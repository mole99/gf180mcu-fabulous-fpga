module gf180mcu_ws_ip__logo_fabulous;
endmodule
