magic
tech gf180mcuD
magscale 1 10
timestamp 1764324262
<< metal1 >>
rect 672 13354 52080 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 52080 13354
rect 672 13268 52080 13302
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 17390 13186 17442 13198
rect 17390 13122 17442 13134
rect 21198 13186 21250 13198
rect 37998 13186 38050 13198
rect 35746 13134 35758 13186
rect 35810 13134 35822 13186
rect 21198 13122 21250 13134
rect 37998 13122 38050 13134
rect 41246 13186 41298 13198
rect 41246 13122 41298 13134
rect 45054 13186 45106 13198
rect 45054 13122 45106 13134
rect 10322 13022 10334 13074
rect 10386 13022 10398 13074
rect 13346 13022 13358 13074
rect 13410 13022 13422 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 15698 13022 15710 13074
rect 15762 13022 15774 13074
rect 22866 13022 22878 13074
rect 22930 13022 22942 13074
rect 37314 13022 37326 13074
rect 37378 13022 37390 13074
rect 43698 13022 43710 13074
rect 43762 13022 43774 13074
rect 35422 12962 35474 12974
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 14130 12910 14142 12962
rect 14194 12910 14206 12962
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 18386 12910 18398 12962
rect 18450 12910 18462 12962
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 39106 12910 39118 12962
rect 39170 12910 39182 12962
rect 40674 12910 40686 12962
rect 40738 12910 40750 12962
rect 42914 12910 42926 12962
rect 42978 12910 42990 12962
rect 44482 12910 44494 12962
rect 44546 12910 44558 12962
rect 47170 12910 47182 12962
rect 47234 12910 47246 12962
rect 48962 12910 48974 12962
rect 49026 12910 49038 12962
rect 50866 12910 50878 12962
rect 50930 12910 50942 12962
rect 35422 12898 35474 12910
rect 24222 12850 24274 12862
rect 19170 12798 19182 12850
rect 19234 12798 19246 12850
rect 24222 12786 24274 12798
rect 36318 12850 36370 12862
rect 38434 12798 38446 12850
rect 38498 12798 38510 12850
rect 39778 12798 39790 12850
rect 39842 12798 39854 12850
rect 51202 12798 51214 12850
rect 51266 12798 51278 12850
rect 36318 12786 36370 12798
rect 48190 12738 48242 12750
rect 48190 12674 48242 12686
rect 49758 12738 49810 12750
rect 49758 12674 49810 12686
rect 672 12570 52080 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 52080 12570
rect 672 12484 52080 12518
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 19854 12402 19906 12414
rect 19854 12338 19906 12350
rect 21646 12402 21698 12414
rect 21646 12338 21698 12350
rect 22878 12402 22930 12414
rect 22878 12338 22930 12350
rect 24334 12402 24386 12414
rect 24334 12338 24386 12350
rect 36542 12402 36594 12414
rect 36542 12338 36594 12350
rect 38110 12402 38162 12414
rect 38110 12338 38162 12350
rect 40014 12402 40066 12414
rect 40014 12338 40066 12350
rect 41582 12402 41634 12414
rect 41582 12338 41634 12350
rect 48078 12402 48130 12414
rect 48078 12338 48130 12350
rect 16718 12290 16770 12302
rect 49646 12290 49698 12302
rect 2706 12238 2718 12290
rect 2770 12238 2782 12290
rect 5842 12238 5854 12290
rect 5906 12238 5918 12290
rect 18050 12238 18062 12290
rect 18114 12238 18126 12290
rect 16718 12226 16770 12238
rect 49646 12226 49698 12238
rect 51214 12290 51266 12302
rect 51214 12226 51266 12238
rect 3166 12178 3218 12190
rect 29374 12178 29426 12190
rect 42590 12178 42642 12190
rect 15362 12126 15374 12178
rect 15426 12126 15438 12178
rect 18946 12126 18958 12178
rect 19010 12126 19022 12178
rect 23762 12126 23774 12178
rect 23826 12126 23838 12178
rect 28578 12126 28590 12178
rect 28642 12126 28654 12178
rect 38994 12126 39006 12178
rect 39058 12126 39070 12178
rect 48738 12126 48750 12178
rect 48802 12126 48814 12178
rect 3166 12114 3218 12126
rect 29374 12114 29426 12126
rect 42590 12114 42642 12126
rect 6750 12066 6802 12078
rect 6750 12002 6802 12014
rect 7646 12066 7698 12078
rect 12798 12066 12850 12078
rect 26686 12066 26738 12078
rect 9874 12014 9886 12066
rect 9938 12014 9950 12066
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 12226 12014 12238 12066
rect 12290 12014 12302 12066
rect 15698 12014 15710 12066
rect 15762 12014 15774 12066
rect 17266 12014 17278 12066
rect 17330 12014 17342 12066
rect 20626 12014 20638 12066
rect 20690 12014 20702 12066
rect 23426 12014 23438 12066
rect 23490 12014 23502 12066
rect 7646 12002 7698 12014
rect 12798 12002 12850 12014
rect 26686 12002 26738 12014
rect 27246 12066 27298 12078
rect 27246 12002 27298 12014
rect 29038 12066 29090 12078
rect 29038 12002 29090 12014
rect 29934 12066 29986 12078
rect 29934 12002 29986 12014
rect 31166 12066 31218 12078
rect 43150 12066 43202 12078
rect 37538 12014 37550 12066
rect 37602 12014 37614 12066
rect 39442 12014 39454 12066
rect 39506 12014 39518 12066
rect 41010 12014 41022 12066
rect 41074 12014 41086 12066
rect 47058 12014 47070 12066
rect 47122 12014 47134 12066
rect 50194 12014 50206 12066
rect 50258 12014 50270 12066
rect 31166 12002 31218 12014
rect 43150 12002 43202 12014
rect 6302 11954 6354 11966
rect 6302 11890 6354 11902
rect 7310 11954 7362 11966
rect 7310 11890 7362 11902
rect 8206 11954 8258 11966
rect 8206 11890 8258 11902
rect 13358 11954 13410 11966
rect 13358 11890 13410 11902
rect 30606 11954 30658 11966
rect 30606 11890 30658 11902
rect 672 11786 52080 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 52080 11786
rect 672 11700 52080 11734
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 14030 11618 14082 11630
rect 14030 11554 14082 11566
rect 23326 11618 23378 11630
rect 23326 11554 23378 11566
rect 25118 11618 25170 11630
rect 25118 11554 25170 11566
rect 38670 11618 38722 11630
rect 38670 11554 38722 11566
rect 40798 11618 40850 11630
rect 40798 11554 40850 11566
rect 42366 11618 42418 11630
rect 42366 11554 42418 11566
rect 6190 11506 6242 11518
rect 28478 11506 28530 11518
rect 13010 11454 13022 11506
rect 13074 11454 13086 11506
rect 18050 11454 18062 11506
rect 18114 11454 18126 11506
rect 18834 11454 18846 11506
rect 18898 11454 18910 11506
rect 21186 11454 21198 11506
rect 21250 11454 21262 11506
rect 21970 11454 21982 11506
rect 22034 11454 22046 11506
rect 6190 11442 6242 11454
rect 28478 11442 28530 11454
rect 27918 11394 27970 11406
rect 5730 11342 5742 11394
rect 5794 11342 5806 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 14578 11342 14590 11394
rect 14642 11342 14654 11394
rect 16146 11342 16158 11394
rect 16210 11342 16222 11394
rect 17266 11342 17278 11394
rect 17330 11342 17342 11394
rect 19730 11342 19742 11394
rect 19794 11342 19806 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 37650 11342 37662 11394
rect 37714 11342 37726 11394
rect 38098 11342 38110 11394
rect 38162 11342 38174 11394
rect 40450 11342 40462 11394
rect 40514 11342 40526 11394
rect 41794 11342 41806 11394
rect 41858 11342 41870 11394
rect 48850 11342 48862 11394
rect 48914 11342 48926 11394
rect 50418 11342 50430 11394
rect 50482 11342 50494 11394
rect 27918 11330 27970 11342
rect 17726 11282 17778 11294
rect 5394 11230 5406 11282
rect 5458 11230 5470 11282
rect 12338 11230 12350 11282
rect 12402 11230 12414 11282
rect 15474 11230 15486 11282
rect 15538 11230 15550 11282
rect 17726 11218 17778 11230
rect 20638 11282 20690 11294
rect 36766 11282 36818 11294
rect 24658 11230 24670 11282
rect 24722 11230 24734 11282
rect 20638 11218 20690 11230
rect 36766 11218 36818 11230
rect 49870 11282 49922 11294
rect 49870 11218 49922 11230
rect 51438 11170 51490 11182
rect 51438 11106 51490 11118
rect 672 11002 52080 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 52080 11002
rect 672 10916 52080 10950
rect 10446 10834 10498 10846
rect 10446 10770 10498 10782
rect 11678 10834 11730 10846
rect 11678 10770 11730 10782
rect 14814 10834 14866 10846
rect 14814 10770 14866 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 18286 10834 18338 10846
rect 18286 10770 18338 10782
rect 19854 10834 19906 10846
rect 19854 10770 19906 10782
rect 21870 10834 21922 10846
rect 21870 10770 21922 10782
rect 23438 10834 23490 10846
rect 23438 10770 23490 10782
rect 37774 10834 37826 10846
rect 37774 10770 37826 10782
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 42478 10834 42530 10846
rect 42478 10770 42530 10782
rect 49646 10722 49698 10734
rect 1698 10670 1710 10722
rect 1762 10670 1774 10722
rect 26786 10670 26798 10722
rect 26850 10670 26862 10722
rect 27682 10670 27694 10722
rect 27746 10670 27758 10722
rect 41122 10670 41134 10722
rect 41186 10670 41198 10722
rect 49646 10658 49698 10670
rect 27246 10610 27298 10622
rect 47742 10610 47794 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 12114 10558 12126 10610
rect 12178 10558 12190 10610
rect 15250 10558 15262 10610
rect 15314 10558 15326 10610
rect 21298 10558 21310 10610
rect 21362 10558 21374 10610
rect 40562 10558 40574 10610
rect 40626 10558 40638 10610
rect 42018 10558 42030 10610
rect 42082 10558 42094 10610
rect 48850 10558 48862 10610
rect 48914 10558 48926 10610
rect 50194 10558 50206 10610
rect 50258 10558 50270 10610
rect 27246 10546 27298 10558
rect 47742 10546 47794 10558
rect 48302 10498 48354 10510
rect 16930 10446 16942 10498
rect 16994 10446 17006 10498
rect 17266 10446 17278 10498
rect 17330 10446 17342 10498
rect 18834 10446 18846 10498
rect 18898 10446 18910 10498
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 37202 10446 37214 10498
rect 37266 10446 37278 10498
rect 38770 10446 38782 10498
rect 38834 10446 38846 10498
rect 50978 10446 50990 10498
rect 51042 10446 51054 10498
rect 48302 10434 48354 10446
rect 2158 10386 2210 10398
rect 2158 10322 2210 10334
rect 26350 10386 26402 10398
rect 26350 10322 26402 10334
rect 672 10218 52080 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 52080 10218
rect 672 10132 52080 10166
rect 10670 10050 10722 10062
rect 10670 9986 10722 9998
rect 12462 10050 12514 10062
rect 12462 9986 12514 9998
rect 14030 10050 14082 10062
rect 14030 9986 14082 9998
rect 15598 10050 15650 10062
rect 15598 9986 15650 9998
rect 17614 10050 17666 10062
rect 17614 9986 17666 9998
rect 19294 10050 19346 10062
rect 19294 9986 19346 9998
rect 22318 10050 22370 10062
rect 36206 10050 36258 10062
rect 27682 9998 27694 10050
rect 27746 9998 27758 10050
rect 22318 9986 22370 9998
rect 36206 9986 36258 9998
rect 40798 10050 40850 10062
rect 40798 9986 40850 9998
rect 43934 10050 43986 10062
rect 43934 9986 43986 9998
rect 8878 9938 8930 9950
rect 24558 9938 24610 9950
rect 21410 9886 21422 9938
rect 21474 9886 21486 9938
rect 8878 9874 8930 9886
rect 24558 9874 24610 9886
rect 25118 9938 25170 9950
rect 39106 9886 39118 9938
rect 39170 9886 39182 9938
rect 50418 9886 50430 9938
rect 50482 9886 50494 9938
rect 25118 9874 25170 9886
rect 9438 9826 9490 9838
rect 26798 9826 26850 9838
rect 12786 9774 12798 9826
rect 12850 9774 12862 9826
rect 14466 9774 14478 9826
rect 14530 9774 14542 9826
rect 16146 9774 16158 9826
rect 16210 9774 16222 9826
rect 17042 9774 17054 9826
rect 17106 9774 17118 9826
rect 19842 9774 19854 9826
rect 19906 9774 19918 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 9438 9762 9490 9774
rect 26798 9762 26850 9774
rect 27358 9826 27410 9838
rect 27358 9762 27410 9774
rect 34526 9826 34578 9838
rect 44830 9826 44882 9838
rect 38322 9774 38334 9826
rect 38386 9774 38398 9826
rect 40338 9774 40350 9826
rect 40402 9774 40414 9826
rect 41906 9774 41918 9826
rect 41970 9774 41982 9826
rect 49074 9774 49086 9826
rect 49138 9774 49150 9826
rect 34526 9762 34578 9774
rect 44830 9762 44882 9774
rect 11230 9714 11282 9726
rect 26238 9714 26290 9726
rect 20514 9662 20526 9714
rect 20578 9662 20590 9714
rect 11230 9650 11282 9662
rect 26238 9650 26290 9662
rect 35086 9714 35138 9726
rect 35086 9650 35138 9662
rect 36766 9714 36818 9726
rect 44494 9714 44546 9726
rect 49870 9714 49922 9726
rect 42242 9662 42254 9714
rect 42306 9662 42318 9714
rect 45266 9662 45278 9714
rect 45330 9662 45342 9714
rect 36766 9650 36818 9662
rect 44494 9650 44546 9662
rect 49870 9650 49922 9662
rect 51438 9602 51490 9614
rect 51438 9538 51490 9550
rect 672 9434 52080 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 52080 9434
rect 672 9348 52080 9382
rect 14814 9266 14866 9278
rect 14814 9202 14866 9214
rect 16382 9266 16434 9278
rect 16382 9202 16434 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 20862 9266 20914 9278
rect 20862 9202 20914 9214
rect 40462 9266 40514 9278
rect 40462 9202 40514 9214
rect 49646 9266 49698 9278
rect 49646 9202 49698 9214
rect 22206 9154 22258 9166
rect 8530 9102 8542 9154
rect 8594 9102 8606 9154
rect 11554 9102 11566 9154
rect 11618 9102 11630 9154
rect 22206 9090 22258 9102
rect 13806 9042 13858 9054
rect 24334 9042 24386 9054
rect 39118 9042 39170 9054
rect 12226 8990 12238 9042
rect 12290 8990 12302 9042
rect 16930 8990 16942 9042
rect 16994 8990 17006 9042
rect 22642 8990 22654 9042
rect 22706 8990 22718 9042
rect 38658 8990 38670 9042
rect 38722 8990 38734 9042
rect 13806 8978 13858 8990
rect 24334 8978 24386 8990
rect 39118 8978 39170 8990
rect 13246 8930 13298 8942
rect 24894 8930 24946 8942
rect 15362 8878 15374 8930
rect 15426 8878 15438 8930
rect 17266 8878 17278 8930
rect 17330 8878 17342 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 21858 8878 21870 8930
rect 21922 8878 21934 8930
rect 13246 8866 13298 8878
rect 24894 8866 24946 8878
rect 25790 8930 25842 8942
rect 48302 8930 48354 8942
rect 39890 8878 39902 8930
rect 39954 8878 39966 8930
rect 48626 8878 48638 8930
rect 48690 8878 48702 8930
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 50978 8878 50990 8930
rect 51042 8878 51054 8930
rect 25790 8866 25842 8878
rect 48302 8866 48354 8878
rect 8990 8818 9042 8830
rect 8990 8754 9042 8766
rect 17838 8818 17890 8830
rect 17838 8754 17890 8766
rect 25230 8818 25282 8830
rect 25230 8754 25282 8766
rect 47742 8818 47794 8830
rect 47742 8754 47794 8766
rect 672 8650 52080 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 52080 8650
rect 672 8564 52080 8598
rect 13022 8482 13074 8494
rect 13022 8418 13074 8430
rect 21534 8482 21586 8494
rect 21534 8418 21586 8430
rect 22430 8482 22482 8494
rect 22430 8418 22482 8430
rect 9326 8370 9378 8382
rect 9326 8306 9378 8318
rect 32398 8370 32450 8382
rect 50418 8318 50430 8370
rect 50482 8318 50494 8370
rect 32398 8306 32450 8318
rect 9886 8258 9938 8270
rect 9886 8194 9938 8206
rect 12462 8258 12514 8270
rect 20974 8258 21026 8270
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 19394 8206 19406 8258
rect 19458 8206 19470 8258
rect 12462 8194 12514 8206
rect 20974 8194 21026 8206
rect 24894 8258 24946 8270
rect 24894 8194 24946 8206
rect 29934 8258 29986 8270
rect 29934 8194 29986 8206
rect 48638 8258 48690 8270
rect 48638 8194 48690 8206
rect 49534 8258 49586 8270
rect 49534 8194 49586 8206
rect 13582 8146 13634 8158
rect 13582 8082 13634 8094
rect 15150 8146 15202 8158
rect 21870 8146 21922 8158
rect 18498 8094 18510 8146
rect 18562 8094 18574 8146
rect 15150 8082 15202 8094
rect 21870 8082 21922 8094
rect 25454 8146 25506 8158
rect 32958 8146 33010 8158
rect 29474 8094 29486 8146
rect 29538 8094 29550 8146
rect 49074 8094 49086 8146
rect 49138 8094 49150 8146
rect 49970 8094 49982 8146
rect 50034 8094 50046 8146
rect 25454 8082 25506 8094
rect 32958 8082 33010 8094
rect 51438 8034 51490 8046
rect 51438 7970 51490 7982
rect 672 7866 52080 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 52080 7866
rect 672 7780 52080 7814
rect 13022 7698 13074 7710
rect 13022 7634 13074 7646
rect 14590 7698 14642 7710
rect 14590 7634 14642 7646
rect 50878 7698 50930 7710
rect 50878 7634 50930 7646
rect 23326 7586 23378 7598
rect 18498 7534 18510 7586
rect 18562 7534 18574 7586
rect 23326 7522 23378 7534
rect 29934 7586 29986 7598
rect 29934 7522 29986 7534
rect 49646 7586 49698 7598
rect 49646 7522 49698 7534
rect 23886 7474 23938 7486
rect 14018 7422 14030 7474
rect 14082 7422 14094 7474
rect 48738 7422 48750 7474
rect 48802 7422 48814 7474
rect 51314 7422 51326 7474
rect 51378 7422 51390 7474
rect 23886 7410 23938 7422
rect 15586 7310 15598 7362
rect 15650 7310 15662 7362
rect 18958 7250 19010 7262
rect 18958 7186 19010 7198
rect 29374 7250 29426 7262
rect 29374 7186 29426 7198
rect 672 7082 52080 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 52080 7082
rect 672 6996 52080 7030
rect 19294 6914 19346 6926
rect 19294 6850 19346 6862
rect 6414 6802 6466 6814
rect 6414 6738 6466 6750
rect 8990 6690 9042 6702
rect 18734 6690 18786 6702
rect 5954 6638 5966 6690
rect 6018 6638 6030 6690
rect 9426 6638 9438 6690
rect 9490 6638 9502 6690
rect 8990 6626 9042 6638
rect 18734 6626 18786 6638
rect 22766 6690 22818 6702
rect 22766 6626 22818 6638
rect 23326 6690 23378 6702
rect 23326 6626 23378 6638
rect 29374 6690 29426 6702
rect 29374 6626 29426 6638
rect 44606 6690 44658 6702
rect 48850 6638 48862 6690
rect 48914 6638 48926 6690
rect 50418 6638 50430 6690
rect 50482 6638 50494 6690
rect 44606 6626 44658 6638
rect 29934 6578 29986 6590
rect 51438 6578 51490 6590
rect 45042 6526 45054 6578
rect 45106 6526 45118 6578
rect 49746 6526 49758 6578
rect 49810 6526 49822 6578
rect 29934 6514 29986 6526
rect 51438 6514 51490 6526
rect 672 6298 52080 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 52080 6298
rect 672 6212 52080 6246
rect 51214 6130 51266 6142
rect 51214 6066 51266 6078
rect 9550 6018 9602 6030
rect 5058 5966 5070 6018
rect 5122 5966 5134 6018
rect 9550 5954 9602 5966
rect 23774 6018 23826 6030
rect 49870 6018 49922 6030
rect 48514 5966 48526 6018
rect 48578 5966 48590 6018
rect 23774 5954 23826 5966
rect 49870 5954 49922 5966
rect 5518 5906 5570 5918
rect 24334 5906 24386 5918
rect 9986 5854 9998 5906
rect 10050 5854 10062 5906
rect 5518 5842 5570 5854
rect 24334 5842 24386 5854
rect 38670 5906 38722 5918
rect 38670 5842 38722 5854
rect 49310 5906 49362 5918
rect 49310 5842 49362 5854
rect 6414 5794 6466 5806
rect 6414 5730 6466 5742
rect 10446 5794 10498 5806
rect 10446 5730 10498 5742
rect 38334 5794 38386 5806
rect 38334 5730 38386 5742
rect 39230 5794 39282 5806
rect 50194 5742 50206 5794
rect 50258 5742 50270 5794
rect 39230 5730 39282 5742
rect 5854 5682 5906 5694
rect 5854 5618 5906 5630
rect 11006 5682 11058 5694
rect 11006 5618 11058 5630
rect 37774 5682 37826 5694
rect 37774 5618 37826 5630
rect 48078 5682 48130 5694
rect 48078 5618 48130 5630
rect 672 5514 52080 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 52080 5514
rect 672 5428 52080 5462
rect 14814 5346 14866 5358
rect 14814 5282 14866 5294
rect 17614 5346 17666 5358
rect 17614 5282 17666 5294
rect 23102 5346 23154 5358
rect 23102 5282 23154 5294
rect 6526 5234 6578 5246
rect 6526 5170 6578 5182
rect 14254 5234 14306 5246
rect 14254 5170 14306 5182
rect 17054 5234 17106 5246
rect 17054 5170 17106 5182
rect 22542 5234 22594 5246
rect 22542 5170 22594 5182
rect 25454 5234 25506 5246
rect 51202 5182 51214 5234
rect 51266 5182 51278 5234
rect 25454 5170 25506 5182
rect 24894 5122 24946 5134
rect 24894 5058 24946 5070
rect 38894 5122 38946 5134
rect 38894 5058 38946 5070
rect 39454 5122 39506 5134
rect 48962 5070 48974 5122
rect 49026 5070 49038 5122
rect 49634 5070 49646 5122
rect 49698 5070 49710 5122
rect 50642 5070 50654 5122
rect 50706 5070 50718 5122
rect 39454 5058 39506 5070
rect 6066 4958 6078 5010
rect 6130 4958 6142 5010
rect 672 4730 52080 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 52080 4730
rect 672 4644 52080 4678
rect 51214 4562 51266 4574
rect 51214 4498 51266 4510
rect 10210 4398 10222 4450
rect 10274 4398 10286 4450
rect 14914 4398 14926 4450
rect 14978 4398 14990 4450
rect 33058 4398 33070 4450
rect 33122 4398 33134 4450
rect 48178 4398 48190 4450
rect 48242 4398 48254 4450
rect 32622 4338 32674 4350
rect 48738 4286 48750 4338
rect 48802 4286 48814 4338
rect 50194 4286 50206 4338
rect 50258 4286 50270 4338
rect 32622 4274 32674 4286
rect 27022 4226 27074 4238
rect 27022 4162 27074 4174
rect 42814 4226 42866 4238
rect 42814 4162 42866 4174
rect 44158 4226 44210 4238
rect 44158 4162 44210 4174
rect 44718 4226 44770 4238
rect 44718 4162 44770 4174
rect 46958 4226 47010 4238
rect 49410 4174 49422 4226
rect 49474 4174 49486 4226
rect 46958 4162 47010 4174
rect 10670 4114 10722 4126
rect 10670 4050 10722 4062
rect 15374 4114 15426 4126
rect 15374 4050 15426 4062
rect 26462 4114 26514 4126
rect 26462 4050 26514 4062
rect 42254 4114 42306 4126
rect 42254 4050 42306 4062
rect 46398 4114 46450 4126
rect 46398 4050 46450 4062
rect 47742 4114 47794 4126
rect 47742 4050 47794 4062
rect 672 3946 52080 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 52080 3946
rect 672 3860 52080 3894
rect 2382 3778 2434 3790
rect 2382 3714 2434 3726
rect 20302 3778 20354 3790
rect 20302 3714 20354 3726
rect 27246 3778 27298 3790
rect 27246 3714 27298 3726
rect 29262 3778 29314 3790
rect 29262 3714 29314 3726
rect 32958 3778 33010 3790
rect 32958 3714 33010 3726
rect 45838 3778 45890 3790
rect 45838 3714 45890 3726
rect 46734 3778 46786 3790
rect 46734 3714 46786 3726
rect 19742 3666 19794 3678
rect 19742 3602 19794 3614
rect 27806 3666 27858 3678
rect 27806 3602 27858 3614
rect 33518 3666 33570 3678
rect 33518 3602 33570 3614
rect 45278 3666 45330 3678
rect 45278 3602 45330 3614
rect 47294 3666 47346 3678
rect 48850 3614 48862 3666
rect 48914 3614 48926 3666
rect 47294 3602 47346 3614
rect 25118 3554 25170 3566
rect 25118 3490 25170 3502
rect 29822 3554 29874 3566
rect 29822 3490 29874 3502
rect 44718 3554 44770 3566
rect 50418 3502 50430 3554
rect 50482 3502 50494 3554
rect 44718 3490 44770 3502
rect 46398 3442 46450 3454
rect 1922 3390 1934 3442
rect 1986 3390 1998 3442
rect 24658 3390 24670 3442
rect 24722 3390 24734 3442
rect 46398 3378 46450 3390
rect 49870 3442 49922 3454
rect 49870 3378 49922 3390
rect 51438 3442 51490 3454
rect 51438 3378 51490 3390
rect 672 3162 52080 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 52080 3162
rect 672 3076 52080 3110
rect 51214 2994 51266 3006
rect 51214 2930 51266 2942
rect 2158 2882 2210 2894
rect 16830 2882 16882 2894
rect 48078 2882 48130 2894
rect 3938 2830 3950 2882
rect 4002 2830 4014 2882
rect 10882 2830 10894 2882
rect 10946 2830 10958 2882
rect 11778 2830 11790 2882
rect 11842 2830 11854 2882
rect 39330 2830 39342 2882
rect 39394 2830 39406 2882
rect 2158 2818 2210 2830
rect 16830 2818 16882 2830
rect 48078 2818 48130 2830
rect 11342 2770 11394 2782
rect 1698 2718 1710 2770
rect 1762 2718 1774 2770
rect 11342 2706 11394 2718
rect 12238 2770 12290 2782
rect 12238 2706 12290 2718
rect 17390 2770 17442 2782
rect 17390 2706 17442 2718
rect 37102 2770 37154 2782
rect 37102 2706 37154 2718
rect 38894 2770 38946 2782
rect 38894 2706 38946 2718
rect 45390 2770 45442 2782
rect 47058 2718 47070 2770
rect 47122 2718 47134 2770
rect 48738 2718 48750 2770
rect 48802 2718 48814 2770
rect 50306 2718 50318 2770
rect 50370 2718 50382 2770
rect 45390 2706 45442 2718
rect 4398 2658 4450 2670
rect 4398 2594 4450 2606
rect 37662 2658 37714 2670
rect 37662 2594 37714 2606
rect 45950 2658 46002 2670
rect 49410 2606 49422 2658
rect 49474 2606 49486 2658
rect 45950 2594 46002 2606
rect 672 2378 52080 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 52080 2378
rect 672 2292 52080 2326
rect 13918 2210 13970 2222
rect 13918 2146 13970 2158
rect 20750 2210 20802 2222
rect 20750 2146 20802 2158
rect 32846 2210 32898 2222
rect 32846 2146 32898 2158
rect 43822 2210 43874 2222
rect 43822 2146 43874 2158
rect 18958 2098 19010 2110
rect 18958 2034 19010 2046
rect 20190 2098 20242 2110
rect 20190 2034 20242 2046
rect 33406 2098 33458 2110
rect 33406 2034 33458 2046
rect 39678 2098 39730 2110
rect 39678 2034 39730 2046
rect 47518 2098 47570 2110
rect 48850 2046 48862 2098
rect 48914 2046 48926 2098
rect 50418 2046 50430 2098
rect 50482 2046 50494 2098
rect 47518 2034 47570 2046
rect 39118 1986 39170 1998
rect 19394 1934 19406 1986
rect 19458 1934 19470 1986
rect 47058 1934 47070 1986
rect 47122 1934 47134 1986
rect 39118 1922 39170 1934
rect 14478 1874 14530 1886
rect 49870 1874 49922 1886
rect 44258 1822 44270 1874
rect 44322 1822 44334 1874
rect 14478 1810 14530 1822
rect 49870 1810 49922 1822
rect 51438 1874 51490 1886
rect 51438 1810 51490 1822
rect 672 1594 52080 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 52080 1594
rect 672 1508 52080 1542
rect 49758 1426 49810 1438
rect 49758 1362 49810 1374
rect 48190 1314 48242 1326
rect 20402 1262 20414 1314
rect 20466 1262 20478 1314
rect 48190 1250 48242 1262
rect 51326 1314 51378 1326
rect 51326 1250 51378 1262
rect 20862 1202 20914 1214
rect 48738 1150 48750 1202
rect 48802 1150 48814 1202
rect 20862 1138 20914 1150
rect 47170 1038 47182 1090
rect 47234 1038 47246 1090
rect 50766 978 50818 990
rect 50766 914 50818 926
rect 672 810 52080 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 52080 810
rect 672 724 52080 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 17390 13134 17442 13186
rect 21198 13134 21250 13186
rect 35758 13134 35810 13186
rect 37998 13134 38050 13186
rect 41246 13134 41298 13186
rect 45054 13134 45106 13186
rect 10334 13022 10386 13074
rect 13358 13022 13410 13074
rect 14926 13022 14978 13074
rect 15710 13022 15762 13074
rect 22878 13022 22930 13074
rect 37326 13022 37378 13074
rect 43710 13022 43762 13074
rect 11902 12910 11954 12962
rect 14142 12910 14194 12962
rect 17838 12910 17890 12962
rect 18398 12910 18450 12962
rect 21758 12910 21810 12962
rect 22094 12910 22146 12962
rect 25006 12910 25058 12962
rect 35422 12910 35474 12962
rect 39118 12910 39170 12962
rect 40686 12910 40738 12962
rect 42926 12910 42978 12962
rect 44494 12910 44546 12962
rect 47182 12910 47234 12962
rect 48974 12910 49026 12962
rect 50878 12910 50930 12962
rect 19182 12798 19234 12850
rect 24222 12798 24274 12850
rect 36318 12798 36370 12850
rect 38446 12798 38498 12850
rect 39790 12798 39842 12850
rect 51214 12798 51266 12850
rect 48190 12686 48242 12738
rect 49758 12686 49810 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 11678 12350 11730 12402
rect 14814 12350 14866 12402
rect 19854 12350 19906 12402
rect 21646 12350 21698 12402
rect 22878 12350 22930 12402
rect 24334 12350 24386 12402
rect 36542 12350 36594 12402
rect 38110 12350 38162 12402
rect 40014 12350 40066 12402
rect 41582 12350 41634 12402
rect 48078 12350 48130 12402
rect 2718 12238 2770 12290
rect 5854 12238 5906 12290
rect 16718 12238 16770 12290
rect 18062 12238 18114 12290
rect 49646 12238 49698 12290
rect 51214 12238 51266 12290
rect 3166 12126 3218 12178
rect 15374 12126 15426 12178
rect 18958 12126 19010 12178
rect 23774 12126 23826 12178
rect 28590 12126 28642 12178
rect 29374 12126 29426 12178
rect 39006 12126 39058 12178
rect 42590 12126 42642 12178
rect 48750 12126 48802 12178
rect 6750 12014 6802 12066
rect 7646 12014 7698 12066
rect 9886 12014 9938 12066
rect 10670 12014 10722 12066
rect 12238 12014 12290 12066
rect 12798 12014 12850 12066
rect 15710 12014 15762 12066
rect 17278 12014 17330 12066
rect 20638 12014 20690 12066
rect 23438 12014 23490 12066
rect 26686 12014 26738 12066
rect 27246 12014 27298 12066
rect 29038 12014 29090 12066
rect 29934 12014 29986 12066
rect 31166 12014 31218 12066
rect 37550 12014 37602 12066
rect 39454 12014 39506 12066
rect 41022 12014 41074 12066
rect 43150 12014 43202 12066
rect 47070 12014 47122 12066
rect 50206 12014 50258 12066
rect 6302 11902 6354 11954
rect 7310 11902 7362 11954
rect 8206 11902 8258 11954
rect 13358 11902 13410 11954
rect 30606 11902 30658 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 10894 11566 10946 11618
rect 14030 11566 14082 11618
rect 23326 11566 23378 11618
rect 25118 11566 25170 11618
rect 38670 11566 38722 11618
rect 40798 11566 40850 11618
rect 42366 11566 42418 11618
rect 6190 11454 6242 11506
rect 13022 11454 13074 11506
rect 18062 11454 18114 11506
rect 18846 11454 18898 11506
rect 21198 11454 21250 11506
rect 21982 11454 22034 11506
rect 28478 11454 28530 11506
rect 5742 11342 5794 11394
rect 6638 11342 6690 11394
rect 11454 11342 11506 11394
rect 14590 11342 14642 11394
rect 16158 11342 16210 11394
rect 17278 11342 17330 11394
rect 19742 11342 19794 11394
rect 22766 11342 22818 11394
rect 27918 11342 27970 11394
rect 37662 11342 37714 11394
rect 38110 11342 38162 11394
rect 40462 11342 40514 11394
rect 41806 11342 41858 11394
rect 48862 11342 48914 11394
rect 50430 11342 50482 11394
rect 5406 11230 5458 11282
rect 12350 11230 12402 11282
rect 15486 11230 15538 11282
rect 17726 11230 17778 11282
rect 20638 11230 20690 11282
rect 24670 11230 24722 11282
rect 36766 11230 36818 11282
rect 49870 11230 49922 11282
rect 51438 11118 51490 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 10446 10782 10498 10834
rect 11678 10782 11730 10834
rect 14814 10782 14866 10834
rect 16382 10782 16434 10834
rect 18286 10782 18338 10834
rect 19854 10782 19906 10834
rect 21870 10782 21922 10834
rect 23438 10782 23490 10834
rect 37774 10782 37826 10834
rect 39342 10782 39394 10834
rect 42478 10782 42530 10834
rect 1710 10670 1762 10722
rect 26798 10670 26850 10722
rect 27694 10670 27746 10722
rect 41134 10670 41186 10722
rect 49646 10670 49698 10722
rect 9550 10558 9602 10610
rect 12126 10558 12178 10610
rect 15262 10558 15314 10610
rect 21310 10558 21362 10610
rect 27246 10558 27298 10610
rect 40574 10558 40626 10610
rect 42030 10558 42082 10610
rect 47742 10558 47794 10610
rect 48862 10558 48914 10610
rect 50206 10558 50258 10610
rect 16942 10446 16994 10498
rect 17278 10446 17330 10498
rect 18846 10446 18898 10498
rect 22878 10446 22930 10498
rect 37214 10446 37266 10498
rect 38782 10446 38834 10498
rect 48302 10446 48354 10498
rect 50990 10446 51042 10498
rect 2158 10334 2210 10386
rect 26350 10334 26402 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 10670 9998 10722 10050
rect 12462 9998 12514 10050
rect 14030 9998 14082 10050
rect 15598 9998 15650 10050
rect 17614 9998 17666 10050
rect 19294 9998 19346 10050
rect 22318 9998 22370 10050
rect 27694 9998 27746 10050
rect 36206 9998 36258 10050
rect 40798 9998 40850 10050
rect 43934 9998 43986 10050
rect 8878 9886 8930 9938
rect 21422 9886 21474 9938
rect 24558 9886 24610 9938
rect 25118 9886 25170 9938
rect 39118 9886 39170 9938
rect 50430 9886 50482 9938
rect 9438 9774 9490 9826
rect 12798 9774 12850 9826
rect 14478 9774 14530 9826
rect 16158 9774 16210 9826
rect 17054 9774 17106 9826
rect 19854 9774 19906 9826
rect 21982 9774 22034 9826
rect 26798 9774 26850 9826
rect 27358 9774 27410 9826
rect 34526 9774 34578 9826
rect 38334 9774 38386 9826
rect 40350 9774 40402 9826
rect 41918 9774 41970 9826
rect 44830 9774 44882 9826
rect 49086 9774 49138 9826
rect 11230 9662 11282 9714
rect 20526 9662 20578 9714
rect 26238 9662 26290 9714
rect 35086 9662 35138 9714
rect 36766 9662 36818 9714
rect 42254 9662 42306 9714
rect 44494 9662 44546 9714
rect 45278 9662 45330 9714
rect 49870 9662 49922 9714
rect 51438 9550 51490 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 14814 9214 14866 9266
rect 16382 9214 16434 9266
rect 19070 9214 19122 9266
rect 20862 9214 20914 9266
rect 40462 9214 40514 9266
rect 49646 9214 49698 9266
rect 8542 9102 8594 9154
rect 11566 9102 11618 9154
rect 22206 9102 22258 9154
rect 12238 8990 12290 9042
rect 13806 8990 13858 9042
rect 16942 8990 16994 9042
rect 22654 8990 22706 9042
rect 24334 8990 24386 9042
rect 38670 8990 38722 9042
rect 39118 8990 39170 9042
rect 13246 8878 13298 8930
rect 15374 8878 15426 8930
rect 17278 8878 17330 8930
rect 20078 8878 20130 8930
rect 21870 8878 21922 8930
rect 24894 8878 24946 8930
rect 25790 8878 25842 8930
rect 39902 8878 39954 8930
rect 48302 8878 48354 8930
rect 48638 8878 48690 8930
rect 50206 8878 50258 8930
rect 50990 8878 51042 8930
rect 8990 8766 9042 8818
rect 17838 8766 17890 8818
rect 25230 8766 25282 8818
rect 47742 8766 47794 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 13022 8430 13074 8482
rect 21534 8430 21586 8482
rect 22430 8430 22482 8482
rect 9326 8318 9378 8370
rect 32398 8318 32450 8370
rect 50430 8318 50482 8370
rect 9886 8206 9938 8258
rect 12462 8206 12514 8258
rect 14590 8206 14642 8258
rect 16158 8206 16210 8258
rect 19406 8206 19458 8258
rect 20974 8206 21026 8258
rect 24894 8206 24946 8258
rect 29934 8206 29986 8258
rect 48638 8206 48690 8258
rect 49534 8206 49586 8258
rect 13582 8094 13634 8146
rect 15150 8094 15202 8146
rect 18510 8094 18562 8146
rect 21870 8094 21922 8146
rect 25454 8094 25506 8146
rect 29486 8094 29538 8146
rect 32958 8094 33010 8146
rect 49086 8094 49138 8146
rect 49982 8094 50034 8146
rect 51438 7982 51490 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 13022 7646 13074 7698
rect 14590 7646 14642 7698
rect 50878 7646 50930 7698
rect 18510 7534 18562 7586
rect 23326 7534 23378 7586
rect 29934 7534 29986 7586
rect 49646 7534 49698 7586
rect 14030 7422 14082 7474
rect 23886 7422 23938 7474
rect 48750 7422 48802 7474
rect 51326 7422 51378 7474
rect 15598 7310 15650 7362
rect 18958 7198 19010 7250
rect 29374 7198 29426 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 19294 6862 19346 6914
rect 6414 6750 6466 6802
rect 5966 6638 6018 6690
rect 8990 6638 9042 6690
rect 9438 6638 9490 6690
rect 18734 6638 18786 6690
rect 22766 6638 22818 6690
rect 23326 6638 23378 6690
rect 29374 6638 29426 6690
rect 44606 6638 44658 6690
rect 48862 6638 48914 6690
rect 50430 6638 50482 6690
rect 29934 6526 29986 6578
rect 45054 6526 45106 6578
rect 49758 6526 49810 6578
rect 51438 6526 51490 6578
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 51214 6078 51266 6130
rect 5070 5966 5122 6018
rect 9550 5966 9602 6018
rect 23774 5966 23826 6018
rect 48526 5966 48578 6018
rect 49870 5966 49922 6018
rect 5518 5854 5570 5906
rect 9998 5854 10050 5906
rect 24334 5854 24386 5906
rect 38670 5854 38722 5906
rect 49310 5854 49362 5906
rect 6414 5742 6466 5794
rect 10446 5742 10498 5794
rect 38334 5742 38386 5794
rect 39230 5742 39282 5794
rect 50206 5742 50258 5794
rect 5854 5630 5906 5682
rect 11006 5630 11058 5682
rect 37774 5630 37826 5682
rect 48078 5630 48130 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 14814 5294 14866 5346
rect 17614 5294 17666 5346
rect 23102 5294 23154 5346
rect 6526 5182 6578 5234
rect 14254 5182 14306 5234
rect 17054 5182 17106 5234
rect 22542 5182 22594 5234
rect 25454 5182 25506 5234
rect 51214 5182 51266 5234
rect 24894 5070 24946 5122
rect 38894 5070 38946 5122
rect 39454 5070 39506 5122
rect 48974 5070 49026 5122
rect 49646 5070 49698 5122
rect 50654 5070 50706 5122
rect 6078 4958 6130 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 51214 4510 51266 4562
rect 10222 4398 10274 4450
rect 14926 4398 14978 4450
rect 33070 4398 33122 4450
rect 48190 4398 48242 4450
rect 32622 4286 32674 4338
rect 48750 4286 48802 4338
rect 50206 4286 50258 4338
rect 27022 4174 27074 4226
rect 42814 4174 42866 4226
rect 44158 4174 44210 4226
rect 44718 4174 44770 4226
rect 46958 4174 47010 4226
rect 49422 4174 49474 4226
rect 10670 4062 10722 4114
rect 15374 4062 15426 4114
rect 26462 4062 26514 4114
rect 42254 4062 42306 4114
rect 46398 4062 46450 4114
rect 47742 4062 47794 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 2382 3726 2434 3778
rect 20302 3726 20354 3778
rect 27246 3726 27298 3778
rect 29262 3726 29314 3778
rect 32958 3726 33010 3778
rect 45838 3726 45890 3778
rect 46734 3726 46786 3778
rect 19742 3614 19794 3666
rect 27806 3614 27858 3666
rect 33518 3614 33570 3666
rect 45278 3614 45330 3666
rect 47294 3614 47346 3666
rect 48862 3614 48914 3666
rect 25118 3502 25170 3554
rect 29822 3502 29874 3554
rect 44718 3502 44770 3554
rect 50430 3502 50482 3554
rect 1934 3390 1986 3442
rect 24670 3390 24722 3442
rect 46398 3390 46450 3442
rect 49870 3390 49922 3442
rect 51438 3390 51490 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 51214 2942 51266 2994
rect 2158 2830 2210 2882
rect 3950 2830 4002 2882
rect 10894 2830 10946 2882
rect 11790 2830 11842 2882
rect 16830 2830 16882 2882
rect 39342 2830 39394 2882
rect 48078 2830 48130 2882
rect 1710 2718 1762 2770
rect 11342 2718 11394 2770
rect 12238 2718 12290 2770
rect 17390 2718 17442 2770
rect 37102 2718 37154 2770
rect 38894 2718 38946 2770
rect 45390 2718 45442 2770
rect 47070 2718 47122 2770
rect 48750 2718 48802 2770
rect 50318 2718 50370 2770
rect 4398 2606 4450 2658
rect 37662 2606 37714 2658
rect 45950 2606 46002 2658
rect 49422 2606 49474 2658
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 13918 2158 13970 2210
rect 20750 2158 20802 2210
rect 32846 2158 32898 2210
rect 43822 2158 43874 2210
rect 18958 2046 19010 2098
rect 20190 2046 20242 2098
rect 33406 2046 33458 2098
rect 39678 2046 39730 2098
rect 47518 2046 47570 2098
rect 48862 2046 48914 2098
rect 50430 2046 50482 2098
rect 19406 1934 19458 1986
rect 39118 1934 39170 1986
rect 47070 1934 47122 1986
rect 14478 1822 14530 1874
rect 44270 1822 44322 1874
rect 49870 1822 49922 1874
rect 51438 1822 51490 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 49758 1374 49810 1426
rect 20414 1262 20466 1314
rect 48190 1262 48242 1314
rect 51326 1262 51378 1314
rect 20862 1150 20914 1202
rect 48750 1150 48802 1202
rect 47182 1038 47234 1090
rect 50766 926 50818 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 12320 14112 12432 14224
rect 12544 14112 12656 14224
rect 12768 14112 12880 14224
rect 12992 14112 13104 14224
rect 13216 14112 13328 14224
rect 13440 14112 13552 14224
rect 13664 14112 13776 14224
rect 13888 14112 14000 14224
rect 14112 14112 14224 14224
rect 14336 14112 14448 14224
rect 14560 14112 14672 14224
rect 14784 14112 14896 14224
rect 15008 14112 15120 14224
rect 15232 14112 15344 14224
rect 15456 14112 15568 14224
rect 15680 14112 15792 14224
rect 15904 14112 16016 14224
rect 16128 14112 16240 14224
rect 16352 14112 16464 14224
rect 16576 14112 16688 14224
rect 16800 14112 16912 14224
rect 17024 14112 17136 14224
rect 17248 14112 17360 14224
rect 17472 14112 17584 14224
rect 17696 14112 17808 14224
rect 17920 14112 18032 14224
rect 18144 14112 18256 14224
rect 18368 14112 18480 14224
rect 18592 14112 18704 14224
rect 18816 14112 18928 14224
rect 19040 14112 19152 14224
rect 19264 14112 19376 14224
rect 19488 14112 19600 14224
rect 19712 14112 19824 14224
rect 19936 14112 20048 14224
rect 20160 14112 20272 14224
rect 20384 14112 20496 14224
rect 20608 14112 20720 14224
rect 20832 14112 20944 14224
rect 21056 14112 21168 14224
rect 21280 14112 21392 14224
rect 21504 14112 21616 14224
rect 21728 14112 21840 14224
rect 21952 14112 22064 14224
rect 22176 14112 22288 14224
rect 22400 14112 22512 14224
rect 22624 14112 22736 14224
rect 22848 14112 22960 14224
rect 23072 14112 23184 14224
rect 23296 14112 23408 14224
rect 23520 14112 23632 14224
rect 23744 14112 23856 14224
rect 23968 14112 24080 14224
rect 24192 14112 24304 14224
rect 24416 14112 24528 14224
rect 24640 14112 24752 14224
rect 24864 14112 24976 14224
rect 25088 14112 25200 14224
rect 25312 14112 25424 14224
rect 25536 14112 25648 14224
rect 25760 14112 25872 14224
rect 25984 14112 26096 14224
rect 26208 14112 26320 14224
rect 26432 14112 26544 14224
rect 26656 14112 26768 14224
rect 26880 14112 26992 14224
rect 27104 14112 27216 14224
rect 27328 14112 27440 14224
rect 27552 14112 27664 14224
rect 27776 14112 27888 14224
rect 28000 14112 28112 14224
rect 28224 14112 28336 14224
rect 28448 14112 28560 14224
rect 28672 14112 28784 14224
rect 28896 14112 29008 14224
rect 29120 14112 29232 14224
rect 29344 14112 29456 14224
rect 29568 14112 29680 14224
rect 29792 14112 29904 14224
rect 30016 14112 30128 14224
rect 30240 14112 30352 14224
rect 30464 14112 30576 14224
rect 30688 14112 30800 14224
rect 30912 14112 31024 14224
rect 31136 14112 31248 14224
rect 31360 14112 31472 14224
rect 31584 14112 31696 14224
rect 31808 14112 31920 14224
rect 32032 14112 32144 14224
rect 32256 14112 32368 14224
rect 32480 14112 32592 14224
rect 32704 14112 32816 14224
rect 32928 14112 33040 14224
rect 33152 14112 33264 14224
rect 33376 14112 33488 14224
rect 33600 14112 33712 14224
rect 33824 14112 33936 14224
rect 34048 14112 34160 14224
rect 34272 14112 34384 14224
rect 34496 14112 34608 14224
rect 34720 14112 34832 14224
rect 34944 14112 35056 14224
rect 35168 14112 35280 14224
rect 35392 14112 35504 14224
rect 35616 14112 35728 14224
rect 35840 14112 35952 14224
rect 36064 14112 36176 14224
rect 36288 14112 36400 14224
rect 36512 14112 36624 14224
rect 36736 14112 36848 14224
rect 36960 14112 37072 14224
rect 37184 14112 37296 14224
rect 37408 14112 37520 14224
rect 37632 14112 37744 14224
rect 37856 14112 37968 14224
rect 38080 14112 38192 14224
rect 38304 14112 38416 14224
rect 38528 14112 38640 14224
rect 38752 14112 38864 14224
rect 38976 14112 39088 14224
rect 39200 14112 39312 14224
rect 39424 14112 39536 14224
rect 39648 14112 39760 14224
rect 39872 14112 39984 14224
rect 40096 14112 40208 14224
rect 44156 14196 44212 14206
rect 11564 14084 11620 14094
rect 140 13972 196 13982
rect 140 7476 196 13916
rect 10332 13972 10388 13982
rect 1260 13524 1316 13534
rect 140 7410 196 7420
rect 364 12180 420 12190
rect 364 6916 420 12124
rect 1260 11172 1316 13468
rect 9772 13524 9828 13534
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 7756 13188 7812 13198
rect 1260 11106 1316 11116
rect 2268 13076 2324 13086
rect 1372 10836 1428 10846
rect 1148 9828 1204 9838
rect 364 6850 420 6860
rect 924 8596 980 8606
rect 924 1204 980 8540
rect 1148 7700 1204 9772
rect 1372 9268 1428 10780
rect 2044 10836 2100 10846
rect 1708 10724 1764 10734
rect 1708 10722 1988 10724
rect 1708 10670 1710 10722
rect 1762 10670 1988 10722
rect 1708 10668 1988 10670
rect 1708 10658 1764 10668
rect 1372 9202 1428 9212
rect 1708 9940 1764 9950
rect 1484 9044 1540 9054
rect 1148 7634 1204 7644
rect 1372 8484 1428 8494
rect 1260 7364 1316 7374
rect 1036 4788 1092 4798
rect 1036 2772 1092 4732
rect 1036 2706 1092 2716
rect 1260 2324 1316 7308
rect 1372 6356 1428 8428
rect 1484 6468 1540 8988
rect 1596 8148 1652 8158
rect 1596 6692 1652 8092
rect 1596 6626 1652 6636
rect 1484 6402 1540 6412
rect 1372 6290 1428 6300
rect 1372 5908 1428 5918
rect 1372 2660 1428 5852
rect 1372 2594 1428 2604
rect 1484 4116 1540 4126
rect 1260 2258 1316 2268
rect 1484 2212 1540 4060
rect 1484 2146 1540 2156
rect 1596 3668 1652 3678
rect 1596 1988 1652 3612
rect 1708 2770 1764 9884
rect 1820 6580 1876 6590
rect 1820 4900 1876 6524
rect 1932 6356 1988 10668
rect 1932 6290 1988 6300
rect 1820 4834 1876 4844
rect 1932 3444 1988 3454
rect 2044 3444 2100 10780
rect 2156 10386 2212 10398
rect 2156 10334 2158 10386
rect 2210 10334 2212 10386
rect 2156 8820 2212 10334
rect 2156 8754 2212 8764
rect 2268 7588 2324 13020
rect 2716 12852 2772 12862
rect 2716 12290 2772 12796
rect 6188 12740 6244 12750
rect 3276 12628 3332 12638
rect 2716 12238 2718 12290
rect 2770 12238 2772 12290
rect 2716 12226 2772 12238
rect 3164 12404 3220 12414
rect 3164 12178 3220 12348
rect 3164 12126 3166 12178
rect 3218 12126 3220 12178
rect 3164 12114 3220 12126
rect 3164 11396 3220 11406
rect 3052 10052 3108 10062
rect 2828 8036 2884 8046
rect 2268 7522 2324 7532
rect 2716 7700 2772 7710
rect 2604 6916 2660 6926
rect 2380 4564 2436 4574
rect 1932 3442 2100 3444
rect 1932 3390 1934 3442
rect 1986 3390 2100 3442
rect 1932 3388 2100 3390
rect 2268 4340 2324 4350
rect 1932 3378 1988 3388
rect 2156 2996 2212 3006
rect 2156 2882 2212 2940
rect 2156 2830 2158 2882
rect 2210 2830 2212 2882
rect 2156 2818 2212 2830
rect 1708 2718 1710 2770
rect 1762 2718 1764 2770
rect 1708 2706 1764 2718
rect 2268 2100 2324 4284
rect 2380 3778 2436 4508
rect 2604 4228 2660 6860
rect 2604 4162 2660 4172
rect 2380 3726 2382 3778
rect 2434 3726 2436 3778
rect 2380 3714 2436 3726
rect 2716 3444 2772 7644
rect 2716 3378 2772 3388
rect 2268 2034 2324 2044
rect 1596 1922 1652 1932
rect 924 1138 980 1148
rect 1484 1876 1540 1886
rect 1484 532 1540 1820
rect 1484 466 1540 476
rect 1596 1428 1652 1438
rect 1596 112 1652 1372
rect 1568 0 1680 112
rect 2828 84 2884 7980
rect 2940 5684 2996 5694
rect 2940 980 2996 5628
rect 3052 4788 3108 9996
rect 3164 9828 3220 11340
rect 3276 10724 3332 12572
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 5852 12290 5908 12302
rect 5852 12238 5854 12290
rect 5906 12238 5908 12290
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 5740 11394 5796 11406
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5404 11282 5460 11294
rect 5404 11230 5406 11282
rect 5458 11230 5460 11282
rect 5292 11172 5348 11182
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3276 10658 3332 10668
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 3164 9762 3220 9772
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3612 6356 3668 6366
rect 3388 5796 3444 5806
rect 3052 4722 3108 4732
rect 3164 5460 3220 5470
rect 3164 2772 3220 5404
rect 3276 4676 3332 4686
rect 3388 4676 3444 5740
rect 3332 4620 3444 4676
rect 3276 4610 3332 4620
rect 3612 4452 3668 6300
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 5068 6018 5124 6030
rect 5068 5966 5070 6018
rect 5122 5966 5124 6018
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4172 4788 4228 4798
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 3612 4386 3668 4396
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3948 2884 4004 2894
rect 3948 2790 4004 2828
rect 3164 2706 3220 2716
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 4172 1428 4228 4732
rect 5068 4116 5124 5966
rect 5068 4050 5124 4060
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 4396 2660 4452 2670
rect 4396 2566 4452 2604
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 2940 914 2996 924
rect 4060 1372 4228 1428
rect 4060 112 4116 1372
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 5292 644 5348 11116
rect 5404 6580 5460 11230
rect 5628 9380 5684 9390
rect 5404 6514 5460 6524
rect 5516 9044 5572 9054
rect 5516 5906 5572 8988
rect 5516 5854 5518 5906
rect 5570 5854 5572 5906
rect 5516 5842 5572 5854
rect 5628 4788 5684 9324
rect 5628 4722 5684 4732
rect 5404 4228 5460 4238
rect 5404 980 5460 4172
rect 5404 914 5460 924
rect 5292 578 5348 588
rect 5740 308 5796 11342
rect 5852 8932 5908 12238
rect 6188 11506 6244 12684
rect 6748 12068 6804 12078
rect 6748 11974 6804 12012
rect 7644 12066 7700 12078
rect 7644 12014 7646 12066
rect 7698 12014 7700 12066
rect 6300 11956 6356 11966
rect 6300 11862 6356 11900
rect 7308 11954 7364 11966
rect 7308 11902 7310 11954
rect 7362 11902 7364 11954
rect 6188 11454 6190 11506
rect 6242 11454 6244 11506
rect 6188 11442 6244 11454
rect 6636 11394 6692 11406
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 5852 8866 5908 8876
rect 6524 11172 6580 11182
rect 6524 7364 6580 11116
rect 6636 8372 6692 11342
rect 6636 8306 6692 8316
rect 6524 7298 6580 7308
rect 6636 7252 6692 7262
rect 6412 7140 6468 7150
rect 6412 6802 6468 7084
rect 6412 6750 6414 6802
rect 6466 6750 6468 6802
rect 6412 6738 6468 6750
rect 5964 6690 6020 6702
rect 5964 6638 5966 6690
rect 6018 6638 6020 6690
rect 5852 5684 5908 5694
rect 5852 5590 5908 5628
rect 5964 1316 6020 6638
rect 6412 5794 6468 5806
rect 6412 5742 6414 5794
rect 6466 5742 6468 5794
rect 6412 5348 6468 5742
rect 6412 5282 6468 5292
rect 6524 5236 6580 5246
rect 6524 5142 6580 5180
rect 6076 5010 6132 5022
rect 6076 4958 6078 5010
rect 6130 4958 6132 5010
rect 6076 3220 6132 4958
rect 6636 3892 6692 7196
rect 6860 6580 6916 6590
rect 6636 3826 6692 3836
rect 6748 6244 6804 6254
rect 6076 3154 6132 3164
rect 6636 3220 6692 3230
rect 5964 1250 6020 1260
rect 6412 2660 6468 2670
rect 6412 1092 6468 2604
rect 6636 2660 6692 3164
rect 6636 2594 6692 2604
rect 6748 1652 6804 6188
rect 6412 1026 6468 1036
rect 6524 1596 6804 1652
rect 5740 242 5796 252
rect 6524 112 6580 1596
rect 6860 868 6916 6524
rect 7308 4004 7364 11902
rect 7308 3938 7364 3948
rect 7532 11956 7588 11966
rect 6860 802 6916 812
rect 7532 532 7588 11900
rect 7644 8596 7700 12014
rect 7644 8530 7700 8540
rect 7756 2884 7812 13132
rect 9772 13186 9828 13468
rect 9772 13134 9774 13186
rect 9826 13134 9828 13186
rect 9772 13122 9828 13134
rect 10332 13074 10388 13916
rect 11340 13636 11396 13646
rect 11340 13186 11396 13580
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 10332 13022 10334 13074
rect 10386 13022 10388 13074
rect 10332 13010 10388 13022
rect 10892 12516 10948 12526
rect 8876 12292 8932 12302
rect 8204 11954 8260 11966
rect 8204 11902 8206 11954
rect 8258 11902 8260 11954
rect 7980 11620 8036 11630
rect 7980 6580 8036 11564
rect 8092 9604 8148 9614
rect 8092 8260 8148 9548
rect 8092 8194 8148 8204
rect 7980 6514 8036 6524
rect 7756 2818 7812 2828
rect 8204 2100 8260 11902
rect 8316 10500 8372 10510
rect 8316 7700 8372 10444
rect 8540 10388 8596 10398
rect 8316 7634 8372 7644
rect 8428 9268 8484 9278
rect 8316 6356 8372 6366
rect 8316 4340 8372 6300
rect 8316 4274 8372 4284
rect 8428 3444 8484 9212
rect 8540 9154 8596 10332
rect 8876 9938 8932 12236
rect 9772 12068 9828 12078
rect 8876 9886 8878 9938
rect 8930 9886 8932 9938
rect 8876 9874 8932 9886
rect 8988 11508 9044 11518
rect 8540 9102 8542 9154
rect 8594 9102 8596 9154
rect 8540 9090 8596 9102
rect 8988 9044 9044 11452
rect 9548 10610 9604 10622
rect 9548 10558 9550 10610
rect 9602 10558 9604 10610
rect 9436 9826 9492 9838
rect 9436 9774 9438 9826
rect 9490 9774 9492 9826
rect 8876 8988 9044 9044
rect 9324 9156 9380 9166
rect 8876 6692 8932 8988
rect 8988 8820 9044 8830
rect 8988 8818 9156 8820
rect 8988 8766 8990 8818
rect 9042 8766 9156 8818
rect 8988 8764 9156 8766
rect 8988 8754 9044 8764
rect 8988 6692 9044 6702
rect 8876 6690 9044 6692
rect 8876 6638 8990 6690
rect 9042 6638 9044 6690
rect 8876 6636 9044 6638
rect 8988 6626 9044 6636
rect 9100 5572 9156 8764
rect 9212 8484 9268 8494
rect 9212 6468 9268 8428
rect 9324 8370 9380 9100
rect 9324 8318 9326 8370
rect 9378 8318 9380 8370
rect 9324 8306 9380 8318
rect 9436 7924 9492 9774
rect 9436 7858 9492 7868
rect 9212 6402 9268 6412
rect 9436 6690 9492 6702
rect 9436 6638 9438 6690
rect 9490 6638 9492 6690
rect 9100 5506 9156 5516
rect 8988 5460 9044 5470
rect 8540 5124 8596 5134
rect 8540 4564 8596 5068
rect 8540 4498 8596 4508
rect 8428 3378 8484 3388
rect 8204 2034 8260 2044
rect 7532 466 7588 476
rect 8988 112 9044 5404
rect 9436 3388 9492 6638
rect 9548 6018 9604 10558
rect 9772 8148 9828 12012
rect 9884 12066 9940 12078
rect 9884 12014 9886 12066
rect 9938 12014 9940 12066
rect 9884 11732 9940 12014
rect 10668 12066 10724 12078
rect 10668 12014 10670 12066
rect 10722 12014 10724 12066
rect 9884 11666 9940 11676
rect 10444 11844 10500 11854
rect 10108 10836 10164 10846
rect 10108 10500 10164 10780
rect 10444 10834 10500 11788
rect 10444 10782 10446 10834
rect 10498 10782 10500 10834
rect 10444 10770 10500 10782
rect 10108 10434 10164 10444
rect 10668 10500 10724 12014
rect 10892 11618 10948 12460
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 11340 11620 11396 11630
rect 10668 10434 10724 10444
rect 10556 10164 10612 10174
rect 10556 9044 10612 10108
rect 10668 10052 10724 10062
rect 10668 9958 10724 9996
rect 10556 8978 10612 8988
rect 11228 9714 11284 9726
rect 11228 9662 11230 9714
rect 11282 9662 11284 9714
rect 9996 8596 10052 8606
rect 9772 8082 9828 8092
rect 9884 8258 9940 8270
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 9884 6468 9940 8206
rect 9996 7812 10052 8540
rect 9996 7746 10052 7756
rect 10332 8596 10388 8606
rect 9884 6402 9940 6412
rect 9548 5966 9550 6018
rect 9602 5966 9604 6018
rect 9548 5954 9604 5966
rect 10220 6020 10276 6030
rect 9996 5906 10052 5918
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9996 3388 10052 5854
rect 10220 4450 10276 5964
rect 10332 5796 10388 8540
rect 10332 5730 10388 5740
rect 10444 5794 10500 5806
rect 10444 5742 10446 5794
rect 10498 5742 10500 5794
rect 10444 5012 10500 5742
rect 11004 5684 11060 5694
rect 11004 5590 11060 5628
rect 10444 4946 10500 4956
rect 10220 4398 10222 4450
rect 10274 4398 10276 4450
rect 10220 4386 10276 4398
rect 9436 3332 9604 3388
rect 9548 1316 9604 3332
rect 9548 1250 9604 1260
rect 9884 3332 10052 3388
rect 10668 4114 10724 4126
rect 10668 4062 10670 4114
rect 10722 4062 10724 4114
rect 9884 756 9940 3332
rect 10220 2436 10276 2446
rect 10108 1876 10164 1886
rect 10108 1652 10164 1820
rect 10108 1586 10164 1596
rect 10220 1204 10276 2380
rect 10668 1540 10724 4062
rect 11228 3780 11284 9662
rect 11228 3714 11284 3724
rect 11340 3388 11396 11564
rect 11452 11394 11508 11406
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 7700 11508 11342
rect 11564 9154 11620 14028
rect 12348 14084 12404 14112
rect 12348 14018 12404 14028
rect 11676 13076 11732 13086
rect 11676 12402 11732 13020
rect 11900 12962 11956 12974
rect 11900 12910 11902 12962
rect 11954 12910 11956 12962
rect 11900 12852 11956 12910
rect 11900 12786 11956 12796
rect 12348 12740 12404 12750
rect 11676 12350 11678 12402
rect 11730 12350 11732 12402
rect 11676 12338 11732 12350
rect 11788 12404 11844 12414
rect 11788 11818 11844 12348
rect 12236 12068 12292 12078
rect 12236 11974 12292 12012
rect 11676 11762 11844 11818
rect 11676 10834 11732 11762
rect 12348 11282 12404 12684
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 11218 12404 11230
rect 12460 11956 12516 11966
rect 11676 10782 11678 10834
rect 11730 10782 11732 10834
rect 11676 10770 11732 10782
rect 12124 10610 12180 10622
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 11788 10388 11844 10398
rect 11788 9828 11844 10332
rect 11788 9762 11844 9772
rect 11564 9102 11566 9154
rect 11618 9102 11620 9154
rect 11564 9090 11620 9102
rect 11788 9604 11844 9614
rect 11452 7634 11508 7644
rect 11676 8708 11732 8718
rect 11676 4676 11732 8652
rect 11788 8372 11844 9548
rect 11788 8306 11844 8316
rect 12124 7364 12180 10558
rect 12460 10050 12516 11900
rect 12572 11844 12628 14112
rect 12796 12292 12852 14112
rect 13020 12516 13076 14112
rect 13020 12450 13076 12460
rect 13244 12404 13300 14112
rect 13356 13300 13412 13310
rect 13356 13074 13412 13244
rect 13356 13022 13358 13074
rect 13410 13022 13412 13074
rect 13356 13010 13412 13022
rect 13244 12338 13300 12348
rect 12796 12236 12964 12292
rect 12572 11778 12628 11788
rect 12796 12066 12852 12078
rect 12796 12014 12798 12066
rect 12850 12014 12852 12066
rect 12796 10612 12852 12014
rect 12796 10546 12852 10556
rect 12460 9998 12462 10050
rect 12514 9998 12516 10050
rect 12460 9986 12516 9998
rect 12796 9826 12852 9838
rect 12796 9774 12798 9826
rect 12850 9774 12852 9826
rect 12236 9044 12292 9054
rect 12236 8950 12292 8988
rect 12460 8260 12516 8270
rect 12460 8166 12516 8204
rect 12124 7298 12180 7308
rect 11676 4610 11732 4620
rect 11788 7140 11844 7150
rect 11788 4340 11844 7084
rect 12236 6804 12292 6814
rect 11900 6692 11956 6702
rect 11900 4900 11956 6636
rect 11900 4834 11956 4844
rect 11788 4274 11844 4284
rect 11340 3332 11508 3388
rect 11340 3220 11396 3230
rect 10892 2884 10948 2894
rect 10892 2790 10948 2828
rect 11340 2770 11396 3164
rect 11340 2718 11342 2770
rect 11394 2718 11396 2770
rect 11340 2706 11396 2718
rect 10668 1474 10724 1484
rect 10220 1138 10276 1148
rect 10444 1204 10500 1214
rect 10444 980 10500 1148
rect 10444 914 10500 924
rect 9884 690 9940 700
rect 11452 112 11508 3332
rect 11788 2996 11844 3006
rect 11788 2882 11844 2940
rect 11788 2830 11790 2882
rect 11842 2830 11844 2882
rect 11788 2818 11844 2830
rect 12236 2770 12292 6748
rect 12796 4564 12852 9774
rect 12908 7700 12964 12236
rect 13020 12180 13076 12190
rect 13020 11506 13076 12124
rect 13020 11454 13022 11506
rect 13074 11454 13076 11506
rect 13020 11442 13076 11454
rect 13356 11954 13412 11966
rect 13356 11902 13358 11954
rect 13410 11902 13412 11954
rect 13244 10948 13300 10958
rect 13244 9604 13300 10892
rect 13020 9548 13300 9604
rect 13020 8482 13076 9548
rect 13020 8430 13022 8482
rect 13074 8430 13076 8482
rect 13020 8418 13076 8430
rect 13244 8930 13300 8942
rect 13244 8878 13246 8930
rect 13298 8878 13300 8930
rect 13020 7700 13076 7710
rect 12908 7698 13076 7700
rect 12908 7646 13022 7698
rect 13074 7646 13076 7698
rect 12908 7644 13076 7646
rect 13020 7634 13076 7644
rect 12796 4498 12852 4508
rect 13020 6916 13076 6926
rect 12236 2718 12238 2770
rect 12290 2718 12292 2770
rect 12236 2706 12292 2718
rect 12796 3332 12852 3342
rect 12796 2212 12852 3276
rect 12796 2146 12852 2156
rect 13020 1988 13076 6860
rect 13020 1922 13076 1932
rect 11788 980 11844 990
rect 11788 644 11844 924
rect 11788 578 11844 588
rect 2828 18 2884 28
rect 4032 0 4144 112
rect 6496 0 6608 112
rect 8960 0 9072 112
rect 11424 0 11536 112
rect 13244 84 13300 8878
rect 13356 2324 13412 11902
rect 13468 8148 13524 14112
rect 13692 11956 13748 14112
rect 13692 11890 13748 11900
rect 13916 11844 13972 14112
rect 14140 13188 14196 14112
rect 14364 13524 14420 14112
rect 14364 13458 14420 13468
rect 14476 13860 14532 13870
rect 14140 13132 14420 13188
rect 14140 12962 14196 12974
rect 14140 12910 14142 12962
rect 14194 12910 14196 12962
rect 13916 11778 13972 11788
rect 14028 11956 14084 11966
rect 14028 11618 14084 11900
rect 14140 11844 14196 12910
rect 14140 11778 14196 11788
rect 14028 11566 14030 11618
rect 14082 11566 14084 11618
rect 14028 11554 14084 11566
rect 13580 11172 13636 11182
rect 13580 9716 13636 11116
rect 13580 9650 13636 9660
rect 13804 10276 13860 10286
rect 13804 9042 13860 10220
rect 14028 10052 14084 10062
rect 14028 9958 14084 9996
rect 13804 8990 13806 9042
rect 13858 8990 13860 9042
rect 13804 8978 13860 8990
rect 13692 8372 13748 8382
rect 13580 8148 13636 8158
rect 13468 8146 13636 8148
rect 13468 8094 13582 8146
rect 13634 8094 13636 8146
rect 13468 8092 13636 8094
rect 13580 8082 13636 8092
rect 13580 7812 13636 7822
rect 13468 5796 13524 5806
rect 13468 2996 13524 5740
rect 13468 2930 13524 2940
rect 13356 2258 13412 2268
rect 13580 644 13636 7756
rect 13692 7476 13748 8316
rect 14364 8218 14420 13132
rect 14476 10164 14532 13804
rect 14588 13076 14644 14112
rect 14588 13010 14644 13020
rect 14812 12740 14868 14112
rect 14924 13524 14980 13534
rect 14924 13074 14980 13468
rect 14924 13022 14926 13074
rect 14978 13022 14980 13074
rect 14924 13010 14980 13022
rect 14812 12674 14868 12684
rect 14812 12404 14868 12414
rect 14812 12310 14868 12348
rect 14812 11732 14868 11742
rect 14588 11394 14644 11406
rect 14588 11342 14590 11394
rect 14642 11342 14644 11394
rect 14588 10388 14644 11342
rect 14812 10834 14868 11676
rect 14812 10782 14814 10834
rect 14866 10782 14868 10834
rect 14812 10770 14868 10782
rect 14924 11172 14980 11182
rect 14588 10322 14644 10332
rect 14476 10098 14532 10108
rect 14476 9826 14532 9838
rect 14476 9774 14478 9826
rect 14530 9774 14532 9826
rect 14476 8372 14532 9774
rect 14812 9268 14868 9278
rect 14812 9174 14868 9212
rect 14476 8306 14532 8316
rect 14588 8260 14644 8270
rect 14588 8258 14756 8260
rect 14364 8162 14532 8218
rect 14588 8206 14590 8258
rect 14642 8206 14756 8258
rect 14588 8204 14756 8206
rect 14588 8194 14644 8204
rect 13692 7410 13748 7420
rect 14028 8148 14084 8158
rect 14028 7474 14084 8092
rect 14476 7700 14532 8162
rect 14588 7700 14644 7710
rect 14476 7698 14644 7700
rect 14476 7646 14590 7698
rect 14642 7646 14644 7698
rect 14476 7644 14644 7646
rect 14588 7634 14644 7644
rect 14028 7422 14030 7474
rect 14082 7422 14084 7474
rect 14028 7410 14084 7422
rect 13804 6580 13860 6590
rect 13692 5908 13748 5918
rect 13692 4004 13748 5852
rect 13692 3938 13748 3948
rect 13804 3556 13860 6524
rect 14252 5236 14308 5246
rect 14252 5142 14308 5180
rect 13804 3490 13860 3500
rect 14476 4004 14532 4014
rect 14476 3444 14532 3948
rect 14476 3378 14532 3388
rect 14700 3444 14756 8204
rect 14812 5348 14868 5358
rect 14924 5348 14980 11116
rect 15036 10164 15092 14112
rect 15260 13300 15316 14112
rect 15148 13244 15316 13300
rect 15148 11732 15204 13244
rect 15260 13076 15316 13086
rect 15260 11956 15316 13020
rect 15372 12852 15428 12862
rect 15372 12178 15428 12796
rect 15484 12740 15540 14112
rect 15708 13636 15764 14112
rect 15708 13570 15764 13580
rect 15708 13412 15764 13422
rect 15708 13074 15764 13356
rect 15708 13022 15710 13074
rect 15762 13022 15764 13074
rect 15708 13010 15764 13022
rect 15932 13076 15988 14112
rect 15932 13010 15988 13020
rect 15484 12684 15876 12740
rect 15372 12126 15374 12178
rect 15426 12126 15428 12178
rect 15372 12114 15428 12126
rect 15484 12292 15540 12302
rect 15260 11890 15316 11900
rect 15148 11676 15428 11732
rect 15260 10610 15316 10622
rect 15260 10558 15262 10610
rect 15314 10558 15316 10610
rect 15036 10098 15092 10108
rect 15148 10164 15204 10174
rect 15148 8146 15204 10108
rect 15260 8820 15316 10558
rect 15372 10052 15428 11676
rect 15484 11282 15540 12236
rect 15708 12066 15764 12078
rect 15708 12014 15710 12066
rect 15762 12014 15764 12066
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15484 11218 15540 11230
rect 15596 11620 15652 11630
rect 15372 9986 15428 9996
rect 15484 10612 15540 10622
rect 15484 9716 15540 10556
rect 15596 10050 15652 11564
rect 15708 11060 15764 12014
rect 15708 10994 15764 11004
rect 15596 9998 15598 10050
rect 15650 9998 15652 10050
rect 15596 9986 15652 9998
rect 15708 10500 15764 10510
rect 15708 10052 15764 10444
rect 15708 9986 15764 9996
rect 15372 9660 15540 9716
rect 15372 9492 15428 9660
rect 15372 9426 15428 9436
rect 15820 9268 15876 12684
rect 16156 11620 16212 14112
rect 16156 11554 16212 11564
rect 16268 13188 16324 13198
rect 16156 11394 16212 11406
rect 16156 11342 16158 11394
rect 16210 11342 16212 11394
rect 16156 11284 16212 11342
rect 16268 11396 16324 13132
rect 16380 11732 16436 14112
rect 16380 11666 16436 11676
rect 16492 12516 16548 12526
rect 16492 11620 16548 12460
rect 16492 11554 16548 11564
rect 16268 11330 16324 11340
rect 16156 11218 16212 11228
rect 16044 11060 16100 11070
rect 15820 9202 15876 9212
rect 15932 10276 15988 10286
rect 15260 8754 15316 8764
rect 15372 8930 15428 8942
rect 15372 8878 15374 8930
rect 15426 8878 15428 8930
rect 15148 8094 15150 8146
rect 15202 8094 15204 8146
rect 15148 8082 15204 8094
rect 15260 8596 15316 8606
rect 15036 7588 15092 7598
rect 15036 7476 15092 7532
rect 15036 7420 15204 7476
rect 15148 6580 15204 7420
rect 15148 6514 15204 6524
rect 14812 5346 14980 5348
rect 14812 5294 14814 5346
rect 14866 5294 14980 5346
rect 14812 5292 14980 5294
rect 15036 5348 15092 5358
rect 14812 5282 14868 5292
rect 14924 4900 14980 4910
rect 14924 4450 14980 4844
rect 14924 4398 14926 4450
rect 14978 4398 14980 4450
rect 14924 4386 14980 4398
rect 15036 4228 15092 5292
rect 15260 5236 15316 8540
rect 15372 7588 15428 8878
rect 15708 8820 15764 8830
rect 15708 8148 15764 8764
rect 15708 8082 15764 8092
rect 15820 8708 15876 8718
rect 15372 7522 15428 7532
rect 15596 7362 15652 7374
rect 15596 7310 15598 7362
rect 15650 7310 15652 7362
rect 15596 5348 15652 7310
rect 15596 5282 15652 5292
rect 15260 5170 15316 5180
rect 15036 4162 15092 4172
rect 15148 4452 15204 4462
rect 14700 3378 14756 3388
rect 15036 3780 15092 3790
rect 13692 3332 13748 3342
rect 13692 2772 13748 3276
rect 13692 2706 13748 2716
rect 13916 3108 13972 3118
rect 13916 2660 13972 3052
rect 13916 2594 13972 2604
rect 13916 2212 13972 2222
rect 13916 2118 13972 2156
rect 13580 578 13636 588
rect 13916 1988 13972 1998
rect 13916 112 13972 1932
rect 14476 1876 14532 1886
rect 15036 1876 15092 3724
rect 15148 2436 15204 4396
rect 15372 4114 15428 4126
rect 15372 4062 15374 4114
rect 15426 4062 15428 4114
rect 15372 3388 15428 4062
rect 15708 3556 15764 3566
rect 15372 3332 15540 3388
rect 15484 2996 15540 3332
rect 15484 2930 15540 2940
rect 15148 2370 15204 2380
rect 15596 2100 15652 2110
rect 15036 1820 15316 1876
rect 14476 1782 14532 1820
rect 15260 420 15316 1820
rect 15596 756 15652 2044
rect 15708 1988 15764 3500
rect 15820 2884 15876 8652
rect 15932 8596 15988 10220
rect 16044 8820 16100 11004
rect 16380 10836 16436 10846
rect 16380 10742 16436 10780
rect 16604 10612 16660 14112
rect 16828 13300 16884 14112
rect 16828 13234 16884 13244
rect 16716 12852 16772 12862
rect 16716 12516 16772 12796
rect 16716 12450 16772 12460
rect 16716 12290 16772 12302
rect 16716 12238 16718 12290
rect 16770 12238 16772 12290
rect 16716 11732 16772 12238
rect 16716 11666 16772 11676
rect 16828 11956 16884 11966
rect 16380 10556 16660 10612
rect 16156 9828 16212 9838
rect 16156 9826 16324 9828
rect 16156 9774 16158 9826
rect 16210 9774 16324 9826
rect 16156 9772 16324 9774
rect 16156 9762 16212 9772
rect 16044 8754 16100 8764
rect 16156 9492 16212 9502
rect 15932 8530 15988 8540
rect 16156 8428 16212 9436
rect 15932 8372 16212 8428
rect 15932 6916 15988 8372
rect 15932 6850 15988 6860
rect 16156 8258 16212 8270
rect 16156 8206 16158 8258
rect 16210 8206 16212 8258
rect 15820 2818 15876 2828
rect 15932 4564 15988 4574
rect 15932 2100 15988 4508
rect 16156 2884 16212 8206
rect 16268 7858 16324 9772
rect 16380 9266 16436 10556
rect 16716 10164 16772 10174
rect 16492 9828 16548 9838
rect 16716 9828 16772 10108
rect 16548 9772 16772 9828
rect 16492 9762 16548 9772
rect 16380 9214 16382 9266
rect 16434 9214 16436 9266
rect 16380 9202 16436 9214
rect 16492 8820 16548 8830
rect 16828 8820 16884 11900
rect 17052 10836 17108 14112
rect 17276 12292 17332 14112
rect 17388 13188 17444 13198
rect 17388 13094 17444 13132
rect 17500 12404 17556 14112
rect 17500 12338 17556 12348
rect 17612 13412 17668 13422
rect 17276 12226 17332 12236
rect 17276 12068 17332 12078
rect 17052 10770 17108 10780
rect 17164 12066 17332 12068
rect 17164 12014 17278 12066
rect 17330 12014 17332 12066
rect 17164 12012 17332 12014
rect 17164 10724 17220 12012
rect 17276 12002 17332 12012
rect 17276 11396 17332 11406
rect 17276 11394 17556 11396
rect 17276 11342 17278 11394
rect 17330 11342 17556 11394
rect 17276 11340 17556 11342
rect 17276 11330 17332 11340
rect 17164 10668 17444 10724
rect 16940 10500 16996 10510
rect 17276 10500 17332 10510
rect 16940 10498 17108 10500
rect 16940 10446 16942 10498
rect 16994 10446 17108 10498
rect 16940 10444 17108 10446
rect 16940 10434 16996 10444
rect 17052 10052 17108 10444
rect 17052 9986 17108 9996
rect 17164 10498 17332 10500
rect 17164 10446 17278 10498
rect 17330 10446 17332 10498
rect 17164 10444 17332 10446
rect 17052 9826 17108 9838
rect 17052 9774 17054 9826
rect 17106 9774 17108 9826
rect 17052 9268 17108 9774
rect 17052 9202 17108 9212
rect 16940 9044 16996 9054
rect 16940 8950 16996 8988
rect 16828 8764 16996 8820
rect 16492 8260 16548 8764
rect 16492 8194 16548 8204
rect 16828 8484 16884 8494
rect 16268 7802 16660 7858
rect 16380 7700 16436 7710
rect 16268 4340 16324 4350
rect 16268 3892 16324 4284
rect 16268 3826 16324 3836
rect 16380 3556 16436 7644
rect 16604 7700 16660 7802
rect 16604 7634 16660 7644
rect 16492 7140 16548 7150
rect 16492 6692 16548 7084
rect 16492 6626 16548 6636
rect 16604 6916 16660 6926
rect 16604 5908 16660 6860
rect 16604 5842 16660 5852
rect 16716 6804 16772 6814
rect 16716 5796 16772 6748
rect 16716 5730 16772 5740
rect 16380 3490 16436 3500
rect 16492 5572 16548 5582
rect 16492 3388 16548 5516
rect 16716 5460 16772 5470
rect 16716 4228 16772 5404
rect 16716 4162 16772 4172
rect 16828 3388 16884 8428
rect 16940 6692 16996 8764
rect 17164 7812 17220 10444
rect 17276 10434 17332 10444
rect 17276 8932 17332 8942
rect 17276 8838 17332 8876
rect 17388 8708 17444 10668
rect 17388 8642 17444 8652
rect 17164 7746 17220 7756
rect 16940 6626 16996 6636
rect 17052 7476 17108 7486
rect 16156 2818 16212 2828
rect 16380 3332 16548 3388
rect 16716 3332 16884 3388
rect 16940 5236 16996 5246
rect 16044 2660 16100 2670
rect 16100 2604 16324 2660
rect 16044 2594 16100 2604
rect 15932 2034 15988 2044
rect 16156 2436 16212 2446
rect 15708 1922 15764 1932
rect 16156 1540 16212 2380
rect 16156 1474 16212 1484
rect 16268 1204 16324 2604
rect 16268 1138 16324 1148
rect 15596 690 15652 700
rect 15820 1092 15876 1102
rect 15820 532 15876 1036
rect 15820 466 15876 476
rect 15260 354 15316 364
rect 16380 112 16436 3332
rect 16492 2772 16548 2782
rect 16492 644 16548 2716
rect 16604 2324 16660 2334
rect 16604 1540 16660 2268
rect 16716 1764 16772 3332
rect 16940 3108 16996 5180
rect 17052 5234 17108 7420
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 16940 3042 16996 3052
rect 17052 4788 17108 4798
rect 16828 2884 16884 2894
rect 16828 2790 16884 2828
rect 16716 1698 16772 1708
rect 16604 1474 16660 1484
rect 17052 1428 17108 4732
rect 17500 4676 17556 11340
rect 17612 10050 17668 13356
rect 17724 11956 17780 14112
rect 17836 12962 17892 12974
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17836 12292 17892 12910
rect 17948 12964 18004 14112
rect 18172 13412 18228 14112
rect 18396 13524 18452 14112
rect 18396 13458 18452 13468
rect 18172 13346 18228 13356
rect 17948 12908 18340 12964
rect 17836 12226 17892 12236
rect 18060 12292 18116 12302
rect 18060 12198 18116 12236
rect 17724 11890 17780 11900
rect 17948 11956 18004 11966
rect 17948 11818 18004 11900
rect 17948 11762 18228 11818
rect 18060 11508 18116 11518
rect 18060 11414 18116 11452
rect 17724 11282 17780 11294
rect 17724 11230 17726 11282
rect 17778 11230 17780 11282
rect 17724 10724 17780 11230
rect 18172 10836 18228 11762
rect 18284 11508 18340 12908
rect 18284 11442 18340 11452
rect 18396 12962 18452 12974
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18284 10836 18340 10846
rect 18172 10834 18340 10836
rect 18172 10782 18286 10834
rect 18338 10782 18340 10834
rect 18172 10780 18340 10782
rect 18284 10770 18340 10780
rect 17724 10658 17780 10668
rect 18396 10612 18452 12910
rect 18620 12964 18676 14112
rect 18620 12898 18676 12908
rect 18844 12516 18900 14112
rect 18732 12460 18900 12516
rect 18620 11956 18676 11966
rect 17612 9998 17614 10050
rect 17666 9998 17668 10050
rect 17612 9986 17668 9998
rect 18060 10556 18452 10612
rect 18508 11508 18564 11518
rect 17724 8932 17780 8942
rect 17724 8820 17780 8876
rect 17948 8932 18004 8942
rect 17836 8820 17892 8830
rect 17724 8818 17892 8820
rect 17724 8766 17838 8818
rect 17890 8766 17892 8818
rect 17724 8764 17892 8766
rect 17836 8754 17892 8764
rect 17724 7700 17780 7710
rect 17612 5908 17668 5918
rect 17612 5346 17668 5852
rect 17612 5294 17614 5346
rect 17666 5294 17668 5346
rect 17612 5282 17668 5294
rect 17500 4610 17556 4620
rect 17724 4340 17780 7644
rect 17948 6244 18004 8876
rect 17948 6178 18004 6188
rect 18060 6020 18116 10556
rect 18172 10388 18228 10398
rect 18228 10332 18452 10388
rect 18172 10322 18228 10332
rect 18284 6804 18340 6814
rect 18396 6804 18452 10332
rect 18508 8146 18564 11452
rect 18620 8820 18676 11900
rect 18732 11732 18788 12460
rect 18732 11666 18788 11676
rect 18956 12178 19012 12190
rect 18956 12126 18958 12178
rect 19010 12126 19012 12178
rect 18844 11508 18900 11518
rect 18844 11414 18900 11452
rect 18844 10498 18900 10510
rect 18844 10446 18846 10498
rect 18898 10446 18900 10498
rect 18844 10276 18900 10446
rect 18844 10210 18900 10220
rect 18620 8754 18676 8764
rect 18508 8094 18510 8146
rect 18562 8094 18564 8146
rect 18508 8082 18564 8094
rect 18508 7700 18564 7710
rect 18508 7586 18564 7644
rect 18508 7534 18510 7586
rect 18562 7534 18564 7586
rect 18508 7522 18564 7534
rect 18956 7476 19012 12126
rect 19068 9266 19124 14112
rect 19180 13524 19236 13534
rect 19180 12850 19236 13468
rect 19180 12798 19182 12850
rect 19234 12798 19236 12850
rect 19180 12786 19236 12798
rect 19068 9214 19070 9266
rect 19122 9214 19124 9266
rect 19068 9202 19124 9214
rect 19180 10276 19236 10286
rect 19180 8932 19236 10220
rect 19292 10050 19348 14112
rect 19292 9998 19294 10050
rect 19346 9998 19348 10050
rect 19292 9986 19348 9998
rect 19404 13748 19460 13758
rect 19404 9828 19460 13692
rect 19516 12292 19572 14112
rect 19516 12226 19572 12236
rect 19628 12068 19684 12078
rect 19180 8866 19236 8876
rect 19292 9772 19460 9828
rect 19516 9828 19572 9838
rect 18844 7420 19012 7476
rect 19180 8708 19236 8718
rect 18396 6748 18564 6804
rect 18060 5954 18116 5964
rect 18172 6356 18228 6366
rect 18172 4676 18228 6300
rect 18172 4610 18228 4620
rect 17724 4274 17780 4284
rect 18284 4116 18340 6748
rect 18396 6356 18452 6366
rect 18396 5908 18452 6300
rect 18508 6020 18564 6748
rect 18732 6692 18788 6702
rect 18732 6598 18788 6636
rect 18508 5954 18564 5964
rect 18396 5842 18452 5852
rect 18732 5908 18788 5918
rect 18396 5684 18452 5694
rect 18396 4564 18452 5628
rect 18396 4498 18452 4508
rect 18508 5348 18564 5358
rect 18284 4050 18340 4060
rect 17052 1362 17108 1372
rect 17164 3780 17220 3790
rect 17164 1316 17220 3724
rect 18508 2996 18564 5292
rect 18732 3220 18788 5852
rect 18844 4900 18900 7420
rect 18844 4834 18900 4844
rect 18956 7250 19012 7262
rect 18956 7198 18958 7250
rect 19010 7198 19012 7250
rect 18956 3388 19012 7198
rect 19180 7140 19236 8652
rect 19180 7074 19236 7084
rect 19292 6914 19348 9772
rect 19404 8258 19460 8270
rect 19404 8206 19406 8258
rect 19458 8206 19460 8258
rect 19404 7140 19460 8206
rect 19404 7074 19460 7084
rect 19292 6862 19294 6914
rect 19346 6862 19348 6914
rect 19292 6850 19348 6862
rect 19404 6692 19460 6702
rect 19292 6356 19348 6366
rect 19180 6244 19236 6254
rect 18956 3332 19124 3388
rect 18732 3154 18788 3164
rect 18956 3220 19012 3230
rect 18956 2996 19012 3164
rect 18508 2940 19012 2996
rect 17388 2772 17444 2782
rect 17388 2678 17444 2716
rect 18620 2212 18676 2222
rect 18620 1428 18676 2156
rect 18956 2100 19012 2110
rect 18956 2006 19012 2044
rect 19068 1764 19124 3332
rect 19068 1698 19124 1708
rect 19180 1540 19236 6188
rect 19292 5348 19348 6300
rect 19292 5282 19348 5292
rect 19404 1986 19460 6636
rect 19516 6356 19572 9772
rect 19628 9716 19684 12012
rect 19740 11620 19796 14112
rect 19852 12740 19908 12750
rect 19852 12402 19908 12684
rect 19852 12350 19854 12402
rect 19906 12350 19908 12402
rect 19852 12338 19908 12350
rect 19740 11564 19908 11620
rect 19628 9650 19684 9660
rect 19740 11394 19796 11406
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19516 6290 19572 6300
rect 19628 8036 19684 8046
rect 19628 2660 19684 7980
rect 19740 3666 19796 11342
rect 19852 10834 19908 11564
rect 19964 11508 20020 14112
rect 20076 13860 20132 13870
rect 20076 12964 20132 13804
rect 20188 13188 20244 14112
rect 20188 13122 20244 13132
rect 20300 13860 20356 13870
rect 20076 12908 20244 12964
rect 20188 12068 20244 12908
rect 20188 12002 20244 12012
rect 19964 11442 20020 11452
rect 20188 11732 20244 11742
rect 20188 11060 20244 11676
rect 20300 11284 20356 13804
rect 20300 11218 20356 11228
rect 20188 11004 20356 11060
rect 19852 10782 19854 10834
rect 19906 10782 19908 10834
rect 19852 10770 19908 10782
rect 20076 10500 20132 10510
rect 20076 9940 20132 10444
rect 20076 9874 20132 9884
rect 20188 10388 20244 10398
rect 19852 9828 19908 9838
rect 19852 9734 19908 9772
rect 19964 9268 20020 9278
rect 19964 8932 20020 9212
rect 20188 9268 20244 10332
rect 20188 9202 20244 9212
rect 20300 9044 20356 11004
rect 20412 9492 20468 14112
rect 20636 12740 20692 14112
rect 20524 12684 20692 12740
rect 20860 12740 20916 14112
rect 20524 9714 20580 12684
rect 20860 12674 20916 12684
rect 21084 12516 21140 14112
rect 21308 13524 21364 14112
rect 21308 13458 21364 13468
rect 21532 13524 21588 14112
rect 21532 13458 21588 13468
rect 21196 13188 21252 13198
rect 21756 13188 21812 14112
rect 21756 13132 21924 13188
rect 21196 13094 21252 13132
rect 21756 12962 21812 12974
rect 21756 12910 21758 12962
rect 21810 12910 21812 12962
rect 21644 12852 21700 12862
rect 21420 12796 21644 12852
rect 20748 12460 21140 12516
rect 21196 12740 21252 12750
rect 20636 12066 20692 12078
rect 20636 12014 20638 12066
rect 20690 12014 20692 12066
rect 20636 11956 20692 12014
rect 20636 11890 20692 11900
rect 20636 11284 20692 11294
rect 20748 11284 20804 12460
rect 21196 11844 21252 12684
rect 20636 11282 20804 11284
rect 20636 11230 20638 11282
rect 20690 11230 20804 11282
rect 20636 11228 20804 11230
rect 20972 11788 21252 11844
rect 20636 11218 20692 11228
rect 20524 9662 20526 9714
rect 20578 9662 20580 9714
rect 20524 9650 20580 9662
rect 20412 9436 20916 9492
rect 20860 9266 20916 9436
rect 20860 9214 20862 9266
rect 20914 9214 20916 9266
rect 20860 9202 20916 9214
rect 20188 8988 20356 9044
rect 19964 8866 20020 8876
rect 20076 8930 20132 8942
rect 20076 8878 20078 8930
rect 20130 8878 20132 8930
rect 20076 8260 20132 8878
rect 20076 8194 20132 8204
rect 20188 8036 20244 8988
rect 20972 8932 21028 11788
rect 21196 11620 21252 11630
rect 21196 11506 21252 11564
rect 21196 11454 21198 11506
rect 21250 11454 21252 11506
rect 21196 11442 21252 11454
rect 21308 11396 21364 11406
rect 21308 10610 21364 11340
rect 21308 10558 21310 10610
rect 21362 10558 21364 10610
rect 21308 10546 21364 10558
rect 21308 10388 21364 10398
rect 20972 8866 21028 8876
rect 21196 8932 21252 8942
rect 20748 8820 20804 8830
rect 20076 7980 20244 8036
rect 20524 8764 20748 8820
rect 19740 3614 19742 3666
rect 19794 3614 19796 3666
rect 19740 3602 19796 3614
rect 19852 6132 19908 6142
rect 19628 2594 19684 2604
rect 19404 1934 19406 1986
rect 19458 1934 19460 1986
rect 19404 1922 19460 1934
rect 19516 2212 19572 2222
rect 19852 2212 19908 6076
rect 20076 5348 20132 7980
rect 20524 6916 20580 8764
rect 20748 8754 20804 8764
rect 20972 8260 21028 8270
rect 20972 8166 21028 8204
rect 20524 6850 20580 6860
rect 20300 5348 20356 5358
rect 20076 5282 20132 5292
rect 20188 5292 20300 5348
rect 20076 4900 20132 4910
rect 20188 4900 20244 5292
rect 20300 5282 20356 5292
rect 20132 4844 20244 4900
rect 20300 4900 20356 4910
rect 20076 4834 20132 4844
rect 19180 1474 19236 1484
rect 18620 1362 18676 1372
rect 17164 1250 17220 1260
rect 16492 578 16548 588
rect 18844 252 19236 308
rect 18844 112 18900 252
rect 13244 18 13300 28
rect 13888 0 14000 112
rect 16352 0 16464 112
rect 18816 0 18928 112
rect 19180 84 19236 252
rect 19516 84 19572 2156
rect 19628 2156 19908 2212
rect 19964 4340 20020 4350
rect 19628 532 19684 2156
rect 19964 2100 20020 4284
rect 20300 3778 20356 4844
rect 20300 3726 20302 3778
rect 20354 3726 20356 3778
rect 20300 3714 20356 3726
rect 21196 3668 21252 8876
rect 21308 5124 21364 10332
rect 21420 9938 21476 12796
rect 21644 12786 21700 12796
rect 21644 12404 21700 12414
rect 21644 12310 21700 12348
rect 21644 12068 21700 12078
rect 21644 11620 21700 12012
rect 21644 11554 21700 11564
rect 21420 9886 21422 9938
rect 21474 9886 21476 9938
rect 21420 9874 21476 9886
rect 21532 11508 21588 11518
rect 21532 8482 21588 11452
rect 21532 8430 21534 8482
rect 21586 8430 21588 8482
rect 21532 8418 21588 8430
rect 21644 9828 21700 9838
rect 21532 7028 21588 7038
rect 21532 6692 21588 6972
rect 21532 6626 21588 6636
rect 21308 5058 21364 5068
rect 21420 6356 21476 6366
rect 20972 3612 21252 3668
rect 21308 4116 21364 4126
rect 21308 3668 21364 4060
rect 20412 3444 20468 3454
rect 20300 3332 20356 3342
rect 20300 2996 20356 3276
rect 20300 2930 20356 2940
rect 19740 2044 20020 2100
rect 20188 2100 20244 2110
rect 19740 1092 19796 2044
rect 20188 2006 20244 2044
rect 19852 1876 19908 1886
rect 19852 1764 19908 1820
rect 19852 1708 20132 1764
rect 19740 1026 19796 1036
rect 19628 466 19684 476
rect 19852 756 19908 766
rect 19852 532 19908 700
rect 20076 756 20132 1708
rect 20412 1314 20468 3388
rect 20972 3108 21028 3612
rect 21308 3602 21364 3612
rect 20972 3042 21028 3052
rect 21084 3444 21140 3454
rect 20748 2996 20804 3006
rect 20748 2210 20804 2940
rect 20748 2158 20750 2210
rect 20802 2158 20804 2210
rect 20748 2146 20804 2158
rect 20524 1988 20580 1998
rect 20524 1764 20580 1932
rect 20524 1698 20580 1708
rect 20860 1988 20916 1998
rect 20412 1262 20414 1314
rect 20466 1262 20468 1314
rect 20412 1250 20468 1262
rect 20076 690 20132 700
rect 20636 1204 20692 1214
rect 19852 466 19908 476
rect 19180 28 19572 84
rect 20636 84 20692 1148
rect 20860 1202 20916 1932
rect 21084 1428 21140 3388
rect 21420 3388 21476 6300
rect 21532 5348 21588 5358
rect 21532 4340 21588 5292
rect 21532 4274 21588 4284
rect 21644 3444 21700 9772
rect 21756 6692 21812 12910
rect 21868 10834 21924 13132
rect 21980 11506 22036 14112
rect 21980 11454 21982 11506
rect 22034 11454 22036 11506
rect 21980 11442 22036 11454
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 21868 10782 21870 10834
rect 21922 10782 21924 10834
rect 21868 10770 21924 10782
rect 21980 10388 22036 10398
rect 22092 10388 22148 12910
rect 22204 12404 22260 14112
rect 22204 12338 22260 12348
rect 22316 13524 22372 13534
rect 22036 10332 22148 10388
rect 22204 10388 22260 10398
rect 21980 10322 22036 10332
rect 21980 9826 22036 9838
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21868 8930 21924 8942
rect 21868 8878 21870 8930
rect 21922 8878 21924 8930
rect 21868 8484 21924 8878
rect 21868 8418 21924 8428
rect 21868 8146 21924 8158
rect 21868 8094 21870 8146
rect 21922 8094 21924 8146
rect 21868 7364 21924 8094
rect 21868 7298 21924 7308
rect 21756 6626 21812 6636
rect 21868 6132 21924 6142
rect 21308 3332 21364 3342
rect 21420 3332 21588 3388
rect 21644 3378 21700 3388
rect 21756 5124 21812 5134
rect 21308 3220 21364 3276
rect 21532 3220 21588 3332
rect 21308 3164 21588 3220
rect 21756 2212 21812 5068
rect 21868 5012 21924 6076
rect 21868 4946 21924 4956
rect 21868 4676 21924 4686
rect 21868 4340 21924 4620
rect 21868 4274 21924 4284
rect 21756 2146 21812 2156
rect 21980 2100 22036 9774
rect 22204 9828 22260 10332
rect 22316 10050 22372 13468
rect 22428 13188 22484 14112
rect 22428 13122 22484 13132
rect 22540 13524 22596 13534
rect 22316 9998 22318 10050
rect 22370 9998 22372 10050
rect 22316 9986 22372 9998
rect 22428 12292 22484 12302
rect 22204 9772 22372 9828
rect 22092 9604 22148 9614
rect 22092 8596 22148 9548
rect 22204 9156 22260 9166
rect 22204 9062 22260 9100
rect 22092 8530 22148 8540
rect 22092 8260 22148 8270
rect 22092 6580 22148 8204
rect 22316 7028 22372 9772
rect 22428 8482 22484 12236
rect 22540 9044 22596 13468
rect 22652 10836 22708 14112
rect 22876 13300 22932 14112
rect 22764 13244 22932 13300
rect 22764 11620 22820 13244
rect 22876 13076 22932 13086
rect 22876 12982 22932 13020
rect 22876 12404 22932 12414
rect 23100 12404 23156 14112
rect 22876 12402 23156 12404
rect 22876 12350 22878 12402
rect 22930 12350 23156 12402
rect 22876 12348 23156 12350
rect 23212 13636 23268 13646
rect 22876 12338 22932 12348
rect 22764 11554 22820 11564
rect 22652 10770 22708 10780
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 10276 22820 11342
rect 22764 10210 22820 10220
rect 22876 10498 22932 10510
rect 22876 10446 22878 10498
rect 22930 10446 22932 10498
rect 22876 10164 22932 10446
rect 22876 10098 22932 10108
rect 22988 9828 23044 9838
rect 22764 9156 22820 9166
rect 22652 9044 22708 9054
rect 22540 9042 22708 9044
rect 22540 8990 22654 9042
rect 22706 8990 22708 9042
rect 22540 8988 22708 8990
rect 22652 8978 22708 8988
rect 22764 8820 22820 9100
rect 22540 8764 22820 8820
rect 22540 8708 22596 8764
rect 22540 8642 22596 8652
rect 22988 8708 23044 9772
rect 22988 8642 23044 8652
rect 23100 9604 23156 9614
rect 22428 8430 22430 8482
rect 22482 8430 22484 8482
rect 22428 8418 22484 8430
rect 22876 8484 22932 8494
rect 22316 6962 22372 6972
rect 22428 7476 22484 7486
rect 22092 6514 22148 6524
rect 22316 6580 22372 6590
rect 22316 6356 22372 6524
rect 22316 6290 22372 6300
rect 22428 3538 22484 7420
rect 22764 6692 22820 6702
rect 22764 6598 22820 6636
rect 22540 5460 22596 5470
rect 22540 5234 22596 5404
rect 22540 5182 22542 5234
rect 22594 5182 22596 5234
rect 22540 5170 22596 5182
rect 21980 2034 22036 2044
rect 22092 3482 22484 3538
rect 21084 1362 21140 1372
rect 21196 1876 21252 1886
rect 20860 1150 20862 1202
rect 20914 1150 20916 1202
rect 20860 1138 20916 1150
rect 21196 980 21252 1820
rect 21756 1876 21812 1886
rect 22092 1876 22148 3482
rect 22876 2212 22932 8428
rect 22988 7140 23044 7150
rect 22988 5012 23044 7084
rect 23100 5346 23156 9548
rect 23100 5294 23102 5346
rect 23154 5294 23156 5346
rect 23100 5282 23156 5294
rect 22988 4946 23044 4956
rect 23212 3388 23268 13580
rect 23324 13076 23380 14112
rect 23324 13010 23380 13020
rect 23548 12404 23604 14112
rect 23548 12338 23604 12348
rect 23660 13300 23716 13310
rect 23660 12180 23716 13244
rect 23772 12852 23828 14112
rect 23996 13748 24052 14112
rect 23996 13682 24052 13692
rect 24220 13076 24276 14112
rect 24444 13636 24500 14112
rect 24444 13570 24500 13580
rect 24668 13524 24724 14112
rect 24892 13860 24948 14112
rect 24892 13794 24948 13804
rect 24668 13458 24724 13468
rect 24892 13524 24948 13534
rect 24332 13412 24388 13422
rect 24332 13188 24388 13356
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24892 13188 24948 13468
rect 24332 13132 24948 13188
rect 24220 13010 24276 13020
rect 25004 12962 25060 12974
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 24220 12852 24276 12862
rect 23772 12850 24276 12852
rect 23772 12798 24222 12850
rect 24274 12798 24276 12850
rect 23772 12796 24276 12798
rect 24220 12786 24276 12796
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 24220 12516 24276 12526
rect 24220 12404 24276 12460
rect 24108 12348 24276 12404
rect 24332 12404 24388 12414
rect 23772 12180 23828 12190
rect 23660 12178 23828 12180
rect 23660 12126 23774 12178
rect 23826 12126 23828 12178
rect 23660 12124 23828 12126
rect 23772 12114 23828 12124
rect 23436 12068 23492 12078
rect 23436 11974 23492 12012
rect 24108 11732 24164 12348
rect 24332 12310 24388 12348
rect 25004 12404 25060 12910
rect 25004 12338 25060 12348
rect 24108 11666 24164 11676
rect 24220 12068 24276 12078
rect 24444 12068 24500 12078
rect 23324 11620 23380 11630
rect 23324 11526 23380 11564
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23436 10836 23492 10846
rect 23436 10742 23492 10780
rect 23324 10724 23380 10734
rect 23324 9828 23380 10668
rect 23548 10724 23604 10734
rect 23548 10612 23604 10668
rect 23324 9762 23380 9772
rect 23436 10556 23604 10612
rect 23436 9492 23492 10556
rect 23436 9426 23492 9436
rect 23548 10388 23604 10398
rect 23548 8428 23604 10332
rect 24220 10052 24276 12012
rect 24332 12012 24444 12068
rect 24332 11844 24388 12012
rect 24444 12002 24500 12012
rect 25116 11844 25172 14112
rect 25340 13972 25396 14112
rect 25564 14084 25620 14112
rect 25564 14018 25620 14028
rect 25340 13916 25508 13972
rect 25340 13748 25396 13758
rect 24332 11778 24388 11788
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 25116 11778 25172 11788
rect 25228 12628 25284 12638
rect 24464 11722 24728 11732
rect 25116 11620 25172 11630
rect 25116 11526 25172 11564
rect 24668 11284 24724 11294
rect 24668 11282 25172 11284
rect 24668 11230 24670 11282
rect 24722 11230 25172 11282
rect 24668 11228 25172 11230
rect 24668 11218 24724 11228
rect 24332 10948 24388 10958
rect 24332 10276 24388 10892
rect 25116 10918 25172 11228
rect 25228 11172 25284 12572
rect 25228 11106 25284 11116
rect 25340 11060 25396 13692
rect 25340 10994 25396 11004
rect 25116 10862 25396 10918
rect 25004 10836 25060 10846
rect 24332 10210 24388 10220
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 24220 9996 24612 10052
rect 24556 9938 24612 9996
rect 24556 9886 24558 9938
rect 24610 9886 24612 9938
rect 24556 9874 24612 9886
rect 24444 9828 24500 9838
rect 23660 9772 24444 9828
rect 23660 9380 23716 9772
rect 24444 9762 24500 9772
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 25004 9380 25060 10780
rect 25340 10836 25396 10862
rect 25340 10770 25396 10780
rect 25228 10724 25284 10734
rect 25116 9940 25172 9950
rect 25116 9846 25172 9884
rect 25228 9716 25284 10668
rect 25452 10164 25508 13916
rect 25788 13860 25844 14112
rect 26012 13972 26068 14112
rect 26012 13916 26180 13972
rect 25564 13804 25844 13860
rect 25564 13636 25620 13804
rect 25788 13636 25844 13646
rect 25564 13580 25788 13636
rect 25788 13570 25844 13580
rect 26124 13524 26180 13916
rect 25900 13468 26180 13524
rect 25452 10098 25508 10108
rect 25676 11508 25732 11518
rect 25676 9828 25732 11452
rect 25900 10948 25956 13468
rect 26236 13412 26292 14112
rect 26124 13356 26292 13412
rect 25900 10882 25956 10892
rect 26012 12516 26068 12526
rect 25676 9762 25732 9772
rect 23660 9314 23716 9324
rect 25004 9314 25060 9324
rect 25116 9660 25284 9716
rect 24332 9268 24388 9278
rect 24332 9042 24388 9212
rect 24332 8990 24334 9042
rect 24386 8990 24388 9042
rect 24332 8978 24388 8990
rect 24892 8932 24948 8942
rect 24892 8930 25060 8932
rect 24892 8878 24894 8930
rect 24946 8878 25060 8930
rect 24892 8876 25060 8878
rect 24892 8866 24948 8876
rect 24108 8764 24836 8820
rect 24108 8708 24164 8764
rect 24780 8758 24836 8764
rect 24780 8708 24948 8758
rect 24780 8702 24892 8708
rect 24108 8642 24164 8652
rect 24464 8652 24728 8662
rect 23436 8372 23604 8428
rect 24332 8596 24388 8606
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24892 8642 24948 8652
rect 24464 8586 24728 8596
rect 23772 8372 23828 8382
rect 23436 7924 23492 8372
rect 23436 7858 23492 7868
rect 23660 8316 23772 8372
rect 23660 7812 23716 8316
rect 23772 8306 23828 8316
rect 24332 7924 24388 8540
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24332 7858 24388 7868
rect 24892 8258 24948 8270
rect 24892 8206 24894 8258
rect 24946 8206 24948 8258
rect 23804 7802 24068 7812
rect 23660 7746 23716 7756
rect 23324 7588 23380 7598
rect 23324 7494 23380 7532
rect 23884 7476 23940 7486
rect 23884 7382 23940 7420
rect 24892 7252 24948 8206
rect 24892 7186 24948 7196
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 25004 6916 25060 8876
rect 25116 8148 25172 9660
rect 25564 9380 25620 9390
rect 25340 9156 25396 9166
rect 25228 8818 25284 8830
rect 25228 8766 25230 8818
rect 25282 8766 25284 8818
rect 25228 8260 25284 8766
rect 25228 8194 25284 8204
rect 25116 8082 25172 8092
rect 25340 7700 25396 9100
rect 25340 7634 25396 7644
rect 25452 8146 25508 8158
rect 25452 8094 25454 8146
rect 25506 8094 25508 8146
rect 25340 7364 25396 7374
rect 25116 6916 25172 6926
rect 25004 6860 25116 6916
rect 25116 6850 25172 6860
rect 23324 6692 23380 6702
rect 23324 6598 23380 6636
rect 23548 6636 24612 6692
rect 23548 6356 23604 6636
rect 24444 6468 24500 6478
rect 23548 6290 23604 6300
rect 23660 6412 24444 6468
rect 23660 6244 23716 6412
rect 24444 6402 24500 6412
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24220 6244 24276 6254
rect 23660 6178 23716 6188
rect 23772 6020 23828 6030
rect 23772 5926 23828 5964
rect 23548 5572 23604 5582
rect 23548 4788 23604 5516
rect 24220 5572 24276 6188
rect 24332 6020 24388 6030
rect 24332 5906 24388 5964
rect 24332 5854 24334 5906
rect 24386 5854 24388 5906
rect 24332 5842 24388 5854
rect 24556 5908 24612 6636
rect 25228 5908 25284 5918
rect 24556 5852 25228 5908
rect 25228 5842 25284 5852
rect 24220 5506 24276 5516
rect 24464 5516 24728 5526
rect 24332 5460 24388 5470
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24892 5460 24948 5470
rect 24332 5348 24388 5404
rect 24892 5348 24948 5404
rect 24332 5292 24948 5348
rect 24892 5124 24948 5134
rect 24892 5030 24948 5068
rect 23548 4722 23604 4732
rect 23804 4732 24068 4742
rect 23436 4676 23492 4686
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24332 4676 24388 4686
rect 22876 2146 22932 2156
rect 23100 3332 23268 3388
rect 23324 4452 23380 4462
rect 23436 4452 23492 4620
rect 23548 4452 23604 4462
rect 23436 4396 23548 4452
rect 21812 1820 22148 1876
rect 21756 1810 21812 1820
rect 22204 1764 22260 1774
rect 21868 1708 22204 1764
rect 21308 1540 21364 1550
rect 21308 1204 21364 1484
rect 21308 1138 21364 1148
rect 21196 914 21252 924
rect 21756 868 21812 878
rect 21868 868 21924 1708
rect 22204 1698 22260 1708
rect 21812 812 21924 868
rect 21980 980 22036 990
rect 21980 868 22036 924
rect 22428 868 22484 878
rect 21980 812 22428 868
rect 21756 802 21812 812
rect 22428 802 22484 812
rect 21084 700 21476 756
rect 21084 644 21140 700
rect 20860 588 21140 644
rect 21420 658 21476 700
rect 21420 602 21588 658
rect 22540 644 22596 654
rect 20860 532 20916 588
rect 21532 532 21588 602
rect 21868 588 22540 644
rect 21532 476 21812 532
rect 20860 466 20916 476
rect 21756 420 21812 476
rect 21868 420 21924 588
rect 22540 578 22596 588
rect 23100 644 23156 3332
rect 23100 578 23156 588
rect 23324 644 23380 4396
rect 23548 4386 23604 4396
rect 24332 4004 24388 4620
rect 25228 4676 25284 4686
rect 24556 4228 24612 4238
rect 24556 4116 24612 4172
rect 24556 4060 25060 4116
rect 25004 4004 25060 4060
rect 25116 4004 25172 4014
rect 24332 3938 24388 3948
rect 24464 3948 24728 3958
rect 25004 3948 25116 4004
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 25116 3938 25172 3948
rect 24464 3882 24728 3892
rect 25228 3780 25284 4620
rect 24668 3724 25284 3780
rect 25340 3780 25396 7308
rect 25452 7028 25508 8094
rect 25452 6962 25508 6972
rect 25452 5236 25508 5246
rect 25564 5236 25620 9324
rect 25788 8930 25844 8942
rect 25788 8878 25790 8930
rect 25842 8878 25844 8930
rect 25452 5234 25620 5236
rect 25452 5182 25454 5234
rect 25506 5182 25620 5234
rect 25452 5180 25620 5182
rect 25676 5236 25732 5246
rect 25452 5170 25508 5180
rect 24556 3444 24612 3454
rect 23660 3276 24276 3332
rect 23660 3108 23716 3276
rect 24220 3220 24276 3276
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24556 3220 24612 3388
rect 24668 3442 24724 3724
rect 25340 3714 25396 3724
rect 24668 3390 24670 3442
rect 24722 3390 24724 3442
rect 24668 3378 24724 3390
rect 25116 3554 25172 3566
rect 25116 3502 25118 3554
rect 25170 3502 25172 3554
rect 25116 3444 25172 3502
rect 25116 3378 25172 3388
rect 24556 3164 25284 3220
rect 24220 3154 24276 3164
rect 23804 3098 24068 3108
rect 24332 3108 24388 3118
rect 23660 3042 23716 3052
rect 23548 2884 23604 2894
rect 23548 1652 23604 2828
rect 24332 2436 24388 3052
rect 24892 2436 24948 2446
rect 24332 2370 24388 2380
rect 24464 2380 24728 2390
rect 23996 2324 24052 2334
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 23996 2212 24052 2268
rect 24892 2212 24948 2380
rect 23996 2156 24948 2212
rect 23548 1586 23604 1596
rect 23804 1596 24068 1606
rect 23660 1540 23716 1550
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 24220 1540 24276 1550
rect 23660 1428 23716 1484
rect 24220 1428 24276 1484
rect 23660 1372 24276 1428
rect 24332 924 24948 980
rect 24332 868 24388 924
rect 24892 868 24948 924
rect 24332 802 24388 812
rect 24464 812 24728 822
rect 24220 756 24276 766
rect 23324 578 23380 588
rect 23548 700 23940 756
rect 21756 364 21924 420
rect 21084 242 21364 298
rect 21084 84 21140 242
rect 21308 112 21364 242
rect 20636 28 21140 84
rect 21280 0 21392 112
rect 23548 84 23604 700
rect 23884 644 23940 700
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24892 802 24948 812
rect 24464 746 24728 756
rect 25228 756 25284 3164
rect 25564 2772 25620 2782
rect 25452 1540 25508 1550
rect 25564 1540 25620 2716
rect 25508 1484 25620 1540
rect 25676 1540 25732 5180
rect 25788 4788 25844 8878
rect 26012 6692 26068 12460
rect 26124 9940 26180 13356
rect 26460 13188 26516 14112
rect 26684 13412 26740 14112
rect 26908 13524 26964 14112
rect 27132 13636 27188 14112
rect 27356 13860 27412 14112
rect 26348 13132 26516 13188
rect 26572 13356 26740 13412
rect 26796 13468 26964 13524
rect 27020 13580 27188 13636
rect 27244 13804 27412 13860
rect 27580 13860 27636 14112
rect 27580 13804 27748 13860
rect 26348 12964 26404 13132
rect 26236 12908 26404 12964
rect 26236 12292 26292 12908
rect 26236 12226 26292 12236
rect 26348 12404 26404 12414
rect 26348 10612 26404 12348
rect 26348 10556 26516 10612
rect 26348 10388 26404 10398
rect 26348 10294 26404 10332
rect 26124 9884 26404 9940
rect 26236 9716 26292 9726
rect 26236 9622 26292 9660
rect 26012 6626 26068 6636
rect 26124 5684 26180 5694
rect 26124 4900 26180 5628
rect 25788 4722 25844 4732
rect 25900 4844 26180 4900
rect 25900 4452 25956 4844
rect 25900 4386 25956 4396
rect 26124 4452 26180 4462
rect 25452 1474 25508 1484
rect 25676 1474 25732 1484
rect 23884 588 24052 644
rect 23660 532 23716 542
rect 23996 532 24052 588
rect 24108 532 24164 542
rect 23716 476 23940 532
rect 23996 476 24108 532
rect 23660 466 23716 476
rect 23884 420 23940 476
rect 24108 466 24164 476
rect 23884 364 24052 420
rect 23772 308 23828 318
rect 23772 112 23828 252
rect 23548 18 23604 28
rect 23744 0 23856 112
rect 23996 84 24052 364
rect 24220 308 24276 700
rect 25228 690 25284 700
rect 24220 242 24276 252
rect 26124 308 26180 4396
rect 26348 1988 26404 9884
rect 26460 7140 26516 10556
rect 26572 8820 26628 13356
rect 26796 13300 26852 13468
rect 27020 13300 27076 13580
rect 26796 13244 26964 13300
rect 27020 13244 27188 13300
rect 26908 13188 26964 13244
rect 26908 13122 26964 13132
rect 27020 12740 27076 12750
rect 26684 12068 26740 12078
rect 27020 12068 27076 12684
rect 26684 12066 27076 12068
rect 26684 12014 26686 12066
rect 26738 12014 27076 12066
rect 26684 12012 27076 12014
rect 26684 12002 26740 12012
rect 26796 10724 26852 10734
rect 26684 10722 26852 10724
rect 26684 10670 26798 10722
rect 26850 10670 26852 10722
rect 26684 10668 26852 10670
rect 26684 10388 26740 10668
rect 26796 10658 26852 10668
rect 26684 10322 26740 10332
rect 26796 10322 27076 10378
rect 26684 10164 26740 10174
rect 26796 10164 26852 10322
rect 26740 10108 26852 10164
rect 26908 10164 26964 10174
rect 26684 10098 26740 10108
rect 26796 9828 26852 9838
rect 26796 9734 26852 9772
rect 26572 8754 26628 8764
rect 26796 8260 26852 8270
rect 26572 8204 26796 8260
rect 26572 8148 26628 8204
rect 26796 8194 26852 8204
rect 26572 8082 26628 8092
rect 26908 8038 26964 10108
rect 27020 8148 27076 10322
rect 27020 8082 27076 8092
rect 26684 7982 26964 8038
rect 26684 7924 26740 7982
rect 26684 7858 26740 7868
rect 26460 7084 26852 7140
rect 26572 6916 26628 6926
rect 26460 4114 26516 4126
rect 26460 4062 26462 4114
rect 26514 4062 26516 4114
rect 26460 2436 26516 4062
rect 26572 3220 26628 6860
rect 26796 6916 26852 7084
rect 26796 6850 26852 6860
rect 27020 4226 27076 4238
rect 27020 4174 27022 4226
rect 27074 4174 27076 4226
rect 27020 3892 27076 4174
rect 27020 3826 27076 3836
rect 27132 3780 27188 13244
rect 27244 12740 27300 13804
rect 27244 12674 27300 12684
rect 27692 12740 27748 13804
rect 27692 12674 27748 12684
rect 27244 12068 27300 12078
rect 27804 12068 27860 14112
rect 27244 12066 27412 12068
rect 27244 12014 27246 12066
rect 27298 12014 27412 12066
rect 27244 12012 27412 12014
rect 27244 12002 27300 12012
rect 27356 11508 27412 12012
rect 27356 11442 27412 11452
rect 27580 12012 27860 12068
rect 27244 10948 27300 10958
rect 27244 10610 27300 10892
rect 27244 10558 27246 10610
rect 27298 10558 27300 10610
rect 27244 10546 27300 10558
rect 27468 10052 27524 10062
rect 27356 9826 27412 9838
rect 27356 9774 27358 9826
rect 27410 9774 27412 9826
rect 27356 8484 27412 9774
rect 27468 9828 27524 9996
rect 27468 9762 27524 9772
rect 27356 8418 27412 8428
rect 27580 7476 27636 12012
rect 27692 11844 27748 11854
rect 27692 11732 27748 11788
rect 28028 11844 28084 14112
rect 28252 12404 28308 14112
rect 28252 12338 28308 12348
rect 28476 12180 28532 14112
rect 28028 11778 28084 11788
rect 28364 12124 28532 12180
rect 28588 12178 28644 12190
rect 28588 12126 28590 12178
rect 28642 12126 28644 12178
rect 27692 11676 27860 11732
rect 27692 10724 27748 10734
rect 27692 10630 27748 10668
rect 27692 10052 27748 10062
rect 27692 9958 27748 9996
rect 27804 9118 27860 11676
rect 27916 11394 27972 11406
rect 27916 11342 27918 11394
rect 27970 11342 27972 11394
rect 27916 9268 27972 11342
rect 28364 9828 28420 12124
rect 28476 11732 28532 11742
rect 28476 11506 28532 11676
rect 28476 11454 28478 11506
rect 28530 11454 28532 11506
rect 28476 11442 28532 11454
rect 28364 9762 28420 9772
rect 27916 9202 27972 9212
rect 27804 9062 27972 9118
rect 27804 8820 27860 8830
rect 27692 8708 27748 8718
rect 27692 8372 27748 8652
rect 27804 8596 27860 8764
rect 27804 8530 27860 8540
rect 27804 8372 27860 8382
rect 27692 8316 27804 8372
rect 27804 8306 27860 8316
rect 27580 7410 27636 7420
rect 27244 6692 27300 6702
rect 27244 4340 27300 6636
rect 27244 4274 27300 4284
rect 27580 6468 27636 6478
rect 27244 3780 27300 3790
rect 27132 3778 27300 3780
rect 27132 3726 27246 3778
rect 27298 3726 27300 3778
rect 27132 3724 27300 3726
rect 27244 3714 27300 3724
rect 27580 3332 27636 6412
rect 27580 3266 27636 3276
rect 27692 5572 27748 5582
rect 26572 3154 26628 3164
rect 26460 2370 26516 2380
rect 26684 2772 26740 2782
rect 26684 2436 26740 2716
rect 26684 2370 26740 2380
rect 26348 1922 26404 1932
rect 26796 2100 26852 2110
rect 26124 242 26180 252
rect 26236 1316 26292 1326
rect 26236 112 26292 1260
rect 26796 196 26852 2044
rect 27692 1988 27748 5516
rect 27804 3668 27860 3678
rect 27916 3668 27972 9062
rect 28476 8036 28532 8046
rect 28588 8036 28644 12126
rect 28700 12180 28756 14112
rect 28924 12628 28980 14112
rect 28924 12562 28980 12572
rect 29036 13188 29092 13198
rect 29036 12358 29092 13132
rect 28924 12302 29092 12358
rect 28700 12124 28868 12180
rect 28700 11956 28756 11966
rect 28700 10164 28756 11900
rect 28700 10098 28756 10108
rect 28532 7980 28644 8036
rect 28476 7970 28532 7980
rect 28812 7364 28868 12124
rect 28924 9716 28980 12302
rect 29036 12066 29092 12078
rect 29036 12014 29038 12066
rect 29090 12014 29092 12066
rect 29036 10388 29092 12014
rect 29036 10322 29092 10332
rect 28924 9650 28980 9660
rect 28812 7298 28868 7308
rect 29036 6804 29092 6814
rect 28476 6580 28532 6590
rect 28028 6244 28084 6254
rect 28028 4228 28084 6188
rect 28476 4564 28532 6524
rect 28476 4498 28532 4508
rect 29036 4564 29092 6748
rect 29148 5796 29204 14112
rect 29372 13972 29428 14112
rect 29372 13916 29540 13972
rect 29260 13860 29316 13870
rect 29260 12180 29316 13804
rect 29372 12180 29428 12190
rect 29260 12178 29428 12180
rect 29260 12126 29374 12178
rect 29426 12126 29428 12178
rect 29260 12124 29428 12126
rect 29372 12114 29428 12124
rect 29484 12068 29540 13916
rect 29484 12002 29540 12012
rect 29596 11620 29652 14112
rect 29820 12404 29876 14112
rect 29596 11554 29652 11564
rect 29708 12348 29876 12404
rect 29148 5730 29204 5740
rect 29260 11060 29316 11070
rect 29036 4498 29092 4508
rect 28028 4162 28084 4172
rect 29260 3778 29316 11004
rect 29708 10724 29764 12348
rect 30044 12292 30100 14112
rect 30268 12628 30324 14112
rect 30268 12562 30324 12572
rect 29372 10668 29764 10724
rect 29820 12236 30100 12292
rect 29372 7924 29428 10668
rect 29820 8820 29876 12236
rect 30380 12180 30436 12190
rect 29932 12068 29988 12078
rect 29932 12066 30324 12068
rect 29932 12014 29934 12066
rect 29986 12014 30324 12066
rect 29932 12012 30324 12014
rect 29932 12002 29988 12012
rect 29820 8754 29876 8764
rect 30044 10164 30100 10174
rect 29932 8260 29988 8270
rect 29932 8166 29988 8204
rect 29484 8148 29540 8158
rect 29484 8054 29540 8092
rect 30044 8036 30100 10108
rect 29932 7980 30100 8036
rect 29372 7868 29540 7924
rect 29372 7250 29428 7262
rect 29372 7198 29374 7250
rect 29426 7198 29428 7250
rect 29372 6916 29428 7198
rect 29372 6850 29428 6860
rect 29372 6690 29428 6702
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 29372 5348 29428 6638
rect 29484 6132 29540 7868
rect 29484 6066 29540 6076
rect 29596 7812 29652 7822
rect 29372 5282 29428 5292
rect 29596 5348 29652 7756
rect 29932 7586 29988 7980
rect 30268 7812 30324 12012
rect 30380 11620 30436 12124
rect 30380 11554 30436 11564
rect 30492 10724 30548 14112
rect 30716 12180 30772 14112
rect 30716 12114 30772 12124
rect 30604 11956 30660 11966
rect 30604 11862 30660 11900
rect 30492 10668 30660 10724
rect 30268 7746 30324 7756
rect 29932 7534 29934 7586
rect 29986 7534 29988 7586
rect 29932 7522 29988 7534
rect 30380 7476 30436 7486
rect 30268 7252 30324 7262
rect 30268 6692 30324 7196
rect 30156 6636 30324 6692
rect 29932 6580 29988 6590
rect 29932 6486 29988 6524
rect 29596 5282 29652 5292
rect 29260 3726 29262 3778
rect 29314 3726 29316 3778
rect 29260 3714 29316 3726
rect 28028 3668 28084 3678
rect 27916 3612 28028 3668
rect 27804 3574 27860 3612
rect 28028 3602 28084 3612
rect 29820 3556 29876 3566
rect 29820 3462 29876 3500
rect 29372 3444 29428 3454
rect 27692 1922 27748 1932
rect 28588 2772 28644 2782
rect 27020 1428 27076 1438
rect 27020 868 27076 1372
rect 28588 1092 28644 2716
rect 28588 1026 28644 1036
rect 28700 1316 28756 1326
rect 27020 802 27076 812
rect 26796 130 26852 140
rect 28700 112 28756 1260
rect 29372 308 29428 3388
rect 30156 2436 30212 6636
rect 30380 4228 30436 7420
rect 30604 6356 30660 10668
rect 30940 7364 30996 14112
rect 31164 12292 31220 14112
rect 31388 13972 31444 14112
rect 31388 13906 31444 13916
rect 31612 13972 31668 14112
rect 31612 13906 31668 13916
rect 31836 13188 31892 14112
rect 31836 13122 31892 13132
rect 31612 12964 31668 12974
rect 31164 12236 31444 12292
rect 31164 12066 31220 12078
rect 31164 12014 31166 12066
rect 31218 12014 31220 12066
rect 31052 11620 31108 11630
rect 31052 11396 31108 11564
rect 31052 11330 31108 11340
rect 31164 10948 31220 12014
rect 31164 10882 31220 10892
rect 31276 11844 31332 11854
rect 31052 10388 31108 10398
rect 31052 7476 31108 10332
rect 31164 9828 31220 9838
rect 31164 9492 31220 9772
rect 31164 9426 31220 9436
rect 31052 7410 31108 7420
rect 31164 8260 31220 8270
rect 30940 7298 30996 7308
rect 30604 6290 30660 6300
rect 30380 4162 30436 4172
rect 30604 5236 30660 5246
rect 30268 4116 30324 4126
rect 30268 2660 30324 4060
rect 30268 2594 30324 2604
rect 30380 3332 30436 3342
rect 30156 2370 30212 2380
rect 30380 1204 30436 3276
rect 30492 2660 30548 2670
rect 30492 2324 30548 2604
rect 30492 2258 30548 2268
rect 30380 1138 30436 1148
rect 30268 980 30324 990
rect 30268 420 30324 924
rect 30268 354 30324 364
rect 29372 242 29428 252
rect 24444 84 24500 94
rect 23996 28 24444 84
rect 24444 18 24500 28
rect 26208 0 26320 112
rect 28672 0 28784 112
rect 30492 84 30548 94
rect 30604 84 30660 5180
rect 31164 112 31220 8204
rect 31276 1204 31332 11788
rect 31388 11620 31444 12236
rect 31388 11554 31444 11564
rect 31388 10388 31444 10398
rect 31388 9268 31444 10332
rect 31612 10164 31668 12908
rect 31948 12740 32004 12750
rect 31948 12292 32004 12684
rect 32060 12292 32116 14112
rect 32284 13748 32340 14112
rect 32284 13682 32340 13692
rect 32060 12236 32340 12292
rect 31948 12226 32004 12236
rect 32172 12068 32228 12078
rect 31612 10108 32004 10164
rect 31388 9212 31556 9268
rect 31500 6916 31556 9212
rect 31948 9156 32004 10108
rect 31948 9100 32116 9156
rect 31948 8820 32004 8830
rect 31500 6850 31556 6860
rect 31724 8484 31780 8494
rect 31724 6020 31780 8428
rect 31724 5954 31780 5964
rect 31836 6692 31892 6702
rect 31836 5908 31892 6636
rect 31836 5842 31892 5852
rect 31948 5684 32004 8764
rect 32060 8484 32116 9100
rect 32172 8708 32228 12012
rect 32284 9156 32340 12236
rect 32508 10388 32564 14112
rect 32732 10612 32788 14112
rect 32956 11788 33012 14112
rect 32732 10546 32788 10556
rect 32844 11732 33012 11788
rect 32508 10322 32564 10332
rect 32284 9100 32676 9156
rect 32172 8642 32228 8652
rect 32060 8418 32116 8428
rect 32396 8372 32452 8382
rect 32396 8278 32452 8316
rect 32060 7924 32116 7934
rect 32060 6916 32116 7868
rect 32060 6850 32116 6860
rect 32284 7812 32340 7822
rect 31836 5628 32004 5684
rect 31836 2996 31892 5628
rect 32172 4452 32228 4462
rect 32172 3220 32228 4396
rect 32172 3154 32228 3164
rect 31836 2930 31892 2940
rect 32284 2212 32340 7756
rect 32620 4338 32676 9100
rect 32732 7924 32788 7934
rect 32732 7140 32788 7868
rect 32732 7074 32788 7084
rect 32844 5684 32900 11732
rect 33068 11396 33124 11406
rect 33068 10612 33124 11340
rect 33068 10546 33124 10556
rect 32956 8146 33012 8158
rect 32956 8094 32958 8146
rect 33010 8094 33012 8146
rect 32956 8036 33012 8094
rect 32956 7970 33012 7980
rect 33180 7588 33236 14112
rect 33292 13412 33348 13422
rect 33292 11060 33348 13356
rect 33404 12516 33460 14112
rect 33628 13524 33684 14112
rect 33404 12450 33460 12460
rect 33516 13468 33684 13524
rect 33516 11284 33572 13468
rect 33628 13300 33684 13310
rect 33628 11732 33684 13244
rect 33628 11666 33684 11676
rect 33516 11218 33572 11228
rect 33628 11396 33684 11406
rect 33292 11004 33572 11060
rect 33180 7522 33236 7532
rect 33404 8484 33460 8494
rect 33516 8484 33572 11004
rect 33628 9268 33684 11340
rect 33852 11172 33908 14112
rect 33852 11106 33908 11116
rect 33964 13860 34020 13870
rect 33628 9202 33684 9212
rect 33852 10276 33908 10286
rect 33628 8484 33684 8494
rect 33516 8428 33628 8484
rect 33404 7588 33460 8428
rect 33628 8418 33684 8428
rect 33628 8260 33684 8270
rect 33404 7522 33460 7532
rect 33516 7812 33572 7822
rect 33516 6356 33572 7756
rect 33628 6580 33684 8204
rect 33852 7812 33908 10220
rect 33964 9044 34020 13804
rect 34076 11620 34132 14112
rect 34076 11554 34132 11564
rect 33964 8978 34020 8988
rect 34076 9268 34132 9278
rect 33852 7746 33908 7756
rect 33628 6514 33684 6524
rect 33852 7588 33908 7598
rect 33852 6580 33908 7532
rect 33852 6514 33908 6524
rect 33516 6300 33684 6356
rect 32844 5618 32900 5628
rect 33404 5684 33460 5694
rect 33068 4564 33124 4574
rect 33068 4450 33124 4508
rect 33068 4398 33070 4450
rect 33122 4398 33124 4450
rect 33068 4386 33124 4398
rect 32620 4286 32622 4338
rect 32674 4286 32676 4338
rect 32620 4274 32676 4286
rect 33180 4340 33236 4350
rect 32956 4228 33012 4238
rect 32956 3778 33012 4172
rect 32956 3726 32958 3778
rect 33010 3726 33012 3778
rect 32956 3714 33012 3726
rect 32284 2146 32340 2156
rect 32396 3220 32452 3230
rect 32396 1540 32452 3164
rect 32844 2548 32900 2558
rect 32844 2210 32900 2492
rect 33180 2436 33236 4284
rect 33404 2884 33460 5628
rect 33516 3668 33572 3678
rect 33516 3574 33572 3612
rect 33404 2818 33460 2828
rect 33180 2370 33236 2380
rect 33404 2548 33460 2558
rect 32844 2158 32846 2210
rect 32898 2158 32900 2210
rect 32844 2146 32900 2158
rect 33404 2098 33460 2492
rect 33404 2046 33406 2098
rect 33458 2046 33460 2098
rect 33404 2034 33460 2046
rect 32396 1474 32452 1484
rect 31276 1138 31332 1148
rect 33628 980 33684 6300
rect 34076 5572 34132 9212
rect 34300 8820 34356 14112
rect 34524 12068 34580 14112
rect 34524 12002 34580 12012
rect 34412 11956 34468 11966
rect 34412 10164 34468 11900
rect 34412 10098 34468 10108
rect 34636 10164 34692 10174
rect 34300 8754 34356 8764
rect 34524 9826 34580 9838
rect 34524 9774 34526 9826
rect 34578 9774 34580 9826
rect 34524 6244 34580 9774
rect 34636 7140 34692 10108
rect 34636 7074 34692 7084
rect 34524 6178 34580 6188
rect 34748 6132 34804 14112
rect 34972 11788 35028 14112
rect 35196 13860 35252 14112
rect 35196 13794 35252 13804
rect 35420 13188 35476 14112
rect 35644 13188 35700 14112
rect 35756 13188 35812 13198
rect 35420 13132 35588 13188
rect 35644 13186 35812 13188
rect 35644 13134 35758 13186
rect 35810 13134 35812 13186
rect 35644 13132 35812 13134
rect 35420 12962 35476 12974
rect 35420 12910 35422 12962
rect 35474 12910 35476 12962
rect 34860 11732 35028 11788
rect 35308 11844 35364 11854
rect 34860 10724 34916 11732
rect 34860 10658 34916 10668
rect 34972 10948 35028 10958
rect 34972 9492 35028 10892
rect 35308 10724 35364 11788
rect 35308 10658 35364 10668
rect 35420 10052 35476 12910
rect 35532 11844 35588 13132
rect 35756 13122 35812 13132
rect 35868 12852 35924 14112
rect 36092 13076 36148 14112
rect 36316 13076 36372 14112
rect 36540 13300 36596 14112
rect 36764 13412 36820 14112
rect 36764 13346 36820 13356
rect 36540 13234 36596 13244
rect 36540 13076 36596 13086
rect 36316 13020 36484 13076
rect 36092 13010 36148 13020
rect 36316 12852 36372 12862
rect 35868 12850 36372 12852
rect 35868 12798 36318 12850
rect 36370 12798 36372 12850
rect 35868 12796 36372 12798
rect 36316 12786 36372 12796
rect 35532 11778 35588 11788
rect 35644 12628 35700 12638
rect 35644 11620 35700 12572
rect 36316 12404 36372 12414
rect 35644 11554 35700 11564
rect 35756 12292 35812 12302
rect 35420 9986 35476 9996
rect 34972 9426 35028 9436
rect 35084 9714 35140 9726
rect 35084 9662 35086 9714
rect 35138 9662 35140 9714
rect 35084 8820 35140 9662
rect 35084 8754 35140 8764
rect 35308 9604 35364 9614
rect 35308 7140 35364 9548
rect 35420 8596 35476 8606
rect 35420 7588 35476 8540
rect 35420 7522 35476 7532
rect 35308 7074 35364 7084
rect 35308 6916 35364 6926
rect 34748 6066 34804 6076
rect 35084 6244 35140 6254
rect 34076 5506 34132 5516
rect 33628 914 33684 924
rect 34524 2884 34580 2894
rect 34524 532 34580 2828
rect 35084 1428 35140 6188
rect 35308 4564 35364 6860
rect 35308 4498 35364 4508
rect 35756 4228 35812 12236
rect 36204 10836 36260 10846
rect 36204 10050 36260 10780
rect 36204 9998 36206 10050
rect 36258 9998 36260 10050
rect 36204 9986 36260 9998
rect 36316 7588 36372 12348
rect 36428 11284 36484 13020
rect 36540 12402 36596 13020
rect 36540 12350 36542 12402
rect 36594 12350 36596 12402
rect 36540 12338 36596 12350
rect 36876 12740 36932 12750
rect 36764 11284 36820 11294
rect 36428 11282 36820 11284
rect 36428 11230 36766 11282
rect 36818 11230 36820 11282
rect 36428 11228 36820 11230
rect 36764 11218 36820 11228
rect 36876 11060 36932 12684
rect 36988 12292 37044 14112
rect 37212 12740 37268 14112
rect 37436 13748 37492 14112
rect 37436 13682 37492 13692
rect 37324 13636 37380 13646
rect 37324 13074 37380 13580
rect 37660 13524 37716 14112
rect 37660 13458 37716 13468
rect 37324 13022 37326 13074
rect 37378 13022 37380 13074
rect 37324 13010 37380 13022
rect 37212 12674 37268 12684
rect 37884 12404 37940 14112
rect 37996 13860 38052 13870
rect 37996 13186 38052 13804
rect 38108 13524 38164 14112
rect 38108 13468 38276 13524
rect 37996 13134 37998 13186
rect 38050 13134 38052 13186
rect 37996 13122 38052 13134
rect 38108 13300 38164 13310
rect 37884 12338 37940 12348
rect 38108 12402 38164 13244
rect 38108 12350 38110 12402
rect 38162 12350 38164 12402
rect 38108 12338 38164 12350
rect 36988 12236 37828 12292
rect 37548 12068 37604 12078
rect 37548 11974 37604 12012
rect 36876 10994 36932 11004
rect 37100 11844 37156 11854
rect 36764 9714 36820 9726
rect 36764 9662 36766 9714
rect 36818 9662 36820 9714
rect 36764 8484 36820 9662
rect 36764 8418 36820 8428
rect 36988 8932 37044 8942
rect 36988 8372 37044 8876
rect 36988 8306 37044 8316
rect 36316 7532 36820 7588
rect 35756 4162 35812 4172
rect 36092 6580 36148 6590
rect 35532 2436 35588 2446
rect 35420 2100 35476 2110
rect 35420 1652 35476 2044
rect 35420 1586 35476 1596
rect 35084 1362 35140 1372
rect 35532 644 35588 2380
rect 35532 578 35588 588
rect 34524 466 34580 476
rect 33628 196 33684 206
rect 33628 112 33684 140
rect 36092 112 36148 6524
rect 36652 3332 36708 3342
rect 36652 2772 36708 3276
rect 36652 2706 36708 2716
rect 36764 196 36820 7532
rect 36988 6804 37044 6814
rect 36988 6356 37044 6748
rect 36988 6290 37044 6300
rect 36988 6132 37044 6142
rect 36876 5572 36932 5582
rect 36876 756 36932 5516
rect 36988 4676 37044 6076
rect 36988 4610 37044 4620
rect 37100 2770 37156 11788
rect 37324 11844 37380 11854
rect 37212 10498 37268 10510
rect 37212 10446 37214 10498
rect 37266 10446 37268 10498
rect 37212 8260 37268 10446
rect 37324 9268 37380 11788
rect 37548 11620 37604 11630
rect 37324 9202 37380 9212
rect 37436 11172 37492 11182
rect 37212 8194 37268 8204
rect 37324 6580 37380 6590
rect 37324 5012 37380 6524
rect 37324 4946 37380 4956
rect 37212 4788 37268 4798
rect 37212 2884 37268 4732
rect 37436 3668 37492 11116
rect 37548 6244 37604 11564
rect 37548 6178 37604 6188
rect 37660 11394 37716 11406
rect 37660 11342 37662 11394
rect 37714 11342 37716 11394
rect 37436 3602 37492 3612
rect 37660 2996 37716 11342
rect 37772 10834 37828 12236
rect 37772 10782 37774 10834
rect 37826 10782 37828 10834
rect 37772 10770 37828 10782
rect 37884 12180 37940 12190
rect 37884 10612 37940 12124
rect 38108 11396 38164 11406
rect 38108 11302 38164 11340
rect 37884 10546 37940 10556
rect 37996 11284 38052 11294
rect 37772 5684 37828 5694
rect 37772 5590 37828 5628
rect 37660 2930 37716 2940
rect 37884 5236 37940 5246
rect 37212 2818 37268 2828
rect 37100 2718 37102 2770
rect 37154 2718 37156 2770
rect 37100 2706 37156 2718
rect 37660 2660 37716 2670
rect 37660 2566 37716 2604
rect 37884 1428 37940 5180
rect 37996 4340 38052 11228
rect 38220 11284 38276 13468
rect 38332 12516 38388 14112
rect 38444 12852 38500 12862
rect 38444 12758 38500 12796
rect 38556 12628 38612 14112
rect 38556 12562 38612 12572
rect 38668 12740 38724 12750
rect 38332 12450 38388 12460
rect 38668 11618 38724 12684
rect 38780 12180 38836 14112
rect 38780 12114 38836 12124
rect 38892 13860 38948 13870
rect 38668 11566 38670 11618
rect 38722 11566 38724 11618
rect 38668 11554 38724 11566
rect 38892 11284 38948 13804
rect 39004 13076 39060 14112
rect 39228 13300 39284 14112
rect 39228 13234 39284 13244
rect 39340 13860 39396 13870
rect 39004 13010 39060 13020
rect 39116 12962 39172 12974
rect 39116 12910 39118 12962
rect 39170 12910 39172 12962
rect 38220 11218 38276 11228
rect 38668 11228 38948 11284
rect 39004 12178 39060 12190
rect 39004 12126 39006 12178
rect 39058 12126 39060 12178
rect 38332 9826 38388 9838
rect 38332 9774 38334 9826
rect 38386 9774 38388 9826
rect 38332 9156 38388 9774
rect 38332 9090 38388 9100
rect 38668 9042 38724 11228
rect 38780 10500 38836 10510
rect 38780 10406 38836 10444
rect 38668 8990 38670 9042
rect 38722 8990 38724 9042
rect 38668 8978 38724 8990
rect 39004 8428 39060 12126
rect 39116 11956 39172 12910
rect 39340 12740 39396 13804
rect 39340 12674 39396 12684
rect 39116 11890 39172 11900
rect 39340 12404 39396 12414
rect 39116 11284 39172 11294
rect 39116 9938 39172 11228
rect 39340 10834 39396 12348
rect 39452 12292 39508 14112
rect 39452 12226 39508 12236
rect 39564 13188 39620 13198
rect 39340 10782 39342 10834
rect 39394 10782 39396 10834
rect 39340 10770 39396 10782
rect 39452 12066 39508 12078
rect 39452 12014 39454 12066
rect 39506 12014 39508 12066
rect 39452 10388 39508 12014
rect 39452 10322 39508 10332
rect 39116 9886 39118 9938
rect 39170 9886 39172 9938
rect 39116 9874 39172 9886
rect 39116 9044 39172 9054
rect 39116 8950 39172 8988
rect 39004 8372 39172 8428
rect 38556 7588 38612 7598
rect 37996 4274 38052 4284
rect 38332 5794 38388 5806
rect 38332 5742 38334 5794
rect 38386 5742 38388 5794
rect 38332 2884 38388 5742
rect 38332 2818 38388 2828
rect 37884 1362 37940 1372
rect 36876 690 36932 700
rect 36764 130 36820 140
rect 38556 112 38612 7532
rect 39004 7476 39060 7486
rect 38668 5908 38724 5918
rect 38668 5814 38724 5852
rect 38892 5124 38948 5134
rect 38892 5030 38948 5068
rect 38780 4004 38836 4014
rect 38780 3668 38836 3948
rect 39004 3780 39060 7420
rect 39116 6804 39172 8372
rect 39116 6738 39172 6748
rect 39340 8372 39396 8382
rect 39228 5796 39284 5806
rect 39228 5702 39284 5740
rect 39004 3714 39060 3724
rect 38780 3602 38836 3612
rect 38892 3332 38948 3342
rect 38892 2770 38948 3276
rect 39340 2882 39396 8316
rect 39452 5124 39508 5134
rect 39452 5030 39508 5068
rect 39564 5012 39620 13132
rect 39676 12964 39732 14112
rect 39676 12898 39732 12908
rect 39788 13412 39844 13422
rect 39788 12850 39844 13356
rect 39788 12798 39790 12850
rect 39842 12798 39844 12850
rect 39788 12786 39844 12798
rect 39676 12740 39732 12750
rect 39676 8428 39732 12684
rect 39900 12404 39956 14112
rect 39900 12338 39956 12348
rect 40012 13748 40068 13758
rect 40012 12402 40068 13692
rect 40124 13188 40180 14112
rect 40124 13122 40180 13132
rect 41244 13524 41300 13534
rect 41244 13186 41300 13468
rect 41244 13134 41246 13186
rect 41298 13134 41300 13186
rect 41244 13122 41300 13134
rect 42364 13300 42420 13310
rect 40012 12350 40014 12402
rect 40066 12350 40068 12402
rect 40012 12338 40068 12350
rect 40348 12964 40404 12974
rect 40236 12068 40292 12078
rect 40236 9828 40292 12012
rect 40348 11172 40404 12908
rect 40684 12962 40740 12974
rect 40684 12910 40686 12962
rect 40738 12910 40740 12962
rect 40684 11620 40740 12910
rect 40684 11554 40740 11564
rect 40796 12628 40852 12638
rect 40796 11618 40852 12572
rect 41580 12516 41636 12526
rect 41580 12402 41636 12460
rect 41580 12350 41582 12402
rect 41634 12350 41636 12402
rect 41580 12338 41636 12350
rect 40796 11566 40798 11618
rect 40850 11566 40852 11618
rect 40796 11554 40852 11566
rect 40908 12292 40964 12302
rect 40460 11396 40516 11406
rect 40460 11394 40740 11396
rect 40460 11342 40462 11394
rect 40514 11342 40740 11394
rect 40460 11340 40740 11342
rect 40460 11330 40516 11340
rect 40348 11116 40516 11172
rect 40236 9762 40292 9772
rect 40348 9826 40404 9838
rect 40348 9774 40350 9826
rect 40402 9774 40404 9826
rect 39900 8930 39956 8942
rect 39900 8878 39902 8930
rect 39954 8878 39956 8930
rect 39676 8372 39844 8428
rect 39564 4946 39620 4956
rect 39676 7252 39732 7262
rect 39676 3556 39732 7196
rect 39676 3490 39732 3500
rect 39340 2830 39342 2882
rect 39394 2830 39396 2882
rect 39340 2818 39396 2830
rect 38892 2718 38894 2770
rect 38946 2718 38948 2770
rect 38892 2706 38948 2718
rect 39676 2100 39732 2110
rect 39676 2006 39732 2044
rect 39116 1986 39172 1998
rect 39116 1934 39118 1986
rect 39170 1934 39172 1986
rect 39116 1652 39172 1934
rect 39116 1586 39172 1596
rect 30548 28 30660 84
rect 30492 18 30548 28
rect 31136 0 31248 112
rect 33600 0 33712 112
rect 36064 0 36176 112
rect 38528 0 38640 112
rect 39788 84 39844 8372
rect 39900 6132 39956 8878
rect 39900 6066 39956 6076
rect 40348 5572 40404 9774
rect 40460 9266 40516 11116
rect 40460 9214 40462 9266
rect 40514 9214 40516 9266
rect 40460 9202 40516 9214
rect 40572 10610 40628 10622
rect 40572 10558 40574 10610
rect 40626 10558 40628 10610
rect 40460 9044 40516 9054
rect 40460 6580 40516 8988
rect 40460 6514 40516 6524
rect 40348 5506 40404 5516
rect 40572 5460 40628 10558
rect 40572 5394 40628 5404
rect 40684 4788 40740 11340
rect 40908 10948 40964 12236
rect 41132 12180 41188 12190
rect 40796 10892 40964 10948
rect 41020 12066 41076 12078
rect 41020 12014 41022 12066
rect 41074 12014 41076 12066
rect 40796 10050 40852 10892
rect 40796 9998 40798 10050
rect 40850 9998 40852 10050
rect 40796 9986 40852 9998
rect 40908 10612 40964 10622
rect 40908 9828 40964 10556
rect 40796 9772 40964 9828
rect 40796 6580 40852 9772
rect 40796 6514 40852 6524
rect 40908 9604 40964 9614
rect 40684 4722 40740 4732
rect 40236 4676 40292 4686
rect 40236 2772 40292 4620
rect 40348 4564 40404 4574
rect 40348 3220 40404 4508
rect 40908 4452 40964 9548
rect 41020 8148 41076 12014
rect 41132 10722 41188 12124
rect 41916 11732 41972 11742
rect 41132 10670 41134 10722
rect 41186 10670 41188 10722
rect 41132 10658 41188 10670
rect 41804 11394 41860 11406
rect 41804 11342 41806 11394
rect 41858 11342 41860 11394
rect 41804 10164 41860 11342
rect 41804 10098 41860 10108
rect 41916 9826 41972 11676
rect 42364 11618 42420 13244
rect 43708 13076 43764 13086
rect 43708 12982 43764 13020
rect 42924 12962 42980 12974
rect 42924 12910 42926 12962
rect 42978 12910 42980 12962
rect 42588 12852 42644 12862
rect 42364 11566 42366 11618
rect 42418 11566 42420 11618
rect 42364 11554 42420 11566
rect 42476 12404 42532 12414
rect 42140 11284 42196 11294
rect 41916 9774 41918 9826
rect 41970 9774 41972 9826
rect 41916 9762 41972 9774
rect 42028 10610 42084 10622
rect 42028 10558 42030 10610
rect 42082 10558 42084 10610
rect 41020 8082 41076 8092
rect 41244 8148 41300 8158
rect 40908 4386 40964 4396
rect 40348 3154 40404 3164
rect 40236 2706 40292 2716
rect 41244 2660 41300 8092
rect 42028 7924 42084 10558
rect 42028 7858 42084 7868
rect 42140 5684 42196 11228
rect 42476 10834 42532 12348
rect 42588 12178 42644 12796
rect 42588 12126 42590 12178
rect 42642 12126 42644 12178
rect 42588 12114 42644 12126
rect 42476 10782 42478 10834
rect 42530 10782 42532 10834
rect 42476 10770 42532 10782
rect 42252 9716 42308 9726
rect 42252 9622 42308 9660
rect 42924 8596 42980 12910
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 42924 8530 42980 8540
rect 43148 12066 43204 12078
rect 43148 12014 43150 12066
rect 43202 12014 43204 12066
rect 43148 6356 43204 12014
rect 43484 11060 43540 11070
rect 43148 6290 43204 6300
rect 43372 10612 43428 10622
rect 42140 5618 42196 5628
rect 42812 4226 42868 4238
rect 42812 4174 42814 4226
rect 42866 4174 42868 4226
rect 41244 2594 41300 2604
rect 42252 4114 42308 4126
rect 42252 4062 42254 4114
rect 42306 4062 42308 4114
rect 42252 1316 42308 4062
rect 42812 4116 42868 4174
rect 42812 4050 42868 4060
rect 43372 2100 43428 10556
rect 43372 2034 43428 2044
rect 42252 1250 42308 1260
rect 41020 980 41076 990
rect 41020 112 41076 924
rect 43484 112 43540 11004
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 43932 10500 43988 10510
rect 43932 10050 43988 10444
rect 43932 9998 43934 10050
rect 43986 9998 43988 10050
rect 43932 9986 43988 9998
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 44156 8428 44212 14140
rect 51100 13972 51156 13982
rect 50540 13524 50596 13534
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 45052 13188 45108 13198
rect 45052 13094 45108 13132
rect 48076 13076 48132 13086
rect 44492 12964 44548 12974
rect 44268 12962 44548 12964
rect 44268 12910 44494 12962
rect 44546 12910 44548 12962
rect 44268 12908 44548 12910
rect 44268 10052 44324 12908
rect 44492 12898 44548 12908
rect 47180 12962 47236 12974
rect 47180 12910 47182 12962
rect 47234 12910 47236 12962
rect 45164 12068 45220 12078
rect 47068 12068 47124 12078
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44268 9986 44324 9996
rect 44828 9826 44884 9838
rect 44828 9774 44830 9826
rect 44882 9774 44884 9826
rect 44492 9716 44548 9726
rect 44492 9622 44548 9660
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44156 8372 44324 8428
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 43596 7140 43652 7150
rect 43596 4564 43652 7084
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 44268 5908 44324 8372
rect 44828 8372 44884 9774
rect 44828 8306 44884 8316
rect 45164 8260 45220 12012
rect 46956 12066 47124 12068
rect 46956 12014 47070 12066
rect 47122 12014 47124 12066
rect 46956 12012 47124 12014
rect 45948 10724 46004 10734
rect 45276 9828 45332 9838
rect 45276 9714 45332 9772
rect 45276 9662 45278 9714
rect 45330 9662 45332 9714
rect 45276 9650 45332 9662
rect 45164 8194 45220 8204
rect 45388 8820 45444 8830
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44604 6690 44660 6702
rect 44604 6638 44606 6690
rect 44658 6638 44660 6690
rect 44604 6580 44660 6638
rect 45388 6692 45444 8764
rect 45388 6626 45444 6636
rect 45500 8484 45556 8494
rect 44604 6514 44660 6524
rect 45052 6578 45108 6590
rect 45052 6526 45054 6578
rect 45106 6526 45108 6578
rect 44268 5842 44324 5852
rect 43932 5684 43988 5694
rect 43932 5012 43988 5628
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 45052 5236 45108 6526
rect 45052 5170 45108 5180
rect 43932 4946 43988 4956
rect 45500 5012 45556 8428
rect 45500 4946 45556 4956
rect 45836 4900 45892 4910
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 43596 4508 43764 4564
rect 43708 3332 43764 4508
rect 44156 4228 44212 4238
rect 44156 4134 44212 4172
rect 44716 4228 44772 4238
rect 44716 4226 44884 4228
rect 44716 4174 44718 4226
rect 44770 4174 44884 4226
rect 44716 4172 44884 4174
rect 44716 4162 44772 4172
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 44716 3556 44772 3566
rect 44716 3462 44772 3500
rect 43652 3276 43764 3332
rect 43652 2996 43708 3276
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 43652 2940 43876 2996
rect 43820 2210 43876 2940
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 43820 2158 43822 2210
rect 43874 2158 43876 2210
rect 43820 2146 43876 2158
rect 44268 1876 44324 1886
rect 44268 1782 44324 1820
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 44828 420 44884 4172
rect 45276 3780 45332 3790
rect 45276 3666 45332 3724
rect 45836 3778 45892 4844
rect 45948 4788 46004 10668
rect 46956 9044 47012 12012
rect 47068 12002 47124 12012
rect 47180 9604 47236 12910
rect 48076 12402 48132 13020
rect 48972 12964 49028 12974
rect 48972 12962 49364 12964
rect 48972 12910 48974 12962
rect 49026 12910 49364 12962
rect 48972 12908 49364 12910
rect 48972 12898 49028 12908
rect 48188 12738 48244 12750
rect 48188 12686 48190 12738
rect 48242 12686 48244 12738
rect 48188 12628 48244 12686
rect 48188 12562 48244 12572
rect 48076 12350 48078 12402
rect 48130 12350 48132 12402
rect 48076 12338 48132 12350
rect 47180 9538 47236 9548
rect 47292 12292 47348 12302
rect 46956 8978 47012 8988
rect 46620 8036 46676 8046
rect 46284 6692 46340 6702
rect 45948 4722 46004 4732
rect 46172 5796 46228 5806
rect 45836 3726 45838 3778
rect 45890 3726 45892 3778
rect 45836 3714 45892 3726
rect 45276 3614 45278 3666
rect 45330 3614 45332 3666
rect 45276 3602 45332 3614
rect 45388 2772 45444 2782
rect 45388 2678 45444 2716
rect 46172 2772 46228 5740
rect 46172 2706 46228 2716
rect 45948 2658 46004 2670
rect 45948 2606 45950 2658
rect 46002 2606 46004 2658
rect 45948 2100 46004 2606
rect 46284 2548 46340 6636
rect 46396 4114 46452 4126
rect 46396 4062 46398 4114
rect 46450 4062 46452 4114
rect 46396 3668 46452 4062
rect 46396 3602 46452 3612
rect 46620 3668 46676 7980
rect 46732 4340 46788 4350
rect 46732 3778 46788 4284
rect 46732 3726 46734 3778
rect 46786 3726 46788 3778
rect 46732 3714 46788 3726
rect 46956 4226 47012 4238
rect 46956 4174 46958 4226
rect 47010 4174 47012 4226
rect 46620 3602 46676 3612
rect 46396 3444 46452 3454
rect 46396 3350 46452 3388
rect 46956 2996 47012 4174
rect 47292 3666 47348 12236
rect 48748 12178 48804 12190
rect 48748 12126 48750 12178
rect 48802 12126 48804 12178
rect 47740 11956 47796 11966
rect 47628 10836 47684 10846
rect 47628 8260 47684 10780
rect 47740 10610 47796 11900
rect 47740 10558 47742 10610
rect 47794 10558 47796 10610
rect 47740 10546 47796 10558
rect 48300 10500 48356 10510
rect 48300 10406 48356 10444
rect 48300 8930 48356 8942
rect 48300 8878 48302 8930
rect 48354 8878 48356 8930
rect 47740 8820 47796 8830
rect 47740 8726 47796 8764
rect 48300 8708 48356 8878
rect 48300 8642 48356 8652
rect 48636 8930 48692 8942
rect 48636 8878 48638 8930
rect 48690 8878 48692 8930
rect 48636 8428 48692 8878
rect 47628 8194 47684 8204
rect 48524 8372 48692 8428
rect 48748 8428 48804 12126
rect 48860 11394 48916 11406
rect 48860 11342 48862 11394
rect 48914 11342 48916 11394
rect 48860 11172 48916 11342
rect 48860 11106 48916 11116
rect 48972 11284 49028 11294
rect 48860 10612 48916 10622
rect 48972 10612 49028 11228
rect 48860 10610 49028 10612
rect 48860 10558 48862 10610
rect 48914 10558 49028 10610
rect 48860 10556 49028 10558
rect 48860 10546 48916 10556
rect 49084 9826 49140 9838
rect 49084 9774 49086 9826
rect 49138 9774 49140 9826
rect 48972 9716 49028 9726
rect 48748 8372 48916 8428
rect 47404 7588 47460 7598
rect 47404 6020 47460 7532
rect 48524 6916 48580 8372
rect 48636 8260 48692 8270
rect 48636 8166 48692 8204
rect 48748 7474 48804 7486
rect 48748 7422 48750 7474
rect 48802 7422 48804 7474
rect 48748 7364 48804 7422
rect 48748 7298 48804 7308
rect 48860 6916 48916 8372
rect 48524 6850 48580 6860
rect 48748 6860 48916 6916
rect 47404 5954 47460 5964
rect 48524 6468 48580 6478
rect 48524 6018 48580 6412
rect 48524 5966 48526 6018
rect 48578 5966 48580 6018
rect 48524 5954 48580 5966
rect 48076 5684 48132 5694
rect 48076 5590 48132 5628
rect 48748 5236 48804 6860
rect 48860 6692 48916 6702
rect 48860 6598 48916 6636
rect 48748 5180 48916 5236
rect 48748 5012 48804 5022
rect 48188 4564 48244 4574
rect 48188 4450 48244 4508
rect 48188 4398 48190 4450
rect 48242 4398 48244 4450
rect 48188 4386 48244 4398
rect 48748 4338 48804 4956
rect 48748 4286 48750 4338
rect 48802 4286 48804 4338
rect 48748 4274 48804 4286
rect 47292 3614 47294 3666
rect 47346 3614 47348 3666
rect 47292 3602 47348 3614
rect 47740 4114 47796 4126
rect 47740 4062 47742 4114
rect 47794 4062 47796 4114
rect 47740 3332 47796 4062
rect 48860 3892 48916 5180
rect 48972 5122 49028 9660
rect 49084 8428 49140 9774
rect 49308 8428 49364 12908
rect 49756 12738 49812 12750
rect 49756 12686 49758 12738
rect 49810 12686 49812 12738
rect 49644 12290 49700 12302
rect 49644 12238 49646 12290
rect 49698 12238 49700 12290
rect 49644 11844 49700 12238
rect 49756 12180 49812 12686
rect 49756 12114 49812 12124
rect 50204 12068 50260 12078
rect 50204 11974 50260 12012
rect 49644 11778 49700 11788
rect 50428 11396 50484 11406
rect 50428 11302 50484 11340
rect 49868 11284 49924 11294
rect 49868 11190 49924 11228
rect 49644 10722 49700 10734
rect 49644 10670 49646 10722
rect 49698 10670 49700 10722
rect 49644 10388 49700 10670
rect 50204 10612 50260 10622
rect 50204 10518 50260 10556
rect 49644 10322 49700 10332
rect 50428 9940 50484 9950
rect 50428 9846 50484 9884
rect 49868 9716 49924 9726
rect 49868 9622 49924 9660
rect 50540 9716 50596 13468
rect 50876 12962 50932 12974
rect 50876 12910 50878 12962
rect 50930 12910 50932 12962
rect 50540 9650 50596 9660
rect 50652 10500 50708 10510
rect 49644 9268 49700 9278
rect 49644 9174 49700 9212
rect 50204 8932 50260 8942
rect 50204 8838 50260 8876
rect 50316 8708 50372 8718
rect 49084 8372 49252 8428
rect 49308 8372 49476 8428
rect 49084 8146 49140 8158
rect 49084 8094 49086 8146
rect 49138 8094 49140 8146
rect 49084 6804 49140 8094
rect 49084 6738 49140 6748
rect 48972 5070 48974 5122
rect 49026 5070 49028 5122
rect 48972 5058 49028 5070
rect 49084 5460 49140 5470
rect 48860 3826 48916 3836
rect 48860 3668 48916 3678
rect 48860 3574 48916 3612
rect 47740 3266 47796 3276
rect 46956 2930 47012 2940
rect 47068 2884 47124 2894
rect 47068 2770 47124 2828
rect 48076 2884 48132 2894
rect 48076 2790 48132 2828
rect 47068 2718 47070 2770
rect 47122 2718 47124 2770
rect 47068 2706 47124 2718
rect 48748 2772 48804 2782
rect 48748 2678 48804 2716
rect 46284 2482 46340 2492
rect 45948 2034 46004 2044
rect 47516 2436 47572 2446
rect 47516 2098 47572 2380
rect 47516 2046 47518 2098
rect 47570 2046 47572 2098
rect 47516 2034 47572 2046
rect 48860 2100 48916 2110
rect 48860 2006 48916 2044
rect 47068 1986 47124 1998
rect 47068 1934 47070 1986
rect 47122 1934 47124 1986
rect 47068 1764 47124 1934
rect 47068 1698 47124 1708
rect 48188 1314 48244 1326
rect 48188 1262 48190 1314
rect 48242 1262 48244 1314
rect 47180 1092 47236 1102
rect 47180 998 47236 1036
rect 48188 980 48244 1262
rect 49084 1316 49140 5404
rect 49196 3444 49252 8372
rect 49308 5908 49364 5918
rect 49308 5814 49364 5852
rect 49420 5236 49476 8372
rect 49532 8258 49588 8270
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 7476 49588 8206
rect 49980 8148 50036 8158
rect 49980 8054 50036 8092
rect 49532 7410 49588 7420
rect 49644 7586 49700 7598
rect 49644 7534 49646 7586
rect 49698 7534 49700 7586
rect 49644 6804 49700 7534
rect 49644 6738 49700 6748
rect 49756 6578 49812 6590
rect 49756 6526 49758 6578
rect 49810 6526 49812 6578
rect 49756 5908 49812 6526
rect 49868 6020 49924 6030
rect 49868 5926 49924 5964
rect 49756 5842 49812 5852
rect 50204 5794 50260 5806
rect 50204 5742 50206 5794
rect 50258 5742 50260 5794
rect 50204 5348 50260 5742
rect 50204 5282 50260 5292
rect 49420 5170 49476 5180
rect 49644 5124 49700 5134
rect 49644 5030 49700 5068
rect 50204 4788 50260 4798
rect 50204 4338 50260 4732
rect 50204 4286 50206 4338
rect 50258 4286 50260 4338
rect 50204 4274 50260 4286
rect 49420 4226 49476 4238
rect 49420 4174 49422 4226
rect 49474 4174 49476 4226
rect 49420 3668 49476 4174
rect 49420 3602 49476 3612
rect 49196 3378 49252 3388
rect 49868 3444 49924 3454
rect 49868 3350 49924 3388
rect 50316 2770 50372 8652
rect 50428 8372 50484 8382
rect 50428 8278 50484 8316
rect 50428 6690 50484 6702
rect 50428 6638 50430 6690
rect 50482 6638 50484 6690
rect 50428 3780 50484 6638
rect 50652 5122 50708 10444
rect 50876 8428 50932 12910
rect 50988 10498 51044 10510
rect 50988 10446 50990 10498
rect 51042 10446 51044 10498
rect 50988 9492 51044 10446
rect 50988 9426 51044 9436
rect 51100 9268 51156 13916
rect 51212 13636 51268 13646
rect 51212 12850 51268 13580
rect 51212 12798 51214 12850
rect 51266 12798 51268 12850
rect 51212 12786 51268 12798
rect 51212 12290 51268 12302
rect 51212 12238 51214 12290
rect 51266 12238 51268 12290
rect 51212 10836 51268 12238
rect 51212 10770 51268 10780
rect 51436 11170 51492 11182
rect 51436 11118 51438 11170
rect 51490 11118 51492 11170
rect 51436 9940 51492 11118
rect 51436 9874 51492 9884
rect 51100 9202 51156 9212
rect 51436 9602 51492 9614
rect 51436 9550 51438 9602
rect 51490 9550 51492 9602
rect 51436 9044 51492 9550
rect 51436 8978 51492 8988
rect 50988 8930 51044 8942
rect 50988 8878 50990 8930
rect 51042 8878 51044 8930
rect 50988 8596 51044 8878
rect 50988 8530 51044 8540
rect 50764 8372 50932 8428
rect 50764 5460 50820 8372
rect 50876 8148 50932 8158
rect 50876 7698 50932 8092
rect 50876 7646 50878 7698
rect 50930 7646 50932 7698
rect 50876 7634 50932 7646
rect 51436 8034 51492 8046
rect 51436 7982 51438 8034
rect 51490 7982 51492 8034
rect 51436 7700 51492 7982
rect 51436 7634 51492 7644
rect 51324 7474 51380 7486
rect 51324 7422 51326 7474
rect 51378 7422 51380 7474
rect 51212 6356 51268 6366
rect 51212 6130 51268 6300
rect 51212 6078 51214 6130
rect 51266 6078 51268 6130
rect 51212 6066 51268 6078
rect 50764 5394 50820 5404
rect 51212 5460 51268 5470
rect 51212 5234 51268 5404
rect 51212 5182 51214 5234
rect 51266 5182 51268 5234
rect 51212 5170 51268 5182
rect 50652 5070 50654 5122
rect 50706 5070 50708 5122
rect 50652 5058 50708 5070
rect 51100 5124 51156 5134
rect 51100 4564 51156 5068
rect 51100 4498 51156 4508
rect 51212 5012 51268 5022
rect 51212 4562 51268 4956
rect 51212 4510 51214 4562
rect 51266 4510 51268 4562
rect 51212 4498 51268 4510
rect 50428 3714 50484 3724
rect 50316 2718 50318 2770
rect 50370 2718 50372 2770
rect 50316 2706 50372 2718
rect 50428 3554 50484 3566
rect 50428 3502 50430 3554
rect 50482 3502 50484 3554
rect 49420 2660 49476 2670
rect 49420 2566 49476 2604
rect 50428 2436 50484 3502
rect 51100 3444 51156 3454
rect 50428 2370 50484 2380
rect 50540 2884 50596 2894
rect 50316 2212 50372 2222
rect 50372 2156 50484 2212
rect 50316 2146 50372 2156
rect 50428 2098 50484 2156
rect 50428 2046 50430 2098
rect 50482 2046 50484 2098
rect 50428 2034 50484 2046
rect 49868 1876 49924 1886
rect 49868 1782 49924 1820
rect 49756 1428 49812 1438
rect 49756 1334 49812 1372
rect 49084 1250 49140 1260
rect 48748 1204 48804 1214
rect 48748 1110 48804 1148
rect 48188 914 48244 924
rect 50540 532 50596 2828
rect 51100 2772 51156 3388
rect 51212 3220 51268 3230
rect 51212 2994 51268 3164
rect 51212 2942 51214 2994
rect 51266 2942 51268 2994
rect 51212 2930 51268 2942
rect 51100 2706 51156 2716
rect 51324 1314 51380 7422
rect 51436 7252 51492 7262
rect 51436 6578 51492 7196
rect 51436 6526 51438 6578
rect 51490 6526 51492 6578
rect 51436 6514 51492 6526
rect 51436 4116 51492 4126
rect 51436 3442 51492 4060
rect 51436 3390 51438 3442
rect 51490 3390 51492 3442
rect 51436 3378 51492 3390
rect 51548 2660 51604 2670
rect 51436 2324 51492 2334
rect 51436 1874 51492 2268
rect 51436 1822 51438 1874
rect 51490 1822 51492 1874
rect 51436 1810 51492 1822
rect 51324 1262 51326 1314
rect 51378 1262 51380 1314
rect 51324 1250 51380 1262
rect 50764 978 50820 990
rect 50764 926 50766 978
rect 50818 926 50820 978
rect 50764 644 50820 926
rect 50764 578 50820 588
rect 50540 466 50596 476
rect 44828 354 44884 364
rect 45948 308 46004 318
rect 45948 112 46004 252
rect 50876 308 50932 318
rect 48412 196 48468 206
rect 48412 112 48468 140
rect 50876 112 50932 252
rect 39788 18 39844 28
rect 40992 0 41104 112
rect 43456 0 43568 112
rect 45920 0 46032 112
rect 48384 0 48496 112
rect 50848 0 50960 112
rect 51548 84 51604 2604
rect 51548 18 51604 28
<< via2 >>
rect 44156 14140 44212 14196
rect 11564 14028 11620 14084
rect 140 13916 196 13972
rect 10332 13916 10388 13972
rect 1260 13468 1316 13524
rect 140 7420 196 7476
rect 364 12124 420 12180
rect 9772 13468 9828 13524
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 7756 13132 7812 13188
rect 1260 11116 1316 11172
rect 2268 13020 2324 13076
rect 1372 10780 1428 10836
rect 1148 9772 1204 9828
rect 364 6860 420 6916
rect 924 8540 980 8596
rect 2044 10780 2100 10836
rect 1372 9212 1428 9268
rect 1708 9884 1764 9940
rect 1484 8988 1540 9044
rect 1148 7644 1204 7700
rect 1372 8428 1428 8484
rect 1260 7308 1316 7364
rect 1036 4732 1092 4788
rect 1036 2716 1092 2772
rect 1596 8092 1652 8148
rect 1596 6636 1652 6692
rect 1484 6412 1540 6468
rect 1372 6300 1428 6356
rect 1372 5852 1428 5908
rect 1372 2604 1428 2660
rect 1484 4060 1540 4116
rect 1260 2268 1316 2324
rect 1484 2156 1540 2212
rect 1596 3612 1652 3668
rect 1820 6524 1876 6580
rect 1932 6300 1988 6356
rect 1820 4844 1876 4900
rect 2156 8764 2212 8820
rect 2716 12796 2772 12852
rect 6188 12684 6244 12740
rect 3276 12572 3332 12628
rect 3164 12348 3220 12404
rect 3164 11340 3220 11396
rect 3052 9996 3108 10052
rect 2828 7980 2884 8036
rect 2268 7532 2324 7588
rect 2716 7644 2772 7700
rect 2604 6860 2660 6916
rect 2380 4508 2436 4564
rect 2268 4284 2324 4340
rect 2156 2940 2212 2996
rect 2604 4172 2660 4228
rect 2716 3388 2772 3444
rect 2268 2044 2324 2100
rect 1596 1932 1652 1988
rect 924 1148 980 1204
rect 1484 1820 1540 1876
rect 1484 476 1540 532
rect 1596 1372 1652 1428
rect 2940 5628 2996 5684
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 5292 11116 5348 11172
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3276 10668 3332 10724
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 3164 9772 3220 9828
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3612 6300 3668 6356
rect 3388 5740 3444 5796
rect 3052 4732 3108 4788
rect 3164 5404 3220 5460
rect 3276 4620 3332 4676
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4172 4732 4228 4788
rect 3612 4396 3668 4452
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 3948 2882 4004 2884
rect 3948 2830 3950 2882
rect 3950 2830 4002 2882
rect 4002 2830 4004 2882
rect 3948 2828 4004 2830
rect 3164 2716 3220 2772
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 5068 4060 5124 4116
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 4396 2658 4452 2660
rect 4396 2606 4398 2658
rect 4398 2606 4450 2658
rect 4450 2606 4452 2658
rect 4396 2604 4452 2606
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 2940 924 2996 980
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 5628 9324 5684 9380
rect 5404 6524 5460 6580
rect 5516 8988 5572 9044
rect 5628 4732 5684 4788
rect 5404 4172 5460 4228
rect 5404 924 5460 980
rect 5292 588 5348 644
rect 6748 12066 6804 12068
rect 6748 12014 6750 12066
rect 6750 12014 6802 12066
rect 6802 12014 6804 12066
rect 6748 12012 6804 12014
rect 6300 11954 6356 11956
rect 6300 11902 6302 11954
rect 6302 11902 6354 11954
rect 6354 11902 6356 11954
rect 6300 11900 6356 11902
rect 5852 8876 5908 8932
rect 6524 11116 6580 11172
rect 6636 8316 6692 8372
rect 6524 7308 6580 7364
rect 6636 7196 6692 7252
rect 6412 7084 6468 7140
rect 5852 5682 5908 5684
rect 5852 5630 5854 5682
rect 5854 5630 5906 5682
rect 5906 5630 5908 5682
rect 5852 5628 5908 5630
rect 6412 5292 6468 5348
rect 6524 5234 6580 5236
rect 6524 5182 6526 5234
rect 6526 5182 6578 5234
rect 6578 5182 6580 5234
rect 6524 5180 6580 5182
rect 6860 6524 6916 6580
rect 6636 3836 6692 3892
rect 6748 6188 6804 6244
rect 6076 3164 6132 3220
rect 6636 3164 6692 3220
rect 5964 1260 6020 1316
rect 6412 2604 6468 2660
rect 6636 2604 6692 2660
rect 6412 1036 6468 1092
rect 5740 252 5796 308
rect 7308 3948 7364 4004
rect 7532 11900 7588 11956
rect 6860 812 6916 868
rect 7644 8540 7700 8596
rect 11340 13580 11396 13636
rect 10892 12460 10948 12516
rect 8876 12236 8932 12292
rect 7980 11564 8036 11620
rect 8092 9548 8148 9604
rect 8092 8204 8148 8260
rect 7980 6524 8036 6580
rect 7756 2828 7812 2884
rect 8316 10444 8372 10500
rect 8540 10332 8596 10388
rect 8316 7644 8372 7700
rect 8428 9212 8484 9268
rect 8316 6300 8372 6356
rect 8316 4284 8372 4340
rect 9772 12012 9828 12068
rect 8988 11452 9044 11508
rect 9324 9100 9380 9156
rect 9212 8428 9268 8484
rect 9436 7868 9492 7924
rect 9212 6412 9268 6468
rect 9100 5516 9156 5572
rect 8988 5404 9044 5460
rect 8540 5068 8596 5124
rect 8540 4508 8596 4564
rect 8428 3388 8484 3444
rect 8204 2044 8260 2100
rect 7532 476 7588 532
rect 9884 11676 9940 11732
rect 10444 11788 10500 11844
rect 10108 10780 10164 10836
rect 10108 10444 10164 10500
rect 11340 11564 11396 11620
rect 10668 10444 10724 10500
rect 10556 10108 10612 10164
rect 10668 10050 10724 10052
rect 10668 9998 10670 10050
rect 10670 9998 10722 10050
rect 10722 9998 10724 10050
rect 10668 9996 10724 9998
rect 10556 8988 10612 9044
rect 9996 8540 10052 8596
rect 9772 8092 9828 8148
rect 9996 7756 10052 7812
rect 10332 8540 10388 8596
rect 9884 6412 9940 6468
rect 10220 5964 10276 6020
rect 10332 5740 10388 5796
rect 11004 5682 11060 5684
rect 11004 5630 11006 5682
rect 11006 5630 11058 5682
rect 11058 5630 11060 5682
rect 11004 5628 11060 5630
rect 10444 4956 10500 5012
rect 9548 1260 9604 1316
rect 10220 2380 10276 2436
rect 10108 1820 10164 1876
rect 10108 1596 10164 1652
rect 11228 3724 11284 3780
rect 12348 14028 12404 14084
rect 11676 13020 11732 13076
rect 11900 12796 11956 12852
rect 12348 12684 12404 12740
rect 11788 12348 11844 12404
rect 12236 12066 12292 12068
rect 12236 12014 12238 12066
rect 12238 12014 12290 12066
rect 12290 12014 12292 12066
rect 12236 12012 12292 12014
rect 12460 11900 12516 11956
rect 11788 10332 11844 10388
rect 11788 9772 11844 9828
rect 11788 9548 11844 9604
rect 11452 7644 11508 7700
rect 11676 8652 11732 8708
rect 11788 8316 11844 8372
rect 13020 12460 13076 12516
rect 13356 13244 13412 13300
rect 13244 12348 13300 12404
rect 12572 11788 12628 11844
rect 12796 10556 12852 10612
rect 12236 9042 12292 9044
rect 12236 8990 12238 9042
rect 12238 8990 12290 9042
rect 12290 8990 12292 9042
rect 12236 8988 12292 8990
rect 12460 8258 12516 8260
rect 12460 8206 12462 8258
rect 12462 8206 12514 8258
rect 12514 8206 12516 8258
rect 12460 8204 12516 8206
rect 12124 7308 12180 7364
rect 11676 4620 11732 4676
rect 11788 7084 11844 7140
rect 12236 6748 12292 6804
rect 11900 6636 11956 6692
rect 11900 4844 11956 4900
rect 11788 4284 11844 4340
rect 11340 3164 11396 3220
rect 10892 2882 10948 2884
rect 10892 2830 10894 2882
rect 10894 2830 10946 2882
rect 10946 2830 10948 2882
rect 10892 2828 10948 2830
rect 10668 1484 10724 1540
rect 10220 1148 10276 1204
rect 10444 1148 10500 1204
rect 10444 924 10500 980
rect 9884 700 9940 756
rect 11788 2940 11844 2996
rect 13020 12124 13076 12180
rect 13244 10892 13300 10948
rect 12796 4508 12852 4564
rect 13020 6860 13076 6916
rect 12796 3276 12852 3332
rect 12796 2156 12852 2212
rect 13020 1932 13076 1988
rect 11788 924 11844 980
rect 11788 588 11844 644
rect 2828 28 2884 84
rect 13692 11900 13748 11956
rect 14364 13468 14420 13524
rect 14476 13804 14532 13860
rect 13916 11788 13972 11844
rect 14028 11900 14084 11956
rect 14140 11788 14196 11844
rect 13580 11116 13636 11172
rect 13580 9660 13636 9716
rect 13804 10220 13860 10276
rect 14028 10050 14084 10052
rect 14028 9998 14030 10050
rect 14030 9998 14082 10050
rect 14082 9998 14084 10050
rect 14028 9996 14084 9998
rect 13692 8316 13748 8372
rect 13580 7756 13636 7812
rect 13468 5740 13524 5796
rect 13468 2940 13524 2996
rect 13356 2268 13412 2324
rect 14588 13020 14644 13076
rect 14924 13468 14980 13524
rect 14812 12684 14868 12740
rect 14812 12402 14868 12404
rect 14812 12350 14814 12402
rect 14814 12350 14866 12402
rect 14866 12350 14868 12402
rect 14812 12348 14868 12350
rect 14812 11676 14868 11732
rect 14924 11116 14980 11172
rect 14588 10332 14644 10388
rect 14476 10108 14532 10164
rect 14812 9266 14868 9268
rect 14812 9214 14814 9266
rect 14814 9214 14866 9266
rect 14866 9214 14868 9266
rect 14812 9212 14868 9214
rect 14476 8316 14532 8372
rect 13692 7420 13748 7476
rect 14028 8092 14084 8148
rect 13804 6524 13860 6580
rect 13692 5852 13748 5908
rect 13692 3948 13748 4004
rect 14252 5234 14308 5236
rect 14252 5182 14254 5234
rect 14254 5182 14306 5234
rect 14306 5182 14308 5234
rect 14252 5180 14308 5182
rect 13804 3500 13860 3556
rect 14476 3948 14532 4004
rect 14476 3388 14532 3444
rect 15260 13020 15316 13076
rect 15372 12796 15428 12852
rect 15708 13580 15764 13636
rect 15708 13356 15764 13412
rect 15932 13020 15988 13076
rect 15484 12236 15540 12292
rect 15260 11900 15316 11956
rect 15036 10108 15092 10164
rect 15148 10108 15204 10164
rect 15596 11564 15652 11620
rect 15372 9996 15428 10052
rect 15484 10556 15540 10612
rect 15708 11004 15764 11060
rect 15708 10444 15764 10500
rect 15708 9996 15764 10052
rect 15372 9436 15428 9492
rect 16156 11564 16212 11620
rect 16268 13132 16324 13188
rect 16380 11676 16436 11732
rect 16492 12460 16548 12516
rect 16492 11564 16548 11620
rect 16268 11340 16324 11396
rect 16156 11228 16212 11284
rect 16044 11004 16100 11060
rect 15820 9212 15876 9268
rect 15932 10220 15988 10276
rect 15260 8764 15316 8820
rect 15260 8540 15316 8596
rect 15036 7532 15092 7588
rect 15148 6524 15204 6580
rect 15036 5292 15092 5348
rect 14924 4844 14980 4900
rect 15708 8764 15764 8820
rect 15708 8092 15764 8148
rect 15820 8652 15876 8708
rect 15372 7532 15428 7588
rect 15596 5292 15652 5348
rect 15260 5180 15316 5236
rect 15036 4172 15092 4228
rect 15148 4396 15204 4452
rect 14700 3388 14756 3444
rect 15036 3724 15092 3780
rect 13692 3276 13748 3332
rect 13692 2716 13748 2772
rect 13916 3052 13972 3108
rect 13916 2604 13972 2660
rect 13916 2210 13972 2212
rect 13916 2158 13918 2210
rect 13918 2158 13970 2210
rect 13970 2158 13972 2210
rect 13916 2156 13972 2158
rect 13580 588 13636 644
rect 13916 1932 13972 1988
rect 14476 1874 14532 1876
rect 14476 1822 14478 1874
rect 14478 1822 14530 1874
rect 14530 1822 14532 1874
rect 14476 1820 14532 1822
rect 15708 3500 15764 3556
rect 15484 2940 15540 2996
rect 15148 2380 15204 2436
rect 15596 2044 15652 2100
rect 16380 10834 16436 10836
rect 16380 10782 16382 10834
rect 16382 10782 16434 10834
rect 16434 10782 16436 10834
rect 16380 10780 16436 10782
rect 16828 13244 16884 13300
rect 16716 12796 16772 12852
rect 16716 12460 16772 12516
rect 16716 11676 16772 11732
rect 16828 11900 16884 11956
rect 16044 8764 16100 8820
rect 16156 9436 16212 9492
rect 15932 8540 15988 8596
rect 15932 6860 15988 6916
rect 15820 2828 15876 2884
rect 15932 4508 15988 4564
rect 16716 10108 16772 10164
rect 16492 9772 16548 9828
rect 16492 8764 16548 8820
rect 17388 13186 17444 13188
rect 17388 13134 17390 13186
rect 17390 13134 17442 13186
rect 17442 13134 17444 13186
rect 17388 13132 17444 13134
rect 17500 12348 17556 12404
rect 17612 13356 17668 13412
rect 17276 12236 17332 12292
rect 17052 10780 17108 10836
rect 17052 9996 17108 10052
rect 17052 9212 17108 9268
rect 16940 9042 16996 9044
rect 16940 8990 16942 9042
rect 16942 8990 16994 9042
rect 16994 8990 16996 9042
rect 16940 8988 16996 8990
rect 16492 8204 16548 8260
rect 16828 8428 16884 8484
rect 16380 7644 16436 7700
rect 16268 4284 16324 4340
rect 16268 3836 16324 3892
rect 16604 7644 16660 7700
rect 16492 7084 16548 7140
rect 16492 6636 16548 6692
rect 16604 6860 16660 6916
rect 16604 5852 16660 5908
rect 16716 6748 16772 6804
rect 16716 5740 16772 5796
rect 16380 3500 16436 3556
rect 16492 5516 16548 5572
rect 16716 5404 16772 5460
rect 16716 4172 16772 4228
rect 17276 8930 17332 8932
rect 17276 8878 17278 8930
rect 17278 8878 17330 8930
rect 17330 8878 17332 8930
rect 17276 8876 17332 8878
rect 17388 8652 17444 8708
rect 17164 7756 17220 7812
rect 16940 6636 16996 6692
rect 17052 7420 17108 7476
rect 16156 2828 16212 2884
rect 16940 5180 16996 5236
rect 16044 2604 16100 2660
rect 15932 2044 15988 2100
rect 16156 2380 16212 2436
rect 15708 1932 15764 1988
rect 16156 1484 16212 1540
rect 16268 1148 16324 1204
rect 15596 700 15652 756
rect 15820 1036 15876 1092
rect 15820 476 15876 532
rect 15260 364 15316 420
rect 16492 2716 16548 2772
rect 16604 2268 16660 2324
rect 16940 3052 16996 3108
rect 17052 4732 17108 4788
rect 16828 2882 16884 2884
rect 16828 2830 16830 2882
rect 16830 2830 16882 2882
rect 16882 2830 16884 2882
rect 16828 2828 16884 2830
rect 16716 1708 16772 1764
rect 16604 1484 16660 1540
rect 18396 13468 18452 13524
rect 18172 13356 18228 13412
rect 17836 12236 17892 12292
rect 18060 12290 18116 12292
rect 18060 12238 18062 12290
rect 18062 12238 18114 12290
rect 18114 12238 18116 12290
rect 18060 12236 18116 12238
rect 17724 11900 17780 11956
rect 17948 11900 18004 11956
rect 18060 11506 18116 11508
rect 18060 11454 18062 11506
rect 18062 11454 18114 11506
rect 18114 11454 18116 11506
rect 18060 11452 18116 11454
rect 18284 11452 18340 11508
rect 17724 10668 17780 10724
rect 18620 12908 18676 12964
rect 18620 11900 18676 11956
rect 18508 11452 18564 11508
rect 17724 8876 17780 8932
rect 17948 8876 18004 8932
rect 17724 7644 17780 7700
rect 17612 5852 17668 5908
rect 17500 4620 17556 4676
rect 17948 6188 18004 6244
rect 18172 10332 18228 10388
rect 18284 6748 18340 6804
rect 18732 11676 18788 11732
rect 18844 11506 18900 11508
rect 18844 11454 18846 11506
rect 18846 11454 18898 11506
rect 18898 11454 18900 11506
rect 18844 11452 18900 11454
rect 18844 10220 18900 10276
rect 18620 8764 18676 8820
rect 18508 7644 18564 7700
rect 19180 13468 19236 13524
rect 19180 10220 19236 10276
rect 19404 13692 19460 13748
rect 19516 12236 19572 12292
rect 19628 12012 19684 12068
rect 19180 8876 19236 8932
rect 19516 9772 19572 9828
rect 19180 8652 19236 8708
rect 18060 5964 18116 6020
rect 18172 6300 18228 6356
rect 18172 4620 18228 4676
rect 17724 4284 17780 4340
rect 18396 6300 18452 6356
rect 18732 6690 18788 6692
rect 18732 6638 18734 6690
rect 18734 6638 18786 6690
rect 18786 6638 18788 6690
rect 18732 6636 18788 6638
rect 18508 5964 18564 6020
rect 18396 5852 18452 5908
rect 18732 5852 18788 5908
rect 18396 5628 18452 5684
rect 18396 4508 18452 4564
rect 18508 5292 18564 5348
rect 18284 4060 18340 4116
rect 17052 1372 17108 1428
rect 17164 3724 17220 3780
rect 18844 4844 18900 4900
rect 19180 7084 19236 7140
rect 19404 7084 19460 7140
rect 19404 6636 19460 6692
rect 19292 6300 19348 6356
rect 19180 6188 19236 6244
rect 18732 3164 18788 3220
rect 18956 3164 19012 3220
rect 17388 2770 17444 2772
rect 17388 2718 17390 2770
rect 17390 2718 17442 2770
rect 17442 2718 17444 2770
rect 17388 2716 17444 2718
rect 18620 2156 18676 2212
rect 18956 2098 19012 2100
rect 18956 2046 18958 2098
rect 18958 2046 19010 2098
rect 19010 2046 19012 2098
rect 18956 2044 19012 2046
rect 19068 1708 19124 1764
rect 19292 5292 19348 5348
rect 19852 12684 19908 12740
rect 19628 9660 19684 9716
rect 19516 6300 19572 6356
rect 19628 7980 19684 8036
rect 20076 13804 20132 13860
rect 20188 13132 20244 13188
rect 20300 13804 20356 13860
rect 20188 12012 20244 12068
rect 19964 11452 20020 11508
rect 20188 11676 20244 11732
rect 20300 11228 20356 11284
rect 20076 10444 20132 10500
rect 20076 9884 20132 9940
rect 20188 10332 20244 10388
rect 19852 9826 19908 9828
rect 19852 9774 19854 9826
rect 19854 9774 19906 9826
rect 19906 9774 19908 9826
rect 19852 9772 19908 9774
rect 19964 9212 20020 9268
rect 20188 9212 20244 9268
rect 20860 12684 20916 12740
rect 21308 13468 21364 13524
rect 21532 13468 21588 13524
rect 21196 13186 21252 13188
rect 21196 13134 21198 13186
rect 21198 13134 21250 13186
rect 21250 13134 21252 13186
rect 21196 13132 21252 13134
rect 21644 12796 21700 12852
rect 21196 12684 21252 12740
rect 20636 11900 20692 11956
rect 19964 8876 20020 8932
rect 20076 8204 20132 8260
rect 21196 11564 21252 11620
rect 21308 11340 21364 11396
rect 21308 10332 21364 10388
rect 20972 8876 21028 8932
rect 21196 8876 21252 8932
rect 20748 8764 20804 8820
rect 19852 6076 19908 6132
rect 19628 2604 19684 2660
rect 20972 8258 21028 8260
rect 20972 8206 20974 8258
rect 20974 8206 21026 8258
rect 21026 8206 21028 8258
rect 20972 8204 21028 8206
rect 20524 6860 20580 6916
rect 20076 5292 20132 5348
rect 20300 5292 20356 5348
rect 20076 4844 20132 4900
rect 20300 4844 20356 4900
rect 19516 2156 19572 2212
rect 19180 1484 19236 1540
rect 18620 1372 18676 1428
rect 17164 1260 17220 1316
rect 16492 588 16548 644
rect 13244 28 13300 84
rect 19964 4284 20020 4340
rect 21644 12402 21700 12404
rect 21644 12350 21646 12402
rect 21646 12350 21698 12402
rect 21698 12350 21700 12402
rect 21644 12348 21700 12350
rect 21644 12012 21700 12068
rect 21644 11564 21700 11620
rect 21532 11452 21588 11508
rect 21644 9772 21700 9828
rect 21532 6972 21588 7028
rect 21532 6636 21588 6692
rect 21308 5068 21364 5124
rect 21420 6300 21476 6356
rect 21308 4060 21364 4116
rect 21308 3612 21364 3668
rect 20412 3388 20468 3444
rect 20300 3276 20356 3332
rect 20300 2940 20356 2996
rect 20188 2098 20244 2100
rect 20188 2046 20190 2098
rect 20190 2046 20242 2098
rect 20242 2046 20244 2098
rect 20188 2044 20244 2046
rect 19852 1820 19908 1876
rect 19740 1036 19796 1092
rect 19628 476 19684 532
rect 19852 700 19908 756
rect 20972 3052 21028 3108
rect 21084 3388 21140 3444
rect 20748 2940 20804 2996
rect 20524 1932 20580 1988
rect 20524 1708 20580 1764
rect 20860 1932 20916 1988
rect 20076 700 20132 756
rect 20636 1148 20692 1204
rect 19852 476 19908 532
rect 21532 5292 21588 5348
rect 21532 4284 21588 4340
rect 22204 12348 22260 12404
rect 22316 13468 22372 13524
rect 21980 10332 22036 10388
rect 22204 10332 22260 10388
rect 21868 8428 21924 8484
rect 21868 7308 21924 7364
rect 21756 6636 21812 6692
rect 21868 6076 21924 6132
rect 21644 3388 21700 3444
rect 21756 5068 21812 5124
rect 21308 3276 21364 3332
rect 21868 4956 21924 5012
rect 21868 4620 21924 4676
rect 21868 4284 21924 4340
rect 21756 2156 21812 2212
rect 22428 13132 22484 13188
rect 22540 13468 22596 13524
rect 22428 12236 22484 12292
rect 22092 9548 22148 9604
rect 22204 9154 22260 9156
rect 22204 9102 22206 9154
rect 22206 9102 22258 9154
rect 22258 9102 22260 9154
rect 22204 9100 22260 9102
rect 22092 8540 22148 8596
rect 22092 8204 22148 8260
rect 22876 13074 22932 13076
rect 22876 13022 22878 13074
rect 22878 13022 22930 13074
rect 22930 13022 22932 13074
rect 22876 13020 22932 13022
rect 23212 13580 23268 13636
rect 22764 11564 22820 11620
rect 22652 10780 22708 10836
rect 22764 10220 22820 10276
rect 22876 10108 22932 10164
rect 22988 9772 23044 9828
rect 22764 9100 22820 9156
rect 22540 8652 22596 8708
rect 22988 8652 23044 8708
rect 23100 9548 23156 9604
rect 22876 8428 22932 8484
rect 22316 6972 22372 7028
rect 22428 7420 22484 7476
rect 22092 6524 22148 6580
rect 22316 6524 22372 6580
rect 22316 6300 22372 6356
rect 22764 6690 22820 6692
rect 22764 6638 22766 6690
rect 22766 6638 22818 6690
rect 22818 6638 22820 6690
rect 22764 6636 22820 6638
rect 22540 5404 22596 5460
rect 21980 2044 22036 2100
rect 21084 1372 21140 1428
rect 21196 1820 21252 1876
rect 22988 7084 23044 7140
rect 22988 4956 23044 5012
rect 23324 13020 23380 13076
rect 23548 12348 23604 12404
rect 23660 13244 23716 13300
rect 23996 13692 24052 13748
rect 24444 13580 24500 13636
rect 24892 13804 24948 13860
rect 24668 13468 24724 13524
rect 24892 13468 24948 13524
rect 24332 13356 24388 13412
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 24220 13020 24276 13076
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 24220 12460 24276 12516
rect 24332 12402 24388 12404
rect 24332 12350 24334 12402
rect 24334 12350 24386 12402
rect 24386 12350 24388 12402
rect 24332 12348 24388 12350
rect 23436 12066 23492 12068
rect 23436 12014 23438 12066
rect 23438 12014 23490 12066
rect 23490 12014 23492 12066
rect 23436 12012 23492 12014
rect 25004 12348 25060 12404
rect 24108 11676 24164 11732
rect 24220 12012 24276 12068
rect 23324 11618 23380 11620
rect 23324 11566 23326 11618
rect 23326 11566 23378 11618
rect 23378 11566 23380 11618
rect 23324 11564 23380 11566
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23436 10834 23492 10836
rect 23436 10782 23438 10834
rect 23438 10782 23490 10834
rect 23490 10782 23492 10834
rect 23436 10780 23492 10782
rect 23324 10668 23380 10724
rect 23548 10668 23604 10724
rect 23324 9772 23380 9828
rect 23436 9436 23492 9492
rect 23548 10332 23604 10388
rect 24444 12012 24500 12068
rect 24332 11788 24388 11844
rect 25564 14028 25620 14084
rect 25340 13692 25396 13748
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 25116 11788 25172 11844
rect 25228 12572 25284 12628
rect 24672 11732 24728 11734
rect 25116 11618 25172 11620
rect 25116 11566 25118 11618
rect 25118 11566 25170 11618
rect 25170 11566 25172 11618
rect 25116 11564 25172 11566
rect 24332 10892 24388 10948
rect 25228 11116 25284 11172
rect 25340 11004 25396 11060
rect 24332 10220 24388 10276
rect 25004 10780 25060 10836
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24444 9772 24500 9828
rect 23660 9324 23716 9380
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 25340 10780 25396 10836
rect 25228 10668 25284 10724
rect 25116 9938 25172 9940
rect 25116 9886 25118 9938
rect 25118 9886 25170 9938
rect 25170 9886 25172 9938
rect 25116 9884 25172 9886
rect 25788 13580 25844 13636
rect 25452 10108 25508 10164
rect 25676 11452 25732 11508
rect 25900 10892 25956 10948
rect 26012 12460 26068 12516
rect 25676 9772 25732 9828
rect 25004 9324 25060 9380
rect 24332 9212 24388 9268
rect 24108 8652 24164 8708
rect 24464 8650 24520 8652
rect 24332 8540 24388 8596
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24892 8652 24948 8708
rect 24672 8596 24728 8598
rect 23436 7868 23492 7924
rect 23772 8316 23828 8372
rect 23660 7756 23716 7812
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24332 7868 24388 7924
rect 24012 7812 24068 7814
rect 23324 7586 23380 7588
rect 23324 7534 23326 7586
rect 23326 7534 23378 7586
rect 23378 7534 23380 7586
rect 23324 7532 23380 7534
rect 23884 7474 23940 7476
rect 23884 7422 23886 7474
rect 23886 7422 23938 7474
rect 23938 7422 23940 7474
rect 23884 7420 23940 7422
rect 24892 7196 24948 7252
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 25564 9324 25620 9380
rect 25340 9100 25396 9156
rect 25228 8204 25284 8260
rect 25116 8092 25172 8148
rect 25340 7644 25396 7700
rect 25340 7308 25396 7364
rect 25116 6860 25172 6916
rect 23324 6690 23380 6692
rect 23324 6638 23326 6690
rect 23326 6638 23378 6690
rect 23378 6638 23380 6690
rect 23324 6636 23380 6638
rect 23548 6300 23604 6356
rect 24444 6412 24500 6468
rect 23660 6188 23716 6244
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24220 6188 24276 6244
rect 23772 6018 23828 6020
rect 23772 5966 23774 6018
rect 23774 5966 23826 6018
rect 23826 5966 23828 6018
rect 23772 5964 23828 5966
rect 23548 5516 23604 5572
rect 24332 5964 24388 6020
rect 25228 5852 25284 5908
rect 24220 5516 24276 5572
rect 24464 5514 24520 5516
rect 24332 5404 24388 5460
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 24892 5404 24948 5460
rect 24892 5122 24948 5124
rect 24892 5070 24894 5122
rect 24894 5070 24946 5122
rect 24946 5070 24948 5122
rect 24892 5068 24948 5070
rect 23548 4732 23604 4788
rect 23804 4730 23860 4732
rect 23436 4620 23492 4676
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 22876 2156 22932 2212
rect 23324 4396 23380 4452
rect 24332 4620 24388 4676
rect 23548 4396 23604 4452
rect 21756 1820 21812 1876
rect 22204 1708 22260 1764
rect 21308 1484 21364 1540
rect 21308 1148 21364 1204
rect 21196 924 21252 980
rect 21756 812 21812 868
rect 21980 924 22036 980
rect 22428 812 22484 868
rect 20860 476 20916 532
rect 22540 588 22596 644
rect 23100 588 23156 644
rect 25228 4620 25284 4676
rect 24556 4172 24612 4228
rect 24332 3948 24388 4004
rect 25116 3948 25172 4004
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 25452 6972 25508 7028
rect 25676 5180 25732 5236
rect 25340 3724 25396 3780
rect 24556 3388 24612 3444
rect 23660 3052 23716 3108
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24220 3164 24276 3220
rect 25116 3388 25172 3444
rect 24012 3108 24068 3110
rect 24332 3052 24388 3108
rect 23548 2828 23604 2884
rect 24332 2380 24388 2436
rect 24464 2378 24520 2380
rect 23996 2268 24052 2324
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24892 2380 24948 2436
rect 23548 1596 23604 1652
rect 23804 1594 23860 1596
rect 23660 1484 23716 1540
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24220 1484 24276 1540
rect 24332 812 24388 868
rect 24464 810 24520 812
rect 23324 588 23380 644
rect 24220 700 24276 756
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24892 812 24948 868
rect 24672 756 24728 758
rect 25564 2716 25620 2772
rect 25452 1484 25508 1540
rect 26236 12236 26292 12292
rect 26348 12348 26404 12404
rect 26348 10386 26404 10388
rect 26348 10334 26350 10386
rect 26350 10334 26402 10386
rect 26402 10334 26404 10386
rect 26348 10332 26404 10334
rect 26236 9714 26292 9716
rect 26236 9662 26238 9714
rect 26238 9662 26290 9714
rect 26290 9662 26292 9714
rect 26236 9660 26292 9662
rect 26012 6636 26068 6692
rect 26124 5628 26180 5684
rect 25788 4732 25844 4788
rect 25900 4396 25956 4452
rect 26124 4396 26180 4452
rect 25676 1484 25732 1540
rect 23660 476 23716 532
rect 24108 476 24164 532
rect 23772 252 23828 308
rect 23548 28 23604 84
rect 25228 700 25284 756
rect 24220 252 24276 308
rect 26908 13132 26964 13188
rect 27020 12684 27076 12740
rect 26684 10332 26740 10388
rect 26684 10108 26740 10164
rect 26908 10108 26964 10164
rect 26796 9826 26852 9828
rect 26796 9774 26798 9826
rect 26798 9774 26850 9826
rect 26850 9774 26852 9826
rect 26796 9772 26852 9774
rect 26572 8764 26628 8820
rect 26796 8204 26852 8260
rect 26572 8092 26628 8148
rect 27020 8092 27076 8148
rect 26684 7868 26740 7924
rect 26572 6860 26628 6916
rect 26796 6860 26852 6916
rect 27020 3836 27076 3892
rect 27244 12684 27300 12740
rect 27692 12684 27748 12740
rect 27356 11452 27412 11508
rect 27244 10892 27300 10948
rect 27468 9996 27524 10052
rect 27468 9772 27524 9828
rect 27356 8428 27412 8484
rect 27692 11788 27748 11844
rect 28252 12348 28308 12404
rect 28028 11788 28084 11844
rect 27692 10722 27748 10724
rect 27692 10670 27694 10722
rect 27694 10670 27746 10722
rect 27746 10670 27748 10722
rect 27692 10668 27748 10670
rect 27692 10050 27748 10052
rect 27692 9998 27694 10050
rect 27694 9998 27746 10050
rect 27746 9998 27748 10050
rect 27692 9996 27748 9998
rect 28476 11676 28532 11732
rect 28364 9772 28420 9828
rect 27916 9212 27972 9268
rect 27804 8764 27860 8820
rect 27692 8652 27748 8708
rect 27804 8540 27860 8596
rect 27804 8316 27860 8372
rect 27580 7420 27636 7476
rect 27244 6636 27300 6692
rect 27244 4284 27300 4340
rect 27580 6412 27636 6468
rect 27580 3276 27636 3332
rect 27692 5516 27748 5572
rect 26572 3164 26628 3220
rect 26460 2380 26516 2436
rect 26684 2716 26740 2772
rect 26684 2380 26740 2436
rect 26348 1932 26404 1988
rect 26796 2044 26852 2100
rect 26124 252 26180 308
rect 26236 1260 26292 1316
rect 27804 3666 27860 3668
rect 27804 3614 27806 3666
rect 27806 3614 27858 3666
rect 27858 3614 27860 3666
rect 27804 3612 27860 3614
rect 28924 12572 28980 12628
rect 29036 13132 29092 13188
rect 28700 11900 28756 11956
rect 28700 10108 28756 10164
rect 28476 7980 28532 8036
rect 29036 10332 29092 10388
rect 28924 9660 28980 9716
rect 28812 7308 28868 7364
rect 29036 6748 29092 6804
rect 28476 6524 28532 6580
rect 28028 6188 28084 6244
rect 28476 4508 28532 4564
rect 29260 13804 29316 13860
rect 29484 12012 29540 12068
rect 29596 11564 29652 11620
rect 29148 5740 29204 5796
rect 29260 11004 29316 11060
rect 29036 4508 29092 4564
rect 28028 4172 28084 4228
rect 30268 12572 30324 12628
rect 30380 12124 30436 12180
rect 29820 8764 29876 8820
rect 30044 10108 30100 10164
rect 29932 8258 29988 8260
rect 29932 8206 29934 8258
rect 29934 8206 29986 8258
rect 29986 8206 29988 8258
rect 29932 8204 29988 8206
rect 29484 8146 29540 8148
rect 29484 8094 29486 8146
rect 29486 8094 29538 8146
rect 29538 8094 29540 8146
rect 29484 8092 29540 8094
rect 29372 6860 29428 6916
rect 29484 6076 29540 6132
rect 29596 7756 29652 7812
rect 29372 5292 29428 5348
rect 30380 11564 30436 11620
rect 30716 12124 30772 12180
rect 30604 11954 30660 11956
rect 30604 11902 30606 11954
rect 30606 11902 30658 11954
rect 30658 11902 30660 11954
rect 30604 11900 30660 11902
rect 30268 7756 30324 7812
rect 30380 7420 30436 7476
rect 30268 7196 30324 7252
rect 29932 6578 29988 6580
rect 29932 6526 29934 6578
rect 29934 6526 29986 6578
rect 29986 6526 29988 6578
rect 29932 6524 29988 6526
rect 29596 5292 29652 5348
rect 28028 3612 28084 3668
rect 29820 3554 29876 3556
rect 29820 3502 29822 3554
rect 29822 3502 29874 3554
rect 29874 3502 29876 3554
rect 29820 3500 29876 3502
rect 29372 3388 29428 3444
rect 27692 1932 27748 1988
rect 28588 2716 28644 2772
rect 27020 1372 27076 1428
rect 28588 1036 28644 1092
rect 28700 1260 28756 1316
rect 27020 812 27076 868
rect 26796 140 26852 196
rect 31388 13916 31444 13972
rect 31612 13916 31668 13972
rect 31836 13132 31892 13188
rect 31612 12908 31668 12964
rect 31052 11564 31108 11620
rect 31052 11340 31108 11396
rect 31164 10892 31220 10948
rect 31276 11788 31332 11844
rect 31052 10332 31108 10388
rect 31164 9772 31220 9828
rect 31164 9436 31220 9492
rect 31052 7420 31108 7476
rect 31164 8204 31220 8260
rect 30940 7308 30996 7364
rect 30604 6300 30660 6356
rect 30380 4172 30436 4228
rect 30604 5180 30660 5236
rect 30268 4060 30324 4116
rect 30268 2604 30324 2660
rect 30380 3276 30436 3332
rect 30156 2380 30212 2436
rect 30492 2604 30548 2660
rect 30492 2268 30548 2324
rect 30380 1148 30436 1204
rect 30268 924 30324 980
rect 30268 364 30324 420
rect 29372 252 29428 308
rect 24444 28 24500 84
rect 31388 11564 31444 11620
rect 31388 10332 31444 10388
rect 31948 12684 32004 12740
rect 31948 12236 32004 12292
rect 32284 13692 32340 13748
rect 32172 12012 32228 12068
rect 31948 8764 32004 8820
rect 31500 6860 31556 6916
rect 31724 8428 31780 8484
rect 31724 5964 31780 6020
rect 31836 6636 31892 6692
rect 31836 5852 31892 5908
rect 32732 10556 32788 10612
rect 32508 10332 32564 10388
rect 32172 8652 32228 8708
rect 32060 8428 32116 8484
rect 32396 8370 32452 8372
rect 32396 8318 32398 8370
rect 32398 8318 32450 8370
rect 32450 8318 32452 8370
rect 32396 8316 32452 8318
rect 32060 7868 32116 7924
rect 32060 6860 32116 6916
rect 32284 7756 32340 7812
rect 32172 4396 32228 4452
rect 32172 3164 32228 3220
rect 31836 2940 31892 2996
rect 32732 7868 32788 7924
rect 32732 7084 32788 7140
rect 33068 11340 33124 11396
rect 33068 10556 33124 10612
rect 32956 7980 33012 8036
rect 33292 13356 33348 13412
rect 33404 12460 33460 12516
rect 33628 13244 33684 13300
rect 33628 11676 33684 11732
rect 33516 11228 33572 11284
rect 33628 11340 33684 11396
rect 33180 7532 33236 7588
rect 33404 8428 33460 8484
rect 33852 11116 33908 11172
rect 33964 13804 34020 13860
rect 33628 9212 33684 9268
rect 33852 10220 33908 10276
rect 33628 8428 33684 8484
rect 33628 8204 33684 8260
rect 33404 7532 33460 7588
rect 33516 7756 33572 7812
rect 34076 11564 34132 11620
rect 33964 8988 34020 9044
rect 34076 9212 34132 9268
rect 33852 7756 33908 7812
rect 33628 6524 33684 6580
rect 33852 7532 33908 7588
rect 33852 6524 33908 6580
rect 32844 5628 32900 5684
rect 33404 5628 33460 5684
rect 33068 4508 33124 4564
rect 33180 4284 33236 4340
rect 32956 4172 33012 4228
rect 32284 2156 32340 2212
rect 32396 3164 32452 3220
rect 32844 2492 32900 2548
rect 33516 3666 33572 3668
rect 33516 3614 33518 3666
rect 33518 3614 33570 3666
rect 33570 3614 33572 3666
rect 33516 3612 33572 3614
rect 33404 2828 33460 2884
rect 33180 2380 33236 2436
rect 33404 2492 33460 2548
rect 32396 1484 32452 1540
rect 31276 1148 31332 1204
rect 34524 12012 34580 12068
rect 34412 11900 34468 11956
rect 34412 10108 34468 10164
rect 34636 10108 34692 10164
rect 34300 8764 34356 8820
rect 34636 7084 34692 7140
rect 34524 6188 34580 6244
rect 35196 13804 35252 13860
rect 35308 11788 35364 11844
rect 34860 10668 34916 10724
rect 34972 10892 35028 10948
rect 35308 10668 35364 10724
rect 36092 13020 36148 13076
rect 36764 13356 36820 13412
rect 36540 13244 36596 13300
rect 35532 11788 35588 11844
rect 35644 12572 35700 12628
rect 36316 12348 36372 12404
rect 35644 11564 35700 11620
rect 35756 12236 35812 12292
rect 35420 9996 35476 10052
rect 34972 9436 35028 9492
rect 35084 8764 35140 8820
rect 35308 9548 35364 9604
rect 35420 8540 35476 8596
rect 35420 7532 35476 7588
rect 35308 7084 35364 7140
rect 35308 6860 35364 6916
rect 34748 6076 34804 6132
rect 35084 6188 35140 6244
rect 34076 5516 34132 5572
rect 33628 924 33684 980
rect 34524 2828 34580 2884
rect 35308 4508 35364 4564
rect 36204 10780 36260 10836
rect 36540 13020 36596 13076
rect 36876 12684 36932 12740
rect 37436 13692 37492 13748
rect 37324 13580 37380 13636
rect 37660 13468 37716 13524
rect 37212 12684 37268 12740
rect 37996 13804 38052 13860
rect 38108 13244 38164 13300
rect 37884 12348 37940 12404
rect 37548 12066 37604 12068
rect 37548 12014 37550 12066
rect 37550 12014 37602 12066
rect 37602 12014 37604 12066
rect 37548 12012 37604 12014
rect 36876 11004 36932 11060
rect 37100 11788 37156 11844
rect 36764 8428 36820 8484
rect 36988 8876 37044 8932
rect 36988 8316 37044 8372
rect 35756 4172 35812 4228
rect 36092 6524 36148 6580
rect 35532 2380 35588 2436
rect 35420 2044 35476 2100
rect 35420 1596 35476 1652
rect 35084 1372 35140 1428
rect 35532 588 35588 644
rect 34524 476 34580 532
rect 33628 140 33684 196
rect 36652 3276 36708 3332
rect 36652 2716 36708 2772
rect 36988 6748 37044 6804
rect 36988 6300 37044 6356
rect 36988 6076 37044 6132
rect 36876 5516 36932 5572
rect 36988 4620 37044 4676
rect 37324 11788 37380 11844
rect 37548 11564 37604 11620
rect 37324 9212 37380 9268
rect 37436 11116 37492 11172
rect 37212 8204 37268 8260
rect 37324 6524 37380 6580
rect 37324 4956 37380 5012
rect 37212 4732 37268 4788
rect 37548 6188 37604 6244
rect 37436 3612 37492 3668
rect 37884 12124 37940 12180
rect 38108 11394 38164 11396
rect 38108 11342 38110 11394
rect 38110 11342 38162 11394
rect 38162 11342 38164 11394
rect 38108 11340 38164 11342
rect 37884 10556 37940 10612
rect 37996 11228 38052 11284
rect 37772 5682 37828 5684
rect 37772 5630 37774 5682
rect 37774 5630 37826 5682
rect 37826 5630 37828 5682
rect 37772 5628 37828 5630
rect 37660 2940 37716 2996
rect 37884 5180 37940 5236
rect 37212 2828 37268 2884
rect 37660 2658 37716 2660
rect 37660 2606 37662 2658
rect 37662 2606 37714 2658
rect 37714 2606 37716 2658
rect 37660 2604 37716 2606
rect 38444 12850 38500 12852
rect 38444 12798 38446 12850
rect 38446 12798 38498 12850
rect 38498 12798 38500 12850
rect 38444 12796 38500 12798
rect 38556 12572 38612 12628
rect 38668 12684 38724 12740
rect 38332 12460 38388 12516
rect 38780 12124 38836 12180
rect 38892 13804 38948 13860
rect 39228 13244 39284 13300
rect 39340 13804 39396 13860
rect 39004 13020 39060 13076
rect 38220 11228 38276 11284
rect 38332 9100 38388 9156
rect 38780 10498 38836 10500
rect 38780 10446 38782 10498
rect 38782 10446 38834 10498
rect 38834 10446 38836 10498
rect 38780 10444 38836 10446
rect 39340 12684 39396 12740
rect 39116 11900 39172 11956
rect 39340 12348 39396 12404
rect 39116 11228 39172 11284
rect 39452 12236 39508 12292
rect 39564 13132 39620 13188
rect 39452 10332 39508 10388
rect 39116 9042 39172 9044
rect 39116 8990 39118 9042
rect 39118 8990 39170 9042
rect 39170 8990 39172 9042
rect 39116 8988 39172 8990
rect 38556 7532 38612 7588
rect 37996 4284 38052 4340
rect 38332 2828 38388 2884
rect 37884 1372 37940 1428
rect 36876 700 36932 756
rect 36764 140 36820 196
rect 39004 7420 39060 7476
rect 38668 5906 38724 5908
rect 38668 5854 38670 5906
rect 38670 5854 38722 5906
rect 38722 5854 38724 5906
rect 38668 5852 38724 5854
rect 38892 5122 38948 5124
rect 38892 5070 38894 5122
rect 38894 5070 38946 5122
rect 38946 5070 38948 5122
rect 38892 5068 38948 5070
rect 38780 3948 38836 4004
rect 39116 6748 39172 6804
rect 39340 8316 39396 8372
rect 39228 5794 39284 5796
rect 39228 5742 39230 5794
rect 39230 5742 39282 5794
rect 39282 5742 39284 5794
rect 39228 5740 39284 5742
rect 39004 3724 39060 3780
rect 38780 3612 38836 3668
rect 38892 3276 38948 3332
rect 39452 5122 39508 5124
rect 39452 5070 39454 5122
rect 39454 5070 39506 5122
rect 39506 5070 39508 5122
rect 39452 5068 39508 5070
rect 39676 12908 39732 12964
rect 39788 13356 39844 13412
rect 39676 12684 39732 12740
rect 39900 12348 39956 12404
rect 40012 13692 40068 13748
rect 40124 13132 40180 13188
rect 41244 13468 41300 13524
rect 42364 13244 42420 13300
rect 40348 12908 40404 12964
rect 40236 12012 40292 12068
rect 40684 11564 40740 11620
rect 40796 12572 40852 12628
rect 41580 12460 41636 12516
rect 40908 12236 40964 12292
rect 40236 9772 40292 9828
rect 39564 4956 39620 5012
rect 39676 7196 39732 7252
rect 39676 3500 39732 3556
rect 39676 2098 39732 2100
rect 39676 2046 39678 2098
rect 39678 2046 39730 2098
rect 39730 2046 39732 2098
rect 39676 2044 39732 2046
rect 39116 1596 39172 1652
rect 30492 28 30548 84
rect 39900 6076 39956 6132
rect 40460 8988 40516 9044
rect 40460 6524 40516 6580
rect 40348 5516 40404 5572
rect 40572 5404 40628 5460
rect 41132 12124 41188 12180
rect 40908 10556 40964 10612
rect 40796 6524 40852 6580
rect 40908 9548 40964 9604
rect 40684 4732 40740 4788
rect 40236 4620 40292 4676
rect 40348 4508 40404 4564
rect 41916 11676 41972 11732
rect 41804 10108 41860 10164
rect 43708 13074 43764 13076
rect 43708 13022 43710 13074
rect 43710 13022 43762 13074
rect 43762 13022 43764 13074
rect 43708 13020 43764 13022
rect 42588 12796 42644 12852
rect 42476 12348 42532 12404
rect 42140 11228 42196 11284
rect 41020 8092 41076 8148
rect 41244 8092 41300 8148
rect 40908 4396 40964 4452
rect 40348 3164 40404 3220
rect 40236 2716 40292 2772
rect 42028 7868 42084 7924
rect 42252 9714 42308 9716
rect 42252 9662 42254 9714
rect 42254 9662 42306 9714
rect 42306 9662 42308 9714
rect 42252 9660 42308 9662
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 42924 8540 42980 8596
rect 43484 11004 43540 11060
rect 43148 6300 43204 6356
rect 43372 10556 43428 10612
rect 42140 5628 42196 5684
rect 41244 2604 41300 2660
rect 42812 4060 42868 4116
rect 43372 2044 43428 2100
rect 42252 1260 42308 1316
rect 41020 924 41076 980
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 43932 10444 43988 10500
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 51100 13916 51156 13972
rect 50540 13468 50596 13524
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 45052 13186 45108 13188
rect 45052 13134 45054 13186
rect 45054 13134 45106 13186
rect 45106 13134 45108 13186
rect 45052 13132 45108 13134
rect 48076 13020 48132 13076
rect 45164 12012 45220 12068
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 44268 9996 44324 10052
rect 44492 9714 44548 9716
rect 44492 9662 44494 9714
rect 44494 9662 44546 9714
rect 44546 9662 44548 9714
rect 44492 9660 44548 9662
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 43596 7084 43652 7140
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 44828 8316 44884 8372
rect 45948 10668 46004 10724
rect 45276 9772 45332 9828
rect 45164 8204 45220 8260
rect 45388 8764 45444 8820
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 45388 6636 45444 6692
rect 45500 8428 45556 8484
rect 44604 6524 44660 6580
rect 44268 5852 44324 5908
rect 43932 5628 43988 5684
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 45052 5180 45108 5236
rect 43932 4956 43988 5012
rect 45500 4956 45556 5012
rect 45836 4844 45892 4900
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 44156 4226 44212 4228
rect 44156 4174 44158 4226
rect 44158 4174 44210 4226
rect 44210 4174 44212 4226
rect 44156 4172 44212 4174
rect 44464 3946 44520 3948
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 44716 3554 44772 3556
rect 44716 3502 44718 3554
rect 44718 3502 44770 3554
rect 44770 3502 44772 3554
rect 44716 3500 44772 3502
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 44268 1874 44324 1876
rect 44268 1822 44270 1874
rect 44270 1822 44322 1874
rect 44322 1822 44324 1874
rect 44268 1820 44324 1822
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 45276 3724 45332 3780
rect 48188 12572 48244 12628
rect 47180 9548 47236 9604
rect 47292 12236 47348 12292
rect 46956 8988 47012 9044
rect 46620 7980 46676 8036
rect 46284 6636 46340 6692
rect 45948 4732 46004 4788
rect 46172 5740 46228 5796
rect 45388 2770 45444 2772
rect 45388 2718 45390 2770
rect 45390 2718 45442 2770
rect 45442 2718 45444 2770
rect 45388 2716 45444 2718
rect 46172 2716 46228 2772
rect 46396 3612 46452 3668
rect 46732 4284 46788 4340
rect 46620 3612 46676 3668
rect 46396 3442 46452 3444
rect 46396 3390 46398 3442
rect 46398 3390 46450 3442
rect 46450 3390 46452 3442
rect 46396 3388 46452 3390
rect 47740 11900 47796 11956
rect 47628 10780 47684 10836
rect 48300 10498 48356 10500
rect 48300 10446 48302 10498
rect 48302 10446 48354 10498
rect 48354 10446 48356 10498
rect 48300 10444 48356 10446
rect 47740 8818 47796 8820
rect 47740 8766 47742 8818
rect 47742 8766 47794 8818
rect 47794 8766 47796 8818
rect 47740 8764 47796 8766
rect 48300 8652 48356 8708
rect 47628 8204 47684 8260
rect 48860 11116 48916 11172
rect 48972 11228 49028 11284
rect 48972 9660 49028 9716
rect 47404 7532 47460 7588
rect 48636 8258 48692 8260
rect 48636 8206 48638 8258
rect 48638 8206 48690 8258
rect 48690 8206 48692 8258
rect 48636 8204 48692 8206
rect 48748 7308 48804 7364
rect 48524 6860 48580 6916
rect 47404 5964 47460 6020
rect 48524 6412 48580 6468
rect 48076 5682 48132 5684
rect 48076 5630 48078 5682
rect 48078 5630 48130 5682
rect 48130 5630 48132 5682
rect 48076 5628 48132 5630
rect 48860 6690 48916 6692
rect 48860 6638 48862 6690
rect 48862 6638 48914 6690
rect 48914 6638 48916 6690
rect 48860 6636 48916 6638
rect 48748 4956 48804 5012
rect 48188 4508 48244 4564
rect 49756 12124 49812 12180
rect 50204 12066 50260 12068
rect 50204 12014 50206 12066
rect 50206 12014 50258 12066
rect 50258 12014 50260 12066
rect 50204 12012 50260 12014
rect 49644 11788 49700 11844
rect 50428 11394 50484 11396
rect 50428 11342 50430 11394
rect 50430 11342 50482 11394
rect 50482 11342 50484 11394
rect 50428 11340 50484 11342
rect 49868 11282 49924 11284
rect 49868 11230 49870 11282
rect 49870 11230 49922 11282
rect 49922 11230 49924 11282
rect 49868 11228 49924 11230
rect 50204 10610 50260 10612
rect 50204 10558 50206 10610
rect 50206 10558 50258 10610
rect 50258 10558 50260 10610
rect 50204 10556 50260 10558
rect 49644 10332 49700 10388
rect 50428 9938 50484 9940
rect 50428 9886 50430 9938
rect 50430 9886 50482 9938
rect 50482 9886 50484 9938
rect 50428 9884 50484 9886
rect 49868 9714 49924 9716
rect 49868 9662 49870 9714
rect 49870 9662 49922 9714
rect 49922 9662 49924 9714
rect 49868 9660 49924 9662
rect 50540 9660 50596 9716
rect 50652 10444 50708 10500
rect 49644 9266 49700 9268
rect 49644 9214 49646 9266
rect 49646 9214 49698 9266
rect 49698 9214 49700 9266
rect 49644 9212 49700 9214
rect 50204 8930 50260 8932
rect 50204 8878 50206 8930
rect 50206 8878 50258 8930
rect 50258 8878 50260 8930
rect 50204 8876 50260 8878
rect 50316 8652 50372 8708
rect 49084 6748 49140 6804
rect 49084 5404 49140 5460
rect 48860 3836 48916 3892
rect 48860 3666 48916 3668
rect 48860 3614 48862 3666
rect 48862 3614 48914 3666
rect 48914 3614 48916 3666
rect 48860 3612 48916 3614
rect 47740 3276 47796 3332
rect 46956 2940 47012 2996
rect 47068 2828 47124 2884
rect 48076 2882 48132 2884
rect 48076 2830 48078 2882
rect 48078 2830 48130 2882
rect 48130 2830 48132 2882
rect 48076 2828 48132 2830
rect 48748 2770 48804 2772
rect 48748 2718 48750 2770
rect 48750 2718 48802 2770
rect 48802 2718 48804 2770
rect 48748 2716 48804 2718
rect 46284 2492 46340 2548
rect 45948 2044 46004 2100
rect 47516 2380 47572 2436
rect 48860 2098 48916 2100
rect 48860 2046 48862 2098
rect 48862 2046 48914 2098
rect 48914 2046 48916 2098
rect 48860 2044 48916 2046
rect 47068 1708 47124 1764
rect 47180 1090 47236 1092
rect 47180 1038 47182 1090
rect 47182 1038 47234 1090
rect 47234 1038 47236 1090
rect 47180 1036 47236 1038
rect 49308 5906 49364 5908
rect 49308 5854 49310 5906
rect 49310 5854 49362 5906
rect 49362 5854 49364 5906
rect 49308 5852 49364 5854
rect 49980 8146 50036 8148
rect 49980 8094 49982 8146
rect 49982 8094 50034 8146
rect 50034 8094 50036 8146
rect 49980 8092 50036 8094
rect 49532 7420 49588 7476
rect 49644 6748 49700 6804
rect 49868 6018 49924 6020
rect 49868 5966 49870 6018
rect 49870 5966 49922 6018
rect 49922 5966 49924 6018
rect 49868 5964 49924 5966
rect 49756 5852 49812 5908
rect 50204 5292 50260 5348
rect 49420 5180 49476 5236
rect 49644 5122 49700 5124
rect 49644 5070 49646 5122
rect 49646 5070 49698 5122
rect 49698 5070 49700 5122
rect 49644 5068 49700 5070
rect 50204 4732 50260 4788
rect 49420 3612 49476 3668
rect 49196 3388 49252 3444
rect 49868 3442 49924 3444
rect 49868 3390 49870 3442
rect 49870 3390 49922 3442
rect 49922 3390 49924 3442
rect 49868 3388 49924 3390
rect 50428 8370 50484 8372
rect 50428 8318 50430 8370
rect 50430 8318 50482 8370
rect 50482 8318 50484 8370
rect 50428 8316 50484 8318
rect 50988 9436 51044 9492
rect 51212 13580 51268 13636
rect 51212 10780 51268 10836
rect 51436 9884 51492 9940
rect 51100 9212 51156 9268
rect 51436 8988 51492 9044
rect 50988 8540 51044 8596
rect 50876 8092 50932 8148
rect 51436 7644 51492 7700
rect 51212 6300 51268 6356
rect 50764 5404 50820 5460
rect 51212 5404 51268 5460
rect 51100 5068 51156 5124
rect 51100 4508 51156 4564
rect 51212 4956 51268 5012
rect 50428 3724 50484 3780
rect 49420 2658 49476 2660
rect 49420 2606 49422 2658
rect 49422 2606 49474 2658
rect 49474 2606 49476 2658
rect 49420 2604 49476 2606
rect 51100 3388 51156 3444
rect 50428 2380 50484 2436
rect 50540 2828 50596 2884
rect 50316 2156 50372 2212
rect 49868 1874 49924 1876
rect 49868 1822 49870 1874
rect 49870 1822 49922 1874
rect 49922 1822 49924 1874
rect 49868 1820 49924 1822
rect 49756 1426 49812 1428
rect 49756 1374 49758 1426
rect 49758 1374 49810 1426
rect 49810 1374 49812 1426
rect 49756 1372 49812 1374
rect 49084 1260 49140 1316
rect 48748 1202 48804 1204
rect 48748 1150 48750 1202
rect 48750 1150 48802 1202
rect 48802 1150 48804 1202
rect 48748 1148 48804 1150
rect 48188 924 48244 980
rect 51212 3164 51268 3220
rect 51100 2716 51156 2772
rect 51436 7196 51492 7252
rect 51436 4060 51492 4116
rect 51548 2604 51604 2660
rect 51436 2268 51492 2324
rect 50764 588 50820 644
rect 50540 476 50596 532
rect 44828 364 44884 420
rect 45948 252 46004 308
rect 50876 252 50932 308
rect 48412 140 48468 196
rect 39788 28 39844 84
rect 51548 28 51604 84
<< metal3 >>
rect 14466 14140 14476 14196
rect 14532 14140 16548 14196
rect 16706 14140 16716 14196
rect 16772 14140 31164 14196
rect 31220 14140 31230 14196
rect 31378 14140 31388 14196
rect 31444 14140 35028 14196
rect 35186 14140 35196 14196
rect 35252 14140 39116 14196
rect 39172 14140 39182 14196
rect 39676 14140 44156 14196
rect 44212 14140 44222 14196
rect 16492 14084 16548 14140
rect 34972 14084 35028 14140
rect 11554 14028 11564 14084
rect 11620 14028 12348 14084
rect 12404 14028 12414 14084
rect 13906 14028 13916 14084
rect 13972 14028 16268 14084
rect 16324 14028 16334 14084
rect 16492 14028 25116 14084
rect 25172 14028 25182 14084
rect 25330 14028 25340 14084
rect 25396 14028 25406 14084
rect 25554 14028 25564 14084
rect 25620 14028 33068 14084
rect 33124 14028 33134 14084
rect 34972 14028 37884 14084
rect 37940 14028 37950 14084
rect 38108 14028 38668 14084
rect 0 13972 112 14000
rect 25340 13972 25396 14028
rect 38108 13972 38164 14028
rect 0 13916 140 13972
rect 196 13916 206 13972
rect 10322 13916 10332 13972
rect 10388 13916 22764 13972
rect 22820 13916 22830 13972
rect 22988 13916 25396 13972
rect 26002 13916 26012 13972
rect 26068 13916 29540 13972
rect 31350 13916 31388 13972
rect 31444 13916 31454 13972
rect 31602 13916 31612 13972
rect 31668 13916 38164 13972
rect 38612 13972 38668 14028
rect 39676 13972 39732 14140
rect 52640 13972 52752 14000
rect 38612 13916 39732 13972
rect 51090 13916 51100 13972
rect 51156 13916 52752 13972
rect 0 13888 112 13916
rect 22988 13860 23044 13916
rect 29484 13860 29540 13916
rect 52640 13888 52752 13916
rect 14438 13804 14476 13860
rect 14532 13804 14542 13860
rect 15474 13804 15484 13860
rect 15540 13804 20076 13860
rect 20132 13804 20142 13860
rect 20290 13804 20300 13860
rect 20356 13804 23044 13860
rect 23772 13804 24892 13860
rect 24948 13804 24958 13860
rect 26114 13804 26124 13860
rect 26180 13804 29260 13860
rect 29316 13804 29326 13860
rect 29484 13804 33964 13860
rect 34020 13804 34030 13860
rect 35186 13804 35196 13860
rect 35252 13804 37996 13860
rect 38052 13804 38062 13860
rect 38210 13804 38220 13860
rect 38276 13804 38892 13860
rect 38948 13804 38958 13860
rect 39106 13804 39116 13860
rect 39172 13804 39340 13860
rect 39396 13804 39406 13860
rect 23772 13748 23828 13804
rect 15138 13692 15148 13748
rect 15204 13692 15988 13748
rect 19394 13692 19404 13748
rect 19460 13692 23828 13748
rect 23986 13692 23996 13748
rect 24052 13692 25340 13748
rect 25396 13692 25406 13748
rect 26338 13692 26348 13748
rect 26404 13692 32284 13748
rect 32340 13692 32350 13748
rect 37426 13692 37436 13748
rect 37492 13692 40012 13748
rect 40068 13692 40078 13748
rect 15932 13636 15988 13692
rect 11330 13580 11340 13636
rect 11396 13580 15708 13636
rect 15764 13580 15774 13636
rect 15932 13580 20972 13636
rect 21028 13580 21038 13636
rect 23202 13580 23212 13636
rect 23268 13580 24444 13636
rect 24500 13580 24510 13636
rect 24892 13580 25564 13636
rect 25620 13580 25630 13636
rect 25778 13580 25788 13636
rect 25844 13580 31836 13636
rect 31892 13580 31902 13636
rect 37314 13580 37324 13636
rect 37380 13580 51212 13636
rect 51268 13580 51278 13636
rect 0 13524 112 13552
rect 24892 13524 24948 13580
rect 52640 13524 52752 13552
rect 0 13468 1260 13524
rect 1316 13468 1326 13524
rect 9762 13468 9772 13524
rect 9828 13468 14364 13524
rect 14420 13468 14430 13524
rect 14914 13468 14924 13524
rect 14980 13468 18396 13524
rect 18452 13468 18462 13524
rect 19170 13468 19180 13524
rect 19236 13468 21308 13524
rect 21364 13468 21374 13524
rect 21522 13468 21532 13524
rect 21588 13468 22316 13524
rect 22372 13468 22382 13524
rect 22530 13468 22540 13524
rect 22596 13468 24668 13524
rect 24724 13468 24734 13524
rect 24882 13468 24892 13524
rect 24948 13468 24958 13524
rect 25218 13468 25228 13524
rect 25284 13468 35196 13524
rect 35252 13468 35262 13524
rect 37650 13468 37660 13524
rect 37716 13468 41244 13524
rect 41300 13468 41310 13524
rect 50530 13468 50540 13524
rect 50596 13468 52752 13524
rect 0 13440 112 13468
rect 52640 13440 52752 13468
rect 7532 13356 15484 13412
rect 15540 13356 15550 13412
rect 15698 13356 15708 13412
rect 15764 13356 16716 13412
rect 16772 13356 16782 13412
rect 17602 13356 17612 13412
rect 17668 13356 18172 13412
rect 18228 13356 18238 13412
rect 18498 13356 18508 13412
rect 18564 13356 24332 13412
rect 24388 13356 24398 13412
rect 24882 13356 24892 13412
rect 24948 13356 30156 13412
rect 30212 13356 30222 13412
rect 31154 13356 31164 13412
rect 31220 13356 33292 13412
rect 33348 13356 33358 13412
rect 36754 13356 36764 13412
rect 36820 13356 39788 13412
rect 39844 13356 39854 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 0 13076 112 13104
rect 0 13020 2268 13076
rect 2324 13020 2334 13076
rect 0 12992 112 13020
rect 7532 12852 7588 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 13346 13244 13356 13300
rect 13412 13244 16828 13300
rect 16884 13244 16894 13300
rect 17164 13244 23660 13300
rect 23716 13244 23726 13300
rect 24892 13244 33628 13300
rect 33684 13244 33694 13300
rect 36530 13244 36540 13300
rect 36596 13244 38108 13300
rect 38164 13244 38174 13300
rect 39218 13244 39228 13300
rect 39284 13244 42364 13300
rect 42420 13244 42430 13300
rect 7746 13132 7756 13188
rect 7812 13132 16268 13188
rect 16324 13132 16334 13188
rect 11666 13020 11676 13076
rect 11732 13020 14588 13076
rect 14644 13020 14654 13076
rect 15250 13020 15260 13076
rect 15316 13020 15932 13076
rect 15988 13020 15998 13076
rect 17164 12964 17220 13244
rect 24892 13188 24948 13244
rect 17378 13132 17388 13188
rect 17444 13132 20188 13188
rect 20244 13132 20254 13188
rect 21186 13132 21196 13188
rect 21252 13132 22428 13188
rect 22484 13132 22494 13188
rect 22652 13132 24948 13188
rect 25106 13132 25116 13188
rect 25172 13132 26740 13188
rect 26898 13132 26908 13188
rect 26964 13132 27244 13188
rect 27300 13132 27310 13188
rect 29026 13132 29036 13188
rect 29092 13132 31836 13188
rect 31892 13132 31902 13188
rect 33058 13132 33068 13188
rect 33124 13132 39564 13188
rect 39620 13132 39630 13188
rect 40114 13132 40124 13188
rect 40180 13132 45052 13188
rect 45108 13132 45118 13188
rect 22652 13076 22708 13132
rect 26684 13076 26740 13132
rect 52640 13076 52752 13104
rect 18956 13020 22708 13076
rect 22866 13020 22876 13076
rect 22932 13020 23324 13076
rect 23380 13020 23390 13076
rect 24210 13020 24220 13076
rect 24276 13020 26460 13076
rect 26516 13020 26526 13076
rect 26684 13020 32620 13076
rect 32676 13020 32686 13076
rect 36082 13020 36092 13076
rect 36148 13020 36540 13076
rect 36596 13020 36606 13076
rect 38994 13020 39004 13076
rect 39060 13020 43708 13076
rect 43764 13020 43774 13076
rect 48066 13020 48076 13076
rect 48132 13020 52752 13076
rect 2706 12796 2716 12852
rect 2772 12796 7588 12852
rect 9548 12908 17220 12964
rect 17938 12908 17948 12964
rect 18004 12908 18620 12964
rect 18676 12908 18686 12964
rect 9548 12740 9604 12908
rect 11890 12796 11900 12852
rect 11956 12796 15148 12852
rect 15204 12796 15214 12852
rect 15362 12796 15372 12852
rect 15428 12796 16716 12852
rect 16772 12796 16782 12852
rect 18956 12740 19012 13020
rect 52640 12992 52752 13020
rect 6178 12684 6188 12740
rect 6244 12684 9604 12740
rect 12338 12684 12348 12740
rect 12404 12684 14812 12740
rect 14868 12684 14878 12740
rect 15026 12684 15036 12740
rect 15092 12684 19012 12740
rect 19628 12908 31612 12964
rect 31668 12908 31678 12964
rect 31826 12908 31836 12964
rect 31892 12908 39508 12964
rect 39666 12908 39676 12964
rect 39732 12908 40348 12964
rect 40404 12908 40414 12964
rect 0 12628 112 12656
rect 19628 12628 19684 12908
rect 39452 12852 39508 12908
rect 21634 12796 21644 12852
rect 21700 12796 38444 12852
rect 38500 12796 38510 12852
rect 39452 12796 42588 12852
rect 42644 12796 42654 12852
rect 19842 12684 19852 12740
rect 19908 12684 20860 12740
rect 20916 12684 20926 12740
rect 21186 12684 21196 12740
rect 21252 12684 26348 12740
rect 26404 12684 26414 12740
rect 27010 12684 27020 12740
rect 27076 12684 27114 12740
rect 27234 12684 27244 12740
rect 27300 12684 27468 12740
rect 27524 12684 27534 12740
rect 27682 12684 27692 12740
rect 27748 12684 31948 12740
rect 32004 12684 32014 12740
rect 32610 12684 32620 12740
rect 32676 12684 36876 12740
rect 36932 12684 36942 12740
rect 37202 12684 37212 12740
rect 37268 12684 38668 12740
rect 38724 12684 38734 12740
rect 39330 12684 39340 12740
rect 39396 12684 39676 12740
rect 39732 12684 39742 12740
rect 52640 12628 52752 12656
rect 0 12572 3276 12628
rect 3332 12572 3342 12628
rect 9212 12572 19684 12628
rect 24210 12572 24220 12628
rect 24276 12572 25004 12628
rect 25060 12572 25070 12628
rect 25218 12572 25228 12628
rect 25284 12572 28924 12628
rect 28980 12572 28990 12628
rect 30258 12572 30268 12628
rect 30324 12572 35644 12628
rect 35700 12572 35710 12628
rect 38546 12572 38556 12628
rect 38612 12572 40796 12628
rect 40852 12572 40862 12628
rect 48178 12572 48188 12628
rect 48244 12572 52752 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 9212 12404 9268 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 52640 12544 52752 12572
rect 10882 12460 10892 12516
rect 10948 12460 13020 12516
rect 13076 12460 13086 12516
rect 13468 12460 16492 12516
rect 16548 12460 16558 12516
rect 16706 12460 16716 12516
rect 16772 12460 20748 12516
rect 20804 12460 20814 12516
rect 20972 12460 23548 12516
rect 23604 12460 23614 12516
rect 24210 12460 24220 12516
rect 24276 12460 25228 12516
rect 25284 12460 25294 12516
rect 26002 12460 26012 12516
rect 26068 12460 33404 12516
rect 33460 12460 33470 12516
rect 38322 12460 38332 12516
rect 38388 12460 41580 12516
rect 41636 12460 41646 12516
rect 3154 12348 3164 12404
rect 3220 12348 9268 12404
rect 11778 12348 11788 12404
rect 11844 12348 13244 12404
rect 13300 12348 13310 12404
rect 13468 12292 13524 12460
rect 20972 12404 21028 12460
rect 14802 12348 14812 12404
rect 14868 12348 17500 12404
rect 17556 12348 17566 12404
rect 18050 12348 18060 12404
rect 18116 12348 21028 12404
rect 21634 12348 21644 12404
rect 21700 12348 22204 12404
rect 22260 12348 22270 12404
rect 23538 12348 23548 12404
rect 23604 12348 24332 12404
rect 24388 12348 24398 12404
rect 24994 12348 25004 12404
rect 25060 12348 26348 12404
rect 26404 12348 26414 12404
rect 26572 12348 28252 12404
rect 28308 12348 28318 12404
rect 28466 12348 28476 12404
rect 28532 12348 36316 12404
rect 36372 12348 36382 12404
rect 37874 12348 37884 12404
rect 37940 12348 39340 12404
rect 39396 12348 39406 12404
rect 39890 12348 39900 12404
rect 39956 12348 42476 12404
rect 42532 12348 42542 12404
rect 8866 12236 8876 12292
rect 8932 12236 13524 12292
rect 13682 12236 13692 12292
rect 13748 12236 15260 12292
rect 15316 12236 15326 12292
rect 15474 12236 15484 12292
rect 15540 12236 17276 12292
rect 17332 12236 17342 12292
rect 17798 12236 17836 12292
rect 17892 12236 17902 12292
rect 18050 12236 18060 12292
rect 18116 12236 19516 12292
rect 19572 12236 19582 12292
rect 22418 12236 22428 12292
rect 22484 12236 26236 12292
rect 26292 12236 26302 12292
rect 0 12180 112 12208
rect 26572 12180 26628 12348
rect 26786 12236 26796 12292
rect 26852 12236 31724 12292
rect 31780 12236 31790 12292
rect 31938 12236 31948 12292
rect 32004 12236 35756 12292
rect 35812 12236 35822 12292
rect 39442 12236 39452 12292
rect 39508 12236 40908 12292
rect 40964 12236 40974 12292
rect 43652 12236 47292 12292
rect 47348 12236 47358 12292
rect 0 12124 364 12180
rect 420 12124 430 12180
rect 13010 12124 13020 12180
rect 13076 12178 13636 12180
rect 13692 12178 14868 12180
rect 14924 12178 15540 12180
rect 13076 12124 15540 12178
rect 15698 12124 15708 12180
rect 15764 12124 24892 12180
rect 24948 12124 24958 12180
rect 25106 12124 25116 12180
rect 25172 12124 26628 12180
rect 29260 12124 30380 12180
rect 30436 12124 30446 12180
rect 30706 12124 30716 12180
rect 30772 12124 37884 12180
rect 37940 12124 37950 12180
rect 38770 12124 38780 12180
rect 38836 12124 41132 12180
rect 41188 12124 41198 12180
rect 0 12096 112 12124
rect 13580 12122 13748 12124
rect 14812 12122 14980 12124
rect 6738 12012 6748 12068
rect 6804 12012 9772 12068
rect 9828 12012 9838 12068
rect 12198 12012 12236 12068
rect 12292 12012 12302 12068
rect 15484 11956 15540 12124
rect 29260 12068 29316 12124
rect 43652 12068 43708 12236
rect 52640 12180 52752 12208
rect 49746 12124 49756 12180
rect 49812 12124 52752 12180
rect 52640 12096 52752 12124
rect 15810 12012 15820 12068
rect 15876 12012 19628 12068
rect 19684 12012 19694 12068
rect 20178 12012 20188 12068
rect 20244 12012 21644 12068
rect 21700 12012 21710 12068
rect 23426 12012 23436 12068
rect 23492 12012 24220 12068
rect 24276 12012 24286 12068
rect 24434 12012 24444 12068
rect 24500 12012 29316 12068
rect 29474 12012 29484 12068
rect 29540 12012 30884 12068
rect 32162 12012 32172 12068
rect 32228 12012 34524 12068
rect 34580 12012 34590 12068
rect 37538 12012 37548 12068
rect 37604 12012 40236 12068
rect 40292 12012 40302 12068
rect 40460 12012 43708 12068
rect 45154 12012 45164 12068
rect 45220 12012 50204 12068
rect 50260 12012 50270 12068
rect 30828 11956 30884 12012
rect 6290 11900 6300 11956
rect 6356 11900 7532 11956
rect 7588 11900 7598 11956
rect 12450 11900 12460 11956
rect 12516 11900 13692 11956
rect 13748 11900 13758 11956
rect 14018 11900 14028 11956
rect 14084 11900 15260 11956
rect 15316 11900 15326 11956
rect 15484 11900 16828 11956
rect 16884 11900 16894 11956
rect 17686 11900 17724 11956
rect 17780 11900 17790 11956
rect 17910 11900 17948 11956
rect 18004 11900 18014 11956
rect 18610 11900 18620 11956
rect 18676 11900 20636 11956
rect 20692 11900 20702 11956
rect 22540 11900 25228 11956
rect 25284 11900 25294 11956
rect 25442 11900 25452 11956
rect 25508 11900 26684 11956
rect 26740 11900 26750 11956
rect 26898 11900 26908 11956
rect 26964 11900 28476 11956
rect 28532 11900 28542 11956
rect 28690 11900 28700 11956
rect 28756 11900 30604 11956
rect 30660 11900 30670 11956
rect 30828 11900 32396 11956
rect 32452 11900 32462 11956
rect 34402 11900 34412 11956
rect 34468 11900 39116 11956
rect 39172 11900 39182 11956
rect 22540 11844 22596 11900
rect 40460 11844 40516 12012
rect 43652 11900 47740 11956
rect 47796 11900 47806 11956
rect 43652 11844 43708 11900
rect 10434 11788 10444 11844
rect 10500 11788 12572 11844
rect 12628 11788 12638 11844
rect 13356 11788 13916 11844
rect 13972 11788 13982 11844
rect 14130 11788 14140 11844
rect 14196 11788 15036 11844
rect 15092 11788 15102 11844
rect 15250 11788 15260 11844
rect 15316 11788 22596 11844
rect 22754 11788 22764 11844
rect 22820 11788 24332 11844
rect 24388 11788 24398 11844
rect 25106 11788 25116 11844
rect 25172 11788 27692 11844
rect 27748 11788 27758 11844
rect 28018 11788 28028 11844
rect 28084 11788 31276 11844
rect 31332 11788 31342 11844
rect 31836 11788 35308 11844
rect 35364 11788 35374 11844
rect 35522 11788 35532 11844
rect 35588 11788 37100 11844
rect 37156 11788 37166 11844
rect 37314 11788 37324 11844
rect 37380 11788 40516 11844
rect 42140 11788 43708 11844
rect 49634 11788 49644 11844
rect 49700 11788 51044 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 13356 11732 13412 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 31836 11732 31892 11788
rect 0 11676 3388 11732
rect 9874 11676 9884 11732
rect 9940 11676 13412 11732
rect 14802 11676 14812 11732
rect 14868 11676 16380 11732
rect 16436 11676 16446 11732
rect 16706 11676 16716 11732
rect 16772 11676 18732 11732
rect 18788 11676 18798 11732
rect 20178 11676 20188 11732
rect 20244 11676 24108 11732
rect 24164 11676 24174 11732
rect 24892 11676 28308 11732
rect 28466 11676 28476 11732
rect 28532 11676 31892 11732
rect 31948 11676 33404 11732
rect 33460 11676 33470 11732
rect 33618 11676 33628 11732
rect 33684 11676 36988 11732
rect 37044 11676 37054 11732
rect 37212 11676 41916 11732
rect 41972 11676 41982 11732
rect 0 11648 112 11676
rect 3332 11620 3388 11676
rect 3332 11564 7980 11620
rect 8036 11564 8046 11620
rect 11330 11564 11340 11620
rect 11396 11564 14924 11620
rect 14980 11564 14990 11620
rect 15586 11564 15596 11620
rect 15652 11564 16156 11620
rect 16212 11564 16222 11620
rect 16482 11564 16492 11620
rect 16548 11564 21196 11620
rect 21252 11564 21262 11620
rect 21634 11564 21644 11620
rect 21700 11564 22540 11620
rect 22596 11564 22606 11620
rect 22754 11564 22764 11620
rect 22820 11564 23324 11620
rect 23380 11564 23390 11620
rect 23538 11564 23548 11620
rect 23604 11564 24220 11620
rect 24276 11564 24286 11620
rect 24892 11508 24948 11676
rect 28252 11620 28308 11676
rect 31948 11620 32004 11676
rect 37212 11620 37268 11676
rect 25106 11564 25116 11620
rect 25172 11564 28028 11620
rect 28084 11564 28094 11620
rect 28252 11564 29596 11620
rect 29652 11564 29662 11620
rect 30370 11564 30380 11620
rect 30436 11564 31052 11620
rect 31108 11564 31118 11620
rect 31378 11564 31388 11620
rect 31444 11564 32004 11620
rect 32162 11564 32172 11620
rect 32228 11564 34076 11620
rect 34132 11564 34142 11620
rect 35634 11564 35644 11620
rect 35700 11564 37268 11620
rect 37538 11564 37548 11620
rect 37604 11564 40684 11620
rect 40740 11564 40750 11620
rect 42140 11508 42196 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 50988 11732 51044 11788
rect 52640 11732 52752 11760
rect 50988 11676 52752 11732
rect 52640 11648 52752 11676
rect 8978 11452 8988 11508
rect 9044 11452 18060 11508
rect 18116 11452 18126 11508
rect 18274 11452 18284 11508
rect 18340 11452 18508 11508
rect 18564 11452 18574 11508
rect 18834 11452 18844 11508
rect 18900 11452 19964 11508
rect 20020 11452 20030 11508
rect 21522 11452 21532 11508
rect 21588 11452 24948 11508
rect 25004 11452 25452 11508
rect 25508 11452 25518 11508
rect 25666 11452 25676 11508
rect 25732 11452 27356 11508
rect 27412 11452 27422 11508
rect 28466 11452 28476 11508
rect 28532 11452 42196 11508
rect 25004 11396 25060 11452
rect 3154 11340 3164 11396
rect 3220 11340 13692 11396
rect 13748 11340 13758 11396
rect 16258 11340 16268 11396
rect 16324 11340 21308 11396
rect 21364 11340 21374 11396
rect 21522 11340 21532 11396
rect 21588 11340 25060 11396
rect 25218 11340 25228 11396
rect 25284 11340 29820 11396
rect 29876 11340 29886 11396
rect 30146 11340 30156 11396
rect 30212 11340 30716 11396
rect 30772 11340 30782 11396
rect 31042 11340 31052 11396
rect 31108 11340 33068 11396
rect 33124 11340 33134 11396
rect 33618 11340 33628 11396
rect 33684 11340 38108 11396
rect 38164 11340 38174 11396
rect 40338 11340 40348 11396
rect 40404 11340 50428 11396
rect 50484 11340 50494 11396
rect 0 11284 112 11312
rect 52640 11284 52752 11312
rect 0 11228 15260 11284
rect 15316 11228 15326 11284
rect 16146 11228 16156 11284
rect 16212 11228 20300 11284
rect 20356 11228 20366 11284
rect 20850 11228 20860 11284
rect 20916 11228 33516 11284
rect 33572 11228 33582 11284
rect 33730 11228 33740 11284
rect 33796 11228 37996 11284
rect 38052 11228 38062 11284
rect 38210 11228 38220 11284
rect 38276 11228 39116 11284
rect 39172 11228 39182 11284
rect 42130 11228 42140 11284
rect 42196 11228 48972 11284
rect 49028 11228 49038 11284
rect 49858 11228 49868 11284
rect 49924 11228 52752 11284
rect 0 11200 112 11228
rect 52640 11200 52752 11228
rect 1250 11116 1260 11172
rect 1316 11116 5292 11172
rect 5348 11116 5358 11172
rect 6514 11116 6524 11172
rect 6580 11116 13580 11172
rect 13636 11116 13646 11172
rect 14914 11116 14924 11172
rect 14980 11116 25228 11172
rect 25284 11116 25294 11172
rect 25442 11116 25452 11172
rect 25508 11116 33852 11172
rect 33908 11116 33918 11172
rect 37426 11116 37436 11172
rect 37492 11116 48860 11172
rect 48916 11116 48926 11172
rect 9212 11004 15708 11060
rect 15764 11004 15774 11060
rect 16034 11004 16044 11060
rect 16100 11004 21532 11060
rect 21588 11004 21598 11060
rect 24210 11004 24220 11060
rect 24276 11004 25116 11060
rect 25172 11004 25182 11060
rect 25330 11004 25340 11060
rect 25396 11004 29260 11060
rect 29316 11004 29326 11060
rect 31714 11004 31724 11060
rect 31780 11004 35252 11060
rect 36866 11004 36876 11060
rect 36932 11004 43484 11060
rect 43540 11004 43550 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 0 10836 112 10864
rect 9212 10836 9268 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 35196 10948 35252 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 13234 10892 13244 10948
rect 13300 10892 20860 10948
rect 20916 10892 20926 10948
rect 21084 10892 23716 10948
rect 24322 10892 24332 10948
rect 24388 10892 25900 10948
rect 25956 10892 25966 10948
rect 26226 10892 26236 10948
rect 26292 10892 26740 10948
rect 27206 10892 27244 10948
rect 27300 10892 27310 10948
rect 31154 10892 31164 10948
rect 31220 10892 34972 10948
rect 35028 10892 35038 10948
rect 35196 10892 40460 10948
rect 40516 10892 40526 10948
rect 21084 10836 21140 10892
rect 23660 10836 23716 10892
rect 26684 10836 26740 10892
rect 52640 10836 52752 10864
rect 0 10780 1372 10836
rect 1428 10780 1438 10836
rect 2034 10780 2044 10836
rect 2100 10780 9268 10836
rect 10098 10780 10108 10836
rect 10164 10780 16212 10836
rect 16370 10780 16380 10836
rect 16436 10780 17052 10836
rect 17108 10780 17118 10836
rect 17276 10780 21140 10836
rect 22642 10780 22652 10836
rect 22708 10780 23436 10836
rect 23492 10780 23502 10836
rect 23660 10780 25004 10836
rect 25060 10780 25070 10836
rect 25330 10780 25340 10836
rect 25396 10780 26460 10836
rect 26516 10780 26526 10836
rect 26684 10780 36204 10836
rect 36260 10780 36270 10836
rect 36978 10780 36988 10836
rect 37044 10780 47628 10836
rect 47684 10780 47694 10836
rect 51202 10780 51212 10836
rect 51268 10780 52752 10836
rect 0 10752 112 10780
rect 3266 10668 3276 10724
rect 3332 10668 16100 10724
rect 12786 10556 12796 10612
rect 12852 10556 15484 10612
rect 15540 10556 15550 10612
rect 16044 10500 16100 10668
rect 16156 10612 16212 10780
rect 17276 10724 17332 10780
rect 52640 10752 52752 10780
rect 16482 10668 16492 10724
rect 16548 10668 17332 10724
rect 17714 10668 17724 10724
rect 17780 10668 23324 10724
rect 23380 10668 23390 10724
rect 23538 10668 23548 10724
rect 23604 10668 25004 10724
rect 25060 10668 25070 10724
rect 25218 10668 25228 10724
rect 25284 10668 27692 10724
rect 27748 10668 27758 10724
rect 28802 10668 28812 10724
rect 28868 10668 34860 10724
rect 34916 10668 34926 10724
rect 35298 10668 35308 10724
rect 35364 10668 45948 10724
rect 46004 10668 46014 10724
rect 16156 10556 26684 10612
rect 26740 10556 26750 10612
rect 27010 10556 27020 10612
rect 27076 10556 32732 10612
rect 32788 10556 32798 10612
rect 33058 10556 33068 10612
rect 33124 10556 36652 10612
rect 36708 10556 36718 10612
rect 37874 10556 37884 10612
rect 37940 10556 40908 10612
rect 40964 10556 40974 10612
rect 43362 10556 43372 10612
rect 43428 10556 50204 10612
rect 50260 10556 50270 10612
rect 8306 10444 8316 10500
rect 8372 10444 10108 10500
rect 10164 10444 10174 10500
rect 10658 10444 10668 10500
rect 10724 10444 15708 10500
rect 15764 10444 15774 10500
rect 16044 10444 18452 10500
rect 20066 10444 20076 10500
rect 20132 10444 29596 10500
rect 29652 10444 29662 10500
rect 29922 10444 29932 10500
rect 29988 10444 38780 10500
rect 38836 10444 38846 10500
rect 43652 10444 43932 10500
rect 43988 10444 43998 10500
rect 48290 10444 48300 10500
rect 48356 10444 50652 10500
rect 50708 10444 50718 10500
rect 0 10388 112 10416
rect 18396 10388 18452 10444
rect 0 10332 7028 10388
rect 8530 10332 8540 10388
rect 8596 10332 11788 10388
rect 11844 10332 11854 10388
rect 14578 10332 14588 10388
rect 14644 10332 18172 10388
rect 18228 10332 18238 10388
rect 18396 10332 20188 10388
rect 20244 10332 20254 10388
rect 21298 10332 21308 10388
rect 21364 10332 21980 10388
rect 22036 10332 22046 10388
rect 22194 10332 22204 10388
rect 22260 10332 23380 10388
rect 23538 10332 23548 10388
rect 23604 10332 26348 10388
rect 26404 10332 26414 10388
rect 26562 10332 26572 10388
rect 26628 10332 26684 10388
rect 26740 10332 26750 10388
rect 27122 10332 27132 10388
rect 27188 10332 28812 10388
rect 28868 10332 28878 10388
rect 29026 10332 29036 10388
rect 29092 10332 31052 10388
rect 31108 10332 31118 10388
rect 31378 10332 31388 10388
rect 31444 10332 32508 10388
rect 32564 10332 32574 10388
rect 32834 10332 32844 10388
rect 32900 10332 39452 10388
rect 39508 10332 39518 10388
rect 0 10304 112 10332
rect 6972 10276 7028 10332
rect 23324 10276 23380 10332
rect 43652 10276 43708 10444
rect 52640 10388 52752 10416
rect 49634 10332 49644 10388
rect 49700 10332 52752 10388
rect 52640 10304 52752 10332
rect 6972 10220 10388 10276
rect 13794 10220 13804 10276
rect 13860 10220 15764 10276
rect 15922 10220 15932 10276
rect 15988 10220 18844 10276
rect 18900 10220 18910 10276
rect 19170 10220 19180 10276
rect 19236 10220 22764 10276
rect 22820 10220 22830 10276
rect 23324 10220 24332 10276
rect 24388 10220 24398 10276
rect 25228 10220 33852 10276
rect 33908 10220 33918 10276
rect 35298 10220 35308 10276
rect 35364 10220 43708 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 6636 10108 10276 10164
rect 6636 10052 6692 10108
rect 3042 9996 3052 10052
rect 3108 9996 6692 10052
rect 0 9940 112 9968
rect 10220 9940 10276 10108
rect 10332 10052 10388 10220
rect 15708 10164 15764 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 10546 10108 10556 10164
rect 10612 10108 14476 10164
rect 14532 10108 14542 10164
rect 15026 10108 15036 10164
rect 15092 10108 15148 10164
rect 15204 10108 15214 10164
rect 15708 10108 16492 10164
rect 16548 10108 16558 10164
rect 16706 10108 16716 10164
rect 16772 10108 22876 10164
rect 22932 10108 22942 10164
rect 23090 10108 23100 10164
rect 23156 10108 24220 10164
rect 24276 10108 24286 10164
rect 25228 10052 25284 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 25442 10108 25452 10164
rect 25508 10108 26684 10164
rect 26740 10108 26750 10164
rect 26898 10108 26908 10164
rect 26964 10108 28700 10164
rect 28756 10108 28766 10164
rect 30034 10108 30044 10164
rect 30100 10108 34412 10164
rect 34468 10108 34478 10164
rect 34626 10108 34636 10164
rect 34692 10108 41804 10164
rect 41860 10108 41870 10164
rect 10332 9996 10668 10052
rect 10724 9996 10734 10052
rect 14018 9996 14028 10052
rect 14084 9996 15372 10052
rect 15428 9996 15438 10052
rect 15698 9996 15708 10052
rect 15764 9996 16828 10052
rect 16884 9996 16894 10052
rect 17042 9996 17052 10052
rect 17108 9996 25284 10052
rect 25442 9996 25452 10052
rect 25508 9996 27468 10052
rect 27524 9996 27534 10052
rect 27682 9996 27692 10052
rect 27748 9996 35420 10052
rect 35476 9996 35486 10052
rect 38612 9996 44268 10052
rect 44324 9996 44334 10052
rect 38612 9940 38668 9996
rect 52640 9940 52752 9968
rect 0 9884 1708 9940
rect 1764 9884 1774 9940
rect 10220 9884 20076 9940
rect 20132 9884 20142 9940
rect 20514 9884 20524 9940
rect 20580 9884 21924 9940
rect 22082 9884 22092 9940
rect 22148 9884 22652 9940
rect 22708 9884 22718 9940
rect 23314 9884 23324 9940
rect 23380 9884 24892 9940
rect 24948 9884 24958 9940
rect 25106 9884 25116 9940
rect 25172 9884 26852 9940
rect 26908 9884 26918 9940
rect 27234 9884 27244 9940
rect 27300 9884 38668 9940
rect 39116 9884 50428 9940
rect 50484 9884 50494 9940
rect 51426 9884 51436 9940
rect 51492 9884 52752 9940
rect 0 9856 112 9884
rect 21868 9828 21924 9884
rect 39116 9828 39172 9884
rect 52640 9856 52752 9884
rect 1138 9772 1148 9828
rect 1204 9772 3164 9828
rect 3220 9772 3230 9828
rect 11778 9772 11788 9828
rect 11844 9772 16492 9828
rect 16548 9772 16558 9828
rect 16818 9772 16828 9828
rect 16884 9772 19516 9828
rect 19572 9772 19582 9828
rect 19842 9772 19852 9828
rect 19908 9772 21644 9828
rect 21700 9772 21710 9828
rect 21868 9772 22988 9828
rect 23044 9772 23054 9828
rect 23314 9772 23324 9828
rect 23380 9772 24220 9828
rect 24276 9772 24286 9828
rect 24434 9772 24444 9828
rect 24500 9772 25676 9828
rect 25732 9772 25742 9828
rect 26786 9772 26796 9828
rect 26852 9772 27300 9828
rect 27458 9772 27468 9828
rect 27524 9772 28364 9828
rect 28420 9772 28430 9828
rect 31154 9772 31164 9828
rect 31220 9772 39172 9828
rect 40226 9772 40236 9828
rect 40292 9772 45276 9828
rect 45332 9772 45342 9828
rect 27244 9716 27300 9772
rect 13570 9660 13580 9716
rect 13636 9660 18508 9716
rect 18564 9660 18574 9716
rect 19618 9660 19628 9716
rect 19684 9660 26236 9716
rect 26292 9660 26302 9716
rect 27244 9660 28924 9716
rect 28980 9660 28990 9716
rect 31490 9660 31500 9716
rect 31556 9660 42252 9716
rect 42308 9660 42318 9716
rect 44482 9660 44492 9716
rect 44548 9660 48972 9716
rect 49028 9660 49038 9716
rect 49858 9660 49868 9716
rect 49924 9660 50540 9716
rect 50596 9660 50606 9716
rect 3332 9548 8092 9604
rect 8148 9548 8158 9604
rect 11778 9548 11788 9604
rect 11844 9548 16492 9604
rect 16548 9548 16558 9604
rect 16706 9548 16716 9604
rect 16772 9548 22092 9604
rect 22148 9548 22158 9604
rect 23090 9548 23100 9604
rect 23156 9548 25452 9604
rect 25508 9548 25518 9604
rect 26674 9548 26684 9604
rect 26740 9548 28028 9604
rect 28084 9548 28094 9604
rect 28802 9548 28812 9604
rect 28868 9548 32172 9604
rect 32228 9548 32238 9604
rect 32386 9548 32396 9604
rect 32452 9548 35308 9604
rect 35364 9548 35374 9604
rect 38658 9548 38668 9604
rect 38724 9548 40348 9604
rect 40404 9548 40414 9604
rect 40898 9548 40908 9604
rect 40964 9548 47180 9604
rect 47236 9548 47246 9604
rect 0 9492 112 9520
rect 3332 9492 3388 9548
rect 52640 9492 52752 9520
rect 0 9436 3388 9492
rect 15362 9436 15372 9492
rect 15428 9436 15932 9492
rect 15988 9436 15998 9492
rect 16146 9436 16156 9492
rect 16212 9436 23436 9492
rect 23492 9436 23502 9492
rect 26450 9436 26460 9492
rect 26516 9436 31164 9492
rect 31220 9436 31230 9492
rect 34962 9436 34972 9492
rect 35028 9436 39396 9492
rect 50978 9436 50988 9492
rect 51044 9436 52752 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 5618 9324 5628 9380
rect 5684 9324 19516 9380
rect 19572 9324 19582 9380
rect 19954 9324 19964 9380
rect 20020 9324 23660 9380
rect 23716 9324 23726 9380
rect 24994 9324 25004 9380
rect 25060 9324 25116 9380
rect 25172 9324 25182 9380
rect 25554 9324 25564 9380
rect 25620 9324 29540 9380
rect 29698 9324 29708 9380
rect 29764 9324 31500 9380
rect 31556 9324 31566 9380
rect 31714 9324 31724 9380
rect 31780 9324 35196 9380
rect 35252 9324 35262 9380
rect 29484 9268 29540 9324
rect 1362 9212 1372 9268
rect 1428 9212 8428 9268
rect 8484 9212 8494 9268
rect 14802 9212 14812 9268
rect 14868 9212 15820 9268
rect 15876 9212 15886 9268
rect 16044 9212 17052 9268
rect 17108 9212 17118 9268
rect 17266 9212 17276 9268
rect 17332 9212 19964 9268
rect 20020 9212 20030 9268
rect 20178 9212 20188 9268
rect 20244 9212 24332 9268
rect 24388 9212 24398 9268
rect 25116 9212 27916 9268
rect 27972 9212 27982 9268
rect 29484 9212 33628 9268
rect 33684 9212 33694 9268
rect 34066 9212 34076 9268
rect 34132 9212 37324 9268
rect 37380 9212 37390 9268
rect 16044 9156 16100 9212
rect 25116 9156 25172 9212
rect 9314 9100 9324 9156
rect 9380 9100 16100 9156
rect 16716 9100 22204 9156
rect 22260 9100 22270 9156
rect 22754 9100 22764 9156
rect 22820 9100 25172 9156
rect 25330 9100 25340 9156
rect 25396 9100 38332 9156
rect 38388 9100 38398 9156
rect 0 9044 112 9072
rect 16716 9044 16772 9100
rect 0 8988 1484 9044
rect 1540 8988 1550 9044
rect 5506 8988 5516 9044
rect 5572 8988 10556 9044
rect 10612 8988 10622 9044
rect 12226 8988 12236 9044
rect 12292 8988 16772 9044
rect 16930 8988 16940 9044
rect 16996 8988 21532 9044
rect 21588 8988 21598 9044
rect 21756 8988 26012 9044
rect 26068 8988 26078 9044
rect 26450 8988 26460 9044
rect 26516 8988 33180 9044
rect 33236 8988 33246 9044
rect 33954 8988 33964 9044
rect 34020 8988 39116 9044
rect 39172 8988 39182 9044
rect 0 8960 112 8988
rect 21756 8932 21812 8988
rect 26124 8932 26404 8938
rect 39340 8932 39396 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 52640 9408 52752 9436
rect 49634 9212 49644 9268
rect 49700 9212 51100 9268
rect 51156 9212 51166 9268
rect 52640 9044 52752 9072
rect 40450 8988 40460 9044
rect 40516 8988 46956 9044
rect 47012 8988 47022 9044
rect 51426 8988 51436 9044
rect 51492 8988 52752 9044
rect 52640 8960 52752 8988
rect 5842 8876 5852 8932
rect 5908 8876 17276 8932
rect 17332 8876 17342 8932
rect 17686 8876 17724 8932
rect 17780 8876 17790 8932
rect 17938 8876 17948 8932
rect 18004 8876 19180 8932
rect 19236 8876 19246 8932
rect 19954 8876 19964 8932
rect 20020 8876 20972 8932
rect 21028 8876 21038 8932
rect 21186 8876 21196 8932
rect 21252 8876 21812 8932
rect 21970 8876 21980 8932
rect 22036 8882 36988 8932
rect 22036 8876 26180 8882
rect 26348 8876 36988 8882
rect 37044 8876 37054 8932
rect 39340 8876 50204 8932
rect 50260 8876 50270 8932
rect 2146 8764 2156 8820
rect 2212 8764 13356 8820
rect 13412 8764 13422 8820
rect 15250 8764 15260 8820
rect 15316 8764 15708 8820
rect 15764 8764 15774 8820
rect 16006 8764 16044 8820
rect 16100 8764 16110 8820
rect 16482 8764 16492 8820
rect 16548 8764 18620 8820
rect 18676 8764 18686 8820
rect 18844 8764 20524 8820
rect 20580 8764 20590 8820
rect 20738 8764 20748 8820
rect 20804 8764 26124 8820
rect 26180 8764 26190 8820
rect 26562 8764 26572 8820
rect 26628 8764 27580 8820
rect 27636 8764 27646 8820
rect 27794 8764 27804 8820
rect 27860 8764 29820 8820
rect 29876 8764 29886 8820
rect 30258 8764 30268 8820
rect 30324 8764 31724 8820
rect 31780 8764 31790 8820
rect 31938 8764 31948 8820
rect 32004 8764 34300 8820
rect 34356 8764 34366 8820
rect 35074 8764 35084 8820
rect 35140 8764 44884 8820
rect 45378 8764 45388 8820
rect 45444 8764 47740 8820
rect 47796 8764 47806 8820
rect 18844 8708 18900 8764
rect 7420 8652 11676 8708
rect 11732 8652 11742 8708
rect 15092 8652 15596 8708
rect 15652 8652 15662 8708
rect 15810 8652 15820 8708
rect 15876 8652 17388 8708
rect 17444 8652 17454 8708
rect 17602 8652 17612 8708
rect 17668 8652 18900 8708
rect 19170 8652 19180 8708
rect 19236 8652 22540 8708
rect 22596 8652 22606 8708
rect 22978 8652 22988 8708
rect 23044 8652 24108 8708
rect 24164 8652 24174 8708
rect 24882 8652 24892 8708
rect 24948 8652 26460 8708
rect 26516 8652 26526 8708
rect 26684 8652 27692 8708
rect 27748 8652 27758 8708
rect 27906 8652 27916 8708
rect 27972 8652 32172 8708
rect 32228 8652 32238 8708
rect 35756 8652 40236 8708
rect 40292 8652 40302 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 0 8540 924 8596
rect 980 8540 990 8596
rect 0 8512 112 8540
rect 7420 8484 7476 8652
rect 15092 8596 15148 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 26684 8596 26740 8652
rect 7634 8540 7644 8596
rect 7700 8540 9996 8596
rect 10052 8540 10062 8596
rect 10322 8540 10332 8596
rect 10388 8540 15148 8596
rect 15250 8540 15260 8596
rect 15316 8540 15932 8596
rect 15988 8540 15998 8596
rect 16594 8540 16604 8596
rect 16660 8540 21868 8596
rect 21924 8540 21934 8596
rect 22082 8540 22092 8596
rect 22148 8540 24332 8596
rect 24388 8540 24398 8596
rect 26338 8540 26348 8596
rect 26404 8540 26740 8596
rect 26898 8540 26908 8596
rect 26964 8540 27804 8596
rect 27860 8540 27870 8596
rect 28018 8540 28028 8596
rect 28084 8540 33852 8596
rect 33908 8540 33918 8596
rect 34076 8540 35420 8596
rect 35476 8540 35486 8596
rect 34076 8484 34132 8540
rect 35756 8484 35812 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 44828 8596 44884 8764
rect 48290 8652 48300 8708
rect 48356 8652 50316 8708
rect 50372 8652 50382 8708
rect 52640 8596 52752 8624
rect 35970 8540 35980 8596
rect 36036 8540 42924 8596
rect 42980 8540 42990 8596
rect 44828 8540 48692 8596
rect 50978 8540 50988 8596
rect 51044 8540 52752 8596
rect 1362 8428 1372 8484
rect 1428 8428 7476 8484
rect 9202 8428 9212 8484
rect 9268 8428 13524 8484
rect 15026 8428 15036 8484
rect 15092 8428 15540 8484
rect 15698 8428 15708 8484
rect 15764 8428 16660 8484
rect 16818 8428 16828 8484
rect 16884 8428 20244 8484
rect 21858 8428 21868 8484
rect 21924 8428 22876 8484
rect 22932 8428 22942 8484
rect 23548 8428 27356 8484
rect 27412 8428 27422 8484
rect 27580 8428 31724 8484
rect 31780 8428 31790 8484
rect 32050 8428 32060 8484
rect 32116 8428 33404 8484
rect 33460 8428 33470 8484
rect 33618 8428 33628 8484
rect 33684 8428 34132 8484
rect 35196 8428 35812 8484
rect 36754 8428 36764 8484
rect 36820 8428 45500 8484
rect 45556 8428 45566 8484
rect 13468 8372 13524 8428
rect 15484 8372 15540 8428
rect 16604 8372 16660 8428
rect 20188 8372 20244 8428
rect 23548 8372 23604 8428
rect 27580 8372 27636 8428
rect 35196 8372 35252 8428
rect 48636 8372 48692 8540
rect 52640 8512 52752 8540
rect 6626 8316 6636 8372
rect 6692 8316 11788 8372
rect 11844 8316 11854 8372
rect 13468 8316 13692 8372
rect 13748 8316 13758 8372
rect 14466 8316 14476 8372
rect 14532 8316 15148 8372
rect 15204 8316 15214 8372
rect 15484 8316 16380 8372
rect 16436 8316 16446 8372
rect 16604 8316 19964 8372
rect 20020 8316 20030 8372
rect 20188 8316 23604 8372
rect 23762 8316 23772 8372
rect 23828 8316 26348 8372
rect 26404 8316 26414 8372
rect 26572 8316 27636 8372
rect 27794 8316 27804 8372
rect 27860 8316 28812 8372
rect 28868 8316 28878 8372
rect 29586 8316 29596 8372
rect 29652 8316 32396 8372
rect 32452 8316 32462 8372
rect 32722 8316 32732 8372
rect 32788 8316 35252 8372
rect 36978 8316 36988 8372
rect 37044 8316 39340 8372
rect 39396 8316 39406 8372
rect 40338 8316 40348 8372
rect 40404 8316 44828 8372
rect 44884 8316 44894 8372
rect 48636 8316 50428 8372
rect 50484 8316 50494 8372
rect 26572 8260 26628 8316
rect 8082 8204 8092 8260
rect 8148 8204 12124 8260
rect 12180 8204 12190 8260
rect 12450 8204 12460 8260
rect 12516 8204 16492 8260
rect 16548 8204 16558 8260
rect 16706 8204 16716 8260
rect 16772 8204 18844 8260
rect 18900 8204 18910 8260
rect 20066 8204 20076 8260
rect 20132 8204 20972 8260
rect 21028 8204 21038 8260
rect 22082 8204 22092 8260
rect 22148 8204 25228 8260
rect 25284 8204 25294 8260
rect 25442 8204 25452 8260
rect 25508 8204 26628 8260
rect 26786 8204 26796 8260
rect 26852 8204 29708 8260
rect 29764 8204 29774 8260
rect 29922 8204 29932 8260
rect 29988 8204 31164 8260
rect 31220 8204 31230 8260
rect 33618 8204 33628 8260
rect 33684 8204 37212 8260
rect 37268 8204 37278 8260
rect 37426 8204 37436 8260
rect 37492 8204 45164 8260
rect 45220 8204 45230 8260
rect 47618 8204 47628 8260
rect 47684 8204 48636 8260
rect 48692 8204 48702 8260
rect 0 8148 112 8176
rect 52640 8148 52752 8176
rect 0 8092 1596 8148
rect 1652 8092 1662 8148
rect 9762 8092 9772 8148
rect 9828 8092 13804 8148
rect 13860 8092 13870 8148
rect 14018 8092 14028 8148
rect 14084 8092 15372 8148
rect 15428 8092 15438 8148
rect 15698 8092 15708 8148
rect 15764 8092 25116 8148
rect 25172 8092 25182 8148
rect 25554 8092 25564 8148
rect 25620 8092 26572 8148
rect 26628 8092 26638 8148
rect 27010 8092 27020 8148
rect 27076 8092 28756 8148
rect 29474 8092 29484 8148
rect 29540 8092 41020 8148
rect 41076 8092 41086 8148
rect 41234 8092 41244 8148
rect 41300 8092 49980 8148
rect 50036 8092 50046 8148
rect 50866 8092 50876 8148
rect 50932 8092 52752 8148
rect 0 8064 112 8092
rect 28700 8036 28756 8092
rect 52640 8064 52752 8092
rect 2818 7980 2828 8036
rect 2884 7980 14924 8036
rect 14980 7980 14990 8036
rect 15250 7980 15260 8036
rect 15316 7980 19628 8036
rect 19684 7980 19694 8036
rect 19842 7980 19852 8036
rect 19908 7980 21644 8036
rect 21700 7980 21710 8036
rect 21858 7980 21868 8036
rect 21924 7980 26908 8036
rect 27010 7980 27020 8036
rect 27076 7980 28476 8036
rect 28532 7980 28542 8036
rect 28700 7980 30380 8036
rect 30436 7980 30446 8036
rect 30706 7980 30716 8036
rect 30772 7980 32564 8036
rect 32946 7980 32956 8036
rect 33012 7980 46620 8036
rect 46676 7980 46686 8036
rect 26852 7924 26908 7980
rect 9426 7868 9436 7924
rect 9492 7868 16044 7924
rect 16100 7868 16110 7924
rect 16818 7868 16828 7924
rect 16884 7868 23436 7924
rect 23492 7868 23502 7924
rect 24322 7868 24332 7924
rect 24388 7868 25452 7924
rect 25508 7868 25518 7924
rect 25666 7868 25676 7924
rect 25732 7868 26684 7924
rect 26740 7868 26750 7924
rect 26852 7868 32060 7924
rect 32116 7868 32126 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 32508 7812 32564 7980
rect 32722 7868 32732 7924
rect 32788 7868 42028 7924
rect 42084 7868 42094 7924
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 9986 7756 9996 7812
rect 10052 7756 13580 7812
rect 13636 7756 13646 7812
rect 13794 7756 13804 7812
rect 13860 7756 17164 7812
rect 17220 7756 17230 7812
rect 19170 7756 19180 7812
rect 19236 7756 19852 7812
rect 19908 7756 19918 7812
rect 20066 7756 20076 7812
rect 20132 7756 23660 7812
rect 23716 7756 23726 7812
rect 24210 7756 24220 7812
rect 24276 7756 29596 7812
rect 29652 7756 29662 7812
rect 30258 7756 30268 7812
rect 30324 7756 32284 7812
rect 32340 7756 32350 7812
rect 32508 7756 33516 7812
rect 33572 7756 33582 7812
rect 33842 7756 33852 7812
rect 33908 7756 43708 7812
rect 0 7700 112 7728
rect 0 7644 1148 7700
rect 1204 7644 1214 7700
rect 2706 7644 2716 7700
rect 2772 7644 8316 7700
rect 8372 7644 8382 7700
rect 11442 7644 11452 7700
rect 11508 7644 16380 7700
rect 16436 7644 16446 7700
rect 16594 7644 16604 7700
rect 16660 7644 17724 7700
rect 17780 7644 17790 7700
rect 18498 7644 18508 7700
rect 18564 7644 25340 7700
rect 25396 7644 25406 7700
rect 26674 7644 26684 7700
rect 26740 7644 38556 7700
rect 38612 7644 38622 7700
rect 0 7616 112 7644
rect 43652 7588 43708 7756
rect 52640 7700 52752 7728
rect 51426 7644 51436 7700
rect 51492 7644 52752 7700
rect 52640 7616 52752 7644
rect 2258 7532 2268 7588
rect 2324 7532 15036 7588
rect 15092 7532 15102 7588
rect 15362 7532 15372 7588
rect 15428 7532 23324 7588
rect 23380 7532 23390 7588
rect 23660 7532 29092 7588
rect 29250 7532 29260 7588
rect 29316 7532 33180 7588
rect 33236 7532 33246 7588
rect 33394 7532 33404 7588
rect 33460 7532 33852 7588
rect 33908 7532 33918 7588
rect 35410 7532 35420 7588
rect 35476 7532 38556 7588
rect 38612 7532 38622 7588
rect 43652 7532 47404 7588
rect 47460 7532 47470 7588
rect 23660 7476 23716 7532
rect 130 7420 140 7476
rect 196 7420 10276 7476
rect 13682 7420 13692 7476
rect 13748 7420 16828 7476
rect 16884 7420 16894 7476
rect 17042 7420 17052 7476
rect 17108 7420 22148 7476
rect 22418 7420 22428 7476
rect 22484 7420 23716 7476
rect 23874 7420 23884 7476
rect 23940 7420 27580 7476
rect 27636 7420 27646 7476
rect 1250 7308 1260 7364
rect 1316 7308 6524 7364
rect 6580 7308 6590 7364
rect 0 7252 112 7280
rect 10220 7252 10276 7420
rect 22092 7364 22148 7420
rect 29036 7364 29092 7532
rect 29810 7420 29820 7476
rect 29876 7420 30380 7476
rect 30436 7420 30446 7476
rect 31042 7420 31052 7476
rect 31108 7420 31668 7476
rect 31826 7420 31836 7476
rect 31892 7420 37436 7476
rect 37492 7420 37502 7476
rect 38994 7420 39004 7476
rect 39060 7420 49532 7476
rect 49588 7420 49598 7476
rect 31612 7364 31668 7420
rect 12114 7308 12124 7364
rect 12180 7308 21868 7364
rect 21924 7308 21934 7364
rect 22092 7308 25172 7364
rect 25330 7308 25340 7364
rect 25396 7308 28812 7364
rect 28868 7308 28878 7364
rect 29036 7308 30940 7364
rect 30996 7308 31006 7364
rect 31612 7308 48748 7364
rect 48804 7308 48814 7364
rect 0 7196 6636 7252
rect 6692 7196 6702 7252
rect 10220 7196 24892 7252
rect 24948 7196 24958 7252
rect 0 7168 112 7196
rect 25116 7140 25172 7308
rect 52640 7252 52752 7280
rect 25330 7196 25340 7252
rect 25396 7196 29932 7252
rect 29988 7196 29998 7252
rect 30258 7196 30268 7252
rect 30324 7196 33012 7252
rect 33170 7196 33180 7252
rect 33236 7196 39676 7252
rect 39732 7196 39742 7252
rect 51426 7196 51436 7252
rect 51492 7196 52752 7252
rect 32956 7140 33012 7196
rect 52640 7168 52752 7196
rect 6402 7084 6412 7140
rect 6468 7084 11788 7140
rect 11844 7084 11854 7140
rect 16482 7084 16492 7140
rect 16548 7084 19180 7140
rect 19236 7084 19246 7140
rect 19394 7084 19404 7140
rect 19460 7084 22988 7140
rect 23044 7084 23054 7140
rect 25116 7084 32732 7140
rect 32788 7084 32798 7140
rect 32956 7084 34636 7140
rect 34692 7084 34702 7140
rect 35298 7084 35308 7140
rect 35364 7084 43596 7140
rect 43652 7084 43662 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 7868 6972 21196 7028
rect 21252 6972 21262 7028
rect 21522 6972 21532 7028
rect 21588 6972 22316 7028
rect 22372 6972 22382 7028
rect 24892 6972 25228 7028
rect 25284 6972 25294 7028
rect 25442 6972 25452 7028
rect 25508 6972 43708 7028
rect 354 6860 364 6916
rect 420 6860 2604 6916
rect 2660 6860 2670 6916
rect 0 6804 112 6832
rect 7868 6804 7924 6972
rect 24892 6916 24948 6972
rect 43652 6916 43708 6972
rect 13010 6860 13020 6916
rect 13076 6860 15932 6916
rect 15988 6860 15998 6916
rect 16594 6860 16604 6916
rect 16660 6860 20524 6916
rect 20580 6860 20590 6916
rect 20748 6860 24948 6916
rect 25106 6860 25116 6916
rect 25172 6860 26572 6916
rect 26628 6860 26638 6916
rect 26786 6860 26796 6916
rect 26852 6860 27188 6916
rect 27346 6860 27356 6916
rect 27412 6860 29372 6916
rect 29428 6860 29438 6916
rect 29586 6860 29596 6916
rect 29652 6860 31500 6916
rect 31556 6860 31566 6916
rect 32050 6860 32060 6916
rect 32116 6860 35308 6916
rect 35364 6860 35374 6916
rect 43652 6860 48524 6916
rect 48580 6860 48590 6916
rect 20748 6804 20804 6860
rect 27132 6804 27188 6860
rect 52640 6804 52752 6832
rect 0 6748 1428 6804
rect 0 6720 112 6748
rect 1372 6580 1428 6748
rect 6636 6748 7924 6804
rect 12226 6748 12236 6804
rect 12292 6748 16716 6804
rect 16772 6748 16782 6804
rect 16930 6748 16940 6804
rect 16996 6748 18060 6804
rect 18116 6748 18126 6804
rect 18274 6748 18284 6804
rect 18340 6748 20804 6804
rect 21186 6748 21196 6804
rect 21252 6748 26964 6804
rect 27132 6748 29036 6804
rect 29092 6748 29102 6804
rect 29372 6748 32844 6804
rect 32900 6748 32910 6804
rect 33628 6748 36988 6804
rect 37044 6748 37054 6804
rect 39106 6748 39116 6804
rect 39172 6748 49084 6804
rect 49140 6748 49150 6804
rect 49634 6748 49644 6804
rect 49700 6748 52752 6804
rect 6636 6692 6692 6748
rect 26908 6692 26964 6748
rect 29372 6692 29428 6748
rect 33628 6692 33684 6748
rect 52640 6720 52752 6748
rect 1586 6636 1596 6692
rect 1652 6636 6692 6692
rect 11890 6636 11900 6692
rect 11956 6636 16492 6692
rect 16548 6636 16558 6692
rect 16930 6636 16940 6692
rect 16996 6636 18732 6692
rect 18788 6636 18798 6692
rect 19394 6636 19404 6692
rect 19460 6636 21532 6692
rect 21588 6636 21598 6692
rect 21746 6636 21756 6692
rect 21812 6636 22764 6692
rect 22820 6636 22830 6692
rect 23314 6636 23324 6692
rect 23380 6636 26012 6692
rect 26068 6636 26078 6692
rect 26908 6636 27244 6692
rect 27300 6636 27310 6692
rect 27468 6636 29428 6692
rect 31826 6636 31836 6692
rect 31892 6636 33684 6692
rect 33842 6636 33852 6692
rect 33908 6636 45388 6692
rect 45444 6636 45454 6692
rect 46274 6636 46284 6692
rect 46340 6636 48860 6692
rect 48916 6636 48926 6692
rect 27468 6580 27524 6636
rect 1372 6524 1820 6580
rect 1876 6524 1886 6580
rect 2044 6524 3388 6580
rect 5394 6524 5404 6580
rect 5460 6524 6860 6580
rect 6916 6524 6926 6580
rect 7970 6524 7980 6580
rect 8036 6524 13804 6580
rect 13860 6524 13870 6580
rect 15138 6524 15148 6580
rect 15204 6524 22092 6580
rect 22148 6524 22158 6580
rect 22306 6524 22316 6580
rect 22372 6524 27132 6580
rect 27188 6524 27198 6580
rect 27356 6524 27524 6580
rect 28466 6524 28476 6580
rect 28532 6524 29596 6580
rect 29652 6524 29662 6580
rect 29922 6524 29932 6580
rect 29988 6524 33628 6580
rect 33684 6524 33694 6580
rect 33842 6524 33852 6580
rect 33908 6524 36092 6580
rect 36148 6524 36158 6580
rect 37314 6524 37324 6580
rect 37380 6524 40460 6580
rect 40516 6524 40526 6580
rect 40786 6524 40796 6580
rect 40852 6524 44604 6580
rect 44660 6524 44670 6580
rect 2044 6468 2100 6524
rect 1474 6412 1484 6468
rect 1540 6412 2100 6468
rect 3332 6468 3388 6524
rect 27356 6468 27412 6524
rect 3332 6412 9212 6468
rect 9268 6412 9278 6468
rect 9874 6412 9884 6468
rect 9940 6412 24276 6468
rect 24434 6412 24444 6468
rect 24500 6412 25676 6468
rect 25732 6412 25742 6468
rect 26002 6412 26012 6468
rect 26068 6412 27412 6468
rect 27570 6412 27580 6468
rect 27636 6412 48524 6468
rect 48580 6412 48590 6468
rect 0 6356 112 6384
rect 24220 6356 24276 6412
rect 52640 6356 52752 6384
rect 0 6300 1372 6356
rect 1428 6300 1438 6356
rect 1922 6300 1932 6356
rect 1988 6300 3612 6356
rect 3668 6300 3678 6356
rect 8306 6300 8316 6356
rect 8372 6300 15036 6356
rect 15092 6300 15102 6356
rect 15810 6300 15820 6356
rect 15876 6300 18172 6356
rect 18228 6300 18238 6356
rect 18386 6300 18396 6356
rect 18452 6300 19292 6356
rect 19348 6300 19358 6356
rect 19506 6300 19516 6356
rect 19572 6300 21196 6356
rect 21252 6300 21262 6356
rect 21410 6300 21420 6356
rect 21476 6300 22316 6356
rect 22372 6300 22382 6356
rect 22530 6300 22540 6356
rect 22596 6300 23548 6356
rect 23604 6300 23614 6356
rect 24220 6300 30604 6356
rect 30660 6300 30670 6356
rect 36978 6300 36988 6356
rect 37044 6300 43148 6356
rect 43204 6300 43214 6356
rect 51202 6300 51212 6356
rect 51268 6300 52752 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 52640 6272 52752 6300
rect 6738 6188 6748 6244
rect 6804 6188 16268 6244
rect 16324 6188 16334 6244
rect 16482 6188 16492 6244
rect 16548 6188 17948 6244
rect 18004 6188 18014 6244
rect 19170 6188 19180 6244
rect 19236 6188 23660 6244
rect 23716 6188 23726 6244
rect 24210 6188 24220 6244
rect 24276 6188 26684 6244
rect 26740 6188 26750 6244
rect 28018 6188 28028 6244
rect 28084 6188 34524 6244
rect 34580 6188 34590 6244
rect 35074 6188 35084 6244
rect 35140 6188 37548 6244
rect 37604 6188 37614 6244
rect 12226 6076 12236 6132
rect 12292 6076 19404 6132
rect 19460 6076 19470 6132
rect 19842 6076 19852 6132
rect 19908 6076 20076 6132
rect 20132 6076 20142 6132
rect 21858 6076 21868 6132
rect 21924 6076 29484 6132
rect 29540 6076 29550 6132
rect 29810 6076 29820 6132
rect 29876 6076 34748 6132
rect 34804 6076 34814 6132
rect 36978 6076 36988 6132
rect 37044 6076 39900 6132
rect 39956 6076 39966 6132
rect 10210 5964 10220 6020
rect 10276 5964 18060 6020
rect 18116 5964 18126 6020
rect 18498 5964 18508 6020
rect 18564 5964 23772 6020
rect 23828 5964 23838 6020
rect 24322 5964 24332 6020
rect 24388 5964 27468 6020
rect 27524 5964 27534 6020
rect 31714 5964 31724 6020
rect 31780 5964 38220 6020
rect 38276 5964 38286 6020
rect 47394 5964 47404 6020
rect 47460 5964 49868 6020
rect 49924 5964 49934 6020
rect 0 5908 112 5936
rect 52640 5908 52752 5936
rect 0 5852 1372 5908
rect 1428 5852 1438 5908
rect 13682 5852 13692 5908
rect 13748 5852 16604 5908
rect 16660 5852 16670 5908
rect 17602 5852 17612 5908
rect 17668 5852 18396 5908
rect 18452 5852 18462 5908
rect 18722 5852 18732 5908
rect 18788 5852 25060 5908
rect 25218 5852 25228 5908
rect 25284 5852 31836 5908
rect 31892 5852 31902 5908
rect 0 5824 112 5852
rect 25004 5796 25060 5852
rect 38612 5796 38668 5908
rect 38724 5852 38734 5908
rect 44258 5852 44268 5908
rect 44324 5852 49308 5908
rect 49364 5852 49374 5908
rect 49746 5852 49756 5908
rect 49812 5852 52752 5908
rect 52640 5824 52752 5852
rect 3378 5740 3388 5796
rect 3444 5740 10332 5796
rect 10388 5740 10398 5796
rect 13458 5740 13468 5796
rect 13524 5740 16492 5796
rect 16548 5740 16558 5796
rect 16706 5740 16716 5796
rect 16772 5740 24948 5796
rect 25004 5740 29148 5796
rect 29204 5740 29214 5796
rect 30146 5740 30156 5796
rect 30212 5740 38668 5796
rect 39218 5740 39228 5796
rect 39284 5740 46172 5796
rect 46228 5740 46238 5796
rect 24892 5684 24948 5740
rect 2930 5628 2940 5684
rect 2996 5628 5852 5684
rect 5908 5628 5918 5684
rect 10994 5628 11004 5684
rect 11060 5628 18396 5684
rect 18452 5628 18462 5684
rect 18620 5628 24220 5684
rect 24276 5628 24286 5684
rect 24892 5628 25060 5684
rect 26114 5628 26124 5684
rect 26180 5628 27020 5684
rect 27076 5628 27086 5684
rect 27468 5628 32844 5684
rect 32900 5628 32910 5684
rect 33394 5628 33404 5684
rect 33460 5628 37772 5684
rect 37828 5628 37838 5684
rect 37996 5628 42140 5684
rect 42196 5628 42206 5684
rect 43922 5628 43932 5684
rect 43988 5628 48076 5684
rect 48132 5628 48142 5684
rect 18620 5572 18676 5628
rect 25004 5572 25060 5628
rect 27468 5572 27524 5628
rect 37996 5572 38052 5628
rect 9090 5516 9100 5572
rect 9156 5516 15036 5572
rect 15092 5516 15102 5572
rect 16482 5516 16492 5572
rect 16548 5516 18676 5572
rect 18834 5516 18844 5572
rect 18900 5516 22820 5572
rect 23538 5516 23548 5572
rect 23604 5516 24220 5572
rect 24276 5516 24286 5572
rect 25004 5516 27524 5572
rect 27682 5516 27692 5572
rect 27748 5516 34076 5572
rect 34132 5516 34142 5572
rect 36866 5516 36876 5572
rect 36932 5516 38052 5572
rect 38210 5516 38220 5572
rect 38276 5516 40348 5572
rect 40404 5516 40414 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 22764 5460 22820 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 52640 5460 52752 5488
rect 0 5404 3164 5460
rect 3220 5404 3230 5460
rect 8978 5404 8988 5460
rect 9044 5404 16716 5460
rect 16772 5404 16782 5460
rect 17826 5404 17836 5460
rect 17892 5404 22540 5460
rect 22596 5404 22606 5460
rect 22764 5404 24332 5460
rect 24388 5404 24398 5460
rect 24882 5404 24892 5460
rect 24948 5404 26012 5460
rect 26068 5404 26078 5460
rect 26338 5404 26348 5460
rect 26404 5404 29260 5460
rect 29316 5404 29326 5460
rect 31938 5404 31948 5460
rect 32004 5404 40572 5460
rect 40628 5404 40638 5460
rect 49074 5404 49084 5460
rect 49140 5404 50764 5460
rect 50820 5404 50830 5460
rect 51202 5404 51212 5460
rect 51268 5404 52752 5460
rect 0 5376 112 5404
rect 52640 5376 52752 5404
rect 6402 5292 6412 5348
rect 6468 5292 15036 5348
rect 15092 5292 15102 5348
rect 15586 5292 15596 5348
rect 15652 5292 18508 5348
rect 18564 5292 18574 5348
rect 19282 5292 19292 5348
rect 19348 5292 20076 5348
rect 20132 5292 20142 5348
rect 20290 5292 20300 5348
rect 20356 5292 21308 5348
rect 21364 5292 21374 5348
rect 21522 5292 21532 5348
rect 21588 5292 25956 5348
rect 26114 5292 26124 5348
rect 26180 5292 29372 5348
rect 29428 5292 29438 5348
rect 29586 5292 29596 5348
rect 29652 5292 50204 5348
rect 50260 5292 50270 5348
rect 25900 5236 25956 5292
rect 6514 5180 6524 5236
rect 6580 5180 13916 5236
rect 13972 5180 13982 5236
rect 14242 5180 14252 5236
rect 14308 5180 15260 5236
rect 15316 5180 15326 5236
rect 15474 5180 15484 5236
rect 15540 5180 16380 5236
rect 16436 5180 16446 5236
rect 16930 5180 16940 5236
rect 16996 5180 25676 5236
rect 25732 5180 25742 5236
rect 25900 5180 30436 5236
rect 30594 5180 30604 5236
rect 30660 5180 37884 5236
rect 37940 5180 37950 5236
rect 39116 5180 45052 5236
rect 45108 5180 45118 5236
rect 45276 5180 49420 5236
rect 49476 5180 49486 5236
rect 8530 5068 8540 5124
rect 8596 5068 16268 5124
rect 16324 5068 16334 5124
rect 16930 5068 16940 5124
rect 16996 5068 21308 5124
rect 21364 5068 21374 5124
rect 21746 5068 21756 5124
rect 21812 5068 24892 5124
rect 24948 5068 24958 5124
rect 25106 5068 25116 5124
rect 25172 5068 29932 5124
rect 29988 5068 29998 5124
rect 0 5012 112 5040
rect 30380 5012 30436 5180
rect 35308 5068 38892 5124
rect 38948 5068 38958 5124
rect 35308 5012 35364 5068
rect 0 4956 9268 5012
rect 10434 4956 10444 5012
rect 10500 4956 16492 5012
rect 16548 4956 16558 5012
rect 17042 4956 17052 5012
rect 17108 4956 21868 5012
rect 21924 4956 21934 5012
rect 22978 4956 22988 5012
rect 23044 4956 30100 5012
rect 30380 4956 35364 5012
rect 35522 4956 35532 5012
rect 35588 4956 37324 5012
rect 37380 4956 37390 5012
rect 0 4928 112 4956
rect 9212 4900 9268 4956
rect 30044 4900 30100 4956
rect 39116 4900 39172 5180
rect 45276 5124 45332 5180
rect 39442 5068 39452 5124
rect 39508 5068 45332 5124
rect 49634 5068 49644 5124
rect 49700 5068 51100 5124
rect 51156 5068 51166 5124
rect 52640 5012 52752 5040
rect 39554 4956 39564 5012
rect 39620 4956 43932 5012
rect 43988 4956 43998 5012
rect 45490 4956 45500 5012
rect 45556 4956 48748 5012
rect 48804 4956 48814 5012
rect 51202 4956 51212 5012
rect 51268 4956 52752 5012
rect 52640 4928 52752 4956
rect 1810 4844 1820 4900
rect 1876 4844 6020 4900
rect 9212 4844 11900 4900
rect 11956 4844 11966 4900
rect 14914 4844 14924 4900
rect 14980 4844 18844 4900
rect 18900 4844 18910 4900
rect 19058 4844 19068 4900
rect 19124 4844 20076 4900
rect 20132 4844 20142 4900
rect 20290 4844 20300 4900
rect 20356 4844 29820 4900
rect 29876 4844 29886 4900
rect 30044 4844 39172 4900
rect 40226 4844 40236 4900
rect 40292 4844 45836 4900
rect 45892 4844 45902 4900
rect 5964 4788 6020 4844
rect 1026 4732 1036 4788
rect 1092 4732 3052 4788
rect 3108 4732 3118 4788
rect 4162 4732 4172 4788
rect 4228 4732 5628 4788
rect 5684 4732 5694 4788
rect 5964 4732 15932 4788
rect 15988 4732 15998 4788
rect 16156 4732 16548 4788
rect 17042 4732 17052 4788
rect 17108 4732 23548 4788
rect 23604 4732 23614 4788
rect 24210 4732 24220 4788
rect 24276 4732 25564 4788
rect 25620 4732 25630 4788
rect 25778 4732 25788 4788
rect 25844 4732 35532 4788
rect 35588 4732 35598 4788
rect 37202 4732 37212 4788
rect 37268 4732 40684 4788
rect 40740 4732 40750 4788
rect 45938 4732 45948 4788
rect 46004 4732 50204 4788
rect 50260 4732 50270 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 16156 4676 16212 4732
rect 2156 4620 3276 4676
rect 3332 4620 3342 4676
rect 11666 4620 11676 4676
rect 11732 4620 16212 4676
rect 16492 4676 16548 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 16492 4620 17500 4676
rect 17556 4620 17566 4676
rect 18162 4620 18172 4676
rect 18228 4620 21868 4676
rect 21924 4620 21934 4676
rect 22082 4620 22092 4676
rect 22148 4620 23436 4676
rect 23492 4620 23502 4676
rect 24322 4620 24332 4676
rect 24388 4620 25004 4676
rect 25060 4620 25070 4676
rect 25218 4620 25228 4676
rect 25284 4620 36988 4676
rect 37044 4620 37054 4676
rect 38612 4620 40236 4676
rect 40292 4620 40302 4676
rect 0 4564 112 4592
rect 2156 4564 2212 4620
rect 38612 4564 38668 4620
rect 52640 4564 52752 4592
rect 0 4508 2212 4564
rect 2370 4508 2380 4564
rect 2436 4508 8540 4564
rect 8596 4508 8606 4564
rect 12786 4508 12796 4564
rect 12852 4508 15932 4564
rect 15988 4508 15998 4564
rect 16146 4508 16156 4564
rect 16212 4508 18172 4564
rect 18228 4508 18238 4564
rect 18386 4508 18396 4564
rect 18452 4508 28476 4564
rect 28532 4508 28542 4564
rect 29026 4508 29036 4564
rect 29092 4508 33068 4564
rect 33124 4508 33134 4564
rect 35298 4508 35308 4564
rect 35364 4508 38668 4564
rect 40338 4508 40348 4564
rect 40404 4508 48188 4564
rect 48244 4508 48254 4564
rect 51090 4508 51100 4564
rect 51156 4508 52752 4564
rect 0 4480 112 4508
rect 52640 4480 52752 4508
rect 3602 4396 3612 4452
rect 3668 4396 15148 4452
rect 15204 4396 15214 4452
rect 16492 4396 23324 4452
rect 23380 4396 23390 4452
rect 23538 4396 23548 4452
rect 23604 4396 25900 4452
rect 25956 4396 25966 4452
rect 26114 4396 26124 4452
rect 26180 4396 30156 4452
rect 30212 4396 30222 4452
rect 32162 4396 32172 4452
rect 32228 4396 40908 4452
rect 40964 4396 40974 4452
rect 2258 4284 2268 4340
rect 2324 4284 8316 4340
rect 8372 4284 8382 4340
rect 11778 4284 11788 4340
rect 11844 4284 16268 4340
rect 16324 4284 16334 4340
rect 16492 4228 16548 4396
rect 17714 4284 17724 4340
rect 17780 4284 19628 4340
rect 19684 4284 19694 4340
rect 19954 4284 19964 4340
rect 20020 4284 21532 4340
rect 21588 4284 21598 4340
rect 21858 4284 21868 4340
rect 21924 4284 27020 4340
rect 27076 4284 27086 4340
rect 27234 4284 27244 4340
rect 27300 4284 33180 4340
rect 33236 4284 33246 4340
rect 37986 4284 37996 4340
rect 38052 4284 46732 4340
rect 46788 4284 46798 4340
rect 2594 4172 2604 4228
rect 2660 4172 5404 4228
rect 5460 4172 5470 4228
rect 15026 4172 15036 4228
rect 15092 4172 16548 4228
rect 16706 4172 16716 4228
rect 16772 4172 18564 4228
rect 0 4116 112 4144
rect 18508 4116 18564 4172
rect 19852 4172 24556 4228
rect 24612 4172 24622 4228
rect 24780 4172 28028 4228
rect 28084 4172 28094 4228
rect 30370 4172 30380 4228
rect 30436 4172 32956 4228
rect 33012 4172 33022 4228
rect 35746 4172 35756 4228
rect 35812 4172 44156 4228
rect 44212 4172 44222 4228
rect 19852 4116 19908 4172
rect 24780 4116 24836 4172
rect 52640 4116 52752 4144
rect 0 4060 1484 4116
rect 1540 4060 1550 4116
rect 5058 4060 5068 4116
rect 5124 4060 18284 4116
rect 18340 4060 18350 4116
rect 18508 4060 19908 4116
rect 20066 4060 20076 4116
rect 20132 4060 21308 4116
rect 21364 4060 21374 4116
rect 21522 4060 21532 4116
rect 21588 4060 24836 4116
rect 27010 4060 27020 4116
rect 27076 4060 30044 4116
rect 30100 4060 30110 4116
rect 30258 4060 30268 4116
rect 30324 4060 42812 4116
rect 42868 4060 42878 4116
rect 51426 4060 51436 4116
rect 51492 4060 52752 4116
rect 0 4032 112 4060
rect 52640 4032 52752 4060
rect 7298 3948 7308 4004
rect 7364 3948 13692 4004
rect 13748 3948 13758 4004
rect 14466 3948 14476 4004
rect 14532 3948 20636 4004
rect 20692 3948 20702 4004
rect 20962 3948 20972 4004
rect 21028 3948 22092 4004
rect 22148 3948 22158 4004
rect 22642 3948 22652 4004
rect 22708 3948 24332 4004
rect 24388 3948 24398 4004
rect 25106 3948 25116 4004
rect 25172 3948 38780 4004
rect 38836 3948 38846 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 6626 3836 6636 3892
rect 6692 3836 16100 3892
rect 16258 3836 16268 3892
rect 16324 3836 24220 3892
rect 24276 3836 24286 3892
rect 24994 3836 25004 3892
rect 25060 3836 25620 3892
rect 27010 3836 27020 3892
rect 27076 3836 43708 3892
rect 16044 3780 16100 3836
rect 25564 3780 25620 3836
rect 43652 3780 43708 3836
rect 45052 3836 48860 3892
rect 48916 3836 48926 3892
rect 45052 3780 45108 3836
rect 11218 3724 11228 3780
rect 11284 3724 15036 3780
rect 15092 3724 15102 3780
rect 16044 3724 16940 3780
rect 16996 3724 17006 3780
rect 17154 3724 17164 3780
rect 17220 3724 25340 3780
rect 25396 3724 25406 3780
rect 25564 3724 31948 3780
rect 32004 3724 32014 3780
rect 32620 3724 39004 3780
rect 39060 3724 39070 3780
rect 43652 3724 45108 3780
rect 45266 3724 45276 3780
rect 45332 3724 50428 3780
rect 50484 3724 50494 3780
rect 0 3668 112 3696
rect 32620 3668 32676 3724
rect 52640 3668 52752 3696
rect 0 3612 1596 3668
rect 1652 3612 1662 3668
rect 13682 3612 13692 3668
rect 13748 3612 21084 3668
rect 21140 3612 21150 3668
rect 21298 3612 21308 3668
rect 21364 3612 27804 3668
rect 27860 3612 27870 3668
rect 28018 3612 28028 3668
rect 28084 3612 32676 3668
rect 33506 3612 33516 3668
rect 33572 3612 37436 3668
rect 37492 3612 37502 3668
rect 38770 3612 38780 3668
rect 38836 3612 46396 3668
rect 46452 3612 46462 3668
rect 46610 3612 46620 3668
rect 46676 3612 48860 3668
rect 48916 3612 48926 3668
rect 49410 3612 49420 3668
rect 49476 3612 52752 3668
rect 0 3584 112 3612
rect 52640 3584 52752 3612
rect 13794 3500 13804 3556
rect 13860 3500 15708 3556
rect 15764 3500 15774 3556
rect 16370 3500 16380 3556
rect 16436 3500 18844 3556
rect 18900 3500 18910 3556
rect 19954 3500 19964 3556
rect 20020 3500 29820 3556
rect 29876 3500 29886 3556
rect 39666 3500 39676 3556
rect 39732 3500 44716 3556
rect 44772 3500 44782 3556
rect 1596 3388 2716 3444
rect 2772 3388 2782 3444
rect 8418 3388 8428 3444
rect 8484 3388 11788 3444
rect 12562 3388 12572 3444
rect 12628 3388 14476 3444
rect 14532 3388 14542 3444
rect 14690 3388 14700 3444
rect 14756 3388 20412 3444
rect 20468 3388 20478 3444
rect 20626 3388 20636 3444
rect 20692 3388 21084 3444
rect 21140 3388 21150 3444
rect 21634 3388 21644 3444
rect 21700 3388 21924 3444
rect 22082 3388 22092 3444
rect 22148 3388 24556 3444
rect 24612 3388 24622 3444
rect 25106 3388 25116 3444
rect 25172 3388 29372 3444
rect 29428 3388 29438 3444
rect 29596 3388 36932 3444
rect 46386 3388 46396 3444
rect 46452 3388 49196 3444
rect 49252 3388 49262 3444
rect 49858 3388 49868 3444
rect 49924 3388 51100 3444
rect 51156 3388 51166 3444
rect 0 3220 112 3248
rect 1596 3220 1652 3388
rect 11732 3332 11788 3388
rect 21868 3332 21924 3388
rect 29596 3332 29652 3388
rect 36876 3332 36932 3388
rect 11732 3276 12796 3332
rect 12852 3276 12862 3332
rect 13682 3276 13692 3332
rect 13748 3276 18508 3332
rect 18564 3276 18574 3332
rect 18834 3276 18844 3332
rect 18900 3276 19964 3332
rect 20020 3276 20030 3332
rect 20290 3276 20300 3332
rect 20356 3276 21308 3332
rect 21364 3276 21374 3332
rect 21868 3276 21980 3332
rect 22036 3276 22046 3332
rect 22204 3276 27580 3332
rect 27636 3276 27646 3332
rect 27794 3276 27804 3332
rect 27860 3276 29652 3332
rect 30370 3276 30380 3332
rect 30436 3276 36652 3332
rect 36708 3276 36718 3332
rect 36876 3276 38892 3332
rect 38948 3276 38958 3332
rect 43652 3276 47740 3332
rect 47796 3276 47806 3332
rect 22204 3220 22260 3276
rect 0 3164 1652 3220
rect 6066 3164 6076 3220
rect 6132 3164 6636 3220
rect 6692 3164 6702 3220
rect 11330 3164 11340 3220
rect 11396 3164 18732 3220
rect 18788 3164 18798 3220
rect 18946 3164 18956 3220
rect 19012 3164 22260 3220
rect 22418 3164 22428 3220
rect 22484 3164 23324 3220
rect 23380 3164 23390 3220
rect 24210 3164 24220 3220
rect 24276 3164 26348 3220
rect 26404 3164 26414 3220
rect 26562 3164 26572 3220
rect 26628 3164 32172 3220
rect 32228 3164 32238 3220
rect 32386 3164 32396 3220
rect 32452 3164 35980 3220
rect 36036 3164 36046 3220
rect 36642 3164 36652 3220
rect 36708 3164 40348 3220
rect 40404 3164 40414 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 43652 3108 43708 3276
rect 52640 3220 52752 3248
rect 51202 3164 51212 3220
rect 51268 3164 52752 3220
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 52640 3136 52752 3164
rect 13906 3052 13916 3108
rect 13972 3052 16940 3108
rect 16996 3052 17006 3108
rect 17164 3052 20972 3108
rect 21028 3052 21038 3108
rect 21186 3052 21196 3108
rect 21252 3052 23660 3108
rect 23716 3052 23726 3108
rect 24322 3052 24332 3108
rect 24388 3052 27916 3108
rect 27972 3052 27982 3108
rect 30370 3052 30380 3108
rect 30436 3052 43708 3108
rect 17164 2996 17220 3052
rect 2146 2940 2156 2996
rect 2212 2940 11564 2996
rect 11620 2940 11630 2996
rect 11778 2940 11788 2996
rect 11844 2940 13468 2996
rect 13524 2940 13534 2996
rect 15474 2940 15484 2996
rect 15540 2940 17220 2996
rect 18274 2940 18284 2996
rect 18340 2940 20300 2996
rect 20356 2940 20366 2996
rect 20738 2940 20748 2996
rect 20804 2940 31836 2996
rect 31892 2940 31902 2996
rect 37650 2940 37660 2996
rect 37716 2940 46956 2996
rect 47012 2940 47022 2996
rect 3938 2828 3948 2884
rect 4004 2828 7756 2884
rect 7812 2828 7822 2884
rect 10882 2828 10892 2884
rect 10948 2828 15820 2884
rect 15876 2828 15886 2884
rect 16146 2828 16156 2884
rect 16212 2828 16828 2884
rect 16884 2828 16894 2884
rect 17052 2828 22596 2884
rect 23538 2828 23548 2884
rect 23604 2828 33404 2884
rect 33460 2828 33470 2884
rect 34514 2828 34524 2884
rect 34580 2828 37212 2884
rect 37268 2828 37278 2884
rect 38322 2828 38332 2884
rect 38388 2828 47068 2884
rect 47124 2828 47134 2884
rect 48066 2828 48076 2884
rect 48132 2828 50540 2884
rect 50596 2828 50606 2884
rect 0 2772 112 2800
rect 17052 2772 17108 2828
rect 22540 2772 22596 2828
rect 52640 2772 52752 2800
rect 0 2716 1036 2772
rect 1092 2716 1102 2772
rect 3154 2716 3164 2772
rect 3220 2716 13692 2772
rect 13748 2716 13758 2772
rect 15474 2716 15484 2772
rect 15540 2716 16324 2772
rect 16482 2716 16492 2772
rect 16548 2716 17108 2772
rect 17378 2716 17388 2772
rect 17444 2716 22316 2772
rect 22372 2716 22382 2772
rect 22540 2716 25340 2772
rect 25396 2716 25406 2772
rect 25554 2716 25564 2772
rect 25620 2716 26684 2772
rect 26740 2716 26750 2772
rect 28578 2716 28588 2772
rect 28644 2716 32732 2772
rect 32788 2716 32798 2772
rect 36642 2716 36652 2772
rect 36708 2716 38836 2772
rect 40226 2716 40236 2772
rect 40292 2716 45388 2772
rect 45444 2716 45454 2772
rect 46162 2716 46172 2772
rect 46228 2716 48748 2772
rect 48804 2716 48814 2772
rect 51090 2716 51100 2772
rect 51156 2716 52752 2772
rect 0 2688 112 2716
rect 16268 2660 16324 2716
rect 38780 2660 38836 2716
rect 52640 2688 52752 2716
rect 1362 2604 1372 2660
rect 1428 2604 3388 2660
rect 4386 2604 4396 2660
rect 4452 2604 6412 2660
rect 6468 2604 6478 2660
rect 6626 2604 6636 2660
rect 6692 2604 13916 2660
rect 13972 2604 13982 2660
rect 14130 2604 14140 2660
rect 14196 2604 16044 2660
rect 16100 2604 16110 2660
rect 16268 2604 18284 2660
rect 18340 2604 18350 2660
rect 19618 2604 19628 2660
rect 19684 2604 30268 2660
rect 30324 2604 30334 2660
rect 30482 2604 30492 2660
rect 30548 2604 37660 2660
rect 37716 2604 37726 2660
rect 38780 2604 41244 2660
rect 41300 2604 41310 2660
rect 49410 2604 49420 2660
rect 49476 2604 51548 2660
rect 51604 2604 51614 2660
rect 3332 2548 3388 2604
rect 3332 2492 32844 2548
rect 32900 2492 32910 2548
rect 33394 2492 33404 2548
rect 33460 2492 46284 2548
rect 46340 2492 46350 2548
rect 10210 2380 10220 2436
rect 10276 2380 14308 2436
rect 15138 2380 15148 2436
rect 15204 2380 15932 2436
rect 15988 2380 15998 2436
rect 16146 2380 16156 2436
rect 16212 2380 24332 2436
rect 24388 2380 24398 2436
rect 24882 2380 24892 2436
rect 24948 2380 26460 2436
rect 26516 2380 26526 2436
rect 26674 2380 26684 2436
rect 26740 2380 30156 2436
rect 30212 2380 30222 2436
rect 33170 2380 33180 2436
rect 33236 2380 35532 2436
rect 35588 2380 35598 2436
rect 47506 2380 47516 2436
rect 47572 2380 50428 2436
rect 50484 2380 50494 2436
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 14252 2324 14308 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 52640 2324 52752 2352
rect 0 2268 1260 2324
rect 1316 2268 1326 2324
rect 13346 2268 13356 2324
rect 13412 2268 14196 2324
rect 14252 2268 16604 2324
rect 16660 2268 16670 2324
rect 16818 2268 16828 2324
rect 16884 2268 21196 2324
rect 21252 2268 21262 2324
rect 21634 2268 21644 2324
rect 21700 2268 22204 2324
rect 22260 2268 22270 2324
rect 22428 2268 23996 2324
rect 24052 2268 24062 2324
rect 24892 2268 30492 2324
rect 30548 2268 30558 2324
rect 51426 2268 51436 2324
rect 51492 2268 52752 2324
rect 0 2240 112 2268
rect 14140 2212 14196 2268
rect 22428 2212 22484 2268
rect 24892 2212 24948 2268
rect 52640 2240 52752 2268
rect 1474 2156 1484 2212
rect 1540 2156 12572 2212
rect 12628 2156 12638 2212
rect 12786 2156 12796 2212
rect 12852 2156 13916 2212
rect 13972 2156 13982 2212
rect 14140 2156 18396 2212
rect 18452 2156 18462 2212
rect 18610 2156 18620 2212
rect 18676 2156 19236 2212
rect 19506 2156 19516 2212
rect 19572 2156 21756 2212
rect 21812 2156 21822 2212
rect 21970 2156 21980 2212
rect 22036 2156 22484 2212
rect 22866 2156 22876 2212
rect 22932 2156 24948 2212
rect 32274 2156 32284 2212
rect 32340 2156 50316 2212
rect 50372 2156 50382 2212
rect 19180 2100 19236 2156
rect 1260 2044 2268 2100
rect 2324 2044 2334 2100
rect 8194 2044 8204 2100
rect 8260 2044 14140 2100
rect 14196 2044 14206 2100
rect 14914 2044 14924 2100
rect 14980 2044 15596 2100
rect 15652 2044 15662 2100
rect 15922 2044 15932 2100
rect 15988 2044 18956 2100
rect 19012 2044 19022 2100
rect 19180 2044 19964 2100
rect 20020 2044 20030 2100
rect 20178 2044 20188 2100
rect 20244 2044 21980 2100
rect 22036 2044 22046 2100
rect 22194 2044 22204 2100
rect 22260 2044 26628 2100
rect 26786 2044 26796 2100
rect 26852 2044 35420 2100
rect 35476 2044 35486 2100
rect 39666 2044 39676 2100
rect 39732 2044 43372 2100
rect 43428 2044 43438 2100
rect 45938 2044 45948 2100
rect 46004 2044 48860 2100
rect 48916 2044 48926 2100
rect 0 1876 112 1904
rect 1260 1876 1316 2044
rect 26572 1988 26628 2044
rect 1586 1932 1596 1988
rect 1652 1932 13020 1988
rect 13076 1932 13086 1988
rect 13906 1932 13916 1988
rect 13972 1932 15484 1988
rect 15540 1932 15550 1988
rect 15698 1932 15708 1988
rect 15764 1932 20524 1988
rect 20580 1932 20590 1988
rect 20850 1932 20860 1988
rect 20916 1932 26348 1988
rect 26404 1932 26414 1988
rect 26572 1932 27692 1988
rect 27748 1932 27758 1988
rect 52640 1876 52752 1904
rect 0 1820 1316 1876
rect 1474 1820 1484 1876
rect 1540 1820 10108 1876
rect 10164 1820 10174 1876
rect 14466 1820 14476 1876
rect 14532 1820 19852 1876
rect 19908 1820 19918 1876
rect 20076 1820 21196 1876
rect 21252 1820 21262 1876
rect 21410 1820 21420 1876
rect 21476 1820 21756 1876
rect 21812 1820 21822 1876
rect 22082 1820 22092 1876
rect 22148 1820 44268 1876
rect 44324 1820 44334 1876
rect 49858 1820 49868 1876
rect 49924 1820 52752 1876
rect 0 1792 112 1820
rect 20076 1764 20132 1820
rect 52640 1792 52752 1820
rect 6636 1708 16716 1764
rect 16772 1708 16782 1764
rect 16930 1708 16940 1764
rect 16996 1708 18844 1764
rect 18900 1708 18910 1764
rect 19058 1708 19068 1764
rect 19124 1708 20132 1764
rect 20514 1708 20524 1764
rect 20580 1708 21980 1764
rect 22036 1708 22046 1764
rect 22194 1708 22204 1764
rect 22260 1708 28476 1764
rect 28532 1708 28542 1764
rect 29036 1708 34412 1764
rect 34468 1708 34478 1764
rect 40348 1708 47068 1764
rect 47124 1708 47134 1764
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 0 1428 112 1456
rect 6636 1428 6692 1708
rect 29036 1652 29092 1708
rect 10098 1596 10108 1652
rect 10164 1596 23548 1652
rect 23604 1596 23614 1652
rect 24210 1596 24220 1652
rect 24276 1596 29092 1652
rect 31938 1596 31948 1652
rect 32004 1596 32676 1652
rect 35410 1596 35420 1652
rect 35476 1596 39116 1652
rect 39172 1596 39182 1652
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 32620 1540 32676 1596
rect 40348 1540 40404 1708
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 10658 1484 10668 1540
rect 10724 1484 16156 1540
rect 16212 1484 16222 1540
rect 16594 1484 16604 1540
rect 16660 1484 19180 1540
rect 19236 1484 19246 1540
rect 19394 1484 19404 1540
rect 19460 1484 21308 1540
rect 21364 1484 21374 1540
rect 21746 1484 21756 1540
rect 21812 1484 23660 1540
rect 23716 1484 23726 1540
rect 24210 1484 24220 1540
rect 24276 1484 25452 1540
rect 25508 1484 25518 1540
rect 25666 1484 25676 1540
rect 25732 1484 32396 1540
rect 32452 1484 32462 1540
rect 32620 1484 40404 1540
rect 52640 1428 52752 1456
rect 0 1372 1428 1428
rect 1586 1372 1596 1428
rect 1652 1372 6692 1428
rect 11778 1372 11788 1428
rect 11844 1372 17052 1428
rect 17108 1372 17118 1428
rect 17266 1372 17276 1428
rect 17332 1372 18620 1428
rect 18676 1372 18686 1428
rect 18834 1372 18844 1428
rect 18900 1372 20860 1428
rect 20916 1372 20926 1428
rect 21074 1372 21084 1428
rect 21140 1372 27020 1428
rect 27076 1372 27086 1428
rect 28466 1372 28476 1428
rect 28532 1372 35084 1428
rect 35140 1372 35150 1428
rect 37874 1372 37884 1428
rect 37940 1372 43708 1428
rect 49746 1372 49756 1428
rect 49812 1372 52752 1428
rect 0 1344 112 1372
rect 1372 1316 1428 1372
rect 43652 1316 43708 1372
rect 52640 1344 52752 1372
rect 1372 1260 5964 1316
rect 6020 1260 6030 1316
rect 9538 1260 9548 1316
rect 9604 1260 17164 1316
rect 17220 1260 17230 1316
rect 18172 1260 26236 1316
rect 26292 1260 26302 1316
rect 26450 1260 26460 1316
rect 26516 1260 28700 1316
rect 28756 1260 28766 1316
rect 30258 1260 30268 1316
rect 30324 1260 31836 1316
rect 31892 1260 31902 1316
rect 34188 1260 42252 1316
rect 42308 1260 42318 1316
rect 43652 1260 49084 1316
rect 49140 1260 49150 1316
rect 18172 1204 18228 1260
rect 34188 1204 34244 1260
rect 914 1148 924 1204
rect 980 1148 10220 1204
rect 10276 1148 10286 1204
rect 10434 1148 10444 1204
rect 10500 1148 16100 1204
rect 16258 1148 16268 1204
rect 16324 1148 18228 1204
rect 18386 1148 18396 1204
rect 18452 1148 20636 1204
rect 20692 1148 20702 1204
rect 21298 1148 21308 1204
rect 21364 1148 30380 1204
rect 30436 1148 30446 1204
rect 31266 1148 31276 1204
rect 31332 1148 34244 1204
rect 34402 1148 34412 1204
rect 34468 1148 48748 1204
rect 48804 1148 48814 1204
rect 16044 1092 16100 1148
rect 6402 1036 6412 1092
rect 6468 1036 15820 1092
rect 15876 1036 15886 1092
rect 16044 1036 19740 1092
rect 19796 1036 19806 1092
rect 20972 1036 28588 1092
rect 28644 1036 28654 1092
rect 28802 1036 28812 1092
rect 28868 1036 47180 1092
rect 47236 1036 47246 1092
rect 0 980 112 1008
rect 20972 980 21028 1036
rect 52640 980 52752 1008
rect 0 924 2940 980
rect 2996 924 3006 980
rect 5394 924 5404 980
rect 5460 924 10444 980
rect 10500 924 10510 980
rect 11778 924 11788 980
rect 11844 924 21028 980
rect 21186 924 21196 980
rect 21252 924 21980 980
rect 22036 924 22046 980
rect 22194 924 22204 980
rect 22260 924 30044 980
rect 30100 924 30110 980
rect 30258 924 30268 980
rect 30324 924 32228 980
rect 33618 924 33628 980
rect 33684 924 41020 980
rect 41076 924 41086 980
rect 48178 924 48188 980
rect 48244 924 52752 980
rect 0 896 112 924
rect 6850 812 6860 868
rect 6916 812 21756 868
rect 21812 812 21822 868
rect 22418 812 22428 868
rect 22484 812 24332 868
rect 24388 812 24398 868
rect 24882 812 24892 868
rect 24948 812 26460 868
rect 26516 812 26526 868
rect 27010 812 27020 868
rect 27076 812 31948 868
rect 32004 812 32014 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 32172 756 32228 924
rect 52640 896 52752 924
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 9874 700 9884 756
rect 9940 700 15372 756
rect 15428 700 15438 756
rect 15586 700 15596 756
rect 15652 700 16772 756
rect 16930 700 16940 756
rect 16996 700 19852 756
rect 19908 700 19918 756
rect 20066 700 20076 756
rect 20132 700 22092 756
rect 22148 700 22158 756
rect 22316 700 24220 756
rect 24276 700 24286 756
rect 25218 700 25228 756
rect 25284 700 31948 756
rect 32172 700 36876 756
rect 36932 700 36942 756
rect 16716 644 16772 700
rect 22316 644 22372 700
rect 31892 644 31948 700
rect 5282 588 5292 644
rect 5348 588 11788 644
rect 11844 588 11854 644
rect 13570 588 13580 644
rect 13636 588 16492 644
rect 16548 588 16558 644
rect 16716 588 22372 644
rect 22530 588 22540 644
rect 22596 588 23100 644
rect 23156 588 23166 644
rect 23314 588 23324 644
rect 23380 588 28812 644
rect 28868 588 28878 644
rect 31892 588 34804 644
rect 35522 588 35532 644
rect 35588 588 50764 644
rect 50820 588 50830 644
rect 0 532 112 560
rect 0 476 1484 532
rect 1540 476 1550 532
rect 7522 476 7532 532
rect 7588 476 15596 532
rect 15652 476 15662 532
rect 15810 476 15820 532
rect 15876 476 19628 532
rect 19684 476 19694 532
rect 19842 476 19852 532
rect 19908 476 20860 532
rect 20916 476 20926 532
rect 21186 476 21196 532
rect 21252 476 23660 532
rect 23716 476 23726 532
rect 24098 476 24108 532
rect 24164 476 34524 532
rect 34580 476 34590 532
rect 0 448 112 476
rect 34748 420 34804 588
rect 52640 532 52752 560
rect 50530 476 50540 532
rect 50596 476 52752 532
rect 52640 448 52752 476
rect 15250 364 15260 420
rect 15316 364 30268 420
rect 30324 364 30334 420
rect 34748 364 44828 420
rect 44884 364 44894 420
rect 5730 252 5740 308
rect 5796 252 23772 308
rect 23828 252 23838 308
rect 24210 252 24220 308
rect 24276 252 26124 308
rect 26180 252 26190 308
rect 29362 252 29372 308
rect 29428 252 45948 308
rect 46004 252 46014 308
rect 47740 252 50876 308
rect 50932 252 50942 308
rect 47740 196 47796 252
rect 12114 140 12124 196
rect 12180 140 21196 196
rect 21252 140 21262 196
rect 21522 140 21532 196
rect 21588 140 26796 196
rect 26852 140 26862 196
rect 29922 140 29932 196
rect 29988 140 33628 196
rect 33684 140 33694 196
rect 36754 140 36764 196
rect 36820 140 47796 196
rect 48402 140 48412 196
rect 48468 140 48478 196
rect 0 84 112 112
rect 48412 84 48468 140
rect 52640 84 52752 112
rect 0 28 2828 84
rect 2884 28 2894 84
rect 13234 28 13244 84
rect 13300 28 23548 84
rect 23604 28 23614 84
rect 24434 28 24444 84
rect 24500 28 30492 84
rect 30548 28 30558 84
rect 39778 28 39788 84
rect 39844 28 48468 84
rect 51538 28 51548 84
rect 51604 28 52752 84
rect 0 0 112 28
rect 52640 0 52752 28
<< via3 >>
rect 14476 14140 14532 14196
rect 16716 14140 16772 14196
rect 31164 14140 31220 14196
rect 31388 14140 31444 14196
rect 35196 14140 35252 14196
rect 39116 14140 39172 14196
rect 13916 14028 13972 14084
rect 16268 14028 16324 14084
rect 25116 14028 25172 14084
rect 25340 14028 25396 14084
rect 33068 14028 33124 14084
rect 37884 14028 37940 14084
rect 22764 13916 22820 13972
rect 26012 13916 26068 13972
rect 31388 13916 31444 13972
rect 14476 13804 14532 13860
rect 15484 13804 15540 13860
rect 26124 13804 26180 13860
rect 38220 13804 38276 13860
rect 39116 13804 39172 13860
rect 15148 13692 15204 13748
rect 26348 13692 26404 13748
rect 20972 13580 21028 13636
rect 25564 13580 25620 13636
rect 31836 13580 31892 13636
rect 25228 13468 25284 13524
rect 35196 13468 35252 13524
rect 15484 13356 15540 13412
rect 16716 13356 16772 13412
rect 18508 13356 18564 13412
rect 24892 13356 24948 13412
rect 30156 13356 30212 13412
rect 31164 13356 31220 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 25116 13132 25172 13188
rect 27244 13132 27300 13188
rect 33068 13132 33124 13188
rect 26460 13020 26516 13076
rect 32620 13020 32676 13076
rect 17948 12908 18004 12964
rect 15148 12796 15204 12852
rect 15036 12684 15092 12740
rect 31836 12908 31892 12964
rect 26348 12684 26404 12740
rect 27020 12684 27076 12740
rect 27468 12684 27524 12740
rect 32620 12684 32676 12740
rect 24220 12572 24276 12628
rect 25004 12572 25060 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 20748 12460 20804 12516
rect 23548 12460 23604 12516
rect 25228 12460 25284 12516
rect 18060 12348 18116 12404
rect 28476 12348 28532 12404
rect 13692 12236 13748 12292
rect 15260 12236 15316 12292
rect 17836 12236 17892 12292
rect 26796 12236 26852 12292
rect 31724 12236 31780 12292
rect 15708 12124 15764 12180
rect 24892 12124 24948 12180
rect 25116 12124 25172 12180
rect 12236 12012 12292 12068
rect 15820 12012 15876 12068
rect 17724 11900 17780 11956
rect 17948 11900 18004 11956
rect 25228 11900 25284 11956
rect 25452 11900 25508 11956
rect 26684 11900 26740 11956
rect 26908 11900 26964 11956
rect 28476 11900 28532 11956
rect 32396 11900 32452 11956
rect 15036 11788 15092 11844
rect 15260 11788 15316 11844
rect 22764 11788 22820 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 33404 11676 33460 11732
rect 36988 11676 37044 11732
rect 14924 11564 14980 11620
rect 22540 11564 22596 11620
rect 23548 11564 23604 11620
rect 24220 11564 24276 11620
rect 28028 11564 28084 11620
rect 32172 11564 32228 11620
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 25452 11452 25508 11508
rect 28476 11452 28532 11508
rect 13692 11340 13748 11396
rect 21532 11340 21588 11396
rect 25228 11340 25284 11396
rect 29820 11340 29876 11396
rect 30156 11340 30212 11396
rect 30716 11340 30772 11396
rect 40348 11340 40404 11396
rect 15260 11228 15316 11284
rect 20860 11228 20916 11284
rect 33740 11228 33796 11284
rect 25452 11116 25508 11172
rect 21532 11004 21588 11060
rect 24220 11004 24276 11060
rect 25116 11004 25172 11060
rect 31724 11004 31780 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 20860 10892 20916 10948
rect 26236 10892 26292 10948
rect 27244 10892 27300 10948
rect 40460 10892 40516 10948
rect 26460 10780 26516 10836
rect 36988 10780 37044 10836
rect 16492 10668 16548 10724
rect 25004 10668 25060 10724
rect 28812 10668 28868 10724
rect 26684 10556 26740 10612
rect 27020 10556 27076 10612
rect 36652 10556 36708 10612
rect 29596 10444 29652 10500
rect 29932 10444 29988 10500
rect 26572 10332 26628 10388
rect 27132 10332 27188 10388
rect 28812 10332 28868 10388
rect 32844 10332 32900 10388
rect 35308 10220 35364 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 16492 10108 16548 10164
rect 23100 10108 23156 10164
rect 24220 10108 24276 10164
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 16828 9996 16884 10052
rect 25452 9996 25508 10052
rect 20524 9884 20580 9940
rect 22092 9884 22148 9940
rect 22652 9884 22708 9940
rect 23324 9884 23380 9940
rect 24892 9884 24948 9940
rect 26852 9884 26908 9940
rect 27244 9884 27300 9940
rect 16828 9772 16884 9828
rect 24220 9772 24276 9828
rect 18508 9660 18564 9716
rect 31500 9660 31556 9716
rect 16492 9548 16548 9604
rect 16716 9548 16772 9604
rect 25452 9548 25508 9604
rect 26684 9548 26740 9604
rect 28028 9548 28084 9604
rect 28812 9548 28868 9604
rect 32172 9548 32228 9604
rect 32396 9548 32452 9604
rect 38668 9548 38724 9604
rect 40348 9548 40404 9604
rect 15932 9436 15988 9492
rect 26460 9436 26516 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 19516 9324 19572 9380
rect 19964 9324 20020 9380
rect 25116 9324 25172 9380
rect 29708 9324 29764 9380
rect 31500 9324 31556 9380
rect 31724 9324 31780 9380
rect 35196 9324 35252 9380
rect 17276 9212 17332 9268
rect 21532 8988 21588 9044
rect 26012 8988 26068 9044
rect 26460 8988 26516 9044
rect 33180 8988 33236 9044
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 17724 8876 17780 8932
rect 21980 8876 22036 8932
rect 13356 8764 13412 8820
rect 16044 8764 16100 8820
rect 20524 8764 20580 8820
rect 26124 8764 26180 8820
rect 27580 8764 27636 8820
rect 30268 8764 30324 8820
rect 31724 8764 31780 8820
rect 15596 8652 15652 8708
rect 17612 8652 17668 8708
rect 26460 8652 26516 8708
rect 27916 8652 27972 8708
rect 40236 8652 40292 8708
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 16604 8540 16660 8596
rect 21868 8540 21924 8596
rect 26348 8540 26404 8596
rect 26908 8540 26964 8596
rect 28028 8540 28084 8596
rect 33852 8540 33908 8596
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 35980 8540 36036 8596
rect 15036 8428 15092 8484
rect 15708 8428 15764 8484
rect 15148 8316 15204 8372
rect 16380 8316 16436 8372
rect 19964 8316 20020 8372
rect 26348 8316 26404 8372
rect 28812 8316 28868 8372
rect 29596 8316 29652 8372
rect 32732 8316 32788 8372
rect 40348 8316 40404 8372
rect 12124 8204 12180 8260
rect 16716 8204 16772 8260
rect 18844 8204 18900 8260
rect 25452 8204 25508 8260
rect 29708 8204 29764 8260
rect 37436 8204 37492 8260
rect 13804 8092 13860 8148
rect 15372 8092 15428 8148
rect 25564 8092 25620 8148
rect 14924 7980 14980 8036
rect 15260 7980 15316 8036
rect 19852 7980 19908 8036
rect 21644 7980 21700 8036
rect 21868 7980 21924 8036
rect 27020 7980 27076 8036
rect 30380 7980 30436 8036
rect 30716 7980 30772 8036
rect 16044 7868 16100 7924
rect 16828 7868 16884 7924
rect 25452 7868 25508 7924
rect 25676 7868 25732 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 13804 7756 13860 7812
rect 19180 7756 19236 7812
rect 19852 7756 19908 7812
rect 20076 7756 20132 7812
rect 24220 7756 24276 7812
rect 26684 7644 26740 7700
rect 38556 7644 38612 7700
rect 29260 7532 29316 7588
rect 16828 7420 16884 7476
rect 29820 7420 29876 7476
rect 31836 7420 31892 7476
rect 37436 7420 37492 7476
rect 25340 7196 25396 7252
rect 29932 7196 29988 7252
rect 33180 7196 33236 7252
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 21196 6972 21252 7028
rect 25228 6972 25284 7028
rect 27356 6860 27412 6916
rect 29596 6860 29652 6916
rect 16940 6748 16996 6804
rect 18060 6748 18116 6804
rect 21196 6748 21252 6804
rect 32844 6748 32900 6804
rect 33852 6636 33908 6692
rect 27132 6524 27188 6580
rect 29596 6524 29652 6580
rect 25676 6412 25732 6468
rect 26012 6412 26068 6468
rect 15036 6300 15092 6356
rect 15820 6300 15876 6356
rect 21196 6300 21252 6356
rect 22540 6300 22596 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 16268 6188 16324 6244
rect 16492 6188 16548 6244
rect 26684 6188 26740 6244
rect 12236 6076 12292 6132
rect 19404 6076 19460 6132
rect 20076 6076 20132 6132
rect 29820 6076 29876 6132
rect 27468 5964 27524 6020
rect 38220 5964 38276 6020
rect 16492 5740 16548 5796
rect 30156 5740 30212 5796
rect 24220 5628 24276 5684
rect 27020 5628 27076 5684
rect 15036 5516 15092 5572
rect 18844 5516 18900 5572
rect 38220 5516 38276 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 17836 5404 17892 5460
rect 26012 5404 26068 5460
rect 26348 5404 26404 5460
rect 29260 5404 29316 5460
rect 31948 5404 32004 5460
rect 21308 5292 21364 5348
rect 26124 5292 26180 5348
rect 13916 5180 13972 5236
rect 15484 5180 15540 5236
rect 16380 5180 16436 5236
rect 16268 5068 16324 5124
rect 16940 5068 16996 5124
rect 25116 5068 25172 5124
rect 29932 5068 29988 5124
rect 16492 4956 16548 5012
rect 17052 4956 17108 5012
rect 35532 4956 35588 5012
rect 19068 4844 19124 4900
rect 29820 4844 29876 4900
rect 40236 4844 40292 4900
rect 15932 4732 15988 4788
rect 24220 4732 24276 4788
rect 25564 4732 25620 4788
rect 35532 4732 35588 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 22092 4620 22148 4676
rect 25004 4620 25060 4676
rect 16156 4508 16212 4564
rect 18172 4508 18228 4564
rect 30156 4396 30212 4452
rect 19628 4284 19684 4340
rect 27020 4284 27076 4340
rect 20076 4060 20132 4116
rect 21532 4060 21588 4116
rect 27020 4060 27076 4116
rect 30044 4060 30100 4116
rect 20636 3948 20692 4004
rect 20972 3948 21028 4004
rect 22092 3948 22148 4004
rect 22652 3948 22708 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 24220 3836 24276 3892
rect 25004 3836 25060 3892
rect 16940 3724 16996 3780
rect 31948 3724 32004 3780
rect 13692 3612 13748 3668
rect 21084 3612 21140 3668
rect 18844 3500 18900 3556
rect 19964 3500 20020 3556
rect 12572 3388 12628 3444
rect 20636 3388 20692 3444
rect 22092 3388 22148 3444
rect 18508 3276 18564 3332
rect 18844 3276 18900 3332
rect 19964 3276 20020 3332
rect 21980 3276 22036 3332
rect 27804 3276 27860 3332
rect 22428 3164 22484 3220
rect 23324 3164 23380 3220
rect 26348 3164 26404 3220
rect 35980 3164 36036 3220
rect 36652 3164 36708 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 21196 3052 21252 3108
rect 27916 3052 27972 3108
rect 30380 3052 30436 3108
rect 11564 2940 11620 2996
rect 18284 2940 18340 2996
rect 15484 2716 15540 2772
rect 22316 2716 22372 2772
rect 25340 2716 25396 2772
rect 32732 2716 32788 2772
rect 14140 2604 14196 2660
rect 18284 2604 18340 2660
rect 15932 2380 15988 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 16828 2268 16884 2324
rect 21196 2268 21252 2324
rect 21644 2268 21700 2324
rect 22204 2268 22260 2324
rect 12572 2156 12628 2212
rect 18396 2156 18452 2212
rect 21980 2156 22036 2212
rect 14140 2044 14196 2100
rect 14924 2044 14980 2100
rect 19964 2044 20020 2100
rect 22204 2044 22260 2100
rect 15484 1932 15540 1988
rect 21420 1820 21476 1876
rect 22092 1820 22148 1876
rect 16940 1708 16996 1764
rect 18844 1708 18900 1764
rect 21980 1708 22036 1764
rect 28476 1708 28532 1764
rect 34412 1708 34468 1764
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 24220 1596 24276 1652
rect 31948 1596 32004 1652
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 19404 1484 19460 1540
rect 21756 1484 21812 1540
rect 11788 1372 11844 1428
rect 17276 1372 17332 1428
rect 18844 1372 18900 1428
rect 20860 1372 20916 1428
rect 28476 1372 28532 1428
rect 26460 1260 26516 1316
rect 30268 1260 30324 1316
rect 31836 1260 31892 1316
rect 18396 1148 18452 1204
rect 34412 1148 34468 1204
rect 28812 1036 28868 1092
rect 22204 924 22260 980
rect 30044 924 30100 980
rect 26460 812 26516 868
rect 31948 812 32004 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 15372 700 15428 756
rect 16940 700 16996 756
rect 22092 700 22148 756
rect 28812 588 28868 644
rect 15596 476 15652 532
rect 21196 476 21252 532
rect 12124 140 12180 196
rect 21196 140 21252 196
rect 21532 140 21588 196
rect 29932 140 29988 196
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14224
rect 14476 14196 14532 14206
rect 16716 14196 16772 14206
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 13916 14084 13972 14094
rect 13692 12292 13748 12302
rect 13692 12178 13748 12236
rect 13356 12122 13748 12178
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 12236 12068 12292 12078
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 12124 8260 12180 8270
rect 11564 2998 11620 3006
rect 11564 2996 11844 2998
rect 11620 2942 11844 2996
rect 11564 2930 11620 2940
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 11788 1428 11844 2942
rect 11788 1362 11844 1372
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 12124 196 12180 8204
rect 12236 6132 12292 12012
rect 13356 8820 13412 12122
rect 13356 8754 13412 8764
rect 13692 11396 13748 11406
rect 12236 6066 12292 6076
rect 13692 3668 13748 11340
rect 13804 8148 13860 8158
rect 13804 7812 13860 8092
rect 13804 7746 13860 7756
rect 13916 5236 13972 14028
rect 14476 13860 14532 14140
rect 16268 14140 16716 14158
rect 16268 14102 16772 14140
rect 16268 14084 16324 14102
rect 16268 14018 16324 14028
rect 22764 13972 22820 13982
rect 14476 13794 14532 13804
rect 15484 13860 15540 13870
rect 15148 13748 15204 13758
rect 15148 12852 15204 13692
rect 15484 13412 15540 13804
rect 20972 13636 21028 13646
rect 15484 13346 15540 13356
rect 16716 13412 16772 13422
rect 15148 12786 15204 12796
rect 15036 12740 15092 12750
rect 15036 11998 15092 12684
rect 15260 12292 15316 12302
rect 15260 12178 15316 12236
rect 15708 12180 15764 12190
rect 15260 12124 15708 12178
rect 15260 12122 15764 12124
rect 15708 12114 15764 12122
rect 15820 12068 15876 12078
rect 15820 11998 15876 12012
rect 14924 11942 15092 11998
rect 15148 11942 15876 11998
rect 14924 11620 14980 11942
rect 15036 11844 15092 11854
rect 15148 11818 15204 11942
rect 15092 11788 15204 11818
rect 15036 11762 15204 11788
rect 15260 11844 15316 11854
rect 14924 11554 14980 11564
rect 15260 11284 15316 11788
rect 15260 11218 15316 11228
rect 16492 10724 16548 10734
rect 16492 10164 16548 10668
rect 16492 10098 16548 10108
rect 16492 9604 16548 9614
rect 15932 9492 15988 9502
rect 15932 9118 15988 9436
rect 16492 9298 16548 9548
rect 16716 9604 16772 13356
rect 18508 13412 18564 13422
rect 17948 12964 18004 12974
rect 17836 12292 17892 12302
rect 17724 11956 17780 11966
rect 16828 10052 16884 10062
rect 16828 9828 16884 9996
rect 16828 9762 16884 9772
rect 16716 9538 16772 9548
rect 16492 9268 17332 9298
rect 16492 9242 17276 9268
rect 17276 9202 17332 9212
rect 15932 9062 16772 9118
rect 16044 8820 16100 8830
rect 15596 8708 15876 8758
rect 15652 8702 15876 8708
rect 15596 8642 15652 8652
rect 15036 8484 15092 8494
rect 13916 5170 13972 5180
rect 14924 8036 14980 8046
rect 13692 3602 13748 3612
rect 12572 3444 12628 3454
rect 12572 2212 12628 3388
rect 12572 2146 12628 2156
rect 14140 2660 14196 2670
rect 14140 2100 14196 2604
rect 14140 2034 14196 2044
rect 14924 2100 14980 7980
rect 15036 6356 15092 8428
rect 15708 8484 15764 8494
rect 15148 8372 15204 8382
rect 15148 8218 15204 8316
rect 15708 8218 15764 8428
rect 15148 8162 15316 8218
rect 15260 8036 15316 8162
rect 15372 8162 15764 8218
rect 15372 8148 15428 8162
rect 15372 8082 15428 8092
rect 15260 7970 15316 7980
rect 15036 6290 15092 6300
rect 15820 6356 15876 8702
rect 16044 7924 16100 8764
rect 16604 8596 16660 8606
rect 16604 8398 16660 8540
rect 16380 8372 16660 8398
rect 16436 8342 16660 8372
rect 16380 8306 16436 8316
rect 16716 8260 16772 9062
rect 17724 8932 17780 11900
rect 17724 8866 17780 8876
rect 16716 8194 16772 8204
rect 17612 8708 17668 8718
rect 16044 7858 16100 7868
rect 16828 7924 16884 7934
rect 16828 7476 16884 7868
rect 16828 7410 16884 7420
rect 16940 6804 16996 6814
rect 16940 6418 16996 6748
rect 15820 6290 15876 6300
rect 16268 6362 16996 6418
rect 16268 6244 16324 6362
rect 16268 6178 16324 6188
rect 16492 6244 16548 6254
rect 16492 5796 16548 6188
rect 16492 5730 16548 5740
rect 15036 5572 15092 5582
rect 15036 5158 15092 5516
rect 16268 5462 16548 5518
rect 15484 5236 15540 5246
rect 15484 5158 15540 5180
rect 15036 5102 15540 5158
rect 16268 5124 16324 5462
rect 16492 5338 16548 5462
rect 16492 5282 17108 5338
rect 16268 5058 16324 5068
rect 16380 5236 16436 5246
rect 15932 4788 15988 4798
rect 15932 4618 15988 4732
rect 16380 4618 16436 5180
rect 16492 5124 16996 5158
rect 16492 5102 16940 5124
rect 16492 5012 16548 5102
rect 16940 5058 16996 5068
rect 16492 4946 16548 4956
rect 17052 5012 17108 5282
rect 17052 4946 17108 4956
rect 15932 4564 16212 4618
rect 15932 4562 16156 4564
rect 16380 4562 16772 4618
rect 16156 4498 16212 4508
rect 16716 3178 16772 4562
rect 17612 3898 17668 8652
rect 17836 5460 17892 12236
rect 17948 11956 18004 12908
rect 17948 11890 18004 11900
rect 18060 12404 18116 12414
rect 18060 6804 18116 12348
rect 18508 9716 18564 13356
rect 20748 12516 20804 12526
rect 18508 9650 18564 9660
rect 20524 9940 20580 9950
rect 19516 9380 19572 9390
rect 18060 6738 18116 6748
rect 18844 8260 18900 8270
rect 18844 5572 18900 8204
rect 18844 5506 18900 5516
rect 19180 7812 19236 7822
rect 17836 5394 17892 5404
rect 19068 4900 19124 4910
rect 19068 4798 19124 4844
rect 18172 4742 19124 4798
rect 18172 4564 18228 4742
rect 19180 4618 19236 7756
rect 18172 4498 18228 4508
rect 18508 4562 19236 4618
rect 19404 6132 19460 6142
rect 16940 3842 17668 3898
rect 16940 3780 16996 3842
rect 16940 3714 16996 3724
rect 18508 3332 18564 4562
rect 18508 3266 18564 3276
rect 18844 3556 18900 3566
rect 18844 3332 18900 3500
rect 18844 3266 18900 3276
rect 16716 3122 16884 3178
rect 14924 2034 14980 2044
rect 15484 2772 15540 2782
rect 15484 1988 15540 2716
rect 15484 1922 15540 1932
rect 15932 2436 15988 2446
rect 15932 1918 15988 2380
rect 16828 2324 16884 3122
rect 18284 2996 18340 3006
rect 18284 2660 18340 2940
rect 18284 2594 18340 2604
rect 16828 2258 16884 2268
rect 18396 2212 18452 2222
rect 15932 1862 16996 1918
rect 16940 1764 16996 1862
rect 16940 1698 16996 1708
rect 17276 1428 17332 1438
rect 15372 782 16996 838
rect 15372 756 15428 782
rect 15372 690 15428 700
rect 16940 756 16996 782
rect 16940 690 16996 700
rect 15596 532 15652 542
rect 17276 478 17332 1372
rect 18396 1204 18452 2156
rect 18844 1764 18900 1774
rect 18844 1428 18900 1708
rect 19404 1540 19460 6076
rect 19516 4078 19572 9324
rect 19964 9380 20020 9390
rect 19964 8372 20020 9324
rect 20524 8820 20580 9884
rect 20524 8754 20580 8764
rect 19964 8306 20020 8316
rect 19852 8036 19908 8046
rect 19852 7812 19908 7980
rect 19852 7746 19908 7756
rect 20076 7812 20132 7822
rect 20076 6132 20132 7756
rect 20076 6066 20132 6076
rect 19628 4340 19684 4350
rect 19628 4258 19684 4284
rect 19628 4202 20132 4258
rect 20076 4116 20132 4202
rect 19516 4022 19796 4078
rect 20076 4050 20132 4060
rect 19404 1474 19460 1484
rect 18844 1362 18900 1372
rect 18396 1138 18452 1148
rect 19740 658 19796 4022
rect 20636 4004 20692 4014
rect 19964 3556 20020 3566
rect 19964 3332 20020 3500
rect 20636 3444 20692 3948
rect 20748 3538 20804 12460
rect 20860 11284 20916 11294
rect 20860 10948 20916 11228
rect 20860 10882 20916 10892
rect 20972 4004 21028 13580
rect 22764 11844 22820 13916
rect 23776 12572 24096 14224
rect 24436 13356 24756 14224
rect 31164 14196 31220 14206
rect 25116 14084 25172 14094
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 22764 11778 22820 11788
rect 23548 12516 23604 12526
rect 22540 11620 22596 11630
rect 21532 11396 21588 11406
rect 21532 11060 21588 11340
rect 21532 10994 21588 11004
rect 22092 9940 22148 9950
rect 21532 9044 21588 9054
rect 21532 8938 21588 8988
rect 21980 8938 22036 8942
rect 21532 8932 22036 8938
rect 21532 8882 21980 8932
rect 21980 8866 22036 8876
rect 21868 8596 21924 8606
rect 21644 8036 21700 8046
rect 21644 7858 21700 7980
rect 21868 8036 21924 8540
rect 21868 7970 21924 7980
rect 22092 7858 22148 9884
rect 22540 9658 22596 11564
rect 23548 11620 23604 12460
rect 23548 11554 23604 11564
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 24220 12628 24276 12638
rect 24220 11620 24276 12572
rect 24220 11554 24276 11564
rect 24436 11788 24756 13300
rect 24892 13412 24948 13422
rect 24892 12180 24948 13356
rect 25116 13188 25172 14028
rect 25340 14084 25396 14094
rect 25340 13978 25396 14028
rect 26012 13978 26068 13982
rect 25340 13972 26068 13978
rect 25340 13922 26012 13972
rect 26012 13906 26068 13916
rect 26124 13860 26180 13870
rect 26124 13798 26180 13804
rect 25564 13742 26180 13798
rect 26348 13748 26404 13758
rect 25564 13636 25620 13742
rect 25564 13570 25620 13580
rect 25116 13122 25172 13132
rect 25228 13524 25284 13534
rect 25004 12628 25060 12638
rect 25004 12358 25060 12572
rect 25228 12516 25284 13468
rect 26348 12740 26404 13692
rect 30156 13412 30212 13422
rect 27244 13188 27300 13198
rect 26460 13076 26516 13086
rect 26460 12898 26516 13020
rect 26460 12842 27076 12898
rect 26348 12674 26404 12684
rect 27020 12740 27076 12842
rect 27020 12674 27076 12684
rect 25228 12450 25284 12460
rect 25004 12302 26852 12358
rect 26796 12292 26852 12302
rect 26796 12226 26852 12236
rect 24892 12114 24948 12124
rect 25116 12180 25172 12190
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23100 10164 23156 10174
rect 23100 10018 23156 10108
rect 22652 9962 23156 10018
rect 22652 9940 22708 9962
rect 22652 9874 22708 9884
rect 23324 9940 23380 9950
rect 22540 9602 22708 9658
rect 21644 7802 22148 7858
rect 21196 7028 21252 7038
rect 21196 6804 21252 6972
rect 21196 6738 21252 6748
rect 21196 6362 22596 6418
rect 21196 6356 21252 6362
rect 21196 6290 21252 6300
rect 22540 6356 22596 6362
rect 22540 6290 22596 6300
rect 21308 5348 21364 5358
rect 21308 4798 21364 5292
rect 21308 4742 22148 4798
rect 22092 4676 22148 4742
rect 22092 4610 22148 4620
rect 20972 3938 21028 3948
rect 21532 4116 21588 4126
rect 21532 3718 21588 4060
rect 21084 3668 21588 3718
rect 21140 3662 21588 3668
rect 22092 4004 22148 4014
rect 21084 3602 21140 3612
rect 20748 3482 21700 3538
rect 20636 3378 20692 3388
rect 19964 3266 20020 3276
rect 21196 3108 21252 3118
rect 21196 2324 21252 3052
rect 21196 2258 21252 2268
rect 21644 2324 21700 3482
rect 22092 3444 22148 3948
rect 22652 4004 22708 9602
rect 22652 3938 22708 3948
rect 22092 3378 22148 3388
rect 21980 3332 22036 3342
rect 21980 2458 22036 3276
rect 22428 3220 22484 3230
rect 22428 2818 22484 3164
rect 23324 3220 23380 9884
rect 23324 3154 23380 3164
rect 23776 9436 24096 10948
rect 24220 11060 24276 11070
rect 24220 10164 24276 11004
rect 24220 10098 24276 10108
rect 24436 10220 24756 11732
rect 25116 11458 25172 12124
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23776 6300 24096 7812
rect 24220 9828 24276 9838
rect 24220 7812 24276 9772
rect 24220 7746 24276 7756
rect 24436 8652 24756 10164
rect 24892 11402 25172 11458
rect 25228 11956 25284 11966
rect 24892 9940 24948 11402
rect 25228 11396 25284 11900
rect 25452 11956 25508 11966
rect 25452 11638 25508 11900
rect 25228 11330 25284 11340
rect 25340 11582 25508 11638
rect 26684 11956 26740 11966
rect 25340 11098 25396 11582
rect 25452 11508 25508 11518
rect 25452 11172 25508 11452
rect 25452 11106 25508 11116
rect 25116 11060 25396 11098
rect 25172 11042 25396 11060
rect 25116 10994 25172 11004
rect 26236 10948 26292 10958
rect 25004 10892 26236 10918
rect 25004 10862 26292 10892
rect 26684 10918 26740 11900
rect 26908 11956 26964 11966
rect 26908 10918 26964 11900
rect 26684 10862 26964 10918
rect 27244 10948 27300 13132
rect 27244 10882 27300 10892
rect 27468 12740 27524 12750
rect 25004 10724 25060 10862
rect 26460 10836 26516 10846
rect 26460 10738 26516 10780
rect 26460 10682 27300 10738
rect 25004 10658 25060 10668
rect 26684 10612 26740 10622
rect 26572 10388 26628 10398
rect 26460 10332 26572 10378
rect 26460 10322 26628 10332
rect 24892 9874 24948 9884
rect 25452 10052 25508 10062
rect 25452 9604 25508 9996
rect 25452 9538 25508 9548
rect 26460 9492 26516 10322
rect 26684 9604 26740 10556
rect 27020 10612 27076 10622
rect 27020 10018 27076 10556
rect 26852 9962 27076 10018
rect 27132 10388 27188 10398
rect 26852 9940 26908 9962
rect 26852 9874 26908 9884
rect 26684 9538 26740 9548
rect 26460 9426 26516 9436
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 24436 7084 24756 8596
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 24220 5684 24276 5694
rect 24220 4788 24276 5628
rect 24220 4722 24276 4732
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 23776 3164 24096 4676
rect 24436 3948 24756 5460
rect 25116 9380 25172 9390
rect 25116 5124 25172 9324
rect 27132 9298 27188 10332
rect 27244 9940 27300 10682
rect 27244 9874 27300 9884
rect 26012 9242 27188 9298
rect 26012 9044 26068 9242
rect 26012 8978 26068 8988
rect 26460 9044 26516 9054
rect 26124 8820 26180 8830
rect 25452 8260 25508 8270
rect 25228 8204 25452 8218
rect 25228 8162 25508 8204
rect 26124 8218 26180 8764
rect 26460 8708 26516 8988
rect 26460 8642 26516 8652
rect 26348 8596 26404 8606
rect 26348 8372 26404 8540
rect 26348 8306 26404 8316
rect 26908 8596 26964 8606
rect 26908 8218 26964 8540
rect 26124 8162 26964 8218
rect 25228 7028 25284 8162
rect 25564 8148 25620 8158
rect 25564 8038 25620 8092
rect 25452 7982 25620 8038
rect 27020 8036 27076 8046
rect 25452 7924 25508 7982
rect 25452 7858 25508 7868
rect 25676 7924 25732 7934
rect 25228 6962 25284 6972
rect 25340 7252 25396 7262
rect 25116 5058 25172 5068
rect 22316 2772 22484 2818
rect 22372 2762 22484 2772
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 22316 2706 22372 2716
rect 21980 2402 22148 2458
rect 21644 2258 21700 2268
rect 21980 2212 22036 2222
rect 19964 2100 20020 2110
rect 19964 1918 20020 2044
rect 19964 1876 21476 1918
rect 19964 1862 21420 1876
rect 21420 1810 21476 1820
rect 21980 1764 22036 2156
rect 22092 1876 22148 2402
rect 22204 2324 22260 2334
rect 22204 2100 22260 2268
rect 22204 2034 22260 2044
rect 22092 1810 22148 1820
rect 21980 1698 22036 1708
rect 23776 1596 24096 3108
rect 20860 1540 21812 1558
rect 20860 1502 21756 1540
rect 20860 1428 20916 1502
rect 21756 1474 21812 1484
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 24220 3892 24276 3902
rect 24220 1652 24276 3836
rect 24220 1586 24276 1596
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 25004 4676 25060 4686
rect 25004 3892 25060 4620
rect 25004 3826 25060 3836
rect 25340 2772 25396 7196
rect 25676 6468 25732 7868
rect 26684 7700 26740 7710
rect 25676 6402 25732 6412
rect 26012 6468 26068 6478
rect 26012 5460 26068 6412
rect 26684 6244 26740 7644
rect 26684 6178 26740 6188
rect 27020 5684 27076 7980
rect 27356 6916 27412 6926
rect 27356 6598 27412 6860
rect 27132 6580 27412 6598
rect 27188 6542 27412 6580
rect 27132 6514 27188 6524
rect 27468 6020 27524 12684
rect 28476 12404 28532 12414
rect 28028 12348 28476 12358
rect 28028 12302 28532 12348
rect 28028 11620 28084 12302
rect 28028 11554 28084 11564
rect 28476 11956 28532 11966
rect 28476 11508 28532 11900
rect 28476 11442 28532 11452
rect 29820 11396 29876 11406
rect 28812 10724 28868 10734
rect 28812 10388 28868 10668
rect 28812 10322 28868 10332
rect 29596 10500 29652 10510
rect 28028 9604 28084 9614
rect 27580 8820 27636 8830
rect 27580 8758 27636 8764
rect 27580 8702 27860 8758
rect 27468 5954 27524 5964
rect 27020 5618 27076 5628
rect 26012 5394 26068 5404
rect 26348 5460 26404 5470
rect 26124 5348 26180 5358
rect 26124 4798 26180 5292
rect 25564 4788 26180 4798
rect 25620 4742 26180 4788
rect 25564 4722 25620 4732
rect 26348 3220 26404 5404
rect 27020 4340 27076 4350
rect 27020 4116 27076 4284
rect 27020 4050 27076 4060
rect 27804 3332 27860 8702
rect 27804 3266 27860 3276
rect 27916 8708 27972 8718
rect 26348 3154 26404 3164
rect 27916 3108 27972 8652
rect 28028 8596 28084 9548
rect 28028 8530 28084 8540
rect 28812 9604 28868 9614
rect 28812 8372 28868 9548
rect 28812 8306 28868 8316
rect 29596 8372 29652 10444
rect 29596 8306 29652 8316
rect 29708 9380 29764 9390
rect 29708 8260 29764 9324
rect 29708 8194 29764 8204
rect 29260 7588 29316 7598
rect 29260 5460 29316 7532
rect 29820 7476 29876 11340
rect 30156 11396 30212 13356
rect 31164 13412 31220 14140
rect 31388 14196 31444 14206
rect 31388 13972 31444 14140
rect 35196 14196 35252 14206
rect 31388 13906 31444 13916
rect 33068 14084 33124 14094
rect 31164 13346 31220 13356
rect 31836 13636 31892 13646
rect 31836 12964 31892 13580
rect 33068 13188 33124 14028
rect 35196 13524 35252 14140
rect 39116 14196 39172 14206
rect 37884 14084 37940 14094
rect 37884 13978 37940 14028
rect 37884 13922 38276 13978
rect 38220 13860 38276 13922
rect 38220 13794 38276 13804
rect 39116 13860 39172 14140
rect 39116 13794 39172 13804
rect 35196 13458 35252 13468
rect 33068 13122 33124 13132
rect 31836 12898 31892 12908
rect 32620 13076 32676 13086
rect 32620 12740 32676 13020
rect 32620 12674 32676 12684
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 31724 12292 31780 12302
rect 30156 11330 30212 11340
rect 30716 11396 30772 11406
rect 29820 7410 29876 7420
rect 29932 10500 29988 10510
rect 29932 7252 29988 10444
rect 29932 7186 29988 7196
rect 30268 8820 30324 8830
rect 29596 6916 29652 6926
rect 29596 6580 29652 6860
rect 29596 6514 29652 6524
rect 29260 5394 29316 5404
rect 29820 6132 29876 6142
rect 29820 4900 29876 6076
rect 30156 5796 30212 5806
rect 29820 4834 29876 4844
rect 29932 5124 29988 5134
rect 27916 3042 27972 3052
rect 25340 2706 25396 2716
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 20860 1362 20916 1372
rect 22204 980 22260 990
rect 22204 838 22260 924
rect 22092 782 22260 838
rect 22092 756 22148 782
rect 22092 690 22148 700
rect 19740 602 21252 658
rect 15652 476 17332 478
rect 15596 422 17332 476
rect 21196 532 21252 602
rect 21196 466 21252 476
rect 12124 130 12180 140
rect 21196 242 21588 298
rect 21196 196 21252 242
rect 21196 130 21252 140
rect 21532 196 21588 242
rect 21532 130 21588 140
rect 23776 0 24096 1540
rect 24436 812 24756 2324
rect 28476 1764 28532 1774
rect 28476 1428 28532 1708
rect 28476 1362 28532 1372
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 26460 1316 26516 1326
rect 26460 868 26516 1260
rect 26460 802 26516 812
rect 28812 1092 28868 1102
rect 24436 0 24756 756
rect 28812 644 28868 1036
rect 28812 578 28868 588
rect 29932 196 29988 5068
rect 30156 4452 30212 5740
rect 30156 4386 30212 4396
rect 30268 4258 30324 8764
rect 30044 4202 30324 4258
rect 30380 8036 30436 8046
rect 30044 4116 30100 4202
rect 30044 4050 30100 4060
rect 30380 3108 30436 7980
rect 30716 8036 30772 11340
rect 31724 11060 31780 12236
rect 32396 11956 32452 11966
rect 31724 10994 31780 11004
rect 32172 11620 32228 11630
rect 31500 9716 31556 9726
rect 31500 9380 31556 9660
rect 32172 9604 32228 11564
rect 32172 9538 32228 9548
rect 32396 9604 32452 11900
rect 33404 11732 33460 11742
rect 33404 11458 33460 11676
rect 36988 11732 37044 11742
rect 33404 11402 33796 11458
rect 33740 11284 33796 11402
rect 33740 11218 33796 11228
rect 36988 10836 37044 11676
rect 36988 10770 37044 10780
rect 40348 11396 40404 11406
rect 36652 10612 36708 10622
rect 32396 9538 32452 9548
rect 32844 10388 32900 10398
rect 31500 9314 31556 9324
rect 31724 9380 31780 9390
rect 31724 8820 31780 9324
rect 31724 8754 31780 8764
rect 30716 7970 30772 7980
rect 32732 8372 32788 8382
rect 30380 3042 30436 3052
rect 31836 7476 31892 7486
rect 30268 1316 30324 1326
rect 30268 1018 30324 1260
rect 31836 1316 31892 7420
rect 31948 5460 32004 5470
rect 31948 3780 32004 5404
rect 31948 3714 32004 3724
rect 32732 2772 32788 8316
rect 32844 6804 32900 10332
rect 35308 10276 35364 10286
rect 35308 9478 35364 10220
rect 35196 9422 35364 9478
rect 35196 9380 35252 9422
rect 35196 9314 35252 9324
rect 33180 9044 33236 9054
rect 33180 7252 33236 8988
rect 33180 7186 33236 7196
rect 33852 8596 33908 8606
rect 32844 6738 32900 6748
rect 33852 6692 33908 8540
rect 33852 6626 33908 6636
rect 35980 8596 36036 8606
rect 35532 5012 35588 5022
rect 35532 4788 35588 4956
rect 35532 4722 35588 4732
rect 35980 3220 36036 8540
rect 35980 3154 36036 3164
rect 36652 3220 36708 10556
rect 38668 9604 38724 9614
rect 37436 8260 37492 8270
rect 37436 7476 37492 8204
rect 38668 7858 38724 9548
rect 40348 9604 40404 11340
rect 43776 11004 44096 12516
rect 40348 9538 40404 9548
rect 40460 10948 40516 10958
rect 40460 9478 40516 10892
rect 40348 9422 40516 9478
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 43776 9436 44096 10948
rect 38556 7802 38724 7858
rect 40236 8708 40292 8718
rect 38556 7700 38612 7802
rect 38556 7634 38612 7644
rect 37436 7410 37492 7420
rect 38220 6020 38276 6030
rect 38220 5572 38276 5964
rect 38220 5506 38276 5516
rect 40236 4900 40292 8652
rect 40348 8372 40404 9422
rect 40348 8306 40404 8316
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 40236 4834 40292 4844
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 43776 6300 44096 7812
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 36652 3154 36708 3164
rect 43776 4732 44096 6244
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 43776 3164 44096 4676
rect 32732 2706 32788 2716
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 34412 1764 34468 1774
rect 31836 1250 31892 1260
rect 31948 1652 32004 1662
rect 30044 980 30324 1018
rect 30100 962 30324 980
rect 30044 914 30100 924
rect 31948 868 32004 1596
rect 34412 1204 34468 1708
rect 34412 1138 34468 1148
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 31948 802 32004 812
rect 29932 130 29988 140
rect 43776 0 44096 1540
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44436 3948 44756 5460
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 38528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 37632 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 5712 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 5712 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 45248 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 29232 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 47600 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 36064 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 46816 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 43792 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 27776 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 47600 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 32704 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 17024 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 44576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 34384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 50624 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 30464 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 26208 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 38976 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 1456 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 10528 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 13776 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 32816 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 26320 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 38752 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 24192 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 25088 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 45696 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 24752 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 50624 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 44688 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform 1 0 46256 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 48496 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 29232 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 29232 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform 1 0 24752 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 13552 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 6048 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 8400 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 19152 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 30128 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 14000 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 3360 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 6720 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 2352 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 5712 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 25312 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 17808 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 25312 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 22960 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform -1 0 10304 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform 1 0 26544 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 29120 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform -1 0 22624 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform -1 0 21056 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform -1 0 19712 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 42448 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 47936 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 47600 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 49392 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform -1 0 19488 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform -1 0 17584 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 42112 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform -1 0 24080 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform -1 0 24528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 27104 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 27104 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 38752 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 26992 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform 1 0 49168 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform 1 0 38416 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform 1 0 46592 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 6496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 44464 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 10080 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 41664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 7504 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform -1 0 2576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 21728 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 43680 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 11536 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 15008 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 9744 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 23296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 36960 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 37856 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 15568 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 20496 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 10864 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 20944 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 4592 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 9632 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 13216 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 23520 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 9184 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 12432 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 25312 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 11200 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform 1 0 32480 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform 1 0 27216 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_182
timestamp 1486834041
transform 1 0 21056 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_198
timestamp 1486834041
transform 1 0 22848 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_202
timestamp 1486834041
transform 1 0 23296 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_444
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_454
timestamp 1486834041
transform 1 0 51520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_456
timestamp 1486834041
transform 1 0 51744 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1486834041
transform 1 0 12320 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_112
timestamp 1486834041
transform 1 0 13216 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_116
timestamp 1486834041
transform 1 0 13664 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_125
timestamp 1486834041
transform 1 0 14672 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_133
timestamp 1486834041
transform 1 0 15568 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1486834041
transform 1 0 16016 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_158
timestamp 1486834041
transform 1 0 18368 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_170
timestamp 1486834041
transform 1 0 19712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_172
timestamp 1486834041
transform 1 0 19936 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_181
timestamp 1486834041
transform 1 0 20944 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_197
timestamp 1486834041
transform 1 0 22736 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_205
timestamp 1486834041
transform 1 0 23632 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 24080 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_276
timestamp 1486834041
transform 1 0 31584 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_282
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_294
timestamp 1486834041
transform 1 0 33600 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_326
timestamp 1486834041
transform 1 0 37184 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_392
timestamp 1486834041
transform 1 0 44576 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_408
timestamp 1486834041
transform 1 0 46368 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_426
timestamp 1486834041
transform 1 0 48384 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1486834041
transform 1 0 48608 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_6
timestamp 1486834041
transform 1 0 1344 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_15
timestamp 1486834041
transform 1 0 2352 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_23
timestamp 1486834041
transform 1 0 3248 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_69
timestamp 1486834041
transform 1 0 8400 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_85
timestamp 1486834041
transform 1 0 10192 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_139
timestamp 1486834041
transform 1 0 16240 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_151
timestamp 1486834041
transform 1 0 17584 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_167
timestamp 1486834041
transform 1 0 19376 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 27664 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_247
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1486834041
transform 1 0 35504 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_321
timestamp 1486834041
transform 1 0 36624 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_323
timestamp 1486834041
transform 1 0 36848 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_332
timestamp 1486834041
transform 1 0 37856 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_348
timestamp 1486834041
transform 1 0 39648 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_380
timestamp 1486834041
transform 1 0 43232 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_384
timestamp 1486834041
transform 1 0 43680 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_395
timestamp 1486834041
transform 1 0 44912 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_397
timestamp 1486834041
transform 1 0 45136 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_406
timestamp 1486834041
transform 1 0 46144 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_410
timestamp 1486834041
transform 1 0 46592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_412
timestamp 1486834041
transform 1 0 46816 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_6
timestamp 1486834041
transform 1 0 1344 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_8
timestamp 1486834041
transform 1 0 1568 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_17
timestamp 1486834041
transform 1 0 2576 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_49
timestamp 1486834041
transform 1 0 6160 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_65
timestamp 1486834041
transform 1 0 7952 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_69
timestamp 1486834041
transform 1 0 8400 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_158
timestamp 1486834041
transform 1 0 18368 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_166
timestamp 1486834041
transform 1 0 19264 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_168
timestamp 1486834041
transform 1 0 19488 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_177
timestamp 1486834041
transform 1 0 20496 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_220
timestamp 1486834041
transform 1 0 25312 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_244
timestamp 1486834041
transform 1 0 28000 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_252
timestamp 1486834041
transform 1 0 28896 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_262
timestamp 1486834041
transform 1 0 30016 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_278
timestamp 1486834041
transform 1 0 31808 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_282
timestamp 1486834041
transform 1 0 32256 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1486834041
transform 1 0 32704 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_295
timestamp 1486834041
transform 1 0 33712 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_327
timestamp 1486834041
transform 1 0 37296 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_343
timestamp 1486834041
transform 1 0 39088 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_347
timestamp 1486834041
transform 1 0 39536 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 39760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_384
timestamp 1486834041
transform 1 0 43680 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_400
timestamp 1486834041
transform 1 0 45472 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_418
timestamp 1486834041
transform 1 0 47488 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_426
timestamp 1486834041
transform 1 0 48384 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1486834041
transform 1 0 48608 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_77
timestamp 1486834041
transform 1 0 9296 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_81
timestamp 1486834041
transform 1 0 9744 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_91
timestamp 1486834041
transform 1 0 10864 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_99
timestamp 1486834041
transform 1 0 11760 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1486834041
transform 1 0 12208 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_123
timestamp 1486834041
transform 1 0 14448 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_133
timestamp 1486834041
transform 1 0 15568 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_165
timestamp 1486834041
transform 1 0 19152 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_173
timestamp 1486834041
transform 1 0 20048 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_209
timestamp 1486834041
transform 1 0 24080 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_225
timestamp 1486834041
transform 1 0 25872 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_237
timestamp 1486834041
transform 1 0 27216 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_279
timestamp 1486834041
transform 1 0 31920 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_283
timestamp 1486834041
transform 1 0 32368 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_292
timestamp 1486834041
transform 1 0 33376 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_308
timestamp 1486834041
transform 1 0 35168 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_312
timestamp 1486834041
transform 1 0 35616 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_314
timestamp 1486834041
transform 1 0 35840 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_317
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_349
timestamp 1486834041
transform 1 0 39760 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_365
timestamp 1486834041
transform 1 0 41552 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_369
timestamp 1486834041
transform 1 0 42000 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_378
timestamp 1486834041
transform 1 0 43008 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_382
timestamp 1486834041
transform 1 0 43456 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_384
timestamp 1486834041
transform 1 0 43680 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_395
timestamp 1486834041
transform 1 0 44912 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_403
timestamp 1486834041
transform 1 0 45808 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_415
timestamp 1486834041
transform 1 0 47152 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_34
timestamp 1486834041
transform 1 0 4480 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_42
timestamp 1486834041
transform 1 0 5376 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_54
timestamp 1486834041
transform 1 0 6720 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_104
timestamp 1486834041
transform 1 0 12320 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_128
timestamp 1486834041
transform 1 0 15008 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 15904 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1486834041
transform 1 0 16800 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_153
timestamp 1486834041
transform 1 0 17808 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_185
timestamp 1486834041
transform 1 0 21392 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_193
timestamp 1486834041
transform 1 0 22288 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_202
timestamp 1486834041
transform 1 0 23296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_214
timestamp 1486834041
transform 1 0 24640 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_223
timestamp 1486834041
transform 1 0 25648 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_255
timestamp 1486834041
transform 1 0 29232 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_271
timestamp 1486834041
transform 1 0 31024 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 31920 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_314
timestamp 1486834041
transform 1 0 35840 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_330
timestamp 1486834041
transform 1 0 37632 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_338
timestamp 1486834041
transform 1 0 38528 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_348
timestamp 1486834041
transform 1 0 39648 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 47264 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_426
timestamp 1486834041
transform 1 0 48384 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1486834041
transform 1 0 48608 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_53
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_69
timestamp 1486834041
transform 1 0 8400 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_77
timestamp 1486834041
transform 1 0 9296 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_94
timestamp 1486834041
transform 1 0 11200 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_102
timestamp 1486834041
transform 1 0 12096 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_193
timestamp 1486834041
transform 1 0 22288 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_201
timestamp 1486834041
transform 1 0 23184 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_213
timestamp 1486834041
transform 1 0 24528 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_311
timestamp 1486834041
transform 1 0 35504 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_325
timestamp 1486834041
transform 1 0 37072 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_329
timestamp 1486834041
transform 1 0 37520 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_346
timestamp 1486834041
transform 1 0 39424 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_378
timestamp 1486834041
transform 1 0 43008 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_382
timestamp 1486834041
transform 1 0 43456 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 43680 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_419
timestamp 1486834041
transform 1 0 47600 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_421
timestamp 1486834041
transform 1 0 47824 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_430
timestamp 1486834041
transform 1 0 48832 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_432
timestamp 1486834041
transform 1 0 49056 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_34
timestamp 1486834041
transform 1 0 4480 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_42
timestamp 1486834041
transform 1 0 5376 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_44
timestamp 1486834041
transform 1 0 5600 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_53
timestamp 1486834041
transform 1 0 6608 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_69
timestamp 1486834041
transform 1 0 8400 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_81
timestamp 1486834041
transform 1 0 9744 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_113
timestamp 1486834041
transform 1 0 13328 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_129
timestamp 1486834041
transform 1 0 15120 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_137
timestamp 1486834041
transform 1 0 16016 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 16240 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_158
timestamp 1486834041
transform 1 0 18368 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_168
timestamp 1486834041
transform 1 0 19488 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_184
timestamp 1486834041
transform 1 0 21280 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_192
timestamp 1486834041
transform 1 0 22176 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_204
timestamp 1486834041
transform 1 0 23520 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_208
timestamp 1486834041
transform 1 0 23968 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_244
timestamp 1486834041
transform 1 0 28000 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_252
timestamp 1486834041
transform 1 0 28896 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_254
timestamp 1486834041
transform 1 0 29120 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_263
timestamp 1486834041
transform 1 0 30128 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_279
timestamp 1486834041
transform 1 0 31920 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_384
timestamp 1486834041
transform 1 0 43680 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_388
timestamp 1486834041
transform 1 0 44128 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_390
timestamp 1486834041
transform 1 0 44352 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_399
timestamp 1486834041
transform 1 0 45360 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_415
timestamp 1486834041
transform 1 0 47152 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1486834041
transform 1 0 47600 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_426
timestamp 1486834041
transform 1 0 48384 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1486834041
transform 1 0 48608 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 11984 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_135
timestamp 1486834041
transform 1 0 15792 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_151
timestamp 1486834041
transform 1 0 17584 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_165
timestamp 1486834041
transform 1 0 19152 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_173
timestamp 1486834041
transform 1 0 20048 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_193
timestamp 1486834041
transform 1 0 22288 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_209
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_263
timestamp 1486834041
transform 1 0 30128 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_295
timestamp 1486834041
transform 1 0 33712 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_311
timestamp 1486834041
transform 1 0 35504 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 8064 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_84
timestamp 1486834041
transform 1 0 10080 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_100
timestamp 1486834041
transform 1 0 11872 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_150
timestamp 1486834041
transform 1 0 17472 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_169
timestamp 1486834041
transform 1 0 19600 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_177
timestamp 1486834041
transform 1 0 20496 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_179
timestamp 1486834041
transform 1 0 20720 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_196
timestamp 1486834041
transform 1 0 22624 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_204
timestamp 1486834041
transform 1 0 23520 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_208
timestamp 1486834041
transform 1 0 23968 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_214
timestamp 1486834041
transform 1 0 24640 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_223
timestamp 1486834041
transform 1 0 25648 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_263
timestamp 1486834041
transform 1 0 30128 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 31920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_290
timestamp 1486834041
transform 1 0 33152 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_322
timestamp 1486834041
transform 1 0 36736 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_338
timestamp 1486834041
transform 1 0 38528 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 39424 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 47264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_426
timestamp 1486834041
transform 1 0 48384 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_61
timestamp 1486834041
transform 1 0 7504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_65
timestamp 1486834041
transform 1 0 7952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_67
timestamp 1486834041
transform 1 0 8176 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_76
timestamp 1486834041
transform 1 0 9184 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_84
timestamp 1486834041
transform 1 0 10080 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_88
timestamp 1486834041
transform 1 0 10528 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_90
timestamp 1486834041
transform 1 0 10752 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_199
timestamp 1486834041
transform 1 0 22960 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_207
timestamp 1486834041
transform 1 0 23856 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_209
timestamp 1486834041
transform 1 0 24080 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_226
timestamp 1486834041
transform 1 0 25984 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_242
timestamp 1486834041
transform 1 0 27776 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_244
timestamp 1486834041
transform 1 0 28000 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_333
timestamp 1486834041
transform 1 0 37968 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_345
timestamp 1486834041
transform 1 0 39312 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_363
timestamp 1486834041
transform 1 0 41328 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_379
timestamp 1486834041
transform 1 0 43120 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_383
timestamp 1486834041
transform 1 0 43568 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 8064 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_80
timestamp 1486834041
transform 1 0 9632 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_96
timestamp 1486834041
transform 1 0 11424 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1486834041
transform 1 0 16800 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 24080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_220
timestamp 1486834041
transform 1 0 25312 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_224
timestamp 1486834041
transform 1 0 25760 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_226
timestamp 1486834041
transform 1 0 25984 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_235
timestamp 1486834041
transform 1 0 26992 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_243
timestamp 1486834041
transform 1 0 27888 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_275
timestamp 1486834041
transform 1 0 31472 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_298
timestamp 1486834041
transform 1 0 34048 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_300
timestamp 1486834041
transform 1 0 34272 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_309
timestamp 1486834041
transform 1 0 35280 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_313
timestamp 1486834041
transform 1 0 35728 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_315
timestamp 1486834041
transform 1 0 35952 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_324
timestamp 1486834041
transform 1 0 36960 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_332
timestamp 1486834041
transform 1 0 37856 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_334
timestamp 1486834041
transform 1 0 38080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_349
timestamp 1486834041
transform 1 0 39760 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_374
timestamp 1486834041
transform 1 0 42560 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_382
timestamp 1486834041
transform 1 0 43456 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_384
timestamp 1486834041
transform 1 0 43680 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_401
timestamp 1486834041
transform 1 0 45584 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_417
timestamp 1486834041
transform 1 0 47376 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_426
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1486834041
transform 1 0 48608 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_15
timestamp 1486834041
transform 1 0 2352 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_31
timestamp 1486834041
transform 1 0 4144 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_69
timestamp 1486834041
transform 1 0 8400 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_115
timestamp 1486834041
transform 1 0 13552 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_181
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_211
timestamp 1486834041
transform 1 0 24304 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_227
timestamp 1486834041
transform 1 0 26096 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_244
timestamp 1486834041
transform 1 0 28000 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 35504 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_381
timestamp 1486834041
transform 1 0 43344 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_34
timestamp 1486834041
transform 1 0 4480 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_38
timestamp 1486834041
transform 1 0 4928 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_56
timestamp 1486834041
transform 1 0 6944 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_64
timestamp 1486834041
transform 1 0 7840 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_68
timestamp 1486834041
transform 1 0 8288 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_236
timestamp 1486834041
transform 1 0 27104 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_240
timestamp 1486834041
transform 1 0 27552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_250
timestamp 1486834041
transform 1 0 28672 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_266
timestamp 1486834041
transform 1 0 30464 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_274
timestamp 1486834041
transform 1 0 31360 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_278
timestamp 1486834041
transform 1 0 31808 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_314
timestamp 1486834041
transform 1 0 35840 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_318
timestamp 1486834041
transform 1 0 36288 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_347
timestamp 1486834041
transform 1 0 39536 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_349
timestamp 1486834041
transform 1 0 39760 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_380
timestamp 1486834041
transform 1 0 43232 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_412
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_426
timestamp 1486834041
transform 1 0 48384 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1486834041
transform 1 0 48608 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_10
timestamp 1486834041
transform 1 0 1792 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_14
timestamp 1486834041
transform 1 0 2240 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_24
timestamp 1486834041
transform 1 0 3360 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_32
timestamp 1486834041
transform 1 0 4256 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 4480 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_41
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_43
timestamp 1486834041
transform 1 0 5488 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_52
timestamp 1486834041
transform 1 0 6496 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_69
timestamp 1486834041
transform 1 0 8400 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_115
timestamp 1486834041
transform 1 0 13552 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_219
timestamp 1486834041
transform 1 0 25200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_227
timestamp 1486834041
transform 1 0 26096 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_239
timestamp 1486834041
transform 1 0 27440 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_243
timestamp 1486834041
transform 1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_263
timestamp 1486834041
transform 1 0 30128 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_265
timestamp 1486834041
transform 1 0 30352 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_274
timestamp 1486834041
transform 1 0 31360 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_306
timestamp 1486834041
transform 1 0 34944 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_314
timestamp 1486834041
transform 1 0 35840 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_381
timestamp 1486834041
transform 1 0 43344 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_403
timestamp 1486834041
transform 1 0 45808 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_411
timestamp 1486834041
transform 1 0 46704 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_206
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_221
timestamp 1486834041
transform 1 0 25424 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_237
timestamp 1486834041
transform 1 0 27216 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_329
timestamp 1486834041
transform 1 0 37520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_331
timestamp 1486834041
transform 1 0 37744 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_370
timestamp 1486834041
transform 1 0 42112 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_404
timestamp 1486834041
transform 1 0 45920 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_444
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_454
timestamp 1486834041
transform 1 0 51520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_456
timestamp 1486834041
transform 1 0 51744 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 48496 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 48720 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 50064 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 50288 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 48720 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 50064 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 48496 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 50288 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 50288 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform -1 0 51632 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 46928 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 50288 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 50064 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 50288 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 50064 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 48720 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 48496 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 48608 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 47040 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 46928 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 47040 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 48720 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 48496 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 48608 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 48720 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 50288 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 48720 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 50064 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 48496 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 50288 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 37520 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 38192 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 40880 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 40208 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 41664 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 39760 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 41776 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 44352 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 37744 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 37968 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 39312 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 37072 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 37968 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 39312 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 40544 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 38640 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 12432 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 9296 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 14224 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 12432 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 14784 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 13216 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 15792 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 12432 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 16352 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 14784 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 15568 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 16352 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 15568 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 17136 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 14336 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 20272 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 20048 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 18704 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 17920 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 17136 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 16352 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 17136 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 19600 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 16912 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 17136 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 22064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 22736 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 22624 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 23632 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 23632 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 25424 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 21616 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 19488 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 21616 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 21168 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 21056 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform 1 0 35280 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 52080 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 52080 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 52080 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 52080 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 52080 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 52080 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 52080 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 52080 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 52080 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 52080 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 52080 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 52080 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 52080 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 52080 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 52080 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 52080 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_45
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_51
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_52
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_58
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_59
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_64
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_65
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_66
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_71
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_72
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_73
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_77
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_78
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_79
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_80
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_84
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_91
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_92
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_93
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_94
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_97
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_98
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_99
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_100
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_101
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_103
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_104
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_105
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_106
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_107
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_108
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_110
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_111
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_112
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_113
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_114
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_115
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_116
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_117
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_118
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_119
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_120
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_121
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_122
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_123
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_124
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_125
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_126
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_127
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_128
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_129
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_130
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_131
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_132
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_133
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_136
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_137
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_140
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_141
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_142
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_143
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 52640 0 52752 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 52640 4480 52752 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 52640 4928 52752 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 52640 5376 52752 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 52640 5824 52752 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 52640 6272 52752 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 52640 6720 52752 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 52640 7168 52752 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 52640 7616 52752 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 52640 8064 52752 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 52640 8512 52752 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 52640 448 52752 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 52640 8960 52752 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 52640 9408 52752 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 52640 9856 52752 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 52640 10304 52752 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 52640 10752 52752 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 52640 11200 52752 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 52640 11648 52752 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 52640 12096 52752 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 52640 12544 52752 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 52640 12992 52752 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 52640 896 52752 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 52640 13440 52752 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 52640 13888 52752 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 52640 1344 52752 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 52640 1792 52752 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 52640 2240 52752 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 52640 2688 52752 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 52640 3136 52752 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 52640 3584 52752 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 52640 4032 52752 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 4032 0 4144 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 28672 0 28784 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 31136 0 31248 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 33600 0 33712 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 36064 0 36176 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 38528 0 38640 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 40992 0 41104 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 43456 0 43568 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 45920 0 46032 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 48384 0 48496 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 50848 0 50960 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 6496 0 6608 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 8960 0 9072 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 13888 0 14000 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 16352 0 16464 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 18816 0 18928 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 21280 0 21392 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 23744 0 23856 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 35840 14112 35952 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 38080 14112 38192 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 38528 14112 38640 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 38976 14112 39088 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 39424 14112 39536 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 39872 14112 39984 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 36288 14112 36400 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 36736 14112 36848 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 37184 14112 37296 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 37632 14112 37744 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 12544 14112 12656 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 12992 14112 13104 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 13440 14112 13552 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 13888 14112 14000 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 14336 14112 14448 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 14784 14112 14896 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 15232 14112 15344 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 15680 14112 15792 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 16128 14112 16240 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 16576 14112 16688 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 19264 14112 19376 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 19712 14112 19824 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 20160 14112 20272 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 17024 14112 17136 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 17472 14112 17584 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 17920 14112 18032 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 18368 14112 18480 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 18816 14112 18928 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 22848 14112 22960 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 23296 14112 23408 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 23744 14112 23856 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 20608 14112 20720 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 21056 14112 21168 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 21504 14112 21616 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 21952 14112 22064 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 22400 14112 22512 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 24192 14112 24304 14224 0 FreeSans 448 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 24640 14112 24752 14224 0 FreeSans 448 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 26880 14112 26992 14224 0 FreeSans 448 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 27328 14112 27440 14224 0 FreeSans 448 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 27776 14112 27888 14224 0 FreeSans 448 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 28224 14112 28336 14224 0 FreeSans 448 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 25088 14112 25200 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 25536 14112 25648 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 25984 14112 26096 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 26432 14112 26544 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 30912 14112 31024 14224 0 FreeSans 448 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 31360 14112 31472 14224 0 FreeSans 448 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 31808 14112 31920 14224 0 FreeSans 448 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 28672 14112 28784 14224 0 FreeSans 448 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 29120 14112 29232 14224 0 FreeSans 448 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 29568 14112 29680 14224 0 FreeSans 448 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 30016 14112 30128 14224 0 FreeSans 448 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 30464 14112 30576 14224 0 FreeSans 448 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 34496 14112 34608 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 34944 14112 35056 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 35392 14112 35504 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 32256 14112 32368 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 32704 14112 32816 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 33152 14112 33264 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 33600 14112 33712 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 34048 14112 34160 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1568 0 1680 112 0 FreeSans 448 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 26376 12544 26376 12544 0 VDD
rlabel metal1 26376 13328 26376 13328 0 VSS
rlabel metal3 1470 56 1470 56 0 FrameData[0]
rlabel metal3 1134 4536 1134 4536 0 FrameData[10]
rlabel metal2 16520 6888 16520 6888 0 FrameData[11]
rlabel metal3 1638 5432 1638 5432 0 FrameData[12]
rlabel metal3 742 5880 742 5880 0 FrameData[13]
rlabel metal3 742 6328 742 6328 0 FrameData[14]
rlabel metal3 742 6776 742 6776 0 FrameData[15]
rlabel metal2 39704 5376 39704 5376 0 FrameData[16]
rlabel metal3 630 7672 630 7672 0 FrameData[17]
rlabel metal3 854 8120 854 8120 0 FrameData[18]
rlabel metal3 518 8568 518 8568 0 FrameData[19]
rlabel metal3 798 504 798 504 0 FrameData[1]
rlabel metal3 1792 6440 1792 6440 0 FrameData[20]
rlabel metal2 35448 1848 35448 1848 0 FrameData[21]
rlabel metal3 910 9912 910 9912 0 FrameData[22]
rlabel metal3 7000 10304 7000 10304 0 FrameData[23]
rlabel metal3 742 10808 742 10808 0 FrameData[24]
rlabel metal4 15288 11536 15288 11536 0 FrameData[25]
rlabel metal3 18144 1960 18144 1960 0 FrameData[26]
rlabel metal3 1512 6888 1512 6888 0 FrameData[27]
rlabel metal3 1694 12600 1694 12600 0 FrameData[28]
rlabel metal3 1190 13048 1190 13048 0 FrameData[29]
rlabel metal3 1526 952 1526 952 0 FrameData[2]
rlabel metal2 28616 1904 28616 1904 0 FrameData[30]
rlabel metal3 126 13944 126 13944 0 FrameData[31]
rlabel metal3 742 1400 742 1400 0 FrameData[3]
rlabel metal3 686 1848 686 1848 0 FrameData[4]
rlabel metal3 686 2296 686 2296 0 FrameData[5]
rlabel metal3 574 2744 574 2744 0 FrameData[6]
rlabel metal3 854 3192 854 3192 0 FrameData[7]
rlabel metal3 854 3640 854 3640 0 FrameData[8]
rlabel metal3 798 4088 798 4088 0 FrameData[9]
rlabel metal3 52122 56 52122 56 0 FrameData_O[0]
rlabel metal3 51898 4536 51898 4536 0 FrameData_O[10]
rlabel metal2 51240 4760 51240 4760 0 FrameData_O[11]
rlabel metal2 51240 5320 51240 5320 0 FrameData_O[12]
rlabel metal3 51226 5880 51226 5880 0 FrameData_O[13]
rlabel metal2 51240 6216 51240 6216 0 FrameData_O[14]
rlabel metal3 51170 6776 51170 6776 0 FrameData_O[15]
rlabel metal2 51464 6888 51464 6888 0 FrameData_O[16]
rlabel metal3 52066 7672 52066 7672 0 FrameData_O[17]
rlabel metal3 51786 8120 51786 8120 0 FrameData_O[18]
rlabel metal3 51842 8568 51842 8568 0 FrameData_O[19]
rlabel metal3 51618 504 51618 504 0 FrameData_O[1]
rlabel metal3 52066 9016 52066 9016 0 FrameData_O[20]
rlabel metal3 51842 9464 51842 9464 0 FrameData_O[21]
rlabel metal3 52066 9912 52066 9912 0 FrameData_O[22]
rlabel metal3 51170 10360 51170 10360 0 FrameData_O[23]
rlabel metal3 51954 10808 51954 10808 0 FrameData_O[24]
rlabel metal3 51282 11256 51282 11256 0 FrameData_O[25]
rlabel metal3 51842 11704 51842 11704 0 FrameData_O[26]
rlabel metal3 51226 12152 51226 12152 0 FrameData_O[27]
rlabel metal3 50442 12600 50442 12600 0 FrameData_O[28]
rlabel metal2 48104 12712 48104 12712 0 FrameData_O[29]
rlabel metal3 50442 952 50442 952 0 FrameData_O[2]
rlabel metal3 50232 9688 50232 9688 0 FrameData_O[30]
rlabel metal3 50400 9240 50400 9240 0 FrameData_O[31]
rlabel metal3 51226 1400 51226 1400 0 FrameData_O[3]
rlabel metal3 51282 1848 51282 1848 0 FrameData_O[4]
rlabel metal2 51464 2072 51464 2072 0 FrameData_O[5]
rlabel metal3 51898 2744 51898 2744 0 FrameData_O[6]
rlabel metal2 51240 3080 51240 3080 0 FrameData_O[7]
rlabel metal3 51058 3640 51058 3640 0 FrameData_O[8]
rlabel metal2 51464 3752 51464 3752 0 FrameData_O[9]
rlabel metal2 30576 56 30576 56 0 FrameStrobe[0]
rlabel metal2 28728 686 28728 686 0 FrameStrobe[10]
rlabel metal3 30576 8232 30576 8232 0 FrameStrobe[11]
rlabel metal3 15736 10192 15736 10192 0 FrameStrobe[12]
rlabel metal2 3192 12264 3192 12264 0 FrameStrobe[13]
rlabel metal4 16296 14093 16296 14093 0 FrameStrobe[14]
rlabel metal2 2184 9576 2184 9576 0 FrameStrobe[15]
rlabel metal2 43512 5558 43512 5558 0 FrameStrobe[16]
rlabel metal2 45976 182 45976 182 0 FrameStrobe[17]
rlabel metal2 48440 126 48440 126 0 FrameStrobe[18]
rlabel metal2 50904 182 50904 182 0 FrameStrobe[19]
rlabel metal2 44856 9072 44856 9072 0 FrameStrobe[1]
rlabel metal2 46424 3864 46424 3864 0 FrameStrobe[2]
rlabel metal3 48160 8232 48160 8232 0 FrameStrobe[3]
rlabel metal4 15512 2352 15512 2352 0 FrameStrobe[4]
rlabel metal2 16408 1722 16408 1722 0 FrameStrobe[5]
rlabel metal2 18872 182 18872 182 0 FrameStrobe[6]
rlabel metal2 21336 177 21336 177 0 FrameStrobe[7]
rlabel metal2 23800 182 23800 182 0 FrameStrobe[8]
rlabel metal2 26264 686 26264 686 0 FrameStrobe[9]
rlabel metal2 35896 13482 35896 13482 0 FrameStrobe_O[0]
rlabel metal2 39144 10584 39144 10584 0 FrameStrobe_O[10]
rlabel metal2 41608 12432 41608 12432 0 FrameStrobe_O[11]
rlabel metal2 40824 12096 40824 12096 0 FrameStrobe_O[12]
rlabel metal2 38808 13146 38808 13146 0 FrameStrobe_O[13]
rlabel metal2 39032 13594 39032 13594 0 FrameStrobe_O[14]
rlabel metal2 39256 13706 39256 13706 0 FrameStrobe_O[15]
rlabel metal2 39480 13202 39480 13202 0 FrameStrobe_O[16]
rlabel metal2 39704 13538 39704 13538 0 FrameStrobe_O[17]
rlabel metal2 39928 13258 39928 13258 0 FrameStrobe_O[18]
rlabel metal2 40152 13650 40152 13650 0 FrameStrobe_O[19]
rlabel metal2 36568 12712 36568 12712 0 FrameStrobe_O[1]
rlabel metal2 36344 13594 36344 13594 0 FrameStrobe_O[2]
rlabel metal2 38136 12824 38136 12824 0 FrameStrobe_O[3]
rlabel metal2 39816 13104 39816 13104 0 FrameStrobe_O[4]
rlabel metal2 37016 13202 37016 13202 0 FrameStrobe_O[5]
rlabel metal2 38696 12152 38696 12152 0 FrameStrobe_O[6]
rlabel metal2 40040 13048 40040 13048 0 FrameStrobe_O[7]
rlabel metal2 41272 13328 41272 13328 0 FrameStrobe_O[8]
rlabel metal2 39368 11592 39368 11592 0 FrameStrobe_O[9]
rlabel metal2 12376 14098 12376 14098 0 N1BEG[0]
rlabel metal2 10472 11312 10472 11312 0 N1BEG[1]
rlabel metal2 12992 7672 12992 7672 0 N1BEG[2]
rlabel metal2 10920 12040 10920 12040 0 N1BEG[3]
rlabel metal2 13272 13258 13272 13258 0 N2BEG[0]
rlabel metal2 13496 11130 13496 11130 0 N2BEG[1]
rlabel metal2 12488 10976 12488 10976 0 N2BEG[2]
rlabel metal2 13944 12978 13944 12978 0 N2BEG[3]
rlabel metal2 14560 7672 14560 7672 0 N2BEG[4]
rlabel metal2 9800 13328 9800 13328 0 N2BEG[5]
rlabel metal2 14616 13594 14616 13594 0 N2BEG[6]
rlabel metal2 12376 11984 12376 11984 0 N2BEG[7]
rlabel metal2 15176 9128 15176 9128 0 N2BEGb[0]
rlabel metal2 15288 13706 15288 13706 0 N2BEGb[1]
rlabel metal2 15512 13426 15512 13426 0 N2BEGb[2]
rlabel metal2 15736 13874 15736 13874 0 N2BEGb[3]
rlabel metal2 15960 13594 15960 13594 0 N2BEGb[4]
rlabel metal2 15624 10808 15624 10808 0 N2BEGb[5]
rlabel metal2 16408 12922 16408 12922 0 N2BEGb[6]
rlabel metal2 16632 12362 16632 12362 0 N2BEGb[7]
rlabel metal2 16856 13706 16856 13706 0 N4BEG[0]
rlabel metal2 19096 11690 19096 11690 0 N4BEG[10]
rlabel metal2 19320 12082 19320 12082 0 N4BEG[11]
rlabel metal3 18816 12264 18816 12264 0 N4BEG[12]
rlabel metal2 19880 11200 19880 11200 0 N4BEG[13]
rlabel metal3 19432 11480 19432 11480 0 N4BEG[14]
rlabel metal3 18816 13160 18816 13160 0 N4BEG[15]
rlabel metal2 17080 12474 17080 12474 0 N4BEG[1]
rlabel metal2 15512 11760 15512 11760 0 N4BEG[2]
rlabel metal2 17528 13258 17528 13258 0 N4BEG[3]
rlabel metal2 17752 13034 17752 13034 0 N4BEG[4]
rlabel metal3 18424 11480 18424 11480 0 N4BEG[5]
rlabel metal2 17640 11704 17640 11704 0 N4BEG[6]
rlabel metal2 18424 13818 18424 13818 0 N4BEG[7]
rlabel metal2 18256 10808 18256 10808 0 N4BEG[8]
rlabel metal2 16744 11984 16744 11984 0 N4BEG[9]
rlabel metal2 20888 9352 20888 9352 0 NN4BEG[0]
rlabel metal2 22680 12474 22680 12474 0 NN4BEG[10]
rlabel metal2 22904 13706 22904 13706 0 NN4BEG[11]
rlabel metal2 23128 13258 23128 13258 0 NN4BEG[12]
rlabel metal3 23128 13048 23128 13048 0 NN4BEG[13]
rlabel metal2 23576 13258 23576 13258 0 NN4BEG[14]
rlabel metal2 23800 13482 23800 13482 0 NN4BEG[15]
rlabel metal2 20664 13426 20664 13426 0 NN4BEG[1]
rlabel metal2 19880 12544 19880 12544 0 NN4BEG[2]
rlabel metal2 20720 11256 20720 11256 0 NN4BEG[3]
rlabel metal2 19208 13160 19208 13160 0 NN4BEG[4]
rlabel metal2 21560 13818 21560 13818 0 NN4BEG[5]
rlabel metal2 21784 13650 21784 13650 0 NN4BEG[6]
rlabel metal2 22008 12810 22008 12810 0 NN4BEG[7]
rlabel metal3 21952 12376 21952 12376 0 NN4BEG[8]
rlabel metal3 21840 13160 21840 13160 0 NN4BEG[9]
rlabel metal2 24024 13930 24024 13930 0 S1END[0]
rlabel metal2 24248 13594 24248 13594 0 S1END[1]
rlabel metal2 21896 504 21896 504 0 S1END[2]
rlabel metal2 22624 9016 22624 9016 0 S1END[3]
rlabel metal2 38920 3024 38920 3024 0 S2END[0]
rlabel metal2 27272 10752 27272 10752 0 S2END[1]
rlabel metal2 27216 3752 27216 3752 0 S2END[2]
rlabel metal2 24360 5936 24360 5936 0 S2END[3]
rlabel metal2 35784 8232 35784 8232 0 S2END[4]
rlabel metal2 27832 13090 27832 13090 0 S2END[5]
rlabel metal3 34216 1232 34216 1232 0 S2END[6]
rlabel metal4 25032 11430 25032 11430 0 S2END[7]
rlabel metal2 24920 13986 24920 13986 0 S2MID[0]
rlabel metal2 49560 7840 49560 7840 0 S2MID[1]
rlabel metal2 47768 3696 47768 3696 0 S2MID[2]
rlabel metal2 43960 5320 43960 5320 0 S2MID[3]
rlabel metal2 42616 12488 42616 12488 0 S2MID[4]
rlabel metal2 24360 10584 24360 10584 0 S2MID[5]
rlabel metal2 20888 1568 20888 1568 0 S2MID[6]
rlabel metal2 22456 10360 22456 10360 0 S2MID[7]
rlabel metal4 25480 9800 25480 9800 0 S4END[0]
rlabel metal2 44632 6608 44632 6608 0 S4END[10]
rlabel via3 15624 477 15624 477 0 S4END[11]
rlabel metal2 46760 4032 46760 4032 0 S4END[12]
rlabel metal2 38696 10136 38696 10136 0 S4END[13]
rlabel metal3 46816 5880 46816 5880 0 S4END[14]
rlabel metal2 31864 13650 31864 13650 0 S4END[15]
rlabel metal3 21280 3752 21280 3752 0 S4END[1]
rlabel metal2 25256 11872 25256 11872 0 S4END[2]
rlabel metal3 21896 5880 21896 5880 0 S4END[3]
rlabel metal2 43848 2576 43848 2576 0 S4END[4]
rlabel metal3 24920 11592 24920 11592 0 S4END[5]
rlabel metal2 2408 4144 2408 4144 0 S4END[6]
rlabel metal2 16632 6384 16632 6384 0 S4END[7]
rlabel metal2 41944 10752 41944 10752 0 S4END[8]
rlabel metal3 24248 6384 24248 6384 0 S4END[9]
rlabel metal2 32648 6720 32648 6720 0 SS4END[0]
rlabel metal2 20776 2576 20776 2576 0 SS4END[10]
rlabel metal2 16184 1960 16184 1960 0 SS4END[11]
rlabel metal2 20328 4312 20328 4312 0 SS4END[12]
rlabel metal3 16352 2968 16352 2968 0 SS4END[13]
rlabel metal2 35224 13986 35224 13986 0 SS4END[14]
rlabel metal2 35448 13650 35448 13650 0 SS4END[15]
rlabel metal4 16520 9423 16520 9423 0 SS4END[1]
rlabel metal2 18424 5096 18424 5096 0 SS4END[2]
rlabel metal3 26012 9912 26012 9912 0 SS4END[3]
rlabel metal2 16744 6272 16744 6272 0 SS4END[4]
rlabel metal4 16800 3150 16800 3150 0 SS4END[5]
rlabel metal2 33432 13314 33432 13314 0 SS4END[6]
rlabel metal4 20888 11088 20888 11088 0 SS4END[7]
rlabel metal4 16072 8344 16072 8344 0 SS4END[8]
rlabel metal2 6440 1848 6440 1848 0 SS4END[9]
rlabel metal2 1624 742 1624 742 0 UserCLK
rlabel metal2 35728 13160 35728 13160 0 UserCLKo
rlabel metal2 46200 4256 46200 4256 0 net1
rlabel metal2 51352 4368 51352 4368 0 net10
rlabel metal3 21112 2072 21112 2072 0 net100
rlabel metal2 16296 12264 16296 12264 0 net101
rlabel metal2 16520 12040 16520 12040 0 net102
rlabel metal2 16520 8512 16520 8512 0 net103
rlabel metal3 22288 6664 22288 6664 0 net104
rlabel metal3 31584 10024 31584 10024 0 net105
rlabel metal3 39368 9184 39368 9184 0 net11
rlabel metal2 47096 2800 47096 2800 0 net12
rlabel metal3 39144 9856 39144 9856 0 net13
rlabel metal3 41552 2072 41552 2072 0 net14
rlabel metal2 2184 2912 2184 2912 0 net15
rlabel metal2 30296 672 30296 672 0 net16
rlabel via3 30072 971 30072 971 0 net17
rlabel metal2 48888 11256 48888 11256 0 net18
rlabel metal3 45080 3808 45080 3808 0 net19
rlabel metal3 46760 9688 46760 9688 0 net2
rlabel metal3 45304 5152 45304 5152 0 net20
rlabel metal2 47208 11256 47208 11256 0 net21
rlabel metal2 46984 10528 46984 10528 0 net22
rlabel metal4 28840 840 28840 840 0 net23
rlabel metal3 47824 3416 47824 3416 0 net24
rlabel metal2 48552 7644 48552 7644 0 net25
rlabel metal2 16296 4088 16296 4088 0 net26
rlabel metal3 47432 2072 47432 2072 0 net27
rlabel metal2 50400 2184 50400 2184 0 net28
rlabel metal2 46648 5824 46648 5824 0 net29
rlabel metal3 48104 4760 48104 4760 0 net3
rlabel metal3 49336 8680 49336 8680 0 net30
rlabel metal3 47152 4984 47152 4984 0 net31
rlabel metal2 47544 2240 47544 2240 0 net32
rlabel metal2 51240 13216 51240 13216 0 net33
rlabel metal2 18536 7616 18536 7616 0 net34
rlabel metal2 41048 10080 41048 10080 0 net35
rlabel metal2 34552 1680 34552 1680 0 net36
rlabel metal2 2744 12544 2744 12544 0 net37
rlabel metal2 32424 2352 32424 2352 0 net38
rlabel metal2 1848 10696 1848 10696 0 net39
rlabel metal3 49504 10472 49504 10472 0 net4
rlabel metal2 40376 7672 40376 7672 0 net40
rlabel metal2 39928 7504 39928 7504 0 net41
rlabel metal2 42056 9240 42056 9240 0 net42
rlabel metal2 44296 11480 44296 11480 0 net43
rlabel metal2 45304 9744 45304 9744 0 net44
rlabel metal2 46984 3584 46984 3584 0 net45
rlabel metal2 49112 7448 49112 7448 0 net46
rlabel metal2 39144 12432 39144 12432 0 net47
rlabel metal3 31808 6552 31808 6552 0 net48
rlabel metal2 25592 7280 25592 7280 0 net49
rlabel metal2 46312 4592 46312 4592 0 net5
rlabel metal2 39480 11200 39480 11200 0 net50
rlabel metal4 28504 1568 28504 1568 0 net51
rlabel metal2 16520 1680 16520 1680 0 net52
rlabel metal3 16744 9072 16744 9072 0 net53
rlabel metal2 9576 8288 9576 8288 0 net54
rlabel metal4 15400 8155 15400 8155 0 net55
rlabel metal3 19432 3304 19432 3304 0 net56
rlabel metal2 21896 7728 21896 7728 0 net57
rlabel metal2 20440 2352 20440 2352 0 net58
rlabel metal3 17472 2072 17472 2072 0 net59
rlabel metal2 50232 5544 50232 5544 0 net6
rlabel metal2 43176 9184 43176 9184 0 net60
rlabel metal2 48552 6216 48552 6216 0 net61
rlabel metal2 48216 4480 48216 4480 0 net62
rlabel metal2 30408 2240 30408 2240 0 net63
rlabel metal3 15512 12040 15512 12040 0 net64
rlabel metal3 16520 2856 16520 2856 0 net65
rlabel metal2 42840 4144 42840 4144 0 net66
rlabel metal3 19376 7560 19376 7560 0 net67
rlabel metal2 44856 2296 44856 2296 0 net68
rlabel metal3 21168 5992 21168 5992 0 net69
rlabel metal2 48776 7392 48776 7392 0 net7
rlabel metal2 21336 3864 21336 3864 0 net70
rlabel metal2 25256 10192 25256 10192 0 net71
rlabel metal2 39368 5600 39368 5600 0 net72
rlabel metal4 15176 11880 15176 11880 0 net73
rlabel metal3 20552 8232 20552 8232 0 net74
rlabel metal3 21952 3304 21952 3304 0 net75
rlabel metal3 16632 8680 16632 8680 0 net76
rlabel metal3 17416 10248 17416 10248 0 net77
rlabel metal2 8960 6664 8960 6664 0 net78
rlabel metal2 22568 5320 22568 5320 0 net79
rlabel metal2 45304 3696 45304 3696 0 net8
rlabel metal3 48664 5992 48664 5992 0 net80
rlabel metal3 23016 13888 23016 13888 0 net81
rlabel metal2 47320 7952 47320 7952 0 net82
rlabel metal2 5880 10584 5880 10584 0 net83
rlabel metal2 45080 5880 45080 5880 0 net84
rlabel metal3 16072 9184 16072 9184 0 net85
rlabel metal2 22120 9072 22120 9072 0 net86
rlabel metal2 17192 9128 17192 9128 0 net87
rlabel metal2 2016 3416 2016 3416 0 net88
rlabel metal2 30520 2464 30520 2464 0 net89
rlabel metal3 49560 8344 49560 8344 0 net9
rlabel metal2 16632 9800 16632 9800 0 net90
rlabel metal4 16520 5992 16520 5992 0 net91
rlabel metal2 24584 9968 24584 9968 0 net92
rlabel metal3 21672 10360 21672 10360 0 net93
rlabel metal3 17192 13104 17192 13104 0 net94
rlabel metal2 26824 7000 26824 7000 0 net95
rlabel metal2 21560 12824 21560 12824 0 net96
rlabel metal2 18872 6160 18872 6160 0 net97
rlabel metal2 19768 7504 19768 7504 0 net98
rlabel metal2 18088 8288 18088 8288 0 net99
<< properties >>
string FIXED_BBOX 0 0 52752 14224
<< end >>
