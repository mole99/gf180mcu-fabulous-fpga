* NGSPICE file created from W_IO4.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

.subckt W_IO4 A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 C_I_top C_O_top C_T_top C_config_C_bit0 C_config_C_bit1 C_config_C_bit2
+ C_config_C_bit3 D_I_top D_O_top D_T_top D_config_C_bit0 D_config_C_bit1 D_config_C_bit2
+ D_config_C_bit3 E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3]
+ E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4]
+ E2BEGb[5] E2BEGb[6] E2BEGb[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3]
+ E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] EE4BEG[0] EE4BEG[10] EE4BEG[11]
+ EE4BEG[12] EE4BEG[13] EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4]
+ EE4BEG[5] EE4BEG[6] EE4BEG[7] EE4BEG[8] EE4BEG[9] FrameData[0] FrameData[10] FrameData[11]
+ FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17]
+ FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22]
+ FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28]
+ FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4]
+ FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] UserCLK UserCLKo VDD VSS W1END[0] W1END[1] W1END[2] W1END[3] W2END[0]
+ W2END[1] W2END[2] W2END[3] W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1]
+ W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6] W2MID[7] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XTAP_TAPCELL_ROW_49_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_432_ FrameData[28] net111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_363_ Inst_W_IO4_switch_matrix.E2BEG3 net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_39_Left_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_294_ FrameData[6] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_346_ FrameData[26] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_415_ FrameData[11] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_277_ FrameData[21] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_24_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_200_ W2END[1] WW4END[1] WW4END[9] W6END[1] Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q Inst_W_IO4_switch_matrix.E2BEGb6 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_25_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_131_ W2END[4] W2END[5] W2END[6] W2END[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q _042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_329_ FrameData[9] net53 Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_24_Left_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_114_ _003_ Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q
+ _026_ _027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_46_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Left_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput7 net144 B_I_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput20 net20 D_T_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput31 net31 E2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput42 net60 E2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput64 net82 EE4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput53 net71 E6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput75 net93 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput86 net104 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput97 net115 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_31_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_431_ FrameData[27] net110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_362_ Inst_W_IO4_switch_matrix.E2BEG2 net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_293_ FrameData[5] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_414_ FrameData[10] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_345_ FrameData[25] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_276_ FrameData[20] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_58_Left_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Left_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q _040_ _041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_328_ FrameData[8] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_259_ FrameData[3] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_54_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_113_ W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q _026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput87 net105 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput10 net10 B_config_C_bit1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput8 net8 B_T_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput21 net21 D_config_C_bit0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput32 net32 E2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput65 net83 EE4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput43 net61 E2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput54 net72 E6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput98 net116 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput76 net94 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_430_ FrameData[26] net109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_361_ Inst_W_IO4_switch_matrix.E2BEG1 net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_292_ FrameData[4] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_67_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_413_ FrameData[9] net122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_344_ FrameData[24] net53 Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_275_ FrameData[19] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_327_ FrameData[7] net54 Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_189_ W6END[3] W6END[7] W6END[5] D_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q Inst_W_IO4_switch_matrix.EE4BEG9 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_258_ FrameData[2] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_112_ Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q _020_ _021_ _022_ _025_ net8 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_46_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput88 net106 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput9 net9 B_config_C_bit0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput11 net11 B_config_C_bit2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput22 net22 D_config_C_bit1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput33 net33 E2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput44 net62 E2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput66 net84 EE4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput55 net73 E6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput99 net117 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput77 net95 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_31_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_360_ Inst_W_IO4_switch_matrix.E2BEG0 net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_291_ FrameData[3] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_412_ FrameData[8] net121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_343_ FrameData[23] net53 Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_274_ FrameData[18] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_68_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_326_ FrameData[6] net54 Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_257_ FrameData[1] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_188_ W6END[0] W6END[2] W6END[4] A_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q Inst_W_IO4_switch_matrix.EE4BEG10 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_62_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_111_ Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q _023_ _024_ _025_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_28_Left_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_309_ FrameData[21] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput12 net12 B_config_C_bit3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput23 net23 D_config_C_bit2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput34 net34 E2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput89 net107 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput67 net85 EE4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput45 net63 E6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput56 net74 E6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput78 net96 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_15_Left_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_290_ FrameData[2] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_342_ FrameData[22] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_411_ FrameData[7] net120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_273_ FrameData[17] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_68_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Left_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Left_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_325_ FrameData[5] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_54_Left_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_256_ FrameData[0] net46 Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_187_ W6END[6] W6END[8] W6END[10] B_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q Inst_W_IO4_switch_matrix.EE4BEG11 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_63_Left_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_110_ W2END[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q _024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire126 net7 net144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_3_Left_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_239_ FrameData[15] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_308_ FrameData[20] net50 Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net145 C_I_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput24 net24 D_config_C_bit3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput35 net35 E2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput57 net75 EE4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput46 net64 E6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput68 net86 EE4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput79 net97 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_341_ FrameData[21] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_410_ FrameData[6] net119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_272_ FrameData[16] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_255_ FrameData[31] net41 Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_324_ FrameData[4] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_186_ W6END[1] W6END[3] W6END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q Inst_W_IO4_switch_matrix.EE4BEG12 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_62_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire127 net13 net145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_238_ FrameData[14] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_169_ Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q _074_ _076_ _011_ _077_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_307_ FrameData[19] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput14 net14 C_T_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput25 net25 E1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput36 net36 E2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput69 net87 EE4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput58 net76 EE4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput47 net65 E6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_54_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_340_ FrameData[20] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_271_ FrameData[15] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_19_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_254_ FrameData[30] net41 Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_185_ W6END[7] W6END[9] W6END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q Inst_W_IO4_switch_matrix.EE4BEG13 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_323_ FrameData[3] net55 Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_306_ FrameData[18] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_168_ _000_ Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q
+ _075_ _076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_237_ FrameData[13] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_099_ _004_ W2END[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q _014_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 C_config_C_bit0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput26 net26 E1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput37 net37 E2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput59 net77 EE4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput48 net66 E6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_270_ FrameData[14] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_19_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_399_ Inst_W_IO4_switch_matrix.EE4BEG11 net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_322_ FrameData[2] net55 Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_64_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_184_ W2MID[2] W2MID[4] W2MID[6] Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q Inst_W_IO4_switch_matrix.EE4BEG14 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_253_ FrameData[29] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfanout50 FrameStrobe[1] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_32_Left_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_50_Left_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_305_ FrameData[17] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_098_ _003_ Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q
+ _012_ _013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_236_ FrameData[12] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_167_ W2MID[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q _075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_219_ FrameData[27] net38 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput16 net16 C_config_C_bit1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput27 net27 E1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput38 net56 E2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput49 net67 E6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_17_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_398_ Inst_W_IO4_switch_matrix.EE4BEG10 net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout51 net52 net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_24_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_252_ FrameData[28] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfanout40 FrameStrobe[3] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_321_ FrameData[1] net55 Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_183_ W2MID[3] W2MID[7] W2MID[5] Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q Inst_W_IO4_switch_matrix.EE4BEG15 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_304_ FrameData[16] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_235_ FrameData[11] net42 Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_097_ W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q _012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_166_ W2MID[6] W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q _074_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_23_Left_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_149_ W2END[0] W2END[2] W2END[1] W2END[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q _058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_218_ FrameData[26] net38 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput17 net17 C_config_C_bit2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput28 net28 E1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput39 net57 E2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_10_Left_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_397_ Inst_W_IO4_switch_matrix.EE4BEG9 net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout52 net53 net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_251_ FrameData[27] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfanout41 FrameStrobe[3] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_182_ W1END[2] A_O_top WW4END[11] C_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q Inst_W_IO4_switch_matrix.E6BEG0 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_320_ FrameData[0] net55 Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_13_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_449_ FrameStrobe[13] net127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_165_ Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q _072_ _073_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_234_ FrameData[10] net41 Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_303_ FrameData[15] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_096_ W1END[2] A_O_top W1END[3] C_O_top Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q
+ Inst_W_IO4_switch_matrix.E1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_217_ FrameData[25] net38 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_148_ Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q _055_ _057_ _051_ _053_ net13 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_51_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_079_ W2MID[7] _001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_29_Left_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput18 net18 C_config_C_bit3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput29 net29 E2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_396_ Inst_W_IO4_switch_matrix.EE4BEG8 net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_250_ FrameData[26] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfanout53 net54 net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout42 FrameStrobe[3] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_181_ W1END[3] Inst_A_IO_1_bidirectional_frame_config_pass.Q WW4END[10] Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q
+ Inst_W_IO4_switch_matrix.E6BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_448_ FrameStrobe[12] net126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_30_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_379_ Inst_W_IO4_switch_matrix.E6BEG3 net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_302_ FrameData[14] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_164_ W2MID[0] W2MID[1] W2MID[2] W2MID[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q _072_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_233_ FrameData[9] net42 Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_095_ W1END[1] W1END[2] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q
+ Inst_W_IO4_switch_matrix.E1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ FrameData[24] net38 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_147_ Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q _056_ _057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_078_ W2MID[5] _000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput19 net19 D_I_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_15_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_57_Left_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_66_Left_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_395_ Inst_W_IO4_switch_matrix.EE4BEG7 net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout43 net46 net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_180_ WW4END[7] WW4END[15] A_O_top C_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q Inst_W_IO4_switch_matrix.E6BEG2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout54 net55 net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_70_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_447_ FrameStrobe[11] net125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_378_ Inst_W_IO4_switch_matrix.E6BEG2 net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_232_ FrameData[8] net41 Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_301_ FrameData[13] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_163_ _011_ _070_ Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q _071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_094_ W1END[0] W1END[1] B_O_top D_O_top Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q
+ Inst_W_IO4_switch_matrix.E1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_60_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_215_ FrameData[23] net38 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_146_ W2MID[0] W2MID[1] W2MID[2] W2MID[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q _056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_129_ W2END[0] W2END[2] W2END[1] W2END[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q _040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Left_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_394_ Inst_W_IO4_switch_matrix.EE4BEG6 net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout44 net45 net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout55 FrameStrobe[0] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_446_ FrameStrobe[10] net124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_30_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_377_ Inst_W_IO4_switch_matrix.E6BEG1 net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_61_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_162_ W2END[4] W2END[5] W2END[6] W2END[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q _070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_300_ FrameData[12] net50 Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_231_ FrameData[7] net42 Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_093_ W1END[0] W1END[3] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q
+ Inst_W_IO4_switch_matrix.E1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_429_ FrameData[25] net108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_214_ FrameData[22] net38 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_145_ _009_ _054_ _055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_128_ Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q _034_ _035_ _036_ _039_ net20 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_7_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_393_ Inst_W_IO4_switch_matrix.EE4BEG5 net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_10_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout45 net46 net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_445_ FrameStrobe[9] net142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_376_ Inst_W_IO4_switch_matrix.E6BEG0 net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_161_ Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q _068_ _069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_230_ FrameData[6] net42 Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_092_ W2MID[7] WW4END[7] WW4END[15] W6END[7] Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q Inst_W_IO4_switch_matrix.E2BEG0 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_428_ FrameData[24] net107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_359_ Inst_W_IO4_switch_matrix.E1BEG3 net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_213_ FrameData[21] net38 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_144_ W2MID[4] W2MID[6] W2MID[5] W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q _054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_127_ Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q _037_ _038_ _039_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Left_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Left_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_392_ Inst_W_IO4_switch_matrix.EE4BEG4 net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout46 FrameStrobe[2] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_444_ FrameStrobe[8] net141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_375_ Inst_W_IO4_switch_matrix.E2BEGb7 net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_091_ W2MID[6] WW4END[6] WW4END[14] W6END[6] Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q Inst_W_IO4_switch_matrix.E2BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_160_ W2END[0] W2END[2] W2END[1] W2END[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q _068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_358_ Inst_W_IO4_switch_matrix.E1BEG2 net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_427_ FrameData[23] net106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_289_ FrameData[1] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_212_ FrameData[20] net38 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_143_ _009_ _052_ Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q _053_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_126_ W2END[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q _038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_109_ Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q W2END[6] Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q
+ _023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_391_ Inst_W_IO4_switch_matrix.EE4BEG3 net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Left_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout47 net50 net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_1_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_374_ Inst_W_IO4_switch_matrix.E2BEGb6 net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_443_ FrameStrobe[7] net140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_090_ W2MID[5] WW4END[5] WW4END[13] W6END[5] Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q Inst_W_IO4_switch_matrix.E2BEG2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_426_ FrameData[22] net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_357_ Inst_W_IO4_switch_matrix.E1BEG1 net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_288_ FrameData[0] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_142_ W2END[4] W2END[5] W2END[6] W2END[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q _052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_211_ W2MID[4] WW4END[4] WW4END[12] W6END[4] Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q Inst_W_IO4_switch_matrix.E2BEG3 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_409_ FrameData[5] net118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_6_Left_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_125_ W2END[6] Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q
+ _037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_16_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_108_ _001_ Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q
+ _022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_390_ Inst_W_IO4_switch_matrix.EE4BEG2 net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_9_Left_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xfanout48 net50 net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_70_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_442_ FrameStrobe[6] net139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_373_ Inst_W_IO4_switch_matrix.E2BEGb5 net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_59_Left_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_425_ FrameData[21] net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_287_ FrameData[31] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_356_ Inst_W_IO4_switch_matrix.E1BEG0 net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_141_ Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q _050_ _051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_210_ W2MID[3] WW4END[3] WW4END[11] W6END[3] Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q Inst_W_IO4_switch_matrix.E2BEG4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ FrameData[4] net117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_339_ FrameData[19] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_22_Left_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_124_ _001_ Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q
+ _036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_16_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_107_ _005_ W2END[5] Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q _021_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_31_Left_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Left_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout38 FrameStrobe[4] net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_24_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout49 net50 net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_441_ FrameStrobe[5] net138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_57_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_372_ Inst_W_IO4_switch_matrix.E2BEGb4 net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_424_ FrameData[20] net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_286_ FrameData[30] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_355_ D_O_top clknet_1_1__leaf_UserCLK_regs Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_46_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ W2END[0] W2END[2] W2END[1] W2END[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q _050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_338_ FrameData[18] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_407_ FrameData[3] net116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_269_ FrameData[13] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_123_ W2END[5] _007_ Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q _035_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_106_ _002_ Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q
+ _019_ _020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_19_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout39 net40 net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_1_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_440_ net38 net137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_371_ Inst_W_IO4_switch_matrix.E2BEGb3 net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_52_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_423_ FrameData[19] net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_354_ C_O_top clknet_1_0__leaf_UserCLK_regs Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_285_ FrameData[29] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_337_ FrameData[17] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_406_ FrameData[2] net113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_199_ W2END[0] WW4END[0] WW4END[8] W6END[0] Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q Inst_W_IO4_switch_matrix.E2BEGb7 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_268_ FrameData[12] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_70_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_122_ _002_ Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q
+ _033_ _034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ W2MID[6] Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q _019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_370_ Inst_W_IO4_switch_matrix.E2BEGb2 net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_55_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_422_ FrameData[18] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_284_ FrameData[28] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_353_ B_O_top clknet_1_1__leaf_UserCLK_regs Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_51_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_267_ FrameData[11] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_336_ FrameData[16] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_405_ FrameData[1] net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_198_ W6END[0] W6END[2] W6END[4] A_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q Inst_W_IO4_switch_matrix.EE4BEG0 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput120 net138 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_70_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_121_ W2MID[6] Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q _033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_319_ FrameData[31] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_42_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_104_ Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q _013_ _014_ _015_ _018_ net2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_14_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_13_Left_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_421_ FrameData[17] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_283_ FrameData[27] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_352_ A_O_top clknet_1_0__leaf_UserCLK_regs Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_50_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_404_ FrameData[0] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_266_ FrameData[10] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_335_ FrameData[15] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_197_ W6END[6] W6END[8] W6END[10] B_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q Inst_W_IO4_switch_matrix.EE4BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_47_Left_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_Left_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput110 net128 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput121 net139 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_65_Left_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_120_ Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q _027_ _028_ _029_ _032_ net14 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_1_Left_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_249_ FrameData[25] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_318_ FrameData[30] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_103_ Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q _016_ _017_ _018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_351_ FrameData[31] net54 Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_420_ FrameData[16] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_282_ FrameData[26] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_65_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_334_ FrameData[14] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_403_ Inst_W_IO4_switch_matrix.EE4BEG15 net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_265_ FrameData[9] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_196_ W6END[1] W6END[3] W6END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q Inst_W_IO4_switch_matrix.EE4BEG2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput111 net129 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput122 net140 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput100 net118 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_62_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_317_ FrameData[29] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_248_ FrameData[24] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_179_ WW4END[6] WW4END[14] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q
+ Inst_W_IO4_switch_matrix.E6BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_102_ W2END[2] Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q _017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_350_ FrameData[30] net54 Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_281_ FrameData[25] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_30_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_264_ FrameData[8] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_333_ FrameData[13] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_402_ Inst_W_IO4_switch_matrix.EE4BEG14 net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_195_ W6END[7] W6END[9] W6END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q Inst_W_IO4_switch_matrix.EE4BEG3 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput112 net130 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput123 net141 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput101 net119 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_55_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_316_ FrameData[28] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_247_ FrameData[23] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_178_ W1END[2] A_O_top WW4END[3] C_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q Inst_W_IO4_switch_matrix.E6BEG4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_101_ Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q W2END[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q
+ _016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_17_Left_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_280_ FrameData[24] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_401_ Inst_W_IO4_switch_matrix.EE4BEG13 net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_332_ FrameData[12] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_263_ FrameData[7] net44 Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_194_ W2END[2] W2END[4] W2END[6] C_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q Inst_W_IO4_switch_matrix.EE4BEG4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput113 net131 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput124 net142 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_34_Left_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput102 net120 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_43_Left_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Left_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_70_Left_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_246_ FrameData[22] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_315_ FrameData[27] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_177_ W1END[3] Inst_A_IO_1_bidirectional_frame_config_pass.Q WW4END[2] Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q
+ Inst_W_IO4_switch_matrix.E6BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_100_ _002_ Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q
+ _015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Left_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_229_ FrameData[5] net41 Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_331_ FrameData[11] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_400_ Inst_W_IO4_switch_matrix.EE4BEG12 net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_193_ W2END[3] W2END[5] W2END[7] D_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q Inst_W_IO4_switch_matrix.EE4BEG5 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_262_ FrameData[6] net45 Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput125 net143 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput114 net132 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput103 net121 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_63_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_314_ FrameData[26] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_176_ W1END[1] B_O_top WW4END[9] D_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q Inst_W_IO4_switch_matrix.E6BEG6 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_245_ FrameData[21] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Left_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_28_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_159_ Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q _063_ _067_ _059_ _061_ net7 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_228_ FrameData[4] net42 Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_67_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_330_ FrameData[10] net53 Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_192_ W2MID[2] W2MID[4] W2MID[6] Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q Inst_W_IO4_switch_matrix.EE4BEG6 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_261_ FrameData[5] net46 Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput115 net133 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput104 net122 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_313_ FrameData[25] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_244_ FrameData[20] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_175_ W1END[0] Inst_B_IO_1_bidirectional_frame_config_pass.Q WW4END[8] Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q
+ Inst_W_IO4_switch_matrix.E6BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_227_ FrameData[3] net41 net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_158_ Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q _064_ _066_ _010_ _067_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_6_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_089_ Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q _011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_69_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Left_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_260_ FrameData[4] net46 Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_191_ W2MID[3] W2MID[7] W2MID[5] Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q Inst_W_IO4_switch_matrix.EE4BEG7 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_389_ Inst_W_IO4_switch_matrix.EE4BEG1 net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput116 net134 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput105 net123 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_49_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_312_ FrameData[24] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_243_ FrameData[19] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_30_Left_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_174_ WW4END[5] WW4END[13] B_O_top D_O_top Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q Inst_W_IO4_switch_matrix.E6BEG8 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_157_ _000_ Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q
+ _065_ _066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_226_ FrameData[2] net41 net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_088_ Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q _010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_25_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_209_ W2MID[2] WW4END[2] WW4END[10] W6END[2] Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q Inst_W_IO4_switch_matrix.E2BEG5 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_68_Left_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_190_ W6END[6] W6END[8] W6END[10] C_O_top Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q Inst_W_IO4_switch_matrix.EE4BEG8 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_388_ Inst_W_IO4_switch_matrix.EE4BEG0 net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput106 net124 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput117 net135 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_55_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_242_ FrameData[18] net39 Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_311_ FrameData[23] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_173_ WW4END[4] WW4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q
+ Inst_W_IO4_switch_matrix.E6BEG9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_9_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_6_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_156_ W2MID[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q _065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_087_ Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q _009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_225_ FrameData[1] net41 net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Left_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_208_ W2MID[1] WW4END[1] WW4END[9] W6END[1] Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q Inst_W_IO4_switch_matrix.E2BEG6 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_139_ Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q _045_ _049_ _041_ _043_ net19 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_24_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_54_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_456_ clknet_1_0__leaf_UserCLK net143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput107 net125 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_387_ Inst_W_IO4_switch_matrix.E6BEG11 net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput118 net136 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_310_ FrameData[22] net48 Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_241_ FrameData[17] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_172_ W1END[1] B_O_top WW4END[1] D_O_top Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q Inst_W_IO4_switch_matrix.E6BEG10 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_9_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_439_ net41 net136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_224_ FrameData[0] net41 net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_086_ Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q _008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_155_ W2MID[6] W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q _064_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_0_Left_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_207_ W2MID[0] WW4END[0] WW4END[8] W6END[0] Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q Inst_W_IO4_switch_matrix.E2BEG7 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_138_ Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q _046_ _048_ _008_ _049_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_455_ FrameStrobe[19] net133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_386_ Inst_W_IO4_switch_matrix.E6BEG10 net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput108 net126 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput119 net137 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_70_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput90 net108 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_240_ FrameData[16] net40 Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_171_ W1END[0] Inst_B_IO_1_bidirectional_frame_config_pass.Q WW4END[0] Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q
+ Inst_W_IO4_switch_matrix.E6BEG11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_9_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_369_ Inst_W_IO4_switch_matrix.E2BEGb1 net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_438_ net45 net135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_47_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ FrameData[31] net38 net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_085_ Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q _007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_10_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_154_ Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q _062_ _063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_137_ _000_ Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q
+ _047_ _048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_206_ W2END[7] WW4END[15] WW4END[7] W6END[7] Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q Inst_W_IO4_switch_matrix.E2BEGb0 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Left_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Left_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_55_Left_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Left_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_454_ FrameStrobe[18] net132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_385_ Inst_W_IO4_switch_matrix.E6BEG9 net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net127 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput1 net1 A_I_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput91 net109 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput80 net98 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_31_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_170_ Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q _073_ _077_ _069_ _071_ net1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_37_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_299_ FrameData[11] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_368_ Inst_W_IO4_switch_matrix.E2BEGb0 net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_437_ net50 net134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_222_ FrameData[30] FrameStrobe[4] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_153_ W2MID[0] W2MID[1] W2MID[2] W2MID[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q _062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_084_ Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q _006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_136_ Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q W2MID[4] _047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_205_ W2END[6] WW4END[14] WW4END[6] W6END[6] Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q
+ Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q Inst_W_IO4_switch_matrix.E2BEGb1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_119_ Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q _030_ _031_ _032_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Left_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_453_ FrameStrobe[17] net131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_384_ Inst_W_IO4_switch_matrix.E6BEG8 net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput2 net2 A_T_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput70 net88 EE4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput92 net110 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput81 net99 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_31_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_436_ net55 net123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_367_ Inst_W_IO4_switch_matrix.E2BEG7 net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_298_ FrameData[10] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_14_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_083_ Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q _005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_152_ _010_ _060_ Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q _061_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_221_ FrameData[29] FrameStrobe[4] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_419_ FrameData[15] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_204_ W2END[5] WW4END[13] WW4END[5] W6END[5] Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q Inst_W_IO4_switch_matrix.E2BEGb2 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_135_ W2MID[6] W2MID[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q _046_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_40_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_118_ W2END[2] Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q _031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_452_ FrameStrobe[16] net130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_383_ Inst_W_IO4_switch_matrix.E6BEG7 net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net111 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput82 net100 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput3 net3 A_config_C_bit0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput60 net78 EE4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput71 net89 EE4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_22_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_435_ FrameData[31] net115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_366_ Inst_W_IO4_switch_matrix.E2BEG6 net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_297_ FrameData[9] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_220_ FrameData[28] FrameStrobe[4] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_151_ W2END[4] W2END[5] W2END[6] W2END[7] Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q _060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_082_ Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q _004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_349_ FrameData[29] net54 Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_418_ FrameData[14] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_43_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_203_ W2END[4] WW4END[4] WW4END[12] W6END[4] Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q Inst_W_IO4_switch_matrix.E2BEGb3 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_40_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_134_ Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q _044_ _045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_22_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ W2END[4] Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q
+ _030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_451_ FrameStrobe[15] net129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_382_ Inst_W_IO4_switch_matrix.E6BEG6 net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput83 net101 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput4 net4 A_config_C_bit1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput72 net90 EE4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput61 net79 EE4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput50 net68 E6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput94 net112 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_63_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_434_ FrameData[30] net114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_296_ FrameData[8] net47 Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_365_ Inst_W_IO4_switch_matrix.E2BEG5 net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_46_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_150_ Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q _058_ _059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_081_ W2END[1] _003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_348_ FrameData[28] net51 Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_417_ FrameData[13] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_279_ FrameData[23] net46 Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_43_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_133_ W2MID[0] W2MID[1] W2MID[2] W2MID[3] Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q
+ Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q _044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_40_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_202_ W2END[3] WW4END[3] WW4END[11] W6END[3] Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q Inst_W_IO4_switch_matrix.E2BEGb4 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_116_ _002_ Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q
+ _029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_450_ FrameStrobe[14] net128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_381_ Inst_W_IO4_switch_matrix.E6BEG5 net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput5 net5 A_config_C_bit2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput40 net58 E2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput62 net80 EE4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput51 net69 E6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput73 net91 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput95 net113 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput84 net102 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_49_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_433_ FrameData[29] net112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_364_ Inst_W_IO4_switch_matrix.E2BEG4 net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_295_ FrameData[7] net49 Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_46_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_080_ W2END[0] _002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_12_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_416_ FrameData[12] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_28_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_347_ FrameData[27] net52 Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
X_278_ FrameData[22] net43 Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_43_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_132_ _008_ _042_ Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q _043_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_201_ W2END[2] WW4END[2] WW4END[10] W6END[2] Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q
+ Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q Inst_W_IO4_switch_matrix.E2BEGb5 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_115_ W2END[3] _006_ Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q _028_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_380_ Inst_W_IO4_switch_matrix.E6BEG4 net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 A_config_C_bit3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput30 net30 E2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput41 net59 E2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput52 net70 E6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput85 net103 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput96 net114 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput63 net81 EE4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput74 net92 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
.ends

