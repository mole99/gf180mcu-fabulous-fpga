VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO GF_SRAM
  CLASS BLOCK ;
  FOREIGN GF_SRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 158.480 BY 574.560 ;
  PIN A_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 99.680 158.480 100.240 ;
    END
  END A_SRAM0
  PIN A_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 104.160 158.480 104.720 ;
    END
  END A_SRAM1
  PIN A_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 108.640 158.480 109.200 ;
    END
  END A_SRAM2
  PIN A_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 113.120 158.480 113.680 ;
    END
  END A_SRAM3
  PIN A_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 117.600 158.480 118.160 ;
    END
  END A_SRAM4
  PIN A_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 122.080 158.480 122.640 ;
    END
  END A_SRAM5
  PIN A_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 126.560 158.480 127.120 ;
    END
  END A_SRAM6
  PIN A_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 131.040 158.480 131.600 ;
    END
  END A_SRAM7
  PIN A_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 135.520 158.480 136.080 ;
    END
  END A_SRAM8
  PIN CEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 54.880 158.480 55.440 ;
    END
  END CEN_SRAM
  PIN CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 175.840 158.480 176.400 ;
    END
  END CLK_SRAM
  PIN CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 50.400 158.480 50.960 ;
    END
  END CONFIGURED_top
  PIN D_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 140.000 158.480 140.560 ;
    END
  END D_SRAM0
  PIN D_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 144.480 158.480 145.040 ;
    END
  END D_SRAM1
  PIN D_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 148.960 158.480 149.520 ;
    END
  END D_SRAM2
  PIN D_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 153.440 158.480 154.000 ;
    END
  END D_SRAM3
  PIN D_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 157.920 158.480 158.480 ;
    END
  END D_SRAM4
  PIN D_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 162.400 158.480 162.960 ;
    END
  END D_SRAM5
  PIN D_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 166.880 158.480 167.440 ;
    END
  END D_SRAM6
  PIN D_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 171.360 158.480 171.920 ;
    END
  END D_SRAM7
  PIN GWEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 59.360 158.480 59.920 ;
    END
  END GWEN_SRAM
  PIN Q_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 14.560 158.480 15.120 ;
    END
  END Q_SRAM0
  PIN Q_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 19.040 158.480 19.600 ;
    END
  END Q_SRAM1
  PIN Q_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 23.520 158.480 24.080 ;
    END
  END Q_SRAM2
  PIN Q_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 28.000 158.480 28.560 ;
    END
  END Q_SRAM3
  PIN Q_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.531500 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 32.480 158.480 33.040 ;
    END
  END Q_SRAM4
  PIN Q_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.528500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 36.960 158.480 37.520 ;
    END
  END Q_SRAM5
  PIN Q_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 41.440 158.480 42.000 ;
    END
  END Q_SRAM6
  PIN Q_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.030000 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 45.920 158.480 46.480 ;
    END
  END Q_SRAM7
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 395.920 0.560 396.480 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.160 0.560 398.720 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.400 0.560 400.960 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.640 0.560 403.200 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 422.800 0.560 423.360 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.040 0.560 425.600 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 427.280 0.560 427.840 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 429.520 0.560 430.080 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.901000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.760 0.560 432.320 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 434.000 0.560 434.560 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.240 0.560 436.800 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 438.480 0.560 439.040 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.892000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.880 0.560 405.440 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.892000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 407.120 0.560 407.680 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.892000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 409.360 0.560 409.920 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.892000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.600 0.560 412.160 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.892000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.840 0.560 414.400 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.080 0.560 416.640 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 418.320 0.560 418.880 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.560 0.560 421.120 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.560 0.560 477.120 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 498.960 0.560 499.520 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 501.200 0.560 501.760 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.800 0.560 479.360 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.040 0.560 481.600 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.280 0.560 483.840 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 485.520 0.560 486.080 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.760 0.560 488.320 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.000 0.560 490.560 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.240 0.560 492.800 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 494.480 0.560 495.040 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 496.720 0.560 497.280 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 440.720 0.560 441.280 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.120 0.560 463.680 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.360 0.560 465.920 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 467.600 0.560 468.160 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.840 0.560 470.400 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.080 0.560 472.640 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 474.320 0.560 474.880 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.960 0.560 443.520 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 445.200 0.560 445.760 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 447.440 0.560 448.000 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 449.680 0.560 450.240 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 451.920 0.560 452.480 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.160 0.560 454.720 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 456.400 0.560 456.960 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 458.640 0.560 459.200 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.880 0.560 461.440 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 503.440 0.560 504.000 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.840 0.560 526.400 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.080 0.560 528.640 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.320 0.560 530.880 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.560 0.560 533.120 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.800 0.560 535.360 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.040 0.560 537.600 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 539.280 0.560 539.840 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 541.520 0.560 542.080 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.760 0.560 544.320 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.000 0.560 546.560 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 505.680 0.560 506.240 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.240 0.560 548.800 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 550.480 0.560 551.040 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.720 0.560 553.280 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.960 0.560 555.520 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.200 0.560 557.760 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 559.440 0.560 560.000 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.680 0.560 562.240 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 563.920 0.560 564.480 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 566.160 0.560 566.720 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 568.400 0.560 568.960 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 507.920 0.560 508.480 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 570.640 0.560 571.200 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 572.880 0.560 573.440 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.160 0.560 510.720 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 512.400 0.560 512.960 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.640 0.560 515.200 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 516.880 0.560 517.440 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.120 0.560 519.680 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.360 0.560 521.920 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 523.600 0.560 524.160 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 390.880 158.480 391.440 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 446.880 158.480 447.440 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 452.480 158.480 453.040 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 458.080 158.480 458.640 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 463.680 158.480 464.240 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 469.280 158.480 469.840 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 474.880 158.480 475.440 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 480.480 158.480 481.040 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 486.080 158.480 486.640 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 491.680 158.480 492.240 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 497.280 158.480 497.840 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 396.480 158.480 397.040 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 502.880 158.480 503.440 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 508.480 158.480 509.040 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 514.080 158.480 514.640 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 519.680 158.480 520.240 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 525.280 158.480 525.840 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 530.880 158.480 531.440 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 536.480 158.480 537.040 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 542.080 158.480 542.640 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 547.680 158.480 548.240 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 553.280 158.480 553.840 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 402.080 158.480 402.640 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 558.880 158.480 559.440 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 564.480 158.480 565.040 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 407.680 158.480 408.240 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 413.280 158.480 413.840 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 418.880 158.480 419.440 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 424.480 158.480 425.040 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 430.080 158.480 430.640 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 435.680 158.480 436.240 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 441.280 158.480 441.840 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 574.000 109.200 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 574.000 120.400 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 574.000 121.520 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 574.000 122.640 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 574.000 123.760 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 574.000 124.880 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 574.000 126.000 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 574.000 127.120 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 574.000 128.240 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 574.000 129.360 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 574.000 130.480 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 574.000 110.320 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 574.000 111.440 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 574.000 112.560 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 574.000 113.680 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 574.000 114.800 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 574.000 115.920 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 574.000 117.040 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 574.000 118.160 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 574.000 119.280 574.560 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 574.000 27.440 574.560 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 574.000 28.560 574.560 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 574.000 29.680 574.560 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 574.000 30.800 574.560 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 574.000 31.920 574.560 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 574.000 33.040 574.560 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 574.000 34.160 574.560 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 574.000 35.280 574.560 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 574.000 36.400 574.560 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 574.000 37.520 574.560 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 574.000 38.640 574.560 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 574.000 39.760 574.560 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 574.000 40.880 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 574.000 42.000 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 574.000 43.120 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 574.000 44.240 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 574.000 45.360 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 574.000 46.480 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 574.000 47.600 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 574.000 48.720 574.560 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 574.000 49.840 574.560 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 574.000 61.040 574.560 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 574.000 62.160 574.560 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 574.000 63.280 574.560 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 574.000 64.400 574.560 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 574.000 65.520 574.560 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 574.000 66.640 574.560 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 574.000 50.960 574.560 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 574.000 52.080 574.560 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 574.000 53.200 574.560 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 574.000 54.320 574.560 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 574.000 55.440 574.560 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 574.000 56.560 574.560 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 574.000 57.680 574.560 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 574.000 58.800 574.560 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 574.000 59.920 574.560 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.564500 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 574.000 67.760 574.560 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.564500 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 574.000 68.880 574.560 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.564500 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 574.000 70.000 574.560 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.564500 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 574.000 71.120 574.560 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 574.000 81.200 574.560 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 574.000 82.320 574.560 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 574.000 83.440 574.560 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 574.000 84.560 574.560 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 574.000 85.680 574.560 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 574.000 86.800 574.560 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 574.000 87.920 574.560 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 574.000 89.040 574.560 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 574.000 72.240 574.560 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 574.000 73.360 574.560 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.901000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 574.000 74.480 574.560 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.207000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 574.000 75.600 574.560 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 574.000 76.720 574.560 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 574.000 77.840 574.560 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 574.000 78.960 574.560 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 574.000 80.080 574.560 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 574.000 90.160 574.560 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 574.000 101.360 574.560 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 574.000 102.480 574.560 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 574.000 103.600 574.560 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 574.000 104.720 574.560 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 574.000 105.840 574.560 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 574.000 106.960 574.560 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 574.000 91.280 574.560 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 574.000 92.400 574.560 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    ANTENNADIFFAREA 2.462400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 574.000 93.520 574.560 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 574.000 94.640 574.560 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 574.000 95.760 574.560 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 574.000 96.880 574.560 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 574.000 98.000 574.560 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 574.000 99.120 574.560 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 574.000 100.240 574.560 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 574.000 108.080 574.560 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.400 0.560 288.960 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.640 0.560 291.200 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.880 0.560 293.440 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.120 0.560 295.680 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.360 0.560 297.920 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.600 0.560 300.160 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.840 0.560 302.400 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.080 0.560 304.640 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.320 0.560 306.880 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.560 0.560 309.120 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.800 0.560 311.360 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.040 0.560 313.600 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.280 0.560 315.840 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 317.520 0.560 318.080 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.760 0.560 320.320 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.000 0.560 322.560 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.240 0.560 324.800 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.480 0.560 327.040 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.720 0.560 329.280 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.960 0.560 331.520 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.040 0.560 369.600 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 391.440 0.560 392.000 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.680 0.560 394.240 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 371.280 0.560 371.840 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 373.520 0.560 374.080 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.760 0.560 376.320 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 378.000 0.560 378.560 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.240 0.560 380.800 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 382.480 0.560 383.040 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.720 0.560 385.280 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.960 0.560 387.520 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.200 0.560 389.760 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.200 0.560 333.760 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 0.560 356.160 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 357.840 0.560 358.400 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 360.080 0.560 360.640 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.320 0.560 362.880 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.560 0.560 365.120 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 366.800 0.560 367.360 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 335.440 0.560 336.000 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.680 0.560 338.240 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.920 0.560 340.480 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.160 0.560 342.720 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.400 0.560 344.960 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.640 0.560 347.200 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.880 0.560 349.440 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.120 0.560 351.680 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.360 0.560 353.920 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.108000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 108.640 0.560 109.200 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 0.560 111.440 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 0.560 113.680 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 0.560 115.920 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.952000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 0.560 136.080 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.955000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 0.560 138.320 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.955000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 0.560 140.560 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.877500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 0.560 142.800 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.207000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 0.560 145.040 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.117000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 0.560 147.280 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 0.560 149.520 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 0.560 151.760 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.042500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 0.560 118.160 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.952000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 0.560 120.400 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.952000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 0.560 122.640 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.955000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 0.560 124.880 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 0.560 127.120 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 0.560 129.360 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.006000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 0.560 131.600 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 0.560 133.840 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.606500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 0.560 189.840 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 0.560 212.240 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 0.560 214.480 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 0.560 192.080 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 0.560 194.320 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.453500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 0.560 196.560 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.904000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 0.560 198.800 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.480 0.560 201.040 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 0.560 203.280 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 0.560 205.520 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 0.560 207.760 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 209.440 0.560 210.000 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 0.560 154.000 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 175.840 0.560 176.400 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 0.560 178.640 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 0.560 180.880 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 0.560 183.120 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 0.560 185.360 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 0.560 187.600 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 0.560 156.240 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 0.560 158.480 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 0.560 160.720 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 0.560 162.960 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 0.560 165.200 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 0.560 167.440 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 0.560 169.680 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 0.560 171.920 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 0.560 174.160 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 0.560 216.720 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 0.560 239.120 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 0.560 241.360 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.040 0.560 243.600 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 0.560 245.840 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 247.520 0.560 248.080 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 0.560 250.320 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 0.560 252.560 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.240 0.560 254.800 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 0.560 257.040 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 0.560 259.280 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 0.560 218.960 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 0.560 261.520 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 0.560 263.760 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 0.560 266.000 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.680 0.560 268.240 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 0.560 270.480 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 0.560 272.720 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 0.560 274.960 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.640 0.560 277.200 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 0.560 279.440 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.120 0.560 281.680 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.640 0.560 221.200 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.360 0.560 283.920 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.466500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 0.560 286.160 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 0.560 223.440 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 0.560 225.680 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 0.560 227.920 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 0.560 230.160 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.840 0.560 232.400 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 0.560 234.640 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 0.560 236.880 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 199.360 158.480 199.920 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 255.360 158.480 255.920 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 260.960 158.480 261.520 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 266.560 158.480 267.120 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 272.160 158.480 272.720 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 277.760 158.480 278.320 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 283.360 158.480 283.920 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 288.960 158.480 289.520 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 294.560 158.480 295.120 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 300.160 158.480 300.720 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 305.760 158.480 306.320 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 204.960 158.480 205.520 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 311.360 158.480 311.920 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 316.960 158.480 317.520 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 322.560 158.480 323.120 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 328.160 158.480 328.720 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 333.760 158.480 334.320 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 339.360 158.480 339.920 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 344.960 158.480 345.520 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 350.560 158.480 351.120 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 356.160 158.480 356.720 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 361.760 158.480 362.320 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 210.560 158.480 211.120 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 367.360 158.480 367.920 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 372.960 158.480 373.520 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 216.160 158.480 216.720 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 221.760 158.480 222.320 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 227.360 158.480 227.920 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 232.960 158.480 233.520 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 238.560 158.480 239.120 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 244.160 158.480 244.720 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 249.760 158.480 250.320 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 0.000 130.480 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 47.602497 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.858500 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 0.560 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.456500 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 0.560 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.396500 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 0.560 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.396500 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 0.560 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.396500 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 0.560 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 0.560 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 0.560 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.568500 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 0.560 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.399500 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 0.560 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 0.560 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 0.560 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 0.560 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 0.560 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 0.000 31.920 0.560 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 0.560 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 0.560 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 0.560 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 0.560 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 0.560 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.901000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 0.560 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 0.560 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 0.560 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 0.560 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 0.560 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 0.560 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 0.560 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 0.560 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 0.560 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 0.560 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 0.560 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 0.560 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 0.560 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 0.560 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 0.560 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.507500 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 0.560 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 0.560 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 0.560 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 0.560 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 0.560 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 0.560 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 0.560 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 0.560 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 0.560 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 0.560 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 0.560 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 0.560 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 0.560 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 0.560 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 0.560 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 0.560 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 0.560 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 0.560 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 0.560 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 0.560 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 0.560 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 0.560 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 0.560 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 0.560 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 0.560 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 0.560 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 0.560 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 0.560 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 0.560 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 0.560 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 0.560 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 0.560 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 0.560 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.120 0.560 1.680 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.360 0.560 3.920 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 5.600 0.560 6.160 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.840 0.560 8.400 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.080 0.560 10.640 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 0.560 12.880 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 0.560 15.120 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 0.560 17.360 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 0.560 19.600 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 0.560 21.840 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 0.560 24.080 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 0.560 26.320 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 0.560 28.560 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 0.560 30.800 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 0.560 33.040 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 0.560 35.280 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 0.560 37.520 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 0.560 39.760 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 0.560 42.000 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 0.560 44.240 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 0.560 82.320 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 0.560 104.720 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 0.560 106.960 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 0.560 84.560 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.240 0.560 86.800 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 0.560 89.040 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 0.560 91.280 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 0.560 93.520 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 0.560 95.760 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 0.560 98.000 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 0.560 100.240 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 0.560 102.480 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 0.560 46.480 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 0.560 68.880 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 0.560 71.120 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 0.560 73.360 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 0.560 75.600 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 0.560 77.840 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 0.560 80.080 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 0.560 48.720 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 0.560 50.960 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 0.560 53.200 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 0.560 55.440 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 0.560 57.680 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 0.560 59.920 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 0.560 62.160 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 0.560 64.400 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 0.560 66.640 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 0.000 20.480 574.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.880 0.000 120.480 574.560 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 0.000 23.780 574.560 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.180 0.000 123.780 574.560 ;
    END
  END VSS
  PIN WEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 63.840 158.480 64.400 ;
    END
  END WEN_SRAM0
  PIN WEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 68.320 158.480 68.880 ;
    END
  END WEN_SRAM1
  PIN WEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 72.800 158.480 73.360 ;
    END
  END WEN_SRAM2
  PIN WEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 77.280 158.480 77.840 ;
    END
  END WEN_SRAM3
  PIN WEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 81.760 158.480 82.320 ;
    END
  END WEN_SRAM4
  PIN WEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 86.240 158.480 86.800 ;
    END
  END WEN_SRAM5
  PIN WEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 90.720 158.480 91.280 ;
    END
  END WEN_SRAM6
  PIN WEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 157.920 95.200 158.480 95.760 ;
    END
  END WEN_SRAM7
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 155.550 568.830 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 155.120 568.700 ;
      LAYER Metal2 ;
        RECT 0.140 573.700 26.580 574.000 ;
        RECT 130.780 573.700 157.780 574.000 ;
        RECT 0.140 0.860 157.780 573.700 ;
        RECT 0.140 0.090 26.580 0.860 ;
        RECT 130.780 0.090 157.780 0.860 ;
      LAYER Metal3 ;
        RECT 0.090 573.740 158.340 573.860 ;
        RECT 0.860 572.580 158.340 573.740 ;
        RECT 0.090 571.500 158.340 572.580 ;
        RECT 0.860 570.340 158.340 571.500 ;
        RECT 0.090 569.260 158.340 570.340 ;
        RECT 0.860 568.100 158.340 569.260 ;
        RECT 0.090 567.020 158.340 568.100 ;
        RECT 0.860 565.860 158.340 567.020 ;
        RECT 0.090 565.340 158.340 565.860 ;
        RECT 0.090 564.780 157.620 565.340 ;
        RECT 0.860 564.180 157.620 564.780 ;
        RECT 0.860 563.620 158.340 564.180 ;
        RECT 0.090 562.540 158.340 563.620 ;
        RECT 0.860 561.380 158.340 562.540 ;
        RECT 0.090 560.300 158.340 561.380 ;
        RECT 0.860 559.740 158.340 560.300 ;
        RECT 0.860 559.140 157.620 559.740 ;
        RECT 0.090 558.580 157.620 559.140 ;
        RECT 0.090 558.060 158.340 558.580 ;
        RECT 0.860 556.900 158.340 558.060 ;
        RECT 0.090 555.820 158.340 556.900 ;
        RECT 0.860 554.660 158.340 555.820 ;
        RECT 0.090 554.140 158.340 554.660 ;
        RECT 0.090 553.580 157.620 554.140 ;
        RECT 0.860 552.980 157.620 553.580 ;
        RECT 0.860 552.420 158.340 552.980 ;
        RECT 0.090 551.340 158.340 552.420 ;
        RECT 0.860 550.180 158.340 551.340 ;
        RECT 0.090 549.100 158.340 550.180 ;
        RECT 0.860 548.540 158.340 549.100 ;
        RECT 0.860 547.940 157.620 548.540 ;
        RECT 0.090 547.380 157.620 547.940 ;
        RECT 0.090 546.860 158.340 547.380 ;
        RECT 0.860 545.700 158.340 546.860 ;
        RECT 0.090 544.620 158.340 545.700 ;
        RECT 0.860 543.460 158.340 544.620 ;
        RECT 0.090 542.940 158.340 543.460 ;
        RECT 0.090 542.380 157.620 542.940 ;
        RECT 0.860 541.780 157.620 542.380 ;
        RECT 0.860 541.220 158.340 541.780 ;
        RECT 0.090 540.140 158.340 541.220 ;
        RECT 0.860 538.980 158.340 540.140 ;
        RECT 0.090 537.900 158.340 538.980 ;
        RECT 0.860 537.340 158.340 537.900 ;
        RECT 0.860 536.740 157.620 537.340 ;
        RECT 0.090 536.180 157.620 536.740 ;
        RECT 0.090 535.660 158.340 536.180 ;
        RECT 0.860 534.500 158.340 535.660 ;
        RECT 0.090 533.420 158.340 534.500 ;
        RECT 0.860 532.260 158.340 533.420 ;
        RECT 0.090 531.740 158.340 532.260 ;
        RECT 0.090 531.180 157.620 531.740 ;
        RECT 0.860 530.580 157.620 531.180 ;
        RECT 0.860 530.020 158.340 530.580 ;
        RECT 0.090 528.940 158.340 530.020 ;
        RECT 0.860 527.780 158.340 528.940 ;
        RECT 0.090 526.700 158.340 527.780 ;
        RECT 0.860 526.140 158.340 526.700 ;
        RECT 0.860 525.540 157.620 526.140 ;
        RECT 0.090 524.980 157.620 525.540 ;
        RECT 0.090 524.460 158.340 524.980 ;
        RECT 0.860 523.300 158.340 524.460 ;
        RECT 0.090 522.220 158.340 523.300 ;
        RECT 0.860 521.060 158.340 522.220 ;
        RECT 0.090 520.540 158.340 521.060 ;
        RECT 0.090 519.980 157.620 520.540 ;
        RECT 0.860 519.380 157.620 519.980 ;
        RECT 0.860 518.820 158.340 519.380 ;
        RECT 0.090 517.740 158.340 518.820 ;
        RECT 0.860 516.580 158.340 517.740 ;
        RECT 0.090 515.500 158.340 516.580 ;
        RECT 0.860 514.940 158.340 515.500 ;
        RECT 0.860 514.340 157.620 514.940 ;
        RECT 0.090 513.780 157.620 514.340 ;
        RECT 0.090 513.260 158.340 513.780 ;
        RECT 0.860 512.100 158.340 513.260 ;
        RECT 0.090 511.020 158.340 512.100 ;
        RECT 0.860 509.860 158.340 511.020 ;
        RECT 0.090 509.340 158.340 509.860 ;
        RECT 0.090 508.780 157.620 509.340 ;
        RECT 0.860 508.180 157.620 508.780 ;
        RECT 0.860 507.620 158.340 508.180 ;
        RECT 0.090 506.540 158.340 507.620 ;
        RECT 0.860 505.380 158.340 506.540 ;
        RECT 0.090 504.300 158.340 505.380 ;
        RECT 0.860 503.740 158.340 504.300 ;
        RECT 0.860 503.140 157.620 503.740 ;
        RECT 0.090 502.580 157.620 503.140 ;
        RECT 0.090 502.060 158.340 502.580 ;
        RECT 0.860 500.900 158.340 502.060 ;
        RECT 0.090 499.820 158.340 500.900 ;
        RECT 0.860 498.660 158.340 499.820 ;
        RECT 0.090 498.140 158.340 498.660 ;
        RECT 0.090 497.580 157.620 498.140 ;
        RECT 0.860 496.980 157.620 497.580 ;
        RECT 0.860 496.420 158.340 496.980 ;
        RECT 0.090 495.340 158.340 496.420 ;
        RECT 0.860 494.180 158.340 495.340 ;
        RECT 0.090 493.100 158.340 494.180 ;
        RECT 0.860 492.540 158.340 493.100 ;
        RECT 0.860 491.940 157.620 492.540 ;
        RECT 0.090 491.380 157.620 491.940 ;
        RECT 0.090 490.860 158.340 491.380 ;
        RECT 0.860 489.700 158.340 490.860 ;
        RECT 0.090 488.620 158.340 489.700 ;
        RECT 0.860 487.460 158.340 488.620 ;
        RECT 0.090 486.940 158.340 487.460 ;
        RECT 0.090 486.380 157.620 486.940 ;
        RECT 0.860 485.780 157.620 486.380 ;
        RECT 0.860 485.220 158.340 485.780 ;
        RECT 0.090 484.140 158.340 485.220 ;
        RECT 0.860 482.980 158.340 484.140 ;
        RECT 0.090 481.900 158.340 482.980 ;
        RECT 0.860 481.340 158.340 481.900 ;
        RECT 0.860 480.740 157.620 481.340 ;
        RECT 0.090 480.180 157.620 480.740 ;
        RECT 0.090 479.660 158.340 480.180 ;
        RECT 0.860 478.500 158.340 479.660 ;
        RECT 0.090 477.420 158.340 478.500 ;
        RECT 0.860 476.260 158.340 477.420 ;
        RECT 0.090 475.740 158.340 476.260 ;
        RECT 0.090 475.180 157.620 475.740 ;
        RECT 0.860 474.580 157.620 475.180 ;
        RECT 0.860 474.020 158.340 474.580 ;
        RECT 0.090 472.940 158.340 474.020 ;
        RECT 0.860 471.780 158.340 472.940 ;
        RECT 0.090 470.700 158.340 471.780 ;
        RECT 0.860 470.140 158.340 470.700 ;
        RECT 0.860 469.540 157.620 470.140 ;
        RECT 0.090 468.980 157.620 469.540 ;
        RECT 0.090 468.460 158.340 468.980 ;
        RECT 0.860 467.300 158.340 468.460 ;
        RECT 0.090 466.220 158.340 467.300 ;
        RECT 0.860 465.060 158.340 466.220 ;
        RECT 0.090 464.540 158.340 465.060 ;
        RECT 0.090 463.980 157.620 464.540 ;
        RECT 0.860 463.380 157.620 463.980 ;
        RECT 0.860 462.820 158.340 463.380 ;
        RECT 0.090 461.740 158.340 462.820 ;
        RECT 0.860 460.580 158.340 461.740 ;
        RECT 0.090 459.500 158.340 460.580 ;
        RECT 0.860 458.940 158.340 459.500 ;
        RECT 0.860 458.340 157.620 458.940 ;
        RECT 0.090 457.780 157.620 458.340 ;
        RECT 0.090 457.260 158.340 457.780 ;
        RECT 0.860 456.100 158.340 457.260 ;
        RECT 0.090 455.020 158.340 456.100 ;
        RECT 0.860 453.860 158.340 455.020 ;
        RECT 0.090 453.340 158.340 453.860 ;
        RECT 0.090 452.780 157.620 453.340 ;
        RECT 0.860 452.180 157.620 452.780 ;
        RECT 0.860 451.620 158.340 452.180 ;
        RECT 0.090 450.540 158.340 451.620 ;
        RECT 0.860 449.380 158.340 450.540 ;
        RECT 0.090 448.300 158.340 449.380 ;
        RECT 0.860 447.740 158.340 448.300 ;
        RECT 0.860 447.140 157.620 447.740 ;
        RECT 0.090 446.580 157.620 447.140 ;
        RECT 0.090 446.060 158.340 446.580 ;
        RECT 0.860 444.900 158.340 446.060 ;
        RECT 0.090 443.820 158.340 444.900 ;
        RECT 0.860 442.660 158.340 443.820 ;
        RECT 0.090 442.140 158.340 442.660 ;
        RECT 0.090 441.580 157.620 442.140 ;
        RECT 0.860 440.980 157.620 441.580 ;
        RECT 0.860 440.420 158.340 440.980 ;
        RECT 0.090 439.340 158.340 440.420 ;
        RECT 0.860 438.180 158.340 439.340 ;
        RECT 0.090 437.100 158.340 438.180 ;
        RECT 0.860 436.540 158.340 437.100 ;
        RECT 0.860 435.940 157.620 436.540 ;
        RECT 0.090 435.380 157.620 435.940 ;
        RECT 0.090 434.860 158.340 435.380 ;
        RECT 0.860 433.700 158.340 434.860 ;
        RECT 0.090 432.620 158.340 433.700 ;
        RECT 0.860 431.460 158.340 432.620 ;
        RECT 0.090 430.940 158.340 431.460 ;
        RECT 0.090 430.380 157.620 430.940 ;
        RECT 0.860 429.780 157.620 430.380 ;
        RECT 0.860 429.220 158.340 429.780 ;
        RECT 0.090 428.140 158.340 429.220 ;
        RECT 0.860 426.980 158.340 428.140 ;
        RECT 0.090 425.900 158.340 426.980 ;
        RECT 0.860 425.340 158.340 425.900 ;
        RECT 0.860 424.740 157.620 425.340 ;
        RECT 0.090 424.180 157.620 424.740 ;
        RECT 0.090 423.660 158.340 424.180 ;
        RECT 0.860 422.500 158.340 423.660 ;
        RECT 0.090 421.420 158.340 422.500 ;
        RECT 0.860 420.260 158.340 421.420 ;
        RECT 0.090 419.740 158.340 420.260 ;
        RECT 0.090 419.180 157.620 419.740 ;
        RECT 0.860 418.580 157.620 419.180 ;
        RECT 0.860 418.020 158.340 418.580 ;
        RECT 0.090 416.940 158.340 418.020 ;
        RECT 0.860 415.780 158.340 416.940 ;
        RECT 0.090 414.700 158.340 415.780 ;
        RECT 0.860 414.140 158.340 414.700 ;
        RECT 0.860 413.540 157.620 414.140 ;
        RECT 0.090 412.980 157.620 413.540 ;
        RECT 0.090 412.460 158.340 412.980 ;
        RECT 0.860 411.300 158.340 412.460 ;
        RECT 0.090 410.220 158.340 411.300 ;
        RECT 0.860 409.060 158.340 410.220 ;
        RECT 0.090 408.540 158.340 409.060 ;
        RECT 0.090 407.980 157.620 408.540 ;
        RECT 0.860 407.380 157.620 407.980 ;
        RECT 0.860 406.820 158.340 407.380 ;
        RECT 0.090 405.740 158.340 406.820 ;
        RECT 0.860 404.580 158.340 405.740 ;
        RECT 0.090 403.500 158.340 404.580 ;
        RECT 0.860 402.940 158.340 403.500 ;
        RECT 0.860 402.340 157.620 402.940 ;
        RECT 0.090 401.780 157.620 402.340 ;
        RECT 0.090 401.260 158.340 401.780 ;
        RECT 0.860 400.100 158.340 401.260 ;
        RECT 0.090 399.020 158.340 400.100 ;
        RECT 0.860 397.860 158.340 399.020 ;
        RECT 0.090 397.340 158.340 397.860 ;
        RECT 0.090 396.780 157.620 397.340 ;
        RECT 0.860 396.180 157.620 396.780 ;
        RECT 0.860 395.620 158.340 396.180 ;
        RECT 0.090 394.540 158.340 395.620 ;
        RECT 0.860 393.380 158.340 394.540 ;
        RECT 0.090 392.300 158.340 393.380 ;
        RECT 0.860 391.740 158.340 392.300 ;
        RECT 0.860 391.140 157.620 391.740 ;
        RECT 0.090 390.580 157.620 391.140 ;
        RECT 0.090 390.060 158.340 390.580 ;
        RECT 0.860 388.900 158.340 390.060 ;
        RECT 0.090 387.820 158.340 388.900 ;
        RECT 0.860 386.660 158.340 387.820 ;
        RECT 0.090 385.580 158.340 386.660 ;
        RECT 0.860 384.420 158.340 385.580 ;
        RECT 0.090 383.340 158.340 384.420 ;
        RECT 0.860 382.180 158.340 383.340 ;
        RECT 0.090 381.100 158.340 382.180 ;
        RECT 0.860 379.940 158.340 381.100 ;
        RECT 0.090 378.860 158.340 379.940 ;
        RECT 0.860 377.700 158.340 378.860 ;
        RECT 0.090 376.620 158.340 377.700 ;
        RECT 0.860 375.460 158.340 376.620 ;
        RECT 0.090 374.380 158.340 375.460 ;
        RECT 0.860 373.820 158.340 374.380 ;
        RECT 0.860 373.220 157.620 373.820 ;
        RECT 0.090 372.660 157.620 373.220 ;
        RECT 0.090 372.140 158.340 372.660 ;
        RECT 0.860 370.980 158.340 372.140 ;
        RECT 0.090 369.900 158.340 370.980 ;
        RECT 0.860 368.740 158.340 369.900 ;
        RECT 0.090 368.220 158.340 368.740 ;
        RECT 0.090 367.660 157.620 368.220 ;
        RECT 0.860 367.060 157.620 367.660 ;
        RECT 0.860 366.500 158.340 367.060 ;
        RECT 0.090 365.420 158.340 366.500 ;
        RECT 0.860 364.260 158.340 365.420 ;
        RECT 0.090 363.180 158.340 364.260 ;
        RECT 0.860 362.620 158.340 363.180 ;
        RECT 0.860 362.020 157.620 362.620 ;
        RECT 0.090 361.460 157.620 362.020 ;
        RECT 0.090 360.940 158.340 361.460 ;
        RECT 0.860 359.780 158.340 360.940 ;
        RECT 0.090 358.700 158.340 359.780 ;
        RECT 0.860 357.540 158.340 358.700 ;
        RECT 0.090 357.020 158.340 357.540 ;
        RECT 0.090 356.460 157.620 357.020 ;
        RECT 0.860 355.860 157.620 356.460 ;
        RECT 0.860 355.300 158.340 355.860 ;
        RECT 0.090 354.220 158.340 355.300 ;
        RECT 0.860 353.060 158.340 354.220 ;
        RECT 0.090 351.980 158.340 353.060 ;
        RECT 0.860 351.420 158.340 351.980 ;
        RECT 0.860 350.820 157.620 351.420 ;
        RECT 0.090 350.260 157.620 350.820 ;
        RECT 0.090 349.740 158.340 350.260 ;
        RECT 0.860 348.580 158.340 349.740 ;
        RECT 0.090 347.500 158.340 348.580 ;
        RECT 0.860 346.340 158.340 347.500 ;
        RECT 0.090 345.820 158.340 346.340 ;
        RECT 0.090 345.260 157.620 345.820 ;
        RECT 0.860 344.660 157.620 345.260 ;
        RECT 0.860 344.100 158.340 344.660 ;
        RECT 0.090 343.020 158.340 344.100 ;
        RECT 0.860 341.860 158.340 343.020 ;
        RECT 0.090 340.780 158.340 341.860 ;
        RECT 0.860 340.220 158.340 340.780 ;
        RECT 0.860 339.620 157.620 340.220 ;
        RECT 0.090 339.060 157.620 339.620 ;
        RECT 0.090 338.540 158.340 339.060 ;
        RECT 0.860 337.380 158.340 338.540 ;
        RECT 0.090 336.300 158.340 337.380 ;
        RECT 0.860 335.140 158.340 336.300 ;
        RECT 0.090 334.620 158.340 335.140 ;
        RECT 0.090 334.060 157.620 334.620 ;
        RECT 0.860 333.460 157.620 334.060 ;
        RECT 0.860 332.900 158.340 333.460 ;
        RECT 0.090 331.820 158.340 332.900 ;
        RECT 0.860 330.660 158.340 331.820 ;
        RECT 0.090 329.580 158.340 330.660 ;
        RECT 0.860 329.020 158.340 329.580 ;
        RECT 0.860 328.420 157.620 329.020 ;
        RECT 0.090 327.860 157.620 328.420 ;
        RECT 0.090 327.340 158.340 327.860 ;
        RECT 0.860 326.180 158.340 327.340 ;
        RECT 0.090 325.100 158.340 326.180 ;
        RECT 0.860 323.940 158.340 325.100 ;
        RECT 0.090 323.420 158.340 323.940 ;
        RECT 0.090 322.860 157.620 323.420 ;
        RECT 0.860 322.260 157.620 322.860 ;
        RECT 0.860 321.700 158.340 322.260 ;
        RECT 0.090 320.620 158.340 321.700 ;
        RECT 0.860 319.460 158.340 320.620 ;
        RECT 0.090 318.380 158.340 319.460 ;
        RECT 0.860 317.820 158.340 318.380 ;
        RECT 0.860 317.220 157.620 317.820 ;
        RECT 0.090 316.660 157.620 317.220 ;
        RECT 0.090 316.140 158.340 316.660 ;
        RECT 0.860 314.980 158.340 316.140 ;
        RECT 0.090 313.900 158.340 314.980 ;
        RECT 0.860 312.740 158.340 313.900 ;
        RECT 0.090 312.220 158.340 312.740 ;
        RECT 0.090 311.660 157.620 312.220 ;
        RECT 0.860 311.060 157.620 311.660 ;
        RECT 0.860 310.500 158.340 311.060 ;
        RECT 0.090 309.420 158.340 310.500 ;
        RECT 0.860 308.260 158.340 309.420 ;
        RECT 0.090 307.180 158.340 308.260 ;
        RECT 0.860 306.620 158.340 307.180 ;
        RECT 0.860 306.020 157.620 306.620 ;
        RECT 0.090 305.460 157.620 306.020 ;
        RECT 0.090 304.940 158.340 305.460 ;
        RECT 0.860 303.780 158.340 304.940 ;
        RECT 0.090 302.700 158.340 303.780 ;
        RECT 0.860 301.540 158.340 302.700 ;
        RECT 0.090 301.020 158.340 301.540 ;
        RECT 0.090 300.460 157.620 301.020 ;
        RECT 0.860 299.860 157.620 300.460 ;
        RECT 0.860 299.300 158.340 299.860 ;
        RECT 0.090 298.220 158.340 299.300 ;
        RECT 0.860 297.060 158.340 298.220 ;
        RECT 0.090 295.980 158.340 297.060 ;
        RECT 0.860 295.420 158.340 295.980 ;
        RECT 0.860 294.820 157.620 295.420 ;
        RECT 0.090 294.260 157.620 294.820 ;
        RECT 0.090 293.740 158.340 294.260 ;
        RECT 0.860 292.580 158.340 293.740 ;
        RECT 0.090 291.500 158.340 292.580 ;
        RECT 0.860 290.340 158.340 291.500 ;
        RECT 0.090 289.820 158.340 290.340 ;
        RECT 0.090 289.260 157.620 289.820 ;
        RECT 0.860 288.660 157.620 289.260 ;
        RECT 0.860 288.100 158.340 288.660 ;
        RECT 0.090 286.460 158.340 288.100 ;
        RECT 0.860 285.300 158.340 286.460 ;
        RECT 0.090 284.220 158.340 285.300 ;
        RECT 0.860 283.060 157.620 284.220 ;
        RECT 0.090 281.980 158.340 283.060 ;
        RECT 0.860 280.820 158.340 281.980 ;
        RECT 0.090 279.740 158.340 280.820 ;
        RECT 0.860 278.620 158.340 279.740 ;
        RECT 0.860 278.580 157.620 278.620 ;
        RECT 0.090 277.500 157.620 278.580 ;
        RECT 0.860 277.460 157.620 277.500 ;
        RECT 0.860 276.340 158.340 277.460 ;
        RECT 0.090 275.260 158.340 276.340 ;
        RECT 0.860 274.100 158.340 275.260 ;
        RECT 0.090 273.020 158.340 274.100 ;
        RECT 0.860 271.860 157.620 273.020 ;
        RECT 0.090 270.780 158.340 271.860 ;
        RECT 0.860 269.620 158.340 270.780 ;
        RECT 0.090 268.540 158.340 269.620 ;
        RECT 0.860 267.420 158.340 268.540 ;
        RECT 0.860 267.380 157.620 267.420 ;
        RECT 0.090 266.300 157.620 267.380 ;
        RECT 0.860 266.260 157.620 266.300 ;
        RECT 0.860 265.140 158.340 266.260 ;
        RECT 0.090 264.060 158.340 265.140 ;
        RECT 0.860 262.900 158.340 264.060 ;
        RECT 0.090 261.820 158.340 262.900 ;
        RECT 0.860 260.660 157.620 261.820 ;
        RECT 0.090 259.580 158.340 260.660 ;
        RECT 0.860 258.420 158.340 259.580 ;
        RECT 0.090 257.340 158.340 258.420 ;
        RECT 0.860 256.220 158.340 257.340 ;
        RECT 0.860 256.180 157.620 256.220 ;
        RECT 0.090 255.100 157.620 256.180 ;
        RECT 0.860 255.060 157.620 255.100 ;
        RECT 0.860 253.940 158.340 255.060 ;
        RECT 0.090 252.860 158.340 253.940 ;
        RECT 0.860 251.700 158.340 252.860 ;
        RECT 0.090 250.620 158.340 251.700 ;
        RECT 0.860 249.460 157.620 250.620 ;
        RECT 0.090 248.380 158.340 249.460 ;
        RECT 0.860 247.220 158.340 248.380 ;
        RECT 0.090 246.140 158.340 247.220 ;
        RECT 0.860 245.020 158.340 246.140 ;
        RECT 0.860 244.980 157.620 245.020 ;
        RECT 0.090 243.900 157.620 244.980 ;
        RECT 0.860 243.860 157.620 243.900 ;
        RECT 0.860 242.740 158.340 243.860 ;
        RECT 0.090 241.660 158.340 242.740 ;
        RECT 0.860 240.500 158.340 241.660 ;
        RECT 0.090 239.420 158.340 240.500 ;
        RECT 0.860 238.260 157.620 239.420 ;
        RECT 0.090 237.180 158.340 238.260 ;
        RECT 0.860 236.020 158.340 237.180 ;
        RECT 0.090 234.940 158.340 236.020 ;
        RECT 0.860 233.820 158.340 234.940 ;
        RECT 0.860 233.780 157.620 233.820 ;
        RECT 0.090 232.700 157.620 233.780 ;
        RECT 0.860 232.660 157.620 232.700 ;
        RECT 0.860 231.540 158.340 232.660 ;
        RECT 0.090 230.460 158.340 231.540 ;
        RECT 0.860 229.300 158.340 230.460 ;
        RECT 0.090 228.220 158.340 229.300 ;
        RECT 0.860 227.060 157.620 228.220 ;
        RECT 0.090 225.980 158.340 227.060 ;
        RECT 0.860 224.820 158.340 225.980 ;
        RECT 0.090 223.740 158.340 224.820 ;
        RECT 0.860 222.620 158.340 223.740 ;
        RECT 0.860 222.580 157.620 222.620 ;
        RECT 0.090 221.500 157.620 222.580 ;
        RECT 0.860 221.460 157.620 221.500 ;
        RECT 0.860 220.340 158.340 221.460 ;
        RECT 0.090 219.260 158.340 220.340 ;
        RECT 0.860 218.100 158.340 219.260 ;
        RECT 0.090 217.020 158.340 218.100 ;
        RECT 0.860 215.860 157.620 217.020 ;
        RECT 0.090 214.780 158.340 215.860 ;
        RECT 0.860 213.620 158.340 214.780 ;
        RECT 0.090 212.540 158.340 213.620 ;
        RECT 0.860 211.420 158.340 212.540 ;
        RECT 0.860 211.380 157.620 211.420 ;
        RECT 0.090 210.300 157.620 211.380 ;
        RECT 0.860 210.260 157.620 210.300 ;
        RECT 0.860 209.140 158.340 210.260 ;
        RECT 0.090 208.060 158.340 209.140 ;
        RECT 0.860 206.900 158.340 208.060 ;
        RECT 0.090 205.820 158.340 206.900 ;
        RECT 0.860 204.660 157.620 205.820 ;
        RECT 0.090 203.580 158.340 204.660 ;
        RECT 0.860 202.420 158.340 203.580 ;
        RECT 0.090 201.340 158.340 202.420 ;
        RECT 0.860 200.220 158.340 201.340 ;
        RECT 0.860 200.180 157.620 200.220 ;
        RECT 0.090 199.100 157.620 200.180 ;
        RECT 0.860 199.060 157.620 199.100 ;
        RECT 0.860 197.940 158.340 199.060 ;
        RECT 0.090 196.860 158.340 197.940 ;
        RECT 0.860 195.700 158.340 196.860 ;
        RECT 0.090 194.620 158.340 195.700 ;
        RECT 0.860 193.460 158.340 194.620 ;
        RECT 0.090 192.380 158.340 193.460 ;
        RECT 0.860 191.220 158.340 192.380 ;
        RECT 0.090 190.140 158.340 191.220 ;
        RECT 0.860 188.980 158.340 190.140 ;
        RECT 0.090 187.900 158.340 188.980 ;
        RECT 0.860 186.740 158.340 187.900 ;
        RECT 0.090 185.660 158.340 186.740 ;
        RECT 0.860 184.500 158.340 185.660 ;
        RECT 0.090 183.420 158.340 184.500 ;
        RECT 0.860 182.260 158.340 183.420 ;
        RECT 0.090 181.180 158.340 182.260 ;
        RECT 0.860 180.020 158.340 181.180 ;
        RECT 0.090 178.940 158.340 180.020 ;
        RECT 0.860 177.780 158.340 178.940 ;
        RECT 0.090 176.700 158.340 177.780 ;
        RECT 0.860 175.540 157.620 176.700 ;
        RECT 0.090 174.460 158.340 175.540 ;
        RECT 0.860 173.300 158.340 174.460 ;
        RECT 0.090 172.220 158.340 173.300 ;
        RECT 0.860 171.060 157.620 172.220 ;
        RECT 0.090 169.980 158.340 171.060 ;
        RECT 0.860 168.820 158.340 169.980 ;
        RECT 0.090 167.740 158.340 168.820 ;
        RECT 0.860 166.580 157.620 167.740 ;
        RECT 0.090 165.500 158.340 166.580 ;
        RECT 0.860 164.340 158.340 165.500 ;
        RECT 0.090 163.260 158.340 164.340 ;
        RECT 0.860 162.100 157.620 163.260 ;
        RECT 0.090 161.020 158.340 162.100 ;
        RECT 0.860 159.860 158.340 161.020 ;
        RECT 0.090 158.780 158.340 159.860 ;
        RECT 0.860 157.620 157.620 158.780 ;
        RECT 0.090 156.540 158.340 157.620 ;
        RECT 0.860 155.380 158.340 156.540 ;
        RECT 0.090 154.300 158.340 155.380 ;
        RECT 0.860 153.140 157.620 154.300 ;
        RECT 0.090 152.060 158.340 153.140 ;
        RECT 0.860 150.900 158.340 152.060 ;
        RECT 0.090 149.820 158.340 150.900 ;
        RECT 0.860 148.660 157.620 149.820 ;
        RECT 0.090 147.580 158.340 148.660 ;
        RECT 0.860 146.420 158.340 147.580 ;
        RECT 0.090 145.340 158.340 146.420 ;
        RECT 0.860 144.180 157.620 145.340 ;
        RECT 0.090 143.100 158.340 144.180 ;
        RECT 0.860 141.940 158.340 143.100 ;
        RECT 0.090 140.860 158.340 141.940 ;
        RECT 0.860 139.700 157.620 140.860 ;
        RECT 0.090 138.620 158.340 139.700 ;
        RECT 0.860 137.460 158.340 138.620 ;
        RECT 0.090 136.380 158.340 137.460 ;
        RECT 0.860 135.220 157.620 136.380 ;
        RECT 0.090 134.140 158.340 135.220 ;
        RECT 0.860 132.980 158.340 134.140 ;
        RECT 0.090 131.900 158.340 132.980 ;
        RECT 0.860 130.740 157.620 131.900 ;
        RECT 0.090 129.660 158.340 130.740 ;
        RECT 0.860 128.500 158.340 129.660 ;
        RECT 0.090 127.420 158.340 128.500 ;
        RECT 0.860 126.260 157.620 127.420 ;
        RECT 0.090 125.180 158.340 126.260 ;
        RECT 0.860 124.020 158.340 125.180 ;
        RECT 0.090 122.940 158.340 124.020 ;
        RECT 0.860 121.780 157.620 122.940 ;
        RECT 0.090 120.700 158.340 121.780 ;
        RECT 0.860 119.540 158.340 120.700 ;
        RECT 0.090 118.460 158.340 119.540 ;
        RECT 0.860 117.300 157.620 118.460 ;
        RECT 0.090 116.220 158.340 117.300 ;
        RECT 0.860 115.060 158.340 116.220 ;
        RECT 0.090 113.980 158.340 115.060 ;
        RECT 0.860 112.820 157.620 113.980 ;
        RECT 0.090 111.740 158.340 112.820 ;
        RECT 0.860 110.580 158.340 111.740 ;
        RECT 0.090 109.500 158.340 110.580 ;
        RECT 0.860 108.340 157.620 109.500 ;
        RECT 0.090 107.260 158.340 108.340 ;
        RECT 0.860 106.100 158.340 107.260 ;
        RECT 0.090 105.020 158.340 106.100 ;
        RECT 0.860 103.860 157.620 105.020 ;
        RECT 0.090 102.780 158.340 103.860 ;
        RECT 0.860 101.620 158.340 102.780 ;
        RECT 0.090 100.540 158.340 101.620 ;
        RECT 0.860 99.380 157.620 100.540 ;
        RECT 0.090 98.300 158.340 99.380 ;
        RECT 0.860 97.140 158.340 98.300 ;
        RECT 0.090 96.060 158.340 97.140 ;
        RECT 0.860 94.900 157.620 96.060 ;
        RECT 0.090 93.820 158.340 94.900 ;
        RECT 0.860 92.660 158.340 93.820 ;
        RECT 0.090 91.580 158.340 92.660 ;
        RECT 0.860 90.420 157.620 91.580 ;
        RECT 0.090 89.340 158.340 90.420 ;
        RECT 0.860 88.180 158.340 89.340 ;
        RECT 0.090 87.100 158.340 88.180 ;
        RECT 0.860 85.940 157.620 87.100 ;
        RECT 0.090 84.860 158.340 85.940 ;
        RECT 0.860 83.700 158.340 84.860 ;
        RECT 0.090 82.620 158.340 83.700 ;
        RECT 0.860 81.460 157.620 82.620 ;
        RECT 0.090 80.380 158.340 81.460 ;
        RECT 0.860 79.220 158.340 80.380 ;
        RECT 0.090 78.140 158.340 79.220 ;
        RECT 0.860 76.980 157.620 78.140 ;
        RECT 0.090 75.900 158.340 76.980 ;
        RECT 0.860 74.740 158.340 75.900 ;
        RECT 0.090 73.660 158.340 74.740 ;
        RECT 0.860 72.500 157.620 73.660 ;
        RECT 0.090 71.420 158.340 72.500 ;
        RECT 0.860 70.260 158.340 71.420 ;
        RECT 0.090 69.180 158.340 70.260 ;
        RECT 0.860 68.020 157.620 69.180 ;
        RECT 0.090 66.940 158.340 68.020 ;
        RECT 0.860 65.780 158.340 66.940 ;
        RECT 0.090 64.700 158.340 65.780 ;
        RECT 0.860 63.540 157.620 64.700 ;
        RECT 0.090 62.460 158.340 63.540 ;
        RECT 0.860 61.300 158.340 62.460 ;
        RECT 0.090 60.220 158.340 61.300 ;
        RECT 0.860 59.060 157.620 60.220 ;
        RECT 0.090 57.980 158.340 59.060 ;
        RECT 0.860 56.820 158.340 57.980 ;
        RECT 0.090 55.740 158.340 56.820 ;
        RECT 0.860 54.580 157.620 55.740 ;
        RECT 0.090 53.500 158.340 54.580 ;
        RECT 0.860 52.340 158.340 53.500 ;
        RECT 0.090 51.260 158.340 52.340 ;
        RECT 0.860 50.100 157.620 51.260 ;
        RECT 0.090 49.020 158.340 50.100 ;
        RECT 0.860 47.860 158.340 49.020 ;
        RECT 0.090 46.780 158.340 47.860 ;
        RECT 0.860 45.620 157.620 46.780 ;
        RECT 0.090 44.540 158.340 45.620 ;
        RECT 0.860 43.380 158.340 44.540 ;
        RECT 0.090 42.300 158.340 43.380 ;
        RECT 0.860 41.140 157.620 42.300 ;
        RECT 0.090 40.060 158.340 41.140 ;
        RECT 0.860 38.900 158.340 40.060 ;
        RECT 0.090 37.820 158.340 38.900 ;
        RECT 0.860 36.660 157.620 37.820 ;
        RECT 0.090 35.580 158.340 36.660 ;
        RECT 0.860 34.420 158.340 35.580 ;
        RECT 0.090 33.340 158.340 34.420 ;
        RECT 0.860 32.180 157.620 33.340 ;
        RECT 0.090 31.100 158.340 32.180 ;
        RECT 0.860 29.940 158.340 31.100 ;
        RECT 0.090 28.860 158.340 29.940 ;
        RECT 0.860 27.700 157.620 28.860 ;
        RECT 0.090 26.620 158.340 27.700 ;
        RECT 0.860 25.460 158.340 26.620 ;
        RECT 0.090 24.380 158.340 25.460 ;
        RECT 0.860 23.220 157.620 24.380 ;
        RECT 0.090 22.140 158.340 23.220 ;
        RECT 0.860 20.980 158.340 22.140 ;
        RECT 0.090 19.900 158.340 20.980 ;
        RECT 0.860 18.740 157.620 19.900 ;
        RECT 0.090 17.660 158.340 18.740 ;
        RECT 0.860 16.500 158.340 17.660 ;
        RECT 0.090 15.420 158.340 16.500 ;
        RECT 0.860 14.260 157.620 15.420 ;
        RECT 0.090 13.180 158.340 14.260 ;
        RECT 0.860 12.020 158.340 13.180 ;
        RECT 0.090 10.940 158.340 12.020 ;
        RECT 0.860 9.780 158.340 10.940 ;
        RECT 0.090 8.700 158.340 9.780 ;
        RECT 0.860 7.540 158.340 8.700 ;
        RECT 0.090 6.460 158.340 7.540 ;
        RECT 0.860 5.300 158.340 6.460 ;
        RECT 0.090 4.220 158.340 5.300 ;
        RECT 0.860 3.060 158.340 4.220 ;
        RECT 0.090 1.980 158.340 3.060 ;
        RECT 0.860 0.820 158.340 1.980 ;
        RECT 0.090 0.140 158.340 0.820 ;
      LAYER Metal4 ;
        RECT 0.700 0.090 18.580 573.350 ;
        RECT 20.780 0.090 21.880 573.350 ;
        RECT 24.080 0.090 118.580 573.350 ;
        RECT 120.780 0.090 121.880 573.350 ;
        RECT 124.080 0.090 143.220 573.350 ;
  END
END GF_SRAM
END LIBRARY

