magic
tech gf180mcuD
magscale 1 10
timestamp 1764323266
<< metal1 >>
rect 672 56474 56784 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 43806 56474
rect 43858 56422 43910 56474
rect 43962 56422 44014 56474
rect 44066 56422 56784 56474
rect 672 56388 56784 56422
rect 8094 56194 8146 56206
rect 8094 56130 8146 56142
rect 7982 56082 8034 56094
rect 21646 56082 21698 56094
rect 3378 56030 3390 56082
rect 3442 56030 3454 56082
rect 6738 56030 6750 56082
rect 6802 56030 6814 56082
rect 7410 56030 7422 56082
rect 7474 56030 7486 56082
rect 9874 56030 9886 56082
rect 9938 56030 9950 56082
rect 13234 56030 13246 56082
rect 13298 56030 13310 56082
rect 14018 56030 14030 56082
rect 14082 56030 14094 56082
rect 17378 56030 17390 56082
rect 17442 56030 17454 56082
rect 17938 56030 17950 56082
rect 18002 56030 18014 56082
rect 19282 56030 19294 56082
rect 19346 56030 19358 56082
rect 20626 56030 20638 56082
rect 20690 56030 20702 56082
rect 7982 56018 8034 56030
rect 21646 56018 21698 56030
rect 24558 56082 24610 56094
rect 30606 56082 30658 56094
rect 36430 56082 36482 56094
rect 38446 56082 38498 56094
rect 25106 56030 25118 56082
rect 25170 56030 25182 56082
rect 26898 56030 26910 56082
rect 26962 56030 26974 56082
rect 28690 56030 28702 56082
rect 28754 56030 28766 56082
rect 33170 56030 33182 56082
rect 33234 56030 33246 56082
rect 34514 56030 34526 56082
rect 34578 56030 34590 56082
rect 35522 56030 35534 56082
rect 35586 56030 35598 56082
rect 36866 56030 36878 56082
rect 36930 56030 36942 56082
rect 37538 56030 37550 56082
rect 37602 56030 37614 56082
rect 24558 56018 24610 56030
rect 30606 56018 30658 56030
rect 36430 56018 36482 56030
rect 38446 56018 38498 56030
rect 39454 56082 39506 56094
rect 43822 56082 43874 56094
rect 42130 56030 42142 56082
rect 42194 56030 42206 56082
rect 43250 56030 43262 56082
rect 43314 56030 43326 56082
rect 39454 56018 39506 56030
rect 43822 56018 43874 56030
rect 45166 56082 45218 56094
rect 45166 56018 45218 56030
rect 45838 56082 45890 56094
rect 55022 56082 55074 56094
rect 54562 56030 54574 56082
rect 54626 56030 54638 56082
rect 45838 56018 45890 56030
rect 55022 56018 55074 56030
rect 3950 55970 4002 55982
rect 2258 55918 2270 55970
rect 2322 55918 2334 55970
rect 3602 55918 3614 55970
rect 3666 55918 3678 55970
rect 3950 55906 4002 55918
rect 4846 55970 4898 55982
rect 21982 55970 22034 55982
rect 25790 55970 25842 55982
rect 53566 55970 53618 55982
rect 6290 55918 6302 55970
rect 6354 55918 6366 55970
rect 10098 55918 10110 55970
rect 10162 55918 10174 55970
rect 10770 55918 10782 55970
rect 10834 55918 10846 55970
rect 11890 55918 11902 55970
rect 11954 55918 11966 55970
rect 13458 55918 13470 55970
rect 13522 55918 13534 55970
rect 14354 55918 14366 55970
rect 14418 55918 14430 55970
rect 16818 55918 16830 55970
rect 16882 55918 16894 55970
rect 18162 55918 18174 55970
rect 18226 55918 18238 55970
rect 18834 55918 18846 55970
rect 18898 55918 18910 55970
rect 20402 55918 20414 55970
rect 20466 55918 20478 55970
rect 22642 55918 22654 55970
rect 22706 55918 22718 55970
rect 23314 55918 23326 55970
rect 23378 55918 23390 55970
rect 24210 55918 24222 55970
rect 24274 55918 24286 55970
rect 24882 55918 24894 55970
rect 24946 55918 24958 55970
rect 28242 55918 28254 55970
rect 28306 55918 28318 55970
rect 29922 55918 29934 55970
rect 29986 55918 29998 55970
rect 32722 55918 32734 55970
rect 32786 55918 32798 55970
rect 41010 55918 41022 55970
rect 41074 55918 41086 55970
rect 43474 55918 43486 55970
rect 43538 55918 43550 55970
rect 44146 55918 44158 55970
rect 44210 55918 44222 55970
rect 46162 55918 46174 55970
rect 46226 55918 46238 55970
rect 47058 55918 47070 55970
rect 47122 55918 47134 55970
rect 47730 55918 47742 55970
rect 47794 55918 47806 55970
rect 49074 55918 49086 55970
rect 49138 55918 49150 55970
rect 49746 55918 49758 55970
rect 49810 55918 49822 55970
rect 50530 55918 50542 55970
rect 50594 55918 50606 55970
rect 51874 55918 51886 55970
rect 51938 55918 51950 55970
rect 52546 55918 52558 55970
rect 52610 55918 52622 55970
rect 53218 55918 53230 55970
rect 53282 55918 53294 55970
rect 4846 55906 4898 55918
rect 21982 55906 22034 55918
rect 25790 55906 25842 55918
rect 53566 55906 53618 55918
rect 1262 55858 1314 55870
rect 1934 55858 1986 55870
rect 1586 55806 1598 55858
rect 1650 55806 1662 55858
rect 1262 55794 1314 55806
rect 1934 55794 1986 55806
rect 2606 55858 2658 55870
rect 4958 55858 5010 55870
rect 2930 55806 2942 55858
rect 2994 55806 3006 55858
rect 4274 55806 4286 55858
rect 4338 55806 4350 55858
rect 2606 55794 2658 55806
rect 4958 55794 5010 55806
rect 5294 55858 5346 55870
rect 5966 55858 6018 55870
rect 9102 55858 9154 55870
rect 5618 55806 5630 55858
rect 5682 55806 5694 55858
rect 6962 55806 6974 55858
rect 7026 55806 7038 55858
rect 7634 55806 7646 55858
rect 7698 55806 7710 55858
rect 5294 55794 5346 55806
rect 5966 55794 6018 55806
rect 9102 55794 9154 55806
rect 10446 55858 10498 55870
rect 10446 55794 10498 55806
rect 11118 55858 11170 55870
rect 11118 55794 11170 55806
rect 11566 55858 11618 55870
rect 11566 55794 11618 55806
rect 12462 55858 12514 55870
rect 12462 55794 12514 55806
rect 15598 55858 15650 55870
rect 15598 55794 15650 55806
rect 16494 55858 16546 55870
rect 18510 55858 18562 55870
rect 20190 55858 20242 55870
rect 17154 55806 17166 55858
rect 17218 55806 17230 55858
rect 19506 55806 19518 55858
rect 19570 55806 19582 55858
rect 16494 55794 16546 55806
rect 18510 55794 18562 55806
rect 20190 55794 20242 55806
rect 21534 55858 21586 55870
rect 21534 55794 21586 55806
rect 21870 55858 21922 55870
rect 21870 55794 21922 55806
rect 22318 55858 22370 55870
rect 22318 55794 22370 55806
rect 22990 55858 23042 55870
rect 22990 55794 23042 55806
rect 25454 55858 25506 55870
rect 25454 55794 25506 55806
rect 25678 55858 25730 55870
rect 25678 55794 25730 55806
rect 26126 55858 26178 55870
rect 27918 55858 27970 55870
rect 29262 55858 29314 55870
rect 30270 55858 30322 55870
rect 31726 55858 31778 55870
rect 32398 55858 32450 55870
rect 33742 55858 33794 55870
rect 40014 55858 40066 55870
rect 40686 55858 40738 55870
rect 26450 55806 26462 55858
rect 26514 55806 26526 55858
rect 27122 55806 27134 55858
rect 27186 55806 27198 55858
rect 28914 55806 28926 55858
rect 28978 55806 28990 55858
rect 29586 55806 29598 55858
rect 29650 55806 29662 55858
rect 30930 55806 30942 55858
rect 30994 55806 31006 55858
rect 32050 55806 32062 55858
rect 32114 55806 32126 55858
rect 33394 55806 33406 55858
rect 33458 55806 33470 55858
rect 34066 55806 34078 55858
rect 34130 55806 34142 55858
rect 34738 55806 34750 55858
rect 34802 55806 34814 55858
rect 35746 55806 35758 55858
rect 35810 55806 35822 55858
rect 36082 55806 36094 55858
rect 36146 55806 36158 55858
rect 37090 55806 37102 55858
rect 37154 55806 37166 55858
rect 37762 55806 37774 55858
rect 37826 55806 37838 55858
rect 38098 55806 38110 55858
rect 38162 55806 38174 55858
rect 39106 55806 39118 55858
rect 39170 55806 39182 55858
rect 40338 55806 40350 55858
rect 40402 55806 40414 55858
rect 26126 55794 26178 55806
rect 27918 55794 27970 55806
rect 29262 55794 29314 55806
rect 30270 55794 30322 55806
rect 31726 55794 31778 55806
rect 32398 55794 32450 55806
rect 33742 55794 33794 55806
rect 40014 55794 40066 55806
rect 40686 55794 40738 55806
rect 41358 55858 41410 55870
rect 44830 55858 44882 55870
rect 46734 55858 46786 55870
rect 41682 55806 41694 55858
rect 41746 55806 41758 55858
rect 42354 55806 42366 55858
rect 42418 55806 42430 55858
rect 44482 55806 44494 55858
rect 44546 55806 44558 55858
rect 45490 55806 45502 55858
rect 45554 55806 45566 55858
rect 41358 55794 41410 55806
rect 44830 55794 44882 55806
rect 46734 55794 46786 55806
rect 47406 55858 47458 55870
rect 47406 55794 47458 55806
rect 48078 55858 48130 55870
rect 48750 55858 48802 55870
rect 48402 55806 48414 55858
rect 48466 55806 48478 55858
rect 48078 55794 48130 55806
rect 48750 55794 48802 55806
rect 49422 55858 49474 55870
rect 49422 55794 49474 55806
rect 50878 55858 50930 55870
rect 51550 55858 51602 55870
rect 51202 55806 51214 55858
rect 51266 55806 51278 55858
rect 50878 55794 50930 55806
rect 51550 55794 51602 55806
rect 52222 55858 52274 55870
rect 52222 55794 52274 55806
rect 52894 55858 52946 55870
rect 56030 55858 56082 55870
rect 54338 55806 54350 55858
rect 54402 55806 54414 55858
rect 55346 55806 55358 55858
rect 55410 55806 55422 55858
rect 55682 55806 55694 55858
rect 55746 55806 55758 55858
rect 52894 55794 52946 55806
rect 56030 55794 56082 55806
rect 56254 55858 56306 55870
rect 56254 55794 56306 55806
rect 672 55690 56784 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 44466 55690
rect 44518 55638 44570 55690
rect 44622 55638 44674 55690
rect 44726 55638 56784 55690
rect 672 55604 56784 55638
rect 20190 55522 20242 55534
rect 38558 55522 38610 55534
rect 7298 55470 7310 55522
rect 7362 55470 7374 55522
rect 20514 55470 20526 55522
rect 20578 55470 20590 55522
rect 22194 55470 22206 55522
rect 22258 55470 22270 55522
rect 20190 55458 20242 55470
rect 38558 55458 38610 55470
rect 39230 55522 39282 55534
rect 39230 55458 39282 55470
rect 40238 55522 40290 55534
rect 43474 55470 43486 55522
rect 43538 55470 43550 55522
rect 40238 55458 40290 55470
rect 3390 55410 3442 55422
rect 1698 55358 1710 55410
rect 1762 55358 1774 55410
rect 3390 55346 3442 55358
rect 3502 55410 3554 55422
rect 6190 55410 6242 55422
rect 13470 55410 13522 55422
rect 17502 55410 17554 55422
rect 29038 55410 29090 55422
rect 31502 55410 31554 55422
rect 35982 55410 36034 55422
rect 41134 55410 41186 55422
rect 4498 55358 4510 55410
rect 4562 55358 4574 55410
rect 6962 55358 6974 55410
rect 7026 55358 7038 55410
rect 8306 55358 8318 55410
rect 8370 55358 8382 55410
rect 9426 55358 9438 55410
rect 9490 55358 9502 55410
rect 9762 55358 9774 55410
rect 9826 55358 9838 55410
rect 10770 55358 10782 55410
rect 10834 55358 10846 55410
rect 11106 55358 11118 55410
rect 11170 55358 11182 55410
rect 12114 55358 12126 55410
rect 12178 55358 12190 55410
rect 12450 55358 12462 55410
rect 12514 55358 12526 55410
rect 14466 55358 14478 55410
rect 14530 55358 14542 55410
rect 15474 55358 15486 55410
rect 15538 55358 15550 55410
rect 15810 55358 15822 55410
rect 15874 55358 15886 55410
rect 17826 55358 17838 55410
rect 17890 55358 17902 55410
rect 18498 55358 18510 55410
rect 18562 55358 18574 55410
rect 19170 55358 19182 55410
rect 19234 55358 19246 55410
rect 19506 55358 19518 55410
rect 19570 55358 19582 55410
rect 20850 55358 20862 55410
rect 20914 55358 20926 55410
rect 21522 55358 21534 55410
rect 21586 55358 21598 55410
rect 22866 55358 22878 55410
rect 22930 55358 22942 55410
rect 23538 55358 23550 55410
rect 23602 55358 23614 55410
rect 24546 55358 24558 55410
rect 24610 55358 24622 55410
rect 25330 55358 25342 55410
rect 25394 55358 25406 55410
rect 26562 55358 26574 55410
rect 26626 55358 26638 55410
rect 27234 55358 27246 55410
rect 27298 55358 27310 55410
rect 27906 55358 27918 55410
rect 27970 55358 27982 55410
rect 28242 55358 28254 55410
rect 28306 55358 28318 55410
rect 29810 55358 29822 55410
rect 29874 55358 29886 55410
rect 30482 55358 30494 55410
rect 30546 55358 30558 55410
rect 30818 55358 30830 55410
rect 30882 55358 30894 55410
rect 31826 55358 31838 55410
rect 31890 55358 31902 55410
rect 33170 55358 33182 55410
rect 33234 55358 33246 55410
rect 33842 55358 33854 55410
rect 33906 55358 33918 55410
rect 35634 55358 35646 55410
rect 35698 55358 35710 55410
rect 36306 55358 36318 55410
rect 36370 55358 36382 55410
rect 37202 55358 37214 55410
rect 37266 55358 37278 55410
rect 37538 55358 37550 55410
rect 37602 55358 37614 55410
rect 38882 55358 38894 55410
rect 38946 55358 38958 55410
rect 39554 55358 39566 55410
rect 39618 55358 39630 55410
rect 40562 55358 40574 55410
rect 40626 55358 40638 55410
rect 41458 55358 41470 55410
rect 41522 55358 41534 55410
rect 42130 55358 42142 55410
rect 42194 55358 42206 55410
rect 42802 55358 42814 55410
rect 42866 55358 42878 55410
rect 43810 55358 43822 55410
rect 43874 55358 43886 55410
rect 44482 55358 44494 55410
rect 44546 55358 44558 55410
rect 45154 55358 45166 55410
rect 45218 55358 45230 55410
rect 46050 55358 46062 55410
rect 46114 55358 46126 55410
rect 46722 55358 46734 55410
rect 46786 55358 46798 55410
rect 53666 55358 53678 55410
rect 53730 55358 53742 55410
rect 54674 55358 54686 55410
rect 54738 55358 54750 55410
rect 55906 55358 55918 55410
rect 55970 55358 55982 55410
rect 3502 55346 3554 55358
rect 6190 55346 6242 55358
rect 13470 55346 13522 55358
rect 17502 55346 17554 55358
rect 29038 55346 29090 55358
rect 31502 55346 31554 55358
rect 35982 55346 36034 55358
rect 41134 55346 41186 55358
rect 3166 55298 3218 55310
rect 3166 55234 3218 55246
rect 6078 55298 6130 55310
rect 6078 55234 6130 55246
rect 6414 55298 6466 55310
rect 6414 55234 6466 55246
rect 6638 55298 6690 55310
rect 6638 55234 6690 55246
rect 7646 55298 7698 55310
rect 9102 55298 9154 55310
rect 10446 55298 10498 55310
rect 8082 55246 8094 55298
rect 8146 55246 8158 55298
rect 9986 55246 9998 55298
rect 10050 55246 10062 55298
rect 7646 55234 7698 55246
rect 9102 55234 9154 55246
rect 10446 55234 10498 55246
rect 11454 55298 11506 55310
rect 12798 55298 12850 55310
rect 11890 55246 11902 55298
rect 11954 55246 11966 55298
rect 11454 55234 11506 55246
rect 12798 55234 12850 55246
rect 13022 55298 13074 55310
rect 13022 55234 13074 55246
rect 13582 55298 13634 55310
rect 15150 55298 15202 55310
rect 14690 55246 14702 55298
rect 14754 55246 14766 55298
rect 13582 55234 13634 55246
rect 15150 55234 15202 55246
rect 16158 55298 16210 55310
rect 22542 55298 22594 55310
rect 25678 55298 25730 55310
rect 26910 55298 26962 55310
rect 18274 55246 18286 55298
rect 18338 55246 18350 55298
rect 18946 55246 18958 55298
rect 19010 55246 19022 55298
rect 19730 55246 19742 55298
rect 19794 55246 19806 55298
rect 20290 55246 20302 55298
rect 20354 55246 20366 55298
rect 21074 55246 21086 55298
rect 21138 55246 21150 55298
rect 21746 55246 21758 55298
rect 21810 55246 21822 55298
rect 23090 55246 23102 55298
rect 23154 55246 23166 55298
rect 23762 55246 23774 55298
rect 23826 55246 23838 55298
rect 24770 55246 24782 55298
rect 24834 55246 24846 55298
rect 26338 55246 26350 55298
rect 26402 55246 26414 55298
rect 16158 55234 16210 55246
rect 22542 55234 22594 55246
rect 25678 55234 25730 55246
rect 26910 55234 26962 55246
rect 27582 55298 27634 55310
rect 27582 55234 27634 55246
rect 28590 55298 28642 55310
rect 28590 55234 28642 55246
rect 28926 55298 28978 55310
rect 31166 55298 31218 55310
rect 29586 55246 29598 55298
rect 29650 55246 29662 55298
rect 30258 55246 30270 55298
rect 30322 55246 30334 55298
rect 28926 55234 28978 55246
rect 31166 55234 31218 55246
rect 32510 55298 32562 55310
rect 34638 55298 34690 55310
rect 32946 55246 32958 55298
rect 33010 55246 33022 55298
rect 33618 55246 33630 55298
rect 33682 55246 33694 55298
rect 34514 55246 34526 55298
rect 34578 55246 34590 55298
rect 32510 55234 32562 55246
rect 34638 55234 34690 55246
rect 34750 55298 34802 55310
rect 34750 55234 34802 55246
rect 34862 55298 34914 55310
rect 43150 55298 43202 55310
rect 35410 55246 35422 55298
rect 35474 55246 35486 55298
rect 41906 55246 41918 55298
rect 41970 55246 41982 55298
rect 42578 55246 42590 55298
rect 42642 55246 42654 55298
rect 34862 55234 34914 55246
rect 43150 55234 43202 55246
rect 44158 55298 44210 55310
rect 44158 55234 44210 55246
rect 44830 55298 44882 55310
rect 46398 55298 46450 55310
rect 54014 55298 54066 55310
rect 56254 55298 56306 55310
rect 45378 55246 45390 55298
rect 45442 55246 45454 55298
rect 46946 55246 46958 55298
rect 47010 55246 47022 55298
rect 48850 55246 48862 55298
rect 48914 55246 48926 55298
rect 54898 55246 54910 55298
rect 54962 55246 54974 55298
rect 44830 55234 44882 55246
rect 46398 55234 46450 55246
rect 54014 55234 54066 55246
rect 56254 55234 56306 55246
rect 13246 55186 13298 55198
rect 1250 55134 1262 55186
rect 1314 55134 1326 55186
rect 4050 55134 4062 55186
rect 4114 55134 4126 55186
rect 13246 55122 13298 55134
rect 16718 55186 16770 55198
rect 16718 55122 16770 55134
rect 17166 55186 17218 55198
rect 50418 55134 50430 55186
rect 50482 55134 50494 55186
rect 17166 55122 17218 55134
rect 2830 55074 2882 55086
rect 2830 55010 2882 55022
rect 5630 55074 5682 55086
rect 5630 55010 5682 55022
rect 16830 55074 16882 55086
rect 16830 55010 16882 55022
rect 29038 55074 29090 55086
rect 29038 55010 29090 55022
rect 32398 55074 32450 55086
rect 32398 55010 32450 55022
rect 34190 55074 34242 55086
rect 34190 55010 34242 55022
rect 37774 55074 37826 55086
rect 37774 55010 37826 55022
rect 38110 55074 38162 55086
rect 38110 55010 38162 55022
rect 672 54906 56784 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 43806 54906
rect 43858 54854 43910 54906
rect 43962 54854 44014 54906
rect 44066 54854 56784 54906
rect 672 54820 56784 54854
rect 29150 54738 29202 54750
rect 29150 54674 29202 54686
rect 33966 54738 34018 54750
rect 33966 54674 34018 54686
rect 38670 54738 38722 54750
rect 38670 54674 38722 54686
rect 12126 54626 12178 54638
rect 48850 54574 48862 54626
rect 48914 54574 48926 54626
rect 12126 54562 12178 54574
rect 4286 54514 4338 54526
rect 2706 54462 2718 54514
rect 2770 54462 2782 54514
rect 4286 54450 4338 54462
rect 5854 54514 5906 54526
rect 5854 54450 5906 54462
rect 6414 54514 6466 54526
rect 11902 54514 11954 54526
rect 13022 54514 13074 54526
rect 7074 54462 7086 54514
rect 7138 54462 7150 54514
rect 7858 54462 7870 54514
rect 7922 54462 7934 54514
rect 8418 54462 8430 54514
rect 8482 54462 8494 54514
rect 9202 54462 9214 54514
rect 9266 54462 9278 54514
rect 12786 54462 12798 54514
rect 12850 54462 12862 54514
rect 6414 54450 6466 54462
rect 11902 54450 11954 54462
rect 13022 54450 13074 54462
rect 13358 54514 13410 54526
rect 13358 54450 13410 54462
rect 16046 54514 16098 54526
rect 21758 54514 21810 54526
rect 18834 54462 18846 54514
rect 18898 54462 18910 54514
rect 19954 54462 19966 54514
rect 20018 54462 20030 54514
rect 16046 54450 16098 54462
rect 21758 54450 21810 54462
rect 23774 54514 23826 54526
rect 29486 54514 29538 54526
rect 34974 54514 35026 54526
rect 39006 54514 39058 54526
rect 26114 54462 26126 54514
rect 26178 54462 26190 54514
rect 27010 54462 27022 54514
rect 27074 54462 27086 54514
rect 30146 54462 30158 54514
rect 30210 54462 30222 54514
rect 30930 54462 30942 54514
rect 30994 54462 31006 54514
rect 32386 54462 32398 54514
rect 32450 54462 32462 54514
rect 34738 54462 34750 54514
rect 34802 54462 34814 54514
rect 36530 54462 36542 54514
rect 36594 54462 36606 54514
rect 23774 54450 23826 54462
rect 29486 54450 29538 54462
rect 34974 54450 35026 54462
rect 39006 54450 39058 54462
rect 41134 54514 41186 54526
rect 41134 54450 41186 54462
rect 42478 54514 42530 54526
rect 42478 54450 42530 54462
rect 42702 54514 42754 54526
rect 42702 54450 42754 54462
rect 44158 54514 44210 54526
rect 44158 54450 44210 54462
rect 44494 54514 44546 54526
rect 53006 54514 53058 54526
rect 45602 54462 45614 54514
rect 45666 54462 45678 54514
rect 46162 54462 46174 54514
rect 46226 54462 46238 54514
rect 44494 54450 44546 54462
rect 53006 54450 53058 54462
rect 5966 54402 6018 54414
rect 11678 54402 11730 54414
rect 1474 54350 1486 54402
rect 1538 54350 1550 54402
rect 2146 54350 2158 54402
rect 2210 54350 2222 54402
rect 3154 54350 3166 54402
rect 3218 54350 3230 54402
rect 8978 54350 8990 54402
rect 9042 54350 9054 54402
rect 10322 54350 10334 54402
rect 10386 54350 10398 54402
rect 10994 54350 11006 54402
rect 11058 54350 11070 54402
rect 5966 54338 6018 54350
rect 11678 54338 11730 54350
rect 12238 54402 12290 54414
rect 22094 54402 22146 54414
rect 28478 54402 28530 54414
rect 35422 54402 35474 54414
rect 43374 54402 43426 54414
rect 13794 54350 13806 54402
rect 13858 54350 13870 54402
rect 16370 54350 16382 54402
rect 16434 54350 16446 54402
rect 18498 54350 18510 54402
rect 18562 54350 18574 54402
rect 19730 54350 19742 54402
rect 19794 54350 19806 54402
rect 21186 54350 21198 54402
rect 21250 54350 21262 54402
rect 22418 54350 22430 54402
rect 22482 54350 22494 54402
rect 30034 54350 30046 54402
rect 30098 54350 30110 54402
rect 31154 54350 31166 54402
rect 31218 54350 31230 54402
rect 31826 54350 31838 54402
rect 31890 54350 31902 54402
rect 35186 54350 35198 54402
rect 35250 54350 35262 54402
rect 36866 54350 36878 54402
rect 36930 54350 36942 54402
rect 39218 54350 39230 54402
rect 39282 54350 39294 54402
rect 39554 54350 39566 54402
rect 39618 54350 39630 54402
rect 40786 54350 40798 54402
rect 40850 54350 40862 54402
rect 42130 54350 42142 54402
rect 42194 54350 42206 54402
rect 12238 54338 12290 54350
rect 22094 54338 22146 54350
rect 28478 54338 28530 54350
rect 35422 54338 35474 54350
rect 43374 54338 43426 54350
rect 44270 54402 44322 54414
rect 45378 54350 45390 54402
rect 45442 54350 45454 54402
rect 51986 54350 51998 54402
rect 52050 54350 52062 54402
rect 52658 54350 52670 54402
rect 52722 54350 52734 54402
rect 54002 54350 54014 54402
rect 54066 54350 54078 54402
rect 44270 54338 44322 54350
rect 1150 54290 1202 54302
rect 1150 54226 1202 54238
rect 1822 54290 1874 54302
rect 1822 54226 1874 54238
rect 5070 54290 5122 54302
rect 6190 54290 6242 54302
rect 5394 54238 5406 54290
rect 5458 54238 5470 54290
rect 5070 54226 5122 54238
rect 6190 54226 6242 54238
rect 6638 54290 6690 54302
rect 9774 54290 9826 54302
rect 7298 54238 7310 54290
rect 7362 54238 7374 54290
rect 7634 54238 7646 54290
rect 7698 54238 7710 54290
rect 8642 54238 8654 54290
rect 8706 54238 8718 54290
rect 6638 54226 6690 54238
rect 9774 54226 9826 54238
rect 10670 54290 10722 54302
rect 10670 54226 10722 54238
rect 11342 54290 11394 54302
rect 11342 54226 11394 54238
rect 13134 54290 13186 54302
rect 13134 54226 13186 54238
rect 13246 54290 13298 54302
rect 13246 54226 13298 54238
rect 14142 54290 14194 54302
rect 14142 54226 14194 54238
rect 14478 54290 14530 54302
rect 14478 54226 14530 54238
rect 15150 54290 15202 54302
rect 15150 54226 15202 54238
rect 15822 54290 15874 54302
rect 15822 54226 15874 54238
rect 17278 54290 17330 54302
rect 17278 54226 17330 54238
rect 19518 54290 19570 54302
rect 19518 54226 19570 54238
rect 20862 54290 20914 54302
rect 20862 54226 20914 54238
rect 21534 54290 21586 54302
rect 21534 54226 21586 54238
rect 21982 54290 22034 54302
rect 21982 54226 22034 54238
rect 22766 54290 22818 54302
rect 23438 54290 23490 54302
rect 23090 54238 23102 54290
rect 23154 54238 23166 54290
rect 22766 54226 22818 54238
rect 23438 54226 23490 54238
rect 23886 54290 23938 54302
rect 23886 54226 23938 54238
rect 24110 54290 24162 54302
rect 24110 54226 24162 54238
rect 24446 54290 24498 54302
rect 27582 54290 27634 54302
rect 28590 54290 28642 54302
rect 25554 54238 25566 54290
rect 25618 54238 25630 54290
rect 27234 54238 27246 54290
rect 27298 54238 27310 54290
rect 27906 54238 27918 54290
rect 27970 54238 27982 54290
rect 24446 54226 24498 54238
rect 27582 54226 27634 54238
rect 28590 54226 28642 54238
rect 28814 54290 28866 54302
rect 28814 54226 28866 54238
rect 31502 54290 31554 54302
rect 38110 54290 38162 54302
rect 32834 54238 32846 54290
rect 32898 54238 32910 54290
rect 35074 54238 35086 54290
rect 35138 54238 35150 54290
rect 31502 54226 31554 54238
rect 38110 54226 38162 54238
rect 40462 54290 40514 54302
rect 41806 54290 41858 54302
rect 43486 54290 43538 54302
rect 41458 54238 41470 54290
rect 41522 54238 41534 54290
rect 43026 54238 43038 54290
rect 43090 54238 43102 54290
rect 40462 54226 40514 54238
rect 41806 54226 41858 54238
rect 43486 54226 43538 54238
rect 43710 54290 43762 54302
rect 45054 54290 45106 54302
rect 44706 54238 44718 54290
rect 44770 54238 44782 54290
rect 43710 54226 43762 54238
rect 45054 54226 45106 54238
rect 52334 54290 52386 54302
rect 52334 54226 52386 54238
rect 53342 54290 53394 54302
rect 54350 54290 54402 54302
rect 55358 54290 55410 54302
rect 53666 54238 53678 54290
rect 53730 54238 53742 54290
rect 55010 54238 55022 54290
rect 55074 54238 55086 54290
rect 53342 54226 53394 54238
rect 54350 54226 54402 54238
rect 55358 54226 55410 54238
rect 56030 54290 56082 54302
rect 56354 54238 56366 54290
rect 56418 54238 56430 54290
rect 56030 54226 56082 54238
rect 672 54122 56784 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 44466 54122
rect 44518 54070 44570 54122
rect 44622 54070 44674 54122
rect 44726 54070 56784 54122
rect 672 54036 56784 54070
rect 25678 53954 25730 53966
rect 2146 53902 2158 53954
rect 2210 53902 2222 53954
rect 6066 53902 6078 53954
rect 6130 53902 6142 53954
rect 16146 53902 16158 53954
rect 16210 53902 16222 53954
rect 19282 53902 19294 53954
rect 19346 53902 19358 53954
rect 20850 53902 20862 53954
rect 20914 53902 20926 53954
rect 25678 53890 25730 53902
rect 30158 53954 30210 53966
rect 30158 53890 30210 53902
rect 32510 53954 32562 53966
rect 49422 53954 49474 53966
rect 34178 53902 34190 53954
rect 34242 53902 34254 53954
rect 53218 53902 53230 53954
rect 53282 53902 53294 53954
rect 32510 53890 32562 53902
rect 49422 53890 49474 53902
rect 20078 53842 20130 53854
rect 32398 53842 32450 53854
rect 1474 53790 1486 53842
rect 1538 53790 1550 53842
rect 2482 53790 2494 53842
rect 2546 53790 2558 53842
rect 3714 53790 3726 53842
rect 3778 53790 3790 53842
rect 9650 53790 9662 53842
rect 9714 53790 9726 53842
rect 13682 53790 13694 53842
rect 13746 53790 13758 53842
rect 15138 53790 15150 53842
rect 15202 53790 15214 53842
rect 17378 53790 17390 53842
rect 17442 53790 17454 53842
rect 21746 53790 21758 53842
rect 21810 53790 21822 53842
rect 22642 53790 22654 53842
rect 22706 53790 22718 53842
rect 23314 53790 23326 53842
rect 23378 53790 23390 53842
rect 28018 53790 28030 53842
rect 28082 53790 28094 53842
rect 29026 53790 29038 53842
rect 29090 53790 29102 53842
rect 30818 53790 30830 53842
rect 30882 53790 30894 53842
rect 31826 53790 31838 53842
rect 31890 53790 31902 53842
rect 35746 53790 35758 53842
rect 35810 53790 35822 53842
rect 38210 53790 38222 53842
rect 38274 53790 38286 53842
rect 41570 53790 41582 53842
rect 41634 53790 41646 53842
rect 43138 53790 43150 53842
rect 43202 53790 43214 53842
rect 45490 53790 45502 53842
rect 45554 53790 45566 53842
rect 46162 53790 46174 53842
rect 46226 53790 46238 53842
rect 46498 53790 46510 53842
rect 46562 53790 46574 53842
rect 47170 53790 47182 53842
rect 47234 53790 47246 53842
rect 48402 53790 48414 53842
rect 48466 53790 48478 53842
rect 49074 53790 49086 53842
rect 49138 53790 49150 53842
rect 50194 53790 50206 53842
rect 50258 53790 50270 53842
rect 50530 53790 50542 53842
rect 50594 53790 50606 53842
rect 51202 53790 51214 53842
rect 51266 53790 51278 53842
rect 51874 53790 51886 53842
rect 51938 53790 51950 53842
rect 52882 53790 52894 53842
rect 52946 53790 52958 53842
rect 54226 53790 54238 53842
rect 54290 53790 54302 53842
rect 55346 53790 55358 53842
rect 55410 53790 55422 53842
rect 56354 53790 56366 53842
rect 56418 53790 56430 53842
rect 20078 53778 20130 53790
rect 32398 53778 32450 53790
rect 1150 53730 1202 53742
rect 9998 53730 10050 53742
rect 13022 53730 13074 53742
rect 15486 53730 15538 53742
rect 1922 53678 1934 53730
rect 1986 53678 1998 53730
rect 2706 53678 2718 53730
rect 2770 53678 2782 53730
rect 11666 53678 11678 53730
rect 11730 53678 11742 53730
rect 12450 53678 12462 53730
rect 12514 53678 12526 53730
rect 13906 53678 13918 53730
rect 13970 53678 13982 53730
rect 14242 53678 14254 53730
rect 14306 53678 14318 53730
rect 1150 53666 1202 53678
rect 9998 53666 10050 53678
rect 13022 53666 13074 53678
rect 15486 53666 15538 53678
rect 15822 53730 15874 53742
rect 19966 53730 20018 53742
rect 22094 53730 22146 53742
rect 19506 53678 19518 53730
rect 19570 53678 19582 53730
rect 20626 53678 20638 53730
rect 20690 53678 20702 53730
rect 15822 53666 15874 53678
rect 19966 53666 20018 53678
rect 22094 53666 22146 53678
rect 22990 53730 23042 53742
rect 24446 53730 24498 53742
rect 23538 53678 23550 53730
rect 23602 53678 23614 53730
rect 22990 53666 23042 53678
rect 24446 53666 24498 53678
rect 24670 53730 24722 53742
rect 24670 53666 24722 53678
rect 24782 53730 24834 53742
rect 24782 53666 24834 53678
rect 25006 53730 25058 53742
rect 25902 53730 25954 53742
rect 26350 53730 26402 53742
rect 25442 53678 25454 53730
rect 25506 53678 25518 53730
rect 26114 53678 26126 53730
rect 26178 53678 26190 53730
rect 25006 53666 25058 53678
rect 25902 53666 25954 53678
rect 26350 53666 26402 53678
rect 26798 53730 26850 53742
rect 26798 53666 26850 53678
rect 27022 53730 27074 53742
rect 31166 53730 31218 53742
rect 27794 53678 27806 53730
rect 27858 53678 27870 53730
rect 27022 53666 27074 53678
rect 31166 53666 31218 53678
rect 31502 53730 31554 53742
rect 31502 53666 31554 53678
rect 32734 53730 32786 53742
rect 44718 53730 44770 53742
rect 47518 53730 47570 53742
rect 49870 53730 49922 53742
rect 51550 53730 51602 53742
rect 52558 53730 52610 53742
rect 41794 53678 41806 53730
rect 41858 53678 41870 53730
rect 45266 53678 45278 53730
rect 45330 53678 45342 53730
rect 45938 53678 45950 53730
rect 46002 53678 46014 53730
rect 46722 53678 46734 53730
rect 46786 53678 46798 53730
rect 48178 53678 48190 53730
rect 48242 53678 48254 53730
rect 50754 53678 50766 53730
rect 50818 53678 50830 53730
rect 52098 53678 52110 53730
rect 52162 53678 52174 53730
rect 32734 53666 32786 53678
rect 44718 53666 44770 53678
rect 47518 53666 47570 53678
rect 49870 53666 49922 53678
rect 51550 53666 51602 53678
rect 52558 53666 52610 53678
rect 53566 53730 53618 53742
rect 53566 53666 53618 53678
rect 53902 53730 53954 53742
rect 53902 53666 53954 53678
rect 55022 53730 55074 53742
rect 55022 53666 55074 53678
rect 56030 53730 56082 53742
rect 56030 53666 56082 53678
rect 7646 53618 7698 53630
rect 3378 53566 3390 53618
rect 3442 53566 3454 53618
rect 5618 53566 5630 53618
rect 5682 53566 5694 53618
rect 7646 53554 7698 53566
rect 7982 53618 8034 53630
rect 7982 53554 8034 53566
rect 8318 53618 8370 53630
rect 8318 53554 8370 53566
rect 8990 53618 9042 53630
rect 8990 53554 9042 53566
rect 10334 53618 10386 53630
rect 10334 53554 10386 53566
rect 11006 53618 11058 53630
rect 11006 53554 11058 53566
rect 14702 53618 14754 53630
rect 21198 53618 21250 53630
rect 16930 53566 16942 53618
rect 16994 53566 17006 53618
rect 14702 53554 14754 53566
rect 21198 53554 21250 53566
rect 22430 53618 22482 53630
rect 22430 53554 22482 53566
rect 25790 53618 25842 53630
rect 25790 53554 25842 53566
rect 26574 53618 26626 53630
rect 44830 53618 44882 53630
rect 28578 53566 28590 53618
rect 28642 53566 28654 53618
rect 34626 53566 34638 53618
rect 34690 53566 34702 53618
rect 35410 53566 35422 53618
rect 35474 53566 35486 53618
rect 37762 53566 37774 53618
rect 37826 53566 37838 53618
rect 42690 53566 42702 53618
rect 42754 53566 42766 53618
rect 26574 53554 26626 53566
rect 44830 53554 44882 53566
rect 4958 53506 5010 53518
rect 4958 53442 5010 53454
rect 7198 53506 7250 53518
rect 7198 53442 7250 53454
rect 7870 53506 7922 53518
rect 7870 53442 7922 53454
rect 18510 53506 18562 53518
rect 18510 53442 18562 53454
rect 20078 53506 20130 53518
rect 20078 53442 20130 53454
rect 33070 53506 33122 53518
rect 33070 53442 33122 53454
rect 36990 53506 37042 53518
rect 36990 53442 37042 53454
rect 39342 53506 39394 53518
rect 39342 53442 39394 53454
rect 40686 53506 40738 53518
rect 40686 53442 40738 53454
rect 41022 53506 41074 53518
rect 41022 53442 41074 53454
rect 44270 53506 44322 53518
rect 44270 53442 44322 53454
rect 672 53338 56784 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 43806 53338
rect 43858 53286 43910 53338
rect 43962 53286 44014 53338
rect 44066 53286 56784 53338
rect 672 53252 56784 53286
rect 9886 53170 9938 53182
rect 9886 53106 9938 53118
rect 20078 53170 20130 53182
rect 20078 53106 20130 53118
rect 23102 53170 23154 53182
rect 23102 53106 23154 53118
rect 31726 53170 31778 53182
rect 31726 53106 31778 53118
rect 32062 53170 32114 53182
rect 32062 53106 32114 53118
rect 32174 53170 32226 53182
rect 32174 53106 32226 53118
rect 34302 53170 34354 53182
rect 34302 53106 34354 53118
rect 52670 53170 52722 53182
rect 52670 53106 52722 53118
rect 6190 53058 6242 53070
rect 15710 53058 15762 53070
rect 1250 53006 1262 53058
rect 1314 53006 1326 53058
rect 10546 53006 10558 53058
rect 10610 53006 10622 53058
rect 6190 52994 6242 53006
rect 15710 52994 15762 53006
rect 19966 53058 20018 53070
rect 19966 52994 20018 53006
rect 25230 53058 25282 53070
rect 37102 53058 37154 53070
rect 27346 53006 27358 53058
rect 27410 53006 27422 53058
rect 32722 53006 32734 53058
rect 32786 53006 32798 53058
rect 25230 52994 25282 53006
rect 37102 52994 37154 53006
rect 7646 52946 7698 52958
rect 12126 52946 12178 52958
rect 17390 52946 17442 52958
rect 21646 52946 21698 52958
rect 31838 52946 31890 52958
rect 6514 52894 6526 52946
rect 6578 52894 6590 52946
rect 7074 52894 7086 52946
rect 7138 52894 7150 52946
rect 8306 52894 8318 52946
rect 8370 52894 8382 52946
rect 9314 52894 9326 52946
rect 9378 52894 9390 52946
rect 13122 52894 13134 52946
rect 13186 52894 13198 52946
rect 16034 52894 16046 52946
rect 16098 52894 16110 52946
rect 16482 52894 16494 52946
rect 16546 52894 16558 52946
rect 17714 52894 17726 52946
rect 17778 52894 17790 52946
rect 18722 52894 18734 52946
rect 18786 52894 18798 52946
rect 20850 52894 20862 52946
rect 20914 52894 20926 52946
rect 24658 52894 24670 52946
rect 24722 52894 24734 52946
rect 30258 52894 30270 52946
rect 30322 52894 30334 52946
rect 31602 52894 31614 52946
rect 31666 52894 31678 52946
rect 7646 52882 7698 52894
rect 12126 52882 12178 52894
rect 17390 52882 17442 52894
rect 21646 52882 21698 52894
rect 31838 52882 31890 52894
rect 34750 52946 34802 52958
rect 35198 52946 35250 52958
rect 44158 52946 44210 52958
rect 35074 52894 35086 52946
rect 35138 52894 35150 52946
rect 37426 52894 37438 52946
rect 37490 52894 37502 52946
rect 37986 52894 37998 52946
rect 38050 52894 38062 52946
rect 38658 52894 38670 52946
rect 38722 52894 38734 52946
rect 39330 52894 39342 52946
rect 39394 52894 39406 52946
rect 40114 52894 40126 52946
rect 40178 52894 40190 52946
rect 43362 52894 43374 52946
rect 43426 52894 43438 52946
rect 34750 52882 34802 52894
rect 35198 52882 35250 52894
rect 44158 52882 44210 52894
rect 44382 52946 44434 52958
rect 44382 52882 44434 52894
rect 44718 52946 44770 52958
rect 54686 52946 54738 52958
rect 46050 52894 46062 52946
rect 46114 52894 46126 52946
rect 44718 52882 44770 52894
rect 54686 52882 54738 52894
rect 5294 52834 5346 52846
rect 1586 52782 1598 52834
rect 1650 52782 1662 52834
rect 3714 52782 3726 52834
rect 3778 52782 3790 52834
rect 4050 52782 4062 52834
rect 4114 52782 4126 52834
rect 5294 52770 5346 52782
rect 5518 52834 5570 52846
rect 5518 52770 5570 52782
rect 5854 52834 5906 52846
rect 5854 52770 5906 52782
rect 9998 52834 10050 52846
rect 45054 52834 45106 52846
rect 10882 52782 10894 52834
rect 10946 52782 10958 52834
rect 21970 52782 21982 52834
rect 22034 52782 22046 52834
rect 30930 52782 30942 52834
rect 30994 52782 31006 52834
rect 41010 52782 41022 52834
rect 41074 52782 41086 52834
rect 42914 52782 42926 52834
rect 42978 52782 42990 52834
rect 9998 52770 10050 52782
rect 45054 52770 45106 52782
rect 45278 52834 45330 52846
rect 45278 52770 45330 52782
rect 48414 52834 48466 52846
rect 52322 52782 52334 52834
rect 52386 52782 52398 52834
rect 48414 52770 48466 52782
rect 2830 52722 2882 52734
rect 2830 52658 2882 52670
rect 3390 52722 3442 52734
rect 3390 52658 3442 52670
rect 4398 52722 4450 52734
rect 4398 52658 4450 52670
rect 5630 52722 5682 52734
rect 9886 52722 9938 52734
rect 14702 52722 14754 52734
rect 7186 52670 7198 52722
rect 7250 52670 7262 52722
rect 13570 52670 13582 52722
rect 13634 52670 13646 52722
rect 5630 52658 5682 52670
rect 9886 52658 9938 52670
rect 14702 52658 14754 52670
rect 15150 52722 15202 52734
rect 19294 52722 19346 52734
rect 16706 52670 16718 52722
rect 16770 52670 16782 52722
rect 15150 52658 15202 52670
rect 19294 52658 19346 52670
rect 19742 52722 19794 52734
rect 22318 52722 22370 52734
rect 25342 52722 25394 52734
rect 20626 52670 20638 52722
rect 20690 52670 20702 52722
rect 21298 52670 21310 52722
rect 21362 52670 21374 52722
rect 24210 52670 24222 52722
rect 24274 52670 24286 52722
rect 19742 52658 19794 52670
rect 22318 52658 22370 52670
rect 25342 52658 25394 52670
rect 25790 52722 25842 52734
rect 28590 52722 28642 52734
rect 31278 52722 31330 52734
rect 35310 52722 35362 52734
rect 26898 52670 26910 52722
rect 26962 52670 26974 52722
rect 29698 52670 29710 52722
rect 29762 52670 29774 52722
rect 33170 52670 33182 52722
rect 33234 52670 33246 52722
rect 25790 52658 25842 52670
rect 28590 52658 28642 52670
rect 31278 52658 31330 52670
rect 35310 52658 35362 52670
rect 35422 52722 35474 52734
rect 35422 52658 35474 52670
rect 36430 52722 36482 52734
rect 41358 52722 41410 52734
rect 36754 52670 36766 52722
rect 36818 52670 36830 52722
rect 38098 52670 38110 52722
rect 38162 52670 38174 52722
rect 36430 52658 36482 52670
rect 41358 52658 41410 52670
rect 41806 52722 41858 52734
rect 41806 52658 41858 52670
rect 44606 52722 44658 52734
rect 44606 52658 44658 52670
rect 45166 52722 45218 52734
rect 47742 52722 47794 52734
rect 49198 52722 49250 52734
rect 50206 52722 50258 52734
rect 51214 52722 51266 52734
rect 46610 52670 46622 52722
rect 46674 52670 46686 52722
rect 48738 52670 48750 52722
rect 48802 52670 48814 52722
rect 49522 52670 49534 52722
rect 49586 52670 49598 52722
rect 50530 52670 50542 52722
rect 50594 52670 50606 52722
rect 50866 52670 50878 52722
rect 50930 52670 50942 52722
rect 45166 52658 45218 52670
rect 47742 52658 47794 52670
rect 49198 52658 49250 52670
rect 50206 52658 50258 52670
rect 51214 52658 51266 52670
rect 51998 52722 52050 52734
rect 51998 52658 52050 52670
rect 52782 52722 52834 52734
rect 52782 52658 52834 52670
rect 52894 52722 52946 52734
rect 53678 52722 53730 52734
rect 55358 52722 55410 52734
rect 53330 52670 53342 52722
rect 53394 52670 53406 52722
rect 54338 52670 54350 52722
rect 54402 52670 54414 52722
rect 55010 52670 55022 52722
rect 55074 52670 55086 52722
rect 52894 52658 52946 52670
rect 53678 52658 53730 52670
rect 55358 52658 55410 52670
rect 56030 52722 56082 52734
rect 56354 52670 56366 52722
rect 56418 52670 56430 52722
rect 56030 52658 56082 52670
rect 672 52554 56784 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 44466 52554
rect 44518 52502 44570 52554
rect 44622 52502 44674 52554
rect 44726 52502 56784 52554
rect 672 52468 56784 52502
rect 3502 52386 3554 52398
rect 5966 52386 6018 52398
rect 8990 52386 9042 52398
rect 3826 52334 3838 52386
rect 3890 52334 3902 52386
rect 7074 52334 7086 52386
rect 7138 52334 7150 52386
rect 3502 52322 3554 52334
rect 5966 52322 6018 52334
rect 8990 52322 9042 52334
rect 11118 52386 11170 52398
rect 15262 52386 15314 52398
rect 31166 52386 31218 52398
rect 12562 52334 12574 52386
rect 12626 52334 12638 52386
rect 22754 52334 22766 52386
rect 22818 52334 22830 52386
rect 25890 52334 25902 52386
rect 25954 52334 25966 52386
rect 11118 52322 11170 52334
rect 15262 52322 15314 52334
rect 31166 52322 31218 52334
rect 39566 52386 39618 52398
rect 39566 52322 39618 52334
rect 42030 52386 42082 52398
rect 42030 52322 42082 52334
rect 46510 52386 46562 52398
rect 46510 52322 46562 52334
rect 50654 52386 50706 52398
rect 50654 52322 50706 52334
rect 56030 52386 56082 52398
rect 56030 52322 56082 52334
rect 8878 52274 8930 52286
rect 15598 52274 15650 52286
rect 20862 52274 20914 52286
rect 23886 52274 23938 52286
rect 1586 52222 1598 52274
rect 1650 52222 1662 52274
rect 4722 52222 4734 52274
rect 4786 52222 4798 52274
rect 9986 52222 9998 52274
rect 10050 52222 10062 52274
rect 18946 52222 18958 52274
rect 19010 52222 19022 52274
rect 21186 52222 21198 52274
rect 21250 52222 21262 52274
rect 8878 52210 8930 52222
rect 15598 52210 15650 52222
rect 20862 52210 20914 52222
rect 23886 52210 23938 52222
rect 24894 52274 24946 52286
rect 31502 52274 31554 52286
rect 34638 52274 34690 52286
rect 29474 52222 29486 52274
rect 29538 52222 29550 52274
rect 31826 52222 31838 52274
rect 31890 52222 31902 52274
rect 33730 52222 33742 52274
rect 33794 52222 33806 52274
rect 24894 52210 24946 52222
rect 31502 52210 31554 52222
rect 34638 52210 34690 52222
rect 34750 52274 34802 52286
rect 49534 52274 49586 52286
rect 35858 52222 35870 52274
rect 35922 52222 35934 52274
rect 38322 52222 38334 52274
rect 38386 52222 38398 52274
rect 40898 52222 40910 52274
rect 40962 52222 40974 52274
rect 42914 52222 42926 52274
rect 42978 52222 42990 52274
rect 46834 52222 46846 52274
rect 46898 52222 46910 52274
rect 47506 52222 47518 52274
rect 47570 52222 47582 52274
rect 34750 52210 34802 52222
rect 49534 52210 49586 52222
rect 50094 52274 50146 52286
rect 50094 52210 50146 52222
rect 50206 52274 50258 52286
rect 51874 52222 51886 52274
rect 51938 52222 51950 52274
rect 53106 52222 53118 52274
rect 53170 52222 53182 52274
rect 53666 52222 53678 52274
rect 53730 52222 53742 52274
rect 54338 52222 54350 52274
rect 54402 52222 54414 52274
rect 55346 52222 55358 52274
rect 55410 52222 55422 52274
rect 56354 52222 56366 52274
rect 56418 52222 56430 52274
rect 50206 52210 50258 52222
rect 8206 52162 8258 52174
rect 13246 52162 13298 52174
rect 15150 52162 15202 52174
rect 1250 52110 1262 52162
rect 1314 52110 1326 52162
rect 4274 52110 4286 52162
rect 4338 52110 4350 52162
rect 6626 52110 6638 52162
rect 6690 52110 6702 52162
rect 12002 52110 12014 52162
rect 12066 52110 12078 52162
rect 12450 52110 12462 52162
rect 12514 52110 12526 52162
rect 13682 52110 13694 52162
rect 13746 52110 13758 52162
rect 14690 52110 14702 52162
rect 14754 52110 14766 52162
rect 8206 52098 8258 52110
rect 13246 52098 13298 52110
rect 15150 52098 15202 52110
rect 15934 52162 15986 52174
rect 15934 52098 15986 52110
rect 16270 52162 16322 52174
rect 18286 52162 18338 52174
rect 19966 52162 20018 52174
rect 16818 52110 16830 52162
rect 16882 52110 16894 52162
rect 17938 52110 17950 52162
rect 18002 52110 18014 52162
rect 19170 52110 19182 52162
rect 19234 52110 19246 52162
rect 19506 52110 19518 52162
rect 19570 52110 19582 52162
rect 16270 52098 16322 52110
rect 18286 52098 18338 52110
rect 19966 52098 20018 52110
rect 20414 52162 20466 52174
rect 20414 52098 20466 52110
rect 20526 52162 20578 52174
rect 20526 52098 20578 52110
rect 21534 52162 21586 52174
rect 26350 52162 26402 52174
rect 31054 52162 31106 52174
rect 22306 52110 22318 52162
rect 22370 52110 22382 52162
rect 25218 52110 25230 52162
rect 25282 52110 25294 52162
rect 25666 52110 25678 52162
rect 25730 52110 25742 52162
rect 26898 52110 26910 52162
rect 26962 52110 26974 52162
rect 27906 52110 27918 52162
rect 27970 52110 27982 52162
rect 28914 52110 28926 52162
rect 28978 52110 28990 52162
rect 21534 52098 21586 52110
rect 26350 52098 26402 52110
rect 31054 52098 31106 52110
rect 32510 52162 32562 52174
rect 42590 52162 42642 52174
rect 48190 52162 48242 52174
rect 34066 52110 34078 52162
rect 34130 52110 34142 52162
rect 40450 52110 40462 52162
rect 40514 52110 40526 52162
rect 45378 52110 45390 52162
rect 45442 52110 45454 52162
rect 46162 52110 46174 52162
rect 46226 52110 46238 52162
rect 47282 52110 47294 52162
rect 47346 52110 47358 52162
rect 32510 52098 32562 52110
rect 42590 52098 42642 52110
rect 48190 52098 48242 52110
rect 49870 52162 49922 52174
rect 54014 52162 54066 52174
rect 52882 52110 52894 52162
rect 52946 52110 52958 52162
rect 49870 52098 49922 52110
rect 54014 52098 54066 52110
rect 54686 52162 54738 52174
rect 55122 52110 55134 52162
rect 55186 52110 55198 52162
rect 54686 52098 54738 52110
rect 11566 52050 11618 52062
rect 9538 51998 9550 52050
rect 9602 51998 9614 52050
rect 11566 51986 11618 51998
rect 16046 52050 16098 52062
rect 16046 51986 16098 51998
rect 20750 52050 20802 52062
rect 49422 52050 49474 52062
rect 35410 51998 35422 52050
rect 35474 51998 35486 52050
rect 37986 51998 37998 52050
rect 38050 51998 38062 52050
rect 43250 51998 43262 52050
rect 43314 51998 43326 52050
rect 52210 51998 52222 52050
rect 52274 51998 52286 52050
rect 20750 51986 20802 51998
rect 49422 51986 49474 51998
rect 2830 51938 2882 51950
rect 2830 51874 2882 51886
rect 30606 51938 30658 51950
rect 30606 51874 30658 51886
rect 34750 51938 34802 51950
rect 34750 51874 34802 51886
rect 36990 51938 37042 51950
rect 36990 51874 37042 51886
rect 48414 51938 48466 51950
rect 49310 51938 49362 51950
rect 48738 51886 48750 51938
rect 48802 51886 48814 51938
rect 48414 51874 48466 51886
rect 49310 51874 49362 51886
rect 672 51770 56784 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 43806 51770
rect 43858 51718 43910 51770
rect 43962 51718 44014 51770
rect 44066 51718 56784 51770
rect 672 51684 56784 51718
rect 11678 51602 11730 51614
rect 3826 51550 3838 51602
rect 3890 51550 3902 51602
rect 11678 51538 11730 51550
rect 28702 51602 28754 51614
rect 28702 51538 28754 51550
rect 34638 51602 34690 51614
rect 34638 51538 34690 51550
rect 42254 51602 42306 51614
rect 42254 51538 42306 51550
rect 42702 51602 42754 51614
rect 42702 51538 42754 51550
rect 43262 51602 43314 51614
rect 43262 51538 43314 51550
rect 43486 51602 43538 51614
rect 43486 51538 43538 51550
rect 49646 51602 49698 51614
rect 49646 51538 49698 51550
rect 50430 51602 50482 51614
rect 50430 51538 50482 51550
rect 4398 51490 4450 51502
rect 12126 51490 12178 51502
rect 10098 51438 10110 51490
rect 10162 51438 10174 51490
rect 4398 51426 4450 51438
rect 12126 51426 12178 51438
rect 20974 51490 21026 51502
rect 36430 51490 36482 51502
rect 21858 51438 21870 51490
rect 21922 51438 21934 51490
rect 33058 51438 33070 51490
rect 33122 51438 33134 51490
rect 36642 51438 36654 51490
rect 36706 51438 36718 51490
rect 37650 51438 37662 51490
rect 37714 51438 37726 51490
rect 46386 51438 46398 51490
rect 46450 51438 46462 51490
rect 48514 51438 48526 51490
rect 48578 51438 48590 51490
rect 49858 51438 49870 51490
rect 49922 51438 49934 51490
rect 20974 51426 21026 51438
rect 36430 51426 36482 51438
rect 4174 51378 4226 51390
rect 1250 51326 1262 51378
rect 1314 51326 1326 51378
rect 1362 51326 1374 51378
rect 1426 51326 1438 51378
rect 4174 51314 4226 51326
rect 5406 51378 5458 51390
rect 5406 51314 5458 51326
rect 5518 51378 5570 51390
rect 7758 51378 7810 51390
rect 14254 51378 14306 51390
rect 23998 51378 24050 51390
rect 5954 51326 5966 51378
rect 6018 51326 6030 51378
rect 6738 51326 6750 51378
rect 6802 51326 6814 51378
rect 7074 51326 7086 51378
rect 7138 51326 7150 51378
rect 8418 51326 8430 51378
rect 8482 51326 8494 51378
rect 9314 51326 9326 51378
rect 9378 51326 9390 51378
rect 13122 51326 13134 51378
rect 13186 51326 13198 51378
rect 13570 51326 13582 51378
rect 13634 51326 13646 51378
rect 15026 51326 15038 51378
rect 15090 51326 15102 51378
rect 15810 51326 15822 51378
rect 15874 51326 15886 51378
rect 17154 51326 17166 51378
rect 17218 51326 17230 51378
rect 17602 51326 17614 51378
rect 17666 51326 17678 51378
rect 18386 51326 18398 51378
rect 18450 51326 18462 51378
rect 18834 51326 18846 51378
rect 18898 51326 18910 51378
rect 19842 51326 19854 51378
rect 19906 51326 19918 51378
rect 20626 51326 20638 51378
rect 20690 51326 20702 51378
rect 5518 51314 5570 51326
rect 7758 51314 7810 51326
rect 14254 51314 14306 51326
rect 23998 51314 24050 51326
rect 24670 51378 24722 51390
rect 26350 51378 26402 51390
rect 28590 51378 28642 51390
rect 30606 51378 30658 51390
rect 35422 51378 35474 51390
rect 42814 51378 42866 51390
rect 25106 51326 25118 51378
rect 25170 51326 25182 51378
rect 25442 51326 25454 51378
rect 25506 51326 25518 51378
rect 26786 51326 26798 51378
rect 26850 51326 26862 51378
rect 27682 51326 27694 51378
rect 27746 51326 27758 51378
rect 29474 51326 29486 51378
rect 29538 51326 29550 51378
rect 30034 51326 30046 51378
rect 30098 51326 30110 51378
rect 31154 51326 31166 51378
rect 31218 51326 31230 51378
rect 32162 51326 32174 51378
rect 32226 51326 32238 51378
rect 35074 51326 35086 51378
rect 35138 51326 35150 51378
rect 40674 51326 40686 51378
rect 40738 51326 40750 51378
rect 24670 51314 24722 51326
rect 26350 51314 26402 51326
rect 28590 51314 28642 51326
rect 30606 51314 30658 51326
rect 35422 51314 35474 51326
rect 42814 51314 42866 51326
rect 44494 51378 44546 51390
rect 44494 51314 44546 51326
rect 44718 51378 44770 51390
rect 44718 51314 44770 51326
rect 44942 51378 44994 51390
rect 45726 51378 45778 51390
rect 50206 51378 50258 51390
rect 45266 51326 45278 51378
rect 45330 51326 45342 51378
rect 49186 51326 49198 51378
rect 49250 51326 49262 51378
rect 44942 51314 44994 51326
rect 45726 51314 45778 51326
rect 50206 51314 50258 51326
rect 50990 51378 51042 51390
rect 50990 51314 51042 51326
rect 51102 51378 51154 51390
rect 51102 51314 51154 51326
rect 51326 51378 51378 51390
rect 51326 51314 51378 51326
rect 51438 51378 51490 51390
rect 53342 51378 53394 51390
rect 52098 51326 52110 51378
rect 52162 51326 52174 51378
rect 52658 51326 52670 51378
rect 52722 51326 52734 51378
rect 51438 51314 51490 51326
rect 53342 51314 53394 51326
rect 3390 51266 3442 51278
rect 1810 51214 1822 51266
rect 1874 51214 1886 51266
rect 3390 51202 3442 51214
rect 6302 51266 6354 51278
rect 12798 51266 12850 51278
rect 16494 51266 16546 51278
rect 7298 51214 7310 51266
rect 7362 51214 7374 51266
rect 10546 51214 10558 51266
rect 10610 51214 10622 51266
rect 13794 51214 13806 51266
rect 13858 51214 13870 51266
rect 6302 51202 6354 51214
rect 12798 51202 12850 51214
rect 16494 51202 16546 51214
rect 16830 51266 16882 51278
rect 24222 51266 24274 51278
rect 17826 51214 17838 51266
rect 17890 51214 17902 51266
rect 16830 51202 16882 51214
rect 24222 51202 24274 51214
rect 24334 51266 24386 51278
rect 29150 51266 29202 51278
rect 36318 51266 36370 51278
rect 25666 51214 25678 51266
rect 25730 51214 25742 51266
rect 30146 51214 30158 51266
rect 30210 51214 30222 51266
rect 24334 51202 24386 51214
rect 29150 51202 29202 51214
rect 36318 51202 36370 51214
rect 36542 51266 36594 51278
rect 49870 51266 49922 51278
rect 53006 51266 53058 51278
rect 38098 51214 38110 51266
rect 38162 51214 38174 51266
rect 39778 51214 39790 51266
rect 39842 51214 39854 51266
rect 41122 51214 41134 51266
rect 41186 51214 41198 51266
rect 52322 51214 52334 51266
rect 52386 51214 52398 51266
rect 36542 51202 36594 51214
rect 49870 51202 49922 51214
rect 53006 51202 53058 51214
rect 54574 51266 54626 51278
rect 54898 51214 54910 51266
rect 54962 51214 54974 51266
rect 54574 51202 54626 51214
rect 2942 51154 2994 51166
rect 2942 51090 2994 51102
rect 3502 51154 3554 51166
rect 3502 51090 3554 51102
rect 5630 51154 5682 51166
rect 5630 51090 5682 51102
rect 5742 51154 5794 51166
rect 5742 51090 5794 51102
rect 12238 51154 12290 51166
rect 12238 51090 12290 51102
rect 16382 51154 16434 51166
rect 16382 51090 16434 51102
rect 20862 51154 20914 51166
rect 20862 51090 20914 51102
rect 21086 51154 21138 51166
rect 21086 51090 21138 51102
rect 21198 51154 21250 51166
rect 23438 51154 23490 51166
rect 22306 51102 22318 51154
rect 22370 51102 22382 51154
rect 21198 51090 21250 51102
rect 23438 51090 23490 51102
rect 28702 51154 28754 51166
rect 35198 51154 35250 51166
rect 33506 51102 33518 51154
rect 33570 51102 33582 51154
rect 28702 51090 28754 51102
rect 35198 51090 35250 51102
rect 35534 51154 35586 51166
rect 35534 51090 35586 51102
rect 35646 51154 35698 51166
rect 35646 51090 35698 51102
rect 39230 51154 39282 51166
rect 39230 51090 39282 51102
rect 40126 51154 40178 51166
rect 40126 51090 40178 51102
rect 43598 51154 43650 51166
rect 43598 51090 43650 51102
rect 44270 51154 44322 51166
rect 44270 51090 44322 51102
rect 44382 51154 44434 51166
rect 44382 51090 44434 51102
rect 45614 51154 45666 51166
rect 45614 51090 45666 51102
rect 45838 51154 45890 51166
rect 45838 51090 45890 51102
rect 52894 51154 52946 51166
rect 54238 51154 54290 51166
rect 55582 51154 55634 51166
rect 53666 51102 53678 51154
rect 53730 51102 53742 51154
rect 55234 51102 55246 51154
rect 55298 51102 55310 51154
rect 52894 51090 52946 51102
rect 54238 51090 54290 51102
rect 55582 51090 55634 51102
rect 56030 51154 56082 51166
rect 56354 51102 56366 51154
rect 56418 51102 56430 51154
rect 56030 51090 56082 51102
rect 672 50986 56784 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 44466 50986
rect 44518 50934 44570 50986
rect 44622 50934 44674 50986
rect 44726 50934 56784 50986
rect 672 50900 56784 50934
rect 35982 50818 36034 50830
rect 9538 50766 9550 50818
rect 9602 50766 9614 50818
rect 12338 50766 12350 50818
rect 12402 50766 12414 50818
rect 25554 50766 25566 50818
rect 25618 50766 25630 50818
rect 29586 50766 29598 50818
rect 29650 50766 29662 50818
rect 35982 50754 36034 50766
rect 42814 50818 42866 50830
rect 51998 50818 52050 50830
rect 54462 50818 54514 50830
rect 46274 50766 46286 50818
rect 46338 50766 46350 50818
rect 53442 50766 53454 50818
rect 53506 50766 53518 50818
rect 55346 50766 55358 50818
rect 55410 50766 55422 50818
rect 42814 50754 42866 50766
rect 51998 50754 52050 50766
rect 54462 50754 54514 50766
rect 6862 50706 6914 50718
rect 18510 50706 18562 50718
rect 1586 50654 1598 50706
rect 1650 50654 1662 50706
rect 4722 50654 4734 50706
rect 4786 50654 4798 50706
rect 7298 50654 7310 50706
rect 7362 50654 7374 50706
rect 14914 50654 14926 50706
rect 14978 50654 14990 50706
rect 18050 50654 18062 50706
rect 18114 50654 18126 50706
rect 6862 50642 6914 50654
rect 18510 50642 18562 50654
rect 20750 50706 20802 50718
rect 28590 50706 28642 50718
rect 36430 50706 36482 50718
rect 37886 50706 37938 50718
rect 45054 50706 45106 50718
rect 21746 50654 21758 50706
rect 21810 50654 21822 50706
rect 33730 50654 33742 50706
rect 33794 50654 33806 50706
rect 35074 50654 35086 50706
rect 35138 50654 35150 50706
rect 35410 50654 35422 50706
rect 35474 50654 35486 50706
rect 37426 50654 37438 50706
rect 37490 50654 37502 50706
rect 41570 50654 41582 50706
rect 41634 50654 41646 50706
rect 43922 50654 43934 50706
rect 43986 50654 43998 50706
rect 20750 50642 20802 50654
rect 28590 50642 28642 50654
rect 36430 50642 36482 50654
rect 37886 50642 37938 50654
rect 45054 50642 45106 50654
rect 47406 50706 47458 50718
rect 52894 50706 52946 50718
rect 49074 50654 49086 50706
rect 49138 50654 49150 50706
rect 49634 50654 49646 50706
rect 49698 50654 49710 50706
rect 50754 50654 50766 50706
rect 50818 50654 50830 50706
rect 56354 50654 56366 50706
rect 56418 50654 56430 50706
rect 47406 50642 47458 50654
rect 52894 50642 52946 50654
rect 3502 50594 3554 50606
rect 3502 50530 3554 50542
rect 3838 50594 3890 50606
rect 3838 50530 3890 50542
rect 3950 50594 4002 50606
rect 8318 50594 8370 50606
rect 11342 50594 11394 50606
rect 13022 50594 13074 50606
rect 15262 50594 15314 50606
rect 4498 50542 4510 50594
rect 4562 50542 4574 50594
rect 5282 50542 5294 50594
rect 5346 50542 5358 50594
rect 6066 50542 6078 50594
rect 6130 50542 6142 50594
rect 7522 50542 7534 50594
rect 7586 50542 7598 50594
rect 7970 50542 7982 50594
rect 8034 50542 8046 50594
rect 9090 50542 9102 50594
rect 9154 50542 9166 50594
rect 11778 50542 11790 50594
rect 11842 50542 11854 50594
rect 12226 50542 12238 50594
rect 12290 50542 12302 50594
rect 13458 50542 13470 50594
rect 13522 50542 13534 50594
rect 14466 50542 14478 50594
rect 14530 50542 14542 50594
rect 3950 50530 4002 50542
rect 8318 50530 8370 50542
rect 11342 50530 11394 50542
rect 13022 50530 13074 50542
rect 15262 50530 15314 50542
rect 15598 50594 15650 50606
rect 15598 50530 15650 50542
rect 15822 50594 15874 50606
rect 15822 50530 15874 50542
rect 16158 50594 16210 50606
rect 22430 50594 22482 50606
rect 26238 50594 26290 50606
rect 30270 50594 30322 50606
rect 35646 50594 35698 50606
rect 40350 50594 40402 50606
rect 45278 50594 45330 50606
rect 17378 50542 17390 50594
rect 17442 50542 17454 50594
rect 17826 50542 17838 50594
rect 17890 50542 17902 50594
rect 19058 50542 19070 50594
rect 19122 50542 19134 50594
rect 20066 50542 20078 50594
rect 20130 50542 20142 50594
rect 21186 50542 21198 50594
rect 21250 50542 21262 50594
rect 21522 50542 21534 50594
rect 21586 50542 21598 50594
rect 22754 50542 22766 50594
rect 22818 50542 22830 50594
rect 23762 50542 23774 50594
rect 23826 50542 23838 50594
rect 24994 50542 25006 50594
rect 25058 50542 25070 50594
rect 25330 50542 25342 50594
rect 25394 50542 25406 50594
rect 26562 50542 26574 50594
rect 26626 50542 26638 50594
rect 27570 50542 27582 50594
rect 27634 50542 27646 50594
rect 28914 50542 28926 50594
rect 28978 50542 28990 50594
rect 29362 50542 29374 50594
rect 29426 50542 29438 50594
rect 30818 50542 30830 50594
rect 30882 50542 30894 50594
rect 31714 50542 31726 50594
rect 31778 50542 31790 50594
rect 34066 50542 34078 50594
rect 34130 50542 34142 50594
rect 36754 50542 36766 50594
rect 36818 50542 36830 50594
rect 37202 50542 37214 50594
rect 37266 50542 37278 50594
rect 38658 50542 38670 50594
rect 38722 50542 38734 50594
rect 39554 50542 39566 50594
rect 39618 50542 39630 50594
rect 41906 50542 41918 50594
rect 41970 50542 41982 50594
rect 16158 50530 16210 50542
rect 22430 50530 22482 50542
rect 26238 50530 26290 50542
rect 30270 50530 30322 50542
rect 35646 50530 35698 50542
rect 40350 50530 40402 50542
rect 45278 50530 45330 50542
rect 48526 50594 48578 50606
rect 48526 50530 48578 50542
rect 48862 50594 48914 50606
rect 55022 50594 55074 50606
rect 53666 50542 53678 50594
rect 53730 50542 53742 50594
rect 56130 50542 56142 50594
rect 56194 50542 56206 50594
rect 48862 50530 48914 50542
rect 55022 50530 55074 50542
rect 2830 50482 2882 50494
rect 1250 50430 1262 50482
rect 1314 50430 1326 50482
rect 2830 50418 2882 50430
rect 3614 50482 3666 50494
rect 3614 50418 3666 50430
rect 16046 50482 16098 50494
rect 16046 50418 16098 50430
rect 17054 50482 17106 50494
rect 17054 50418 17106 50430
rect 24558 50482 24610 50494
rect 54238 50482 54290 50494
rect 44370 50430 44382 50482
rect 44434 50430 44446 50482
rect 44930 50430 44942 50482
rect 44994 50430 45006 50482
rect 45826 50430 45838 50482
rect 45890 50430 45902 50482
rect 50418 50430 50430 50482
rect 50482 50430 50494 50482
rect 52770 50430 52782 50482
rect 52834 50430 52846 50482
rect 54562 50430 54574 50482
rect 54626 50430 54638 50482
rect 24558 50418 24610 50430
rect 54238 50418 54290 50430
rect 10670 50370 10722 50382
rect 10670 50306 10722 50318
rect 32510 50370 32562 50382
rect 32510 50306 32562 50318
rect 53118 50370 53170 50382
rect 53118 50306 53170 50318
rect 672 50202 56784 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 43806 50202
rect 43858 50150 43910 50202
rect 43962 50150 44014 50202
rect 44066 50150 56784 50202
rect 672 50116 56784 50150
rect 22654 50034 22706 50046
rect 35422 50034 35474 50046
rect 35074 49982 35086 50034
rect 35138 49982 35150 50034
rect 22654 49970 22706 49982
rect 35422 49970 35474 49982
rect 36430 50034 36482 50046
rect 36430 49970 36482 49982
rect 43374 50034 43426 50046
rect 48750 50034 48802 50046
rect 47506 49982 47518 50034
rect 47570 49982 47582 50034
rect 43374 49970 43426 49982
rect 48750 49970 48802 49982
rect 44606 49922 44658 49934
rect 13122 49870 13134 49922
rect 13186 49870 13198 49922
rect 21074 49870 21086 49922
rect 21138 49870 21150 49922
rect 32274 49870 32286 49922
rect 32338 49870 32350 49922
rect 39218 49870 39230 49922
rect 39282 49870 39294 49922
rect 44606 49858 44658 49870
rect 3166 49810 3218 49822
rect 1250 49758 1262 49810
rect 1314 49758 1326 49810
rect 3166 49746 3218 49758
rect 4398 49810 4450 49822
rect 10558 49810 10610 49822
rect 14702 49810 14754 49822
rect 19182 49810 19234 49822
rect 25118 49810 25170 49822
rect 29822 49810 29874 49822
rect 5618 49758 5630 49810
rect 5682 49758 5694 49810
rect 5954 49758 5966 49810
rect 6018 49758 6030 49810
rect 6738 49758 6750 49810
rect 6802 49758 6814 49810
rect 7186 49758 7198 49810
rect 7250 49758 7262 49810
rect 8306 49758 8318 49810
rect 8370 49758 8382 49810
rect 9202 49758 9214 49810
rect 9266 49758 9278 49810
rect 10098 49758 10110 49810
rect 10162 49758 10174 49810
rect 11330 49758 11342 49810
rect 11394 49758 11406 49810
rect 11778 49758 11790 49810
rect 11842 49758 11854 49810
rect 15474 49758 15486 49810
rect 15538 49758 15550 49810
rect 15922 49758 15934 49810
rect 15986 49758 15998 49810
rect 16706 49758 16718 49810
rect 16770 49758 16782 49810
rect 17378 49758 17390 49810
rect 17442 49758 17454 49810
rect 18162 49758 18174 49810
rect 18226 49758 18238 49810
rect 23762 49758 23774 49810
rect 23826 49758 23838 49810
rect 24210 49758 24222 49810
rect 24274 49758 24286 49810
rect 25554 49758 25566 49810
rect 25618 49758 25630 49810
rect 26450 49758 26462 49810
rect 26514 49758 26526 49810
rect 4398 49746 4450 49758
rect 10558 49746 10610 49758
rect 14702 49746 14754 49758
rect 19182 49746 19234 49758
rect 25118 49746 25170 49758
rect 29822 49746 29874 49758
rect 30046 49810 30098 49822
rect 30046 49746 30098 49758
rect 30270 49810 30322 49822
rect 30270 49746 30322 49758
rect 32958 49810 33010 49822
rect 35646 49810 35698 49822
rect 44494 49810 44546 49822
rect 34514 49758 34526 49810
rect 34578 49758 34590 49810
rect 38098 49758 38110 49810
rect 38162 49758 38174 49810
rect 41682 49758 41694 49810
rect 41746 49758 41758 49810
rect 32958 49746 33010 49758
rect 35646 49746 35698 49758
rect 44494 49746 44546 49758
rect 44718 49810 44770 49822
rect 46846 49810 46898 49822
rect 48078 49810 48130 49822
rect 45266 49758 45278 49810
rect 45330 49758 45342 49810
rect 47282 49758 47294 49810
rect 47346 49758 47358 49810
rect 47842 49758 47854 49810
rect 47906 49758 47918 49810
rect 44718 49746 44770 49758
rect 46846 49746 46898 49758
rect 48078 49746 48130 49758
rect 48974 49810 49026 49822
rect 50990 49810 51042 49822
rect 50194 49758 50206 49810
rect 50258 49758 50270 49810
rect 48974 49746 49026 49758
rect 50990 49746 51042 49758
rect 51214 49810 51266 49822
rect 51214 49746 51266 49758
rect 51326 49810 51378 49822
rect 52994 49758 53006 49810
rect 53058 49758 53070 49810
rect 51326 49746 51378 49758
rect 3502 49698 3554 49710
rect 1586 49646 1598 49698
rect 1650 49646 1662 49698
rect 3502 49634 3554 49646
rect 3838 49698 3890 49710
rect 3838 49634 3890 49646
rect 4174 49698 4226 49710
rect 4174 49634 4226 49646
rect 5182 49698 5234 49710
rect 12238 49698 12290 49710
rect 6178 49646 6190 49698
rect 6242 49646 6254 49698
rect 5182 49634 5234 49646
rect 12238 49634 12290 49646
rect 15150 49698 15202 49710
rect 23438 49698 23490 49710
rect 29598 49698 29650 49710
rect 16146 49646 16158 49698
rect 16210 49646 16222 49698
rect 19394 49646 19406 49698
rect 19458 49646 19470 49698
rect 19954 49646 19966 49698
rect 20018 49646 20030 49698
rect 21522 49646 21534 49698
rect 21586 49646 21598 49698
rect 24434 49646 24446 49698
rect 24498 49646 24510 49698
rect 15150 49634 15202 49646
rect 23438 49634 23490 49646
rect 29598 49634 29650 49646
rect 30718 49698 30770 49710
rect 38558 49698 38610 49710
rect 44158 49698 44210 49710
rect 31826 49646 31838 49698
rect 31890 49646 31902 49698
rect 37650 49646 37662 49698
rect 37714 49646 37726 49698
rect 42130 49646 42142 49698
rect 42194 49646 42206 49698
rect 30718 49634 30770 49646
rect 38558 49634 38610 49646
rect 44158 49634 44210 49646
rect 47966 49698 48018 49710
rect 47966 49634 48018 49646
rect 49646 49698 49698 49710
rect 50878 49698 50930 49710
rect 50418 49646 50430 49698
rect 50482 49646 50494 49698
rect 49646 49634 49698 49646
rect 50878 49634 50930 49646
rect 2830 49586 2882 49598
rect 2830 49522 2882 49534
rect 3390 49586 3442 49598
rect 3390 49522 3442 49534
rect 4062 49586 4114 49598
rect 18846 49586 18898 49598
rect 11218 49534 11230 49586
rect 11282 49534 11294 49586
rect 13570 49534 13582 49586
rect 13634 49534 13646 49586
rect 4062 49522 4114 49534
rect 18846 49522 18898 49534
rect 29710 49586 29762 49598
rect 38670 49586 38722 49598
rect 40798 49586 40850 49598
rect 49422 49586 49474 49598
rect 34066 49534 34078 49586
rect 34130 49534 34142 49586
rect 39666 49534 39678 49586
rect 39730 49534 39742 49586
rect 45714 49534 45726 49586
rect 45778 49534 45790 49586
rect 48402 49534 48414 49586
rect 48466 49534 48478 49586
rect 29710 49522 29762 49534
rect 38670 49522 38722 49534
rect 40798 49522 40850 49534
rect 49422 49522 49474 49534
rect 49534 49586 49586 49598
rect 52334 49586 52386 49598
rect 54686 49586 54738 49598
rect 51986 49534 51998 49586
rect 52050 49534 52062 49586
rect 53554 49534 53566 49586
rect 53618 49534 53630 49586
rect 49534 49522 49586 49534
rect 52334 49522 52386 49534
rect 54686 49522 54738 49534
rect 55246 49586 55298 49598
rect 55918 49586 55970 49598
rect 55570 49534 55582 49586
rect 55634 49534 55646 49586
rect 56242 49534 56254 49586
rect 56306 49534 56318 49586
rect 55246 49522 55298 49534
rect 55918 49522 55970 49534
rect 672 49418 56784 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 44466 49418
rect 44518 49366 44570 49418
rect 44622 49366 44674 49418
rect 44726 49366 56784 49418
rect 672 49332 56784 49366
rect 1150 49250 1202 49262
rect 1822 49250 1874 49262
rect 16046 49250 16098 49262
rect 1474 49198 1486 49250
rect 1538 49198 1550 49250
rect 2146 49198 2158 49250
rect 2210 49198 2222 49250
rect 3490 49198 3502 49250
rect 3554 49198 3566 49250
rect 7074 49198 7086 49250
rect 7138 49198 7150 49250
rect 1150 49186 1202 49198
rect 1822 49186 1874 49198
rect 16046 49186 16098 49198
rect 25118 49250 25170 49262
rect 25118 49186 25170 49198
rect 30606 49250 30658 49262
rect 30606 49186 30658 49198
rect 30830 49250 30882 49262
rect 30830 49186 30882 49198
rect 31390 49250 31442 49262
rect 31390 49186 31442 49198
rect 34750 49250 34802 49262
rect 48974 49250 49026 49262
rect 35858 49198 35870 49250
rect 35922 49198 35934 49250
rect 39666 49198 39678 49250
rect 39730 49198 39742 49250
rect 40898 49198 40910 49250
rect 40962 49198 40974 49250
rect 47170 49198 47182 49250
rect 47234 49198 47246 49250
rect 55346 49198 55358 49250
rect 55410 49198 55422 49250
rect 56354 49198 56366 49250
rect 56418 49198 56430 49250
rect 34750 49186 34802 49198
rect 48974 49186 49026 49198
rect 3950 49138 4002 49150
rect 3950 49074 4002 49086
rect 9326 49138 9378 49150
rect 46510 49138 46562 49150
rect 10322 49086 10334 49138
rect 10386 49086 10398 49138
rect 13794 49086 13806 49138
rect 13858 49086 13870 49138
rect 18050 49086 18062 49138
rect 18114 49086 18126 49138
rect 19170 49086 19182 49138
rect 19234 49086 19246 49138
rect 21746 49086 21758 49138
rect 21810 49086 21822 49138
rect 25778 49086 25790 49138
rect 25842 49086 25854 49138
rect 26226 49086 26238 49138
rect 26290 49086 26302 49138
rect 27682 49086 27694 49138
rect 27746 49086 27758 49138
rect 33618 49086 33630 49138
rect 33682 49086 33694 49138
rect 37426 49086 37438 49138
rect 37490 49086 37502 49138
rect 45266 49086 45278 49138
rect 45330 49086 45342 49138
rect 50082 49086 50094 49138
rect 50146 49086 50158 49138
rect 52994 49086 53006 49138
rect 53058 49086 53070 49138
rect 54338 49086 54350 49138
rect 54402 49086 54414 49138
rect 9326 49074 9378 49086
rect 46510 49074 46562 49086
rect 8206 49026 8258 49038
rect 10782 49026 10834 49038
rect 15710 49026 15762 49038
rect 2930 48974 2942 49026
rect 2994 48974 3006 49026
rect 3378 48974 3390 49026
rect 3442 48974 3454 49026
rect 4498 48974 4510 49026
rect 4562 48974 4574 49026
rect 5506 48974 5518 49026
rect 5570 48974 5582 49026
rect 9762 48974 9774 49026
rect 9826 48974 9838 49026
rect 10098 48974 10110 49026
rect 10162 48974 10174 49026
rect 11330 48974 11342 49026
rect 11394 48974 11406 49026
rect 12450 48974 12462 49026
rect 12514 48974 12526 49026
rect 13234 48974 13246 49026
rect 13298 48974 13310 49026
rect 15474 48974 15486 49026
rect 15538 48974 15550 49026
rect 8206 48962 8258 48974
rect 10782 48962 10834 48974
rect 15710 48962 15762 48974
rect 15934 49026 15986 49038
rect 15934 48962 15986 48974
rect 17278 49026 17330 49038
rect 22430 49026 22482 49038
rect 28366 49026 28418 49038
rect 30494 49026 30546 49038
rect 17938 48974 17950 49026
rect 18002 48974 18014 49026
rect 18722 48974 18734 49026
rect 18786 48974 18798 49026
rect 21074 48974 21086 49026
rect 21138 48974 21150 49026
rect 21522 48974 21534 49026
rect 21586 48974 21598 49026
rect 22754 48974 22766 49026
rect 22818 48974 22830 49026
rect 23762 48974 23774 49026
rect 23826 48974 23838 49026
rect 27010 48974 27022 49026
rect 27074 48974 27086 49026
rect 27570 48974 27582 49026
rect 27634 48974 27646 49026
rect 28690 48974 28702 49026
rect 28754 48974 28766 49026
rect 29698 48974 29710 49026
rect 29762 48974 29774 49026
rect 17278 48962 17330 48974
rect 22430 48962 22482 48974
rect 28366 48962 28418 48974
rect 30494 48962 30546 48974
rect 31166 49026 31218 49038
rect 46622 49026 46674 49038
rect 34178 48974 34190 49026
rect 34242 48974 34254 49026
rect 37090 48974 37102 49026
rect 37154 48974 37166 49026
rect 39442 48974 39454 49026
rect 39506 48974 39518 49026
rect 40338 48974 40350 49026
rect 40402 48974 40414 49026
rect 42466 48974 42478 49026
rect 42530 48974 42542 49026
rect 46050 48974 46062 49026
rect 46114 48974 46126 49026
rect 31166 48962 31218 48974
rect 46622 48962 46674 48974
rect 46734 49026 46786 49038
rect 46734 48962 46786 48974
rect 48302 49026 48354 49038
rect 48302 48962 48354 48974
rect 48638 49026 48690 49038
rect 48638 48962 48690 48974
rect 48862 49026 48914 49038
rect 54014 49026 54066 49038
rect 53442 48974 53454 49026
rect 53506 48974 53518 49026
rect 48862 48962 48914 48974
rect 54014 48962 54066 48974
rect 55022 49026 55074 49038
rect 55022 48962 55074 48974
rect 56030 49026 56082 49038
rect 56030 48962 56082 48974
rect 2494 48914 2546 48926
rect 8990 48914 9042 48926
rect 6626 48862 6638 48914
rect 6690 48862 6702 48914
rect 2494 48850 2546 48862
rect 8990 48850 9042 48862
rect 14926 48914 14978 48926
rect 20750 48914 20802 48926
rect 16034 48862 16046 48914
rect 16098 48862 16110 48914
rect 14926 48850 14978 48862
rect 20750 48850 20802 48862
rect 26686 48914 26738 48926
rect 26686 48850 26738 48862
rect 31278 48914 31330 48926
rect 31278 48850 31330 48862
rect 31614 48914 31666 48926
rect 36306 48862 36318 48914
rect 36370 48862 36382 48914
rect 43138 48862 43150 48914
rect 43202 48862 43214 48914
rect 49746 48862 49758 48914
rect 49810 48862 49822 48914
rect 31614 48850 31666 48862
rect 8878 48802 8930 48814
rect 8878 48738 8930 48750
rect 16942 48802 16994 48814
rect 16942 48738 16994 48750
rect 20302 48802 20354 48814
rect 20302 48738 20354 48750
rect 25454 48802 25506 48814
rect 25454 48738 25506 48750
rect 31838 48802 31890 48814
rect 31838 48738 31890 48750
rect 32510 48802 32562 48814
rect 32510 48738 32562 48750
rect 38670 48802 38722 48814
rect 38670 48738 38722 48750
rect 42030 48802 42082 48814
rect 42030 48738 42082 48750
rect 42478 48802 42530 48814
rect 42478 48738 42530 48750
rect 42814 48802 42866 48814
rect 42814 48738 42866 48750
rect 48078 48802 48130 48814
rect 48078 48738 48130 48750
rect 51326 48802 51378 48814
rect 51326 48738 51378 48750
rect 51886 48802 51938 48814
rect 51886 48738 51938 48750
rect 672 48634 56784 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 43806 48634
rect 43858 48582 43910 48634
rect 43962 48582 44014 48634
rect 44066 48582 56784 48634
rect 672 48548 56784 48582
rect 20750 48466 20802 48478
rect 20750 48402 20802 48414
rect 36654 48466 36706 48478
rect 36654 48402 36706 48414
rect 43038 48466 43090 48478
rect 43038 48402 43090 48414
rect 1150 48354 1202 48366
rect 1150 48290 1202 48302
rect 4958 48354 5010 48366
rect 15262 48354 15314 48366
rect 35086 48354 35138 48366
rect 13234 48302 13246 48354
rect 13298 48302 13310 48354
rect 33954 48302 33966 48354
rect 34018 48302 34030 48354
rect 46946 48302 46958 48354
rect 47010 48302 47022 48354
rect 49074 48302 49086 48354
rect 49138 48302 49150 48354
rect 4958 48290 5010 48302
rect 15262 48290 15314 48302
rect 35086 48290 35138 48302
rect 6414 48242 6466 48254
rect 20638 48242 20690 48254
rect 34862 48242 34914 48254
rect 1586 48190 1598 48242
rect 1650 48190 1662 48242
rect 1922 48190 1934 48242
rect 1986 48190 1998 48242
rect 2706 48190 2718 48242
rect 2770 48190 2782 48242
rect 3154 48190 3166 48242
rect 3218 48190 3230 48242
rect 4162 48185 4174 48237
rect 4226 48185 4238 48237
rect 5282 48190 5294 48242
rect 5346 48190 5358 48242
rect 5730 48190 5742 48242
rect 5794 48190 5806 48242
rect 6962 48190 6974 48242
rect 7026 48190 7038 48242
rect 7186 48190 7198 48242
rect 7250 48190 7262 48242
rect 7970 48190 7982 48242
rect 8034 48190 8046 48242
rect 9426 48190 9438 48242
rect 9490 48190 9502 48242
rect 9762 48190 9774 48242
rect 9826 48190 9838 48242
rect 10546 48190 10558 48242
rect 10610 48190 10622 48242
rect 11218 48190 11230 48242
rect 11282 48190 11294 48242
rect 12114 48190 12126 48242
rect 12178 48190 12190 48242
rect 15586 48190 15598 48242
rect 15650 48190 15662 48242
rect 16034 48190 16046 48242
rect 16098 48190 16110 48242
rect 16818 48190 16830 48242
rect 16882 48190 16894 48242
rect 17266 48190 17278 48242
rect 17330 48190 17342 48242
rect 18274 48190 18286 48242
rect 18338 48190 18350 48242
rect 21634 48190 21646 48242
rect 21698 48190 21710 48242
rect 23986 48190 23998 48242
rect 24050 48190 24062 48242
rect 26226 48190 26238 48242
rect 26290 48190 26302 48242
rect 30258 48190 30270 48242
rect 30322 48190 30334 48242
rect 6414 48178 6466 48190
rect 20638 48178 20690 48190
rect 34862 48178 34914 48190
rect 35534 48242 35586 48254
rect 35534 48178 35586 48190
rect 36430 48242 36482 48254
rect 36430 48178 36482 48190
rect 37102 48242 37154 48254
rect 43598 48242 43650 48254
rect 38098 48190 38110 48242
rect 38162 48190 38174 48242
rect 38546 48190 38558 48242
rect 38610 48190 38622 48242
rect 39778 48190 39790 48242
rect 39842 48190 39854 48242
rect 40786 48190 40798 48242
rect 40850 48190 40862 48242
rect 41346 48190 41358 48242
rect 41410 48190 41422 48242
rect 37102 48178 37154 48190
rect 43598 48178 43650 48190
rect 44382 48242 44434 48254
rect 50654 48242 50706 48254
rect 44930 48190 44942 48242
rect 44994 48190 45006 48242
rect 49858 48190 49870 48242
rect 49922 48190 49934 48242
rect 44382 48178 44434 48190
rect 50654 48178 50706 48190
rect 50878 48242 50930 48254
rect 50878 48178 50930 48190
rect 51102 48242 51154 48254
rect 52098 48190 52110 48242
rect 52162 48190 52174 48242
rect 54786 48190 54798 48242
rect 54850 48190 54862 48242
rect 55570 48190 55582 48242
rect 55634 48190 55646 48242
rect 56130 48190 56142 48242
rect 56194 48190 56206 48242
rect 51102 48178 51154 48190
rect 8654 48130 8706 48142
rect 2146 48078 2158 48130
rect 2210 48078 2222 48130
rect 5954 48078 5966 48130
rect 6018 48078 6030 48130
rect 8654 48066 8706 48078
rect 8990 48130 9042 48142
rect 36878 48130 36930 48142
rect 9986 48078 9998 48130
rect 10050 48078 10062 48130
rect 22082 48078 22094 48130
rect 22146 48078 22158 48130
rect 24322 48078 24334 48130
rect 24386 48078 24398 48130
rect 26562 48078 26574 48130
rect 26626 48078 26638 48130
rect 30706 48078 30718 48130
rect 30770 48078 30782 48130
rect 8990 48066 9042 48078
rect 36878 48066 36930 48078
rect 37214 48130 37266 48142
rect 37214 48066 37266 48078
rect 37662 48130 37714 48142
rect 37662 48066 37714 48078
rect 39118 48130 39170 48142
rect 50206 48130 50258 48142
rect 41794 48078 41806 48130
rect 41858 48078 41870 48130
rect 45266 48078 45278 48130
rect 45330 48078 45342 48130
rect 39118 48066 39170 48078
rect 50206 48066 50258 48078
rect 50318 48130 50370 48142
rect 50318 48066 50370 48078
rect 54238 48130 54290 48142
rect 55010 48078 55022 48130
rect 55074 48078 55086 48130
rect 54238 48066 54290 48078
rect 8542 48018 8594 48030
rect 14814 48018 14866 48030
rect 19182 48018 19234 48030
rect 19854 48018 19906 48030
rect 13682 47966 13694 48018
rect 13746 47966 13758 48018
rect 16258 47966 16270 48018
rect 16322 47966 16334 48018
rect 18834 47966 18846 48018
rect 18898 47966 18910 48018
rect 19506 47966 19518 48018
rect 19570 47966 19582 48018
rect 8542 47954 8594 47966
rect 14814 47954 14866 47966
rect 19182 47954 19234 47966
rect 19854 47954 19906 47966
rect 20078 48018 20130 48030
rect 20078 47954 20130 47966
rect 20750 48018 20802 48030
rect 20750 47954 20802 47966
rect 23326 48018 23378 48030
rect 23326 47954 23378 47966
rect 25566 48018 25618 48030
rect 25566 47954 25618 47966
rect 27806 48018 27858 48030
rect 27806 47954 27858 47966
rect 31838 48018 31890 48030
rect 31838 47954 31890 47966
rect 32398 48018 32450 48030
rect 35310 48018 35362 48030
rect 33506 47966 33518 48018
rect 33570 47966 33582 48018
rect 32398 47954 32450 47966
rect 35310 47954 35362 47966
rect 35422 48018 35474 48030
rect 43486 48018 43538 48030
rect 38658 47966 38670 48018
rect 38722 47966 38734 48018
rect 35422 47954 35474 47966
rect 43486 47954 43538 47966
rect 44046 48018 44098 48030
rect 44046 47954 44098 47966
rect 44270 48018 44322 48030
rect 44270 47954 44322 47966
rect 46510 48018 46562 48030
rect 46510 47954 46562 47966
rect 51550 48018 51602 48030
rect 53790 48018 53842 48030
rect 52658 47966 52670 48018
rect 52722 47966 52734 48018
rect 51550 47954 51602 47966
rect 53790 47954 53842 47966
rect 54350 48018 54402 48030
rect 55346 47966 55358 48018
rect 55410 47966 55422 48018
rect 56354 47966 56366 48018
rect 56418 47966 56430 48018
rect 54350 47954 54402 47966
rect 672 47850 56784 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 44466 47850
rect 44518 47798 44570 47850
rect 44622 47798 44674 47850
rect 44726 47798 56784 47850
rect 672 47764 56784 47798
rect 2830 47682 2882 47694
rect 2830 47618 2882 47630
rect 3390 47682 3442 47694
rect 3390 47618 3442 47630
rect 18062 47682 18114 47694
rect 31390 47682 31442 47694
rect 27682 47630 27694 47682
rect 27746 47630 27758 47682
rect 18062 47618 18114 47630
rect 31390 47618 31442 47630
rect 37886 47682 37938 47694
rect 41358 47682 41410 47694
rect 45726 47682 45778 47694
rect 41010 47630 41022 47682
rect 41074 47630 41086 47682
rect 44258 47630 44270 47682
rect 44322 47630 44334 47682
rect 37886 47618 37938 47630
rect 41358 47618 41410 47630
rect 45726 47618 45778 47630
rect 48078 47682 48130 47694
rect 48078 47618 48130 47630
rect 50766 47682 50818 47694
rect 55122 47630 55134 47682
rect 55186 47630 55198 47682
rect 50766 47618 50818 47630
rect 7758 47570 7810 47582
rect 1586 47518 1598 47570
rect 1650 47518 1662 47570
rect 3714 47518 3726 47570
rect 3778 47518 3790 47570
rect 5058 47518 5070 47570
rect 5122 47518 5134 47570
rect 7758 47506 7810 47518
rect 8318 47570 8370 47582
rect 8318 47506 8370 47518
rect 9102 47570 9154 47582
rect 10558 47570 10610 47582
rect 20302 47570 20354 47582
rect 28142 47570 28194 47582
rect 10098 47518 10110 47570
rect 10162 47518 10174 47570
rect 15138 47518 15150 47570
rect 15202 47518 15214 47570
rect 17154 47518 17166 47570
rect 17218 47518 17230 47570
rect 19058 47518 19070 47570
rect 19122 47518 19134 47570
rect 21746 47518 21758 47570
rect 21810 47518 21822 47570
rect 25330 47518 25342 47570
rect 25394 47518 25406 47570
rect 25666 47518 25678 47570
rect 25730 47518 25742 47570
rect 9102 47506 9154 47518
rect 10558 47506 10610 47518
rect 20302 47506 20354 47518
rect 28142 47506 28194 47518
rect 30382 47570 30434 47582
rect 33966 47570 34018 47582
rect 33058 47518 33070 47570
rect 33122 47518 33134 47570
rect 33394 47518 33406 47570
rect 33458 47518 33470 47570
rect 30382 47506 30434 47518
rect 33966 47506 34018 47518
rect 34526 47570 34578 47582
rect 38334 47570 38386 47582
rect 35634 47518 35646 47570
rect 35698 47518 35710 47570
rect 36642 47518 36654 47570
rect 36706 47518 36718 47570
rect 34526 47506 34578 47518
rect 38334 47506 38386 47518
rect 38446 47570 38498 47582
rect 38446 47506 38498 47518
rect 38558 47570 38610 47582
rect 42030 47570 42082 47582
rect 51214 47570 51266 47582
rect 41682 47518 41694 47570
rect 41746 47518 41758 47570
rect 46834 47518 46846 47570
rect 46898 47518 46910 47570
rect 49522 47518 49534 47570
rect 49586 47518 49598 47570
rect 52210 47518 52222 47570
rect 52274 47518 52286 47570
rect 56354 47518 56366 47570
rect 56418 47518 56430 47570
rect 38558 47506 38610 47518
rect 42030 47506 42082 47518
rect 51214 47506 51266 47518
rect 7982 47458 8034 47470
rect 14702 47458 14754 47470
rect 17726 47458 17778 47470
rect 22430 47458 22482 47470
rect 25006 47458 25058 47470
rect 28366 47458 28418 47470
rect 31166 47458 31218 47470
rect 4386 47406 4398 47458
rect 4450 47406 4462 47458
rect 4946 47406 4958 47458
rect 5010 47406 5022 47458
rect 5618 47406 5630 47458
rect 5682 47406 5694 47458
rect 6178 47406 6190 47458
rect 6242 47406 6254 47458
rect 7074 47406 7086 47458
rect 7138 47406 7150 47458
rect 9426 47406 9438 47458
rect 9490 47406 9502 47458
rect 9874 47406 9886 47458
rect 9938 47406 9950 47458
rect 11330 47406 11342 47458
rect 11394 47406 11406 47458
rect 12114 47406 12126 47458
rect 12178 47406 12190 47458
rect 13010 47406 13022 47458
rect 13074 47406 13086 47458
rect 13906 47406 13918 47458
rect 13970 47406 13982 47458
rect 15250 47406 15262 47458
rect 15314 47406 15326 47458
rect 15698 47406 15710 47458
rect 15762 47406 15774 47458
rect 17266 47406 17278 47458
rect 17330 47406 17342 47458
rect 18722 47406 18734 47458
rect 18786 47406 18798 47458
rect 21074 47406 21086 47458
rect 21138 47406 21150 47458
rect 21634 47406 21646 47458
rect 21698 47406 21710 47458
rect 22754 47406 22766 47458
rect 22818 47406 22830 47458
rect 23762 47406 23774 47458
rect 23826 47406 23838 47458
rect 27010 47406 27022 47458
rect 27074 47406 27086 47458
rect 27570 47406 27582 47458
rect 27634 47406 27646 47458
rect 28690 47406 28702 47458
rect 28754 47406 28766 47458
rect 29698 47406 29710 47458
rect 29762 47406 29774 47458
rect 30706 47406 30718 47458
rect 30770 47406 30782 47458
rect 7982 47394 8034 47406
rect 14702 47394 14754 47406
rect 17726 47394 17778 47406
rect 22430 47394 22482 47406
rect 25006 47394 25058 47406
rect 28366 47394 28418 47406
rect 31166 47394 31218 47406
rect 31278 47458 31330 47470
rect 31278 47394 31330 47406
rect 31614 47458 31666 47470
rect 31614 47394 31666 47406
rect 31838 47458 31890 47470
rect 31838 47394 31890 47406
rect 33630 47458 33682 47470
rect 39118 47458 39170 47470
rect 35298 47406 35310 47458
rect 35362 47406 35374 47458
rect 33630 47394 33682 47406
rect 39118 47394 39170 47406
rect 39454 47458 39506 47470
rect 39454 47394 39506 47406
rect 39566 47458 39618 47470
rect 39566 47394 39618 47406
rect 40238 47458 40290 47470
rect 42366 47458 42418 47470
rect 40786 47406 40798 47458
rect 40850 47406 40862 47458
rect 40238 47394 40290 47406
rect 42366 47394 42418 47406
rect 42478 47458 42530 47470
rect 48302 47458 48354 47470
rect 52894 47458 52946 47470
rect 54798 47458 54850 47470
rect 44818 47406 44830 47458
rect 44882 47406 44894 47458
rect 47394 47406 47406 47458
rect 47458 47406 47470 47458
rect 48626 47406 48638 47458
rect 48690 47406 48702 47458
rect 51538 47406 51550 47458
rect 51602 47406 51614 47458
rect 51986 47406 51998 47458
rect 52050 47406 52062 47458
rect 53442 47406 53454 47458
rect 53506 47406 53518 47458
rect 54338 47406 54350 47458
rect 54402 47406 54414 47458
rect 42478 47394 42530 47406
rect 48302 47394 48354 47406
rect 52894 47394 52946 47406
rect 54798 47394 54850 47406
rect 56030 47458 56082 47470
rect 56030 47394 56082 47406
rect 4062 47346 4114 47358
rect 1250 47294 1262 47346
rect 1314 47294 1326 47346
rect 4062 47282 4114 47294
rect 8206 47346 8258 47358
rect 8206 47282 8258 47294
rect 16158 47346 16210 47358
rect 16158 47282 16210 47294
rect 20750 47346 20802 47358
rect 20750 47282 20802 47294
rect 26686 47346 26738 47358
rect 39230 47346 39282 47358
rect 36306 47294 36318 47346
rect 36370 47294 36382 47346
rect 26686 47282 26738 47294
rect 39230 47282 39282 47294
rect 40350 47346 40402 47358
rect 40350 47282 40402 47294
rect 42142 47346 42194 47358
rect 42142 47282 42194 47294
rect 48190 47346 48242 47358
rect 49186 47294 49198 47346
rect 49250 47294 49262 47346
rect 48190 47282 48242 47294
rect 24670 47234 24722 47246
rect 24670 47170 24722 47182
rect 30718 47234 30770 47246
rect 30718 47170 30770 47182
rect 34862 47234 34914 47246
rect 34862 47170 34914 47182
rect 43150 47234 43202 47246
rect 43150 47170 43202 47182
rect 672 47066 56784 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 43806 47066
rect 43858 47014 43910 47066
rect 43962 47014 44014 47066
rect 44066 47014 56784 47066
rect 672 46980 56784 47014
rect 19182 46898 19234 46910
rect 19182 46834 19234 46846
rect 20750 46898 20802 46910
rect 20750 46834 20802 46846
rect 23326 46898 23378 46910
rect 23326 46834 23378 46846
rect 29262 46898 29314 46910
rect 29262 46834 29314 46846
rect 35086 46898 35138 46910
rect 35086 46834 35138 46846
rect 36430 46898 36482 46910
rect 36430 46834 36482 46846
rect 39790 46898 39842 46910
rect 39790 46834 39842 46846
rect 48750 46898 48802 46910
rect 48750 46834 48802 46846
rect 51326 46898 51378 46910
rect 51326 46834 51378 46846
rect 15150 46786 15202 46798
rect 29150 46786 29202 46798
rect 36766 46786 36818 46798
rect 1250 46734 1262 46786
rect 1314 46734 1326 46786
rect 26226 46734 26238 46786
rect 26290 46734 26302 46786
rect 32946 46734 32958 46786
rect 33010 46734 33022 46786
rect 15150 46722 15202 46734
rect 29150 46722 29202 46734
rect 36766 46722 36818 46734
rect 42702 46786 42754 46798
rect 42702 46722 42754 46734
rect 42926 46786 42978 46798
rect 49746 46734 49758 46786
rect 49810 46734 49822 46786
rect 42926 46722 42978 46734
rect 3838 46674 3890 46686
rect 3838 46610 3890 46622
rect 4286 46674 4338 46686
rect 10110 46674 10162 46686
rect 11790 46674 11842 46686
rect 16606 46674 16658 46686
rect 20862 46674 20914 46686
rect 29598 46674 29650 46686
rect 43150 46674 43202 46686
rect 46398 46674 46450 46686
rect 5282 46622 5294 46674
rect 5346 46622 5358 46674
rect 7522 46622 7534 46674
rect 7586 46622 7598 46674
rect 9874 46622 9886 46674
rect 9938 46622 9950 46674
rect 11106 46622 11118 46674
rect 11170 46622 11182 46674
rect 13122 46622 13134 46674
rect 13186 46622 13198 46674
rect 15474 46622 15486 46674
rect 15538 46622 15550 46674
rect 15922 46622 15934 46674
rect 15986 46622 15998 46674
rect 17266 46622 17278 46674
rect 17330 46622 17342 46674
rect 18162 46622 18174 46674
rect 18226 46622 18238 46674
rect 19842 46622 19854 46674
rect 19906 46622 19918 46674
rect 21634 46622 21646 46674
rect 21698 46622 21710 46674
rect 23874 46622 23886 46674
rect 23938 46622 23950 46674
rect 30258 46622 30270 46674
rect 30322 46622 30334 46674
rect 33394 46622 33406 46674
rect 33458 46622 33470 46674
rect 38210 46622 38222 46674
rect 38274 46622 38286 46674
rect 40674 46622 40686 46674
rect 40738 46622 40750 46674
rect 45938 46622 45950 46674
rect 46002 46622 46014 46674
rect 4286 46610 4338 46622
rect 10110 46610 10162 46622
rect 11790 46610 11842 46622
rect 16606 46610 16658 46622
rect 20862 46610 20914 46622
rect 29598 46610 29650 46622
rect 43150 46610 43202 46622
rect 46398 46610 46450 46622
rect 46734 46674 46786 46686
rect 52334 46674 52386 46686
rect 47058 46622 47070 46674
rect 47122 46622 47134 46674
rect 49634 46622 49646 46674
rect 49698 46622 49710 46674
rect 46734 46610 46786 46622
rect 52334 46610 52386 46622
rect 52446 46674 52498 46686
rect 53790 46674 53842 46686
rect 53330 46622 53342 46674
rect 53394 46622 53406 46674
rect 55346 46622 55358 46674
rect 55410 46622 55422 46674
rect 52446 46610 52498 46622
rect 53790 46610 53842 46622
rect 3278 46562 3330 46574
rect 1586 46510 1598 46562
rect 1650 46510 1662 46562
rect 3278 46498 3330 46510
rect 3390 46562 3442 46574
rect 3390 46498 3442 46510
rect 3950 46562 4002 46574
rect 3950 46498 4002 46510
rect 6862 46562 6914 46574
rect 10558 46562 10610 46574
rect 20750 46562 20802 46574
rect 32622 46562 32674 46574
rect 35758 46562 35810 46574
rect 52670 46562 52722 46574
rect 7970 46510 7982 46562
rect 8034 46510 8046 46562
rect 10994 46510 11006 46562
rect 11058 46510 11070 46562
rect 13570 46510 13582 46562
rect 13634 46510 13646 46562
rect 19954 46510 19966 46562
rect 20018 46510 20030 46562
rect 22082 46510 22094 46562
rect 22146 46510 22158 46562
rect 24434 46510 24446 46562
rect 24498 46510 24510 46562
rect 30706 46510 30718 46562
rect 30770 46510 30782 46562
rect 33842 46510 33854 46562
rect 33906 46510 33918 46562
rect 36978 46510 36990 46562
rect 37042 46510 37054 46562
rect 37314 46510 37326 46562
rect 37378 46510 37390 46562
rect 38546 46510 38558 46562
rect 38610 46510 38622 46562
rect 45490 46510 45502 46562
rect 45554 46510 45566 46562
rect 52994 46510 53006 46562
rect 53058 46510 53070 46562
rect 6862 46498 6914 46510
rect 10558 46498 10610 46510
rect 20750 46498 20802 46510
rect 32622 46498 32674 46510
rect 35758 46498 35810 46510
rect 52670 46498 52722 46510
rect 2830 46450 2882 46462
rect 2830 46386 2882 46398
rect 4062 46450 4114 46462
rect 4062 46386 4114 46398
rect 4174 46450 4226 46462
rect 9102 46450 9154 46462
rect 5730 46398 5742 46450
rect 5794 46398 5806 46450
rect 4174 46386 4226 46398
rect 9102 46386 9154 46398
rect 10222 46450 10274 46462
rect 10222 46386 10274 46398
rect 10334 46450 10386 46462
rect 10334 46386 10386 46398
rect 12126 46450 12178 46462
rect 12126 46386 12178 46398
rect 14702 46450 14754 46462
rect 18846 46450 18898 46462
rect 16146 46398 16158 46450
rect 16210 46398 16222 46450
rect 14702 46386 14754 46398
rect 18846 46386 18898 46398
rect 25566 46450 25618 46462
rect 27806 46450 27858 46462
rect 26674 46398 26686 46450
rect 26738 46398 26750 46450
rect 25566 46386 25618 46398
rect 27806 46386 27858 46398
rect 29710 46450 29762 46462
rect 29710 46386 29762 46398
rect 29934 46450 29986 46462
rect 29934 46386 29986 46398
rect 31950 46450 32002 46462
rect 31950 46386 32002 46398
rect 32846 46450 32898 46462
rect 32846 46386 32898 46398
rect 35422 46450 35474 46462
rect 35422 46386 35474 46398
rect 35646 46450 35698 46462
rect 42254 46450 42306 46462
rect 41122 46398 41134 46450
rect 41186 46398 41198 46450
rect 35646 46386 35698 46398
rect 42254 46386 42306 46398
rect 43262 46450 43314 46462
rect 43262 46386 43314 46398
rect 43374 46450 43426 46462
rect 43374 46386 43426 46398
rect 44270 46450 44322 46462
rect 44270 46386 44322 46398
rect 46510 46450 46562 46462
rect 53118 46450 53170 46462
rect 56030 46450 56082 46462
rect 47618 46398 47630 46450
rect 47682 46398 47694 46450
rect 50194 46398 50206 46450
rect 50258 46398 50270 46450
rect 54898 46398 54910 46450
rect 54962 46398 54974 46450
rect 56354 46398 56366 46450
rect 56418 46398 56430 46450
rect 46510 46386 46562 46398
rect 53118 46386 53170 46398
rect 56030 46386 56082 46398
rect 672 46282 56784 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 44466 46282
rect 44518 46230 44570 46282
rect 44622 46230 44674 46282
rect 44726 46230 56784 46282
rect 672 46196 56784 46230
rect 18510 46114 18562 46126
rect 1362 46062 1374 46114
rect 1426 46062 1438 46114
rect 18510 46050 18562 46062
rect 20302 46114 20354 46126
rect 31166 46114 31218 46126
rect 21746 46062 21758 46114
rect 21810 46062 21822 46114
rect 25330 46062 25342 46114
rect 25394 46062 25406 46114
rect 27906 46062 27918 46114
rect 27970 46062 27982 46114
rect 20302 46050 20354 46062
rect 31166 46050 31218 46062
rect 31278 46114 31330 46126
rect 31278 46050 31330 46062
rect 34750 46114 34802 46126
rect 34750 46050 34802 46062
rect 39118 46114 39170 46126
rect 39118 46050 39170 46062
rect 42590 46114 42642 46126
rect 46062 46114 46114 46126
rect 43810 46062 43822 46114
rect 43874 46062 43886 46114
rect 42590 46050 42642 46062
rect 46062 46050 46114 46062
rect 51438 46114 51490 46126
rect 51438 46050 51490 46062
rect 52446 46114 52498 46126
rect 53554 46062 53566 46114
rect 53618 46062 53630 46114
rect 52446 46050 52498 46062
rect 3054 46002 3106 46014
rect 4510 46002 4562 46014
rect 20750 46002 20802 46014
rect 2034 45950 2046 46002
rect 2098 45950 2110 46002
rect 2706 45950 2718 46002
rect 2770 45950 2782 46002
rect 4050 45950 4062 46002
rect 4114 45950 4126 46002
rect 7970 45950 7982 46002
rect 8034 45950 8046 46002
rect 9874 45950 9886 46002
rect 9938 45950 9950 46002
rect 11554 45950 11566 46002
rect 11618 45950 11630 46002
rect 12450 45950 12462 46002
rect 12514 45950 12526 46002
rect 14578 45950 14590 46002
rect 14642 45950 14654 46002
rect 17378 45950 17390 46002
rect 17442 45950 17454 46002
rect 19282 45950 19294 46002
rect 19346 45950 19358 46002
rect 3054 45938 3106 45950
rect 4510 45938 4562 45950
rect 20750 45938 20802 45950
rect 30606 46002 30658 46014
rect 47406 46002 47458 46014
rect 33618 45950 33630 46002
rect 33682 45950 33694 46002
rect 35858 45950 35870 46002
rect 35922 45950 35934 46002
rect 37426 45950 37438 46002
rect 37490 45950 37502 46002
rect 40786 45950 40798 46002
rect 40850 45950 40862 46002
rect 49074 45950 49086 46002
rect 49138 45950 49150 46002
rect 55906 45950 55918 46002
rect 55970 45950 55982 46002
rect 30606 45938 30658 45950
rect 47406 45938 47458 45950
rect 1038 45890 1090 45902
rect 1038 45826 1090 45838
rect 1710 45890 1762 45902
rect 1710 45826 1762 45838
rect 2382 45890 2434 45902
rect 4734 45890 4786 45902
rect 11006 45890 11058 45902
rect 19966 45890 20018 45902
rect 22430 45890 22482 45902
rect 28366 45890 28418 45902
rect 30494 45890 30546 45902
rect 3378 45838 3390 45890
rect 3442 45838 3454 45890
rect 3826 45838 3838 45890
rect 3890 45838 3902 45890
rect 5058 45838 5070 45890
rect 5122 45838 5134 45890
rect 6178 45838 6190 45890
rect 6242 45838 6254 45890
rect 8194 45838 8206 45890
rect 8258 45838 8270 45890
rect 9986 45838 9998 45890
rect 10050 45838 10062 45890
rect 11442 45838 11454 45890
rect 11506 45838 11518 45890
rect 12338 45838 12350 45890
rect 12402 45838 12414 45890
rect 14018 45838 14030 45890
rect 14082 45838 14094 45890
rect 19394 45838 19406 45890
rect 19458 45838 19470 45890
rect 21074 45838 21086 45890
rect 21138 45838 21150 45890
rect 21634 45838 21646 45890
rect 21698 45838 21710 45890
rect 22754 45838 22766 45890
rect 22818 45838 22830 45890
rect 23874 45838 23886 45890
rect 23938 45838 23950 45890
rect 27234 45838 27246 45890
rect 27298 45838 27310 45890
rect 27682 45838 27694 45890
rect 27746 45838 27758 45890
rect 28914 45838 28926 45890
rect 28978 45838 28990 45890
rect 29922 45838 29934 45890
rect 29986 45838 29998 45890
rect 2382 45826 2434 45838
rect 4734 45826 4786 45838
rect 11006 45826 11058 45838
rect 19966 45826 20018 45838
rect 22430 45826 22482 45838
rect 28366 45826 28418 45838
rect 30494 45826 30546 45838
rect 31390 45890 31442 45902
rect 31390 45826 31442 45838
rect 31614 45890 31666 45902
rect 39230 45890 39282 45902
rect 36978 45838 36990 45890
rect 37042 45838 37054 45890
rect 31614 45826 31666 45838
rect 39230 45826 39282 45838
rect 39342 45890 39394 45902
rect 39342 45826 39394 45838
rect 39790 45890 39842 45902
rect 39790 45826 39842 45838
rect 45614 45890 45666 45902
rect 46286 45890 46338 45902
rect 45938 45838 45950 45890
rect 46002 45838 46014 45890
rect 45614 45826 45666 45838
rect 46286 45826 46338 45838
rect 47182 45890 47234 45902
rect 47182 45826 47234 45838
rect 50318 45890 50370 45902
rect 50318 45826 50370 45838
rect 50766 45890 50818 45902
rect 50766 45826 50818 45838
rect 50990 45890 51042 45902
rect 50990 45826 51042 45838
rect 51214 45890 51266 45902
rect 51214 45826 51266 45838
rect 54574 45890 54626 45902
rect 54574 45826 54626 45838
rect 54798 45890 54850 45902
rect 54798 45826 54850 45838
rect 55134 45890 55186 45902
rect 55134 45826 55186 45838
rect 56254 45890 56306 45902
rect 56254 45826 56306 45838
rect 26910 45778 26962 45790
rect 42702 45778 42754 45790
rect 46174 45778 46226 45790
rect 16930 45726 16942 45778
rect 16994 45726 17006 45778
rect 24882 45726 24894 45778
rect 24946 45726 24958 45778
rect 34066 45726 34078 45778
rect 34130 45726 34142 45778
rect 36306 45726 36318 45778
rect 36370 45726 36382 45778
rect 40450 45726 40462 45778
rect 40514 45726 40526 45778
rect 43362 45726 43374 45778
rect 43426 45726 43438 45778
rect 26910 45714 26962 45726
rect 42702 45714 42754 45726
rect 46174 45714 46226 45726
rect 46958 45778 47010 45790
rect 46958 45714 47010 45726
rect 47294 45778 47346 45790
rect 51326 45778 51378 45790
rect 48738 45726 48750 45778
rect 48802 45726 48814 45778
rect 47294 45714 47346 45726
rect 51326 45714 51378 45726
rect 51998 45778 52050 45790
rect 54686 45778 54738 45790
rect 54002 45726 54014 45778
rect 54066 45726 54078 45778
rect 51998 45714 52050 45726
rect 54686 45714 54738 45726
rect 7086 45666 7138 45678
rect 7086 45602 7138 45614
rect 7422 45666 7474 45678
rect 7422 45602 7474 45614
rect 8990 45666 9042 45678
rect 8990 45602 9042 45614
rect 9326 45666 9378 45678
rect 9326 45602 9378 45614
rect 10670 45666 10722 45678
rect 10670 45602 10722 45614
rect 13134 45666 13186 45678
rect 13134 45602 13186 45614
rect 13470 45666 13522 45678
rect 13470 45602 13522 45614
rect 15710 45666 15762 45678
rect 15710 45602 15762 45614
rect 26462 45666 26514 45678
rect 26462 45602 26514 45614
rect 30606 45666 30658 45678
rect 30606 45602 30658 45614
rect 31838 45666 31890 45678
rect 31838 45602 31890 45614
rect 32510 45666 32562 45678
rect 32510 45602 32562 45614
rect 38670 45666 38722 45678
rect 38670 45602 38722 45614
rect 42030 45666 42082 45678
rect 42030 45602 42082 45614
rect 42814 45666 42866 45678
rect 42814 45602 42866 45614
rect 44942 45666 44994 45678
rect 44942 45602 44994 45614
rect 46734 45666 46786 45678
rect 46734 45602 46786 45614
rect 51886 45666 51938 45678
rect 51886 45602 51938 45614
rect 672 45498 56784 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 43806 45498
rect 43858 45446 43910 45498
rect 43962 45446 44014 45498
rect 44066 45446 56784 45498
rect 672 45412 56784 45446
rect 11006 45330 11058 45342
rect 11006 45266 11058 45278
rect 17726 45330 17778 45342
rect 17726 45266 17778 45278
rect 35310 45330 35362 45342
rect 35310 45266 35362 45278
rect 35646 45330 35698 45342
rect 35646 45266 35698 45278
rect 39118 45330 39170 45342
rect 39118 45266 39170 45278
rect 42590 45330 42642 45342
rect 42590 45266 42642 45278
rect 45950 45330 46002 45342
rect 45950 45266 46002 45278
rect 50878 45330 50930 45342
rect 50878 45266 50930 45278
rect 52446 45330 52498 45342
rect 52446 45266 52498 45278
rect 53790 45330 53842 45342
rect 53790 45266 53842 45278
rect 4398 45218 4450 45230
rect 12910 45218 12962 45230
rect 6514 45166 6526 45218
rect 6578 45166 6590 45218
rect 8866 45166 8878 45218
rect 8930 45166 8942 45218
rect 4398 45154 4450 45166
rect 12910 45154 12962 45166
rect 14030 45218 14082 45230
rect 14030 45154 14082 45166
rect 24222 45218 24274 45230
rect 43150 45218 43202 45230
rect 46510 45218 46562 45230
rect 55806 45218 55858 45230
rect 40002 45166 40014 45218
rect 40066 45166 40078 45218
rect 44370 45166 44382 45218
rect 44434 45166 44446 45218
rect 47058 45166 47070 45218
rect 47122 45166 47134 45218
rect 49298 45166 49310 45218
rect 49362 45166 49374 45218
rect 55346 45166 55358 45218
rect 55410 45166 55422 45218
rect 24222 45154 24274 45166
rect 43150 45154 43202 45166
rect 46510 45154 46562 45166
rect 55806 45154 55858 45166
rect 5294 45106 5346 45118
rect 1250 45054 1262 45106
rect 1314 45054 1326 45106
rect 2146 45054 2158 45106
rect 2210 45054 2222 45106
rect 2818 45054 2830 45106
rect 2882 45054 2894 45106
rect 3490 45054 3502 45106
rect 3554 45054 3566 45106
rect 3938 45054 3950 45106
rect 4002 45054 4014 45106
rect 5294 45042 5346 45054
rect 5518 45106 5570 45118
rect 5518 45042 5570 45054
rect 10110 45106 10162 45118
rect 10110 45042 10162 45054
rect 11342 45106 11394 45118
rect 11342 45042 11394 45054
rect 12686 45106 12738 45118
rect 12686 45042 12738 45054
rect 13022 45106 13074 45118
rect 13022 45042 13074 45054
rect 13246 45106 13298 45118
rect 14466 45054 14478 45106
rect 14530 45054 14542 45106
rect 14802 45057 14814 45109
rect 14866 45057 14878 45109
rect 15710 45106 15762 45118
rect 25678 45106 25730 45118
rect 42142 45106 42194 45118
rect 43038 45106 43090 45118
rect 16034 45054 16046 45106
rect 16098 45054 16110 45106
rect 17042 45054 17054 45106
rect 17106 45054 17118 45106
rect 19282 45054 19294 45106
rect 19346 45054 19358 45106
rect 22194 45054 22206 45106
rect 22258 45054 22270 45106
rect 24658 45054 24670 45106
rect 24722 45054 24734 45106
rect 24994 45054 25006 45106
rect 25058 45054 25070 45106
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 27346 45054 27358 45106
rect 27410 45054 27422 45106
rect 30146 45054 30158 45106
rect 30210 45054 30222 45106
rect 30930 45054 30942 45106
rect 30994 45054 31006 45106
rect 33170 45054 33182 45106
rect 33234 45054 33246 45106
rect 37426 45054 37438 45106
rect 37490 45054 37502 45106
rect 40562 45054 40574 45106
rect 40626 45054 40638 45106
rect 42914 45054 42926 45106
rect 42978 45054 42990 45106
rect 13246 45042 13298 45054
rect 15710 45042 15762 45054
rect 25678 45042 25730 45054
rect 42142 45042 42194 45054
rect 43038 45042 43090 45054
rect 46398 45106 46450 45118
rect 56030 45106 56082 45118
rect 49186 45054 49198 45106
rect 49250 45054 49262 45106
rect 52882 45054 52894 45106
rect 52946 45054 52958 45106
rect 46398 45042 46450 45054
rect 56030 45042 56082 45054
rect 4958 44994 5010 45006
rect 3378 44942 3390 44994
rect 3442 44942 3454 44994
rect 4958 44930 5010 44942
rect 5966 44994 6018 45006
rect 8542 44994 8594 45006
rect 6850 44942 6862 44994
rect 6914 44942 6926 44994
rect 5966 44930 6018 44942
rect 8542 44930 8594 44942
rect 8766 44994 8818 45006
rect 39678 44994 39730 45006
rect 9314 44942 9326 44994
rect 9378 44942 9390 44994
rect 9874 44942 9886 44994
rect 9938 44942 9950 44994
rect 11554 44942 11566 44994
rect 11618 44942 11630 44994
rect 12114 44942 12126 44994
rect 12178 44942 12190 44994
rect 22530 44942 22542 44994
rect 22594 44942 22606 44994
rect 29810 44942 29822 44994
rect 29874 44942 29886 44994
rect 33506 44942 33518 44994
rect 33570 44942 33582 44994
rect 37874 44942 37886 44994
rect 37938 44942 37950 44994
rect 8766 44930 8818 44942
rect 39678 44930 39730 44942
rect 39902 44994 39954 45006
rect 39902 44930 39954 44942
rect 51326 44994 51378 45006
rect 56366 44994 56418 45006
rect 53218 44942 53230 44994
rect 53282 44942 53294 44994
rect 51326 44930 51378 44942
rect 56366 44930 56418 44942
rect 5070 44882 5122 44894
rect 5070 44818 5122 44830
rect 5854 44882 5906 44894
rect 5854 44818 5906 44830
rect 8094 44882 8146 44894
rect 8094 44818 8146 44830
rect 10446 44882 10498 44894
rect 23774 44882 23826 44894
rect 28590 44882 28642 44894
rect 32510 44882 32562 44894
rect 15026 44830 15038 44882
rect 15090 44830 15102 44882
rect 18834 44830 18846 44882
rect 18898 44830 18910 44882
rect 25218 44830 25230 44882
rect 25282 44830 25294 44882
rect 31378 44830 31390 44882
rect 31442 44830 31454 44882
rect 10446 44818 10498 44830
rect 23774 44818 23826 44830
rect 28590 44818 28642 44830
rect 32510 44818 32562 44830
rect 34750 44882 34802 44894
rect 34750 44818 34802 44830
rect 35534 44882 35586 44894
rect 35534 44818 35586 44830
rect 36654 44882 36706 44894
rect 43262 44882 43314 44894
rect 48638 44882 48690 44894
rect 51438 44882 51490 44894
rect 36978 44830 36990 44882
rect 37042 44830 37054 44882
rect 41010 44830 41022 44882
rect 41074 44830 41086 44882
rect 44818 44830 44830 44882
rect 44882 44830 44894 44882
rect 47506 44830 47518 44882
rect 47570 44830 47582 44882
rect 49746 44830 49758 44882
rect 49810 44830 49822 44882
rect 36654 44818 36706 44830
rect 43262 44818 43314 44830
rect 48638 44818 48690 44830
rect 51438 44818 51490 44830
rect 52110 44882 52162 44894
rect 56254 44882 56306 44894
rect 54898 44830 54910 44882
rect 54962 44830 54974 44882
rect 52110 44818 52162 44830
rect 56254 44818 56306 44830
rect 672 44714 56784 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 44466 44714
rect 44518 44662 44570 44714
rect 44622 44662 44674 44714
rect 44726 44662 56784 44714
rect 672 44628 56784 44662
rect 16606 44546 16658 44558
rect 5506 44494 5518 44546
rect 5570 44494 5582 44546
rect 16606 44482 16658 44494
rect 16830 44546 16882 44558
rect 19406 44546 19458 44558
rect 18274 44494 18286 44546
rect 18338 44494 18350 44546
rect 16830 44482 16882 44494
rect 19406 44482 19458 44494
rect 21646 44546 21698 44558
rect 31278 44546 31330 44558
rect 27906 44494 27918 44546
rect 27970 44494 27982 44546
rect 21646 44482 21698 44494
rect 31278 44482 31330 44494
rect 31390 44546 31442 44558
rect 31390 44482 31442 44494
rect 37326 44546 37378 44558
rect 37326 44482 37378 44494
rect 37438 44546 37490 44558
rect 42366 44546 42418 44558
rect 38770 44494 38782 44546
rect 38834 44494 38846 44546
rect 37438 44482 37490 44494
rect 42366 44482 42418 44494
rect 50094 44546 50146 44558
rect 50094 44482 50146 44494
rect 50654 44546 50706 44558
rect 50654 44482 50706 44494
rect 4510 44434 4562 44446
rect 1810 44382 1822 44434
rect 1874 44382 1886 44434
rect 4510 44370 4562 44382
rect 8206 44434 8258 44446
rect 16942 44434 16994 44446
rect 23886 44434 23938 44446
rect 30606 44434 30658 44446
rect 9538 44382 9550 44434
rect 9602 44382 9614 44434
rect 12674 44382 12686 44434
rect 12738 44382 12750 44434
rect 14802 44382 14814 44434
rect 14866 44382 14878 44434
rect 20514 44382 20526 44434
rect 20578 44382 20590 44434
rect 22754 44382 22766 44434
rect 22818 44382 22830 44434
rect 25218 44382 25230 44434
rect 25282 44382 25294 44434
rect 8206 44370 8258 44382
rect 16942 44370 16994 44382
rect 23886 44370 23938 44382
rect 30606 44370 30658 44382
rect 31166 44434 31218 44446
rect 37550 44434 37602 44446
rect 33618 44382 33630 44434
rect 33682 44382 33694 44434
rect 35186 44382 35198 44434
rect 35250 44382 35262 44434
rect 31166 44370 31218 44382
rect 37550 44370 37602 44382
rect 38446 44434 38498 44446
rect 42926 44434 42978 44446
rect 38658 44382 38670 44434
rect 38722 44382 38734 44434
rect 41122 44382 41134 44434
rect 41186 44382 41198 44434
rect 43810 44382 43822 44434
rect 43874 44382 43886 44434
rect 46274 44382 46286 44434
rect 46338 44382 46350 44434
rect 48962 44382 48974 44434
rect 49026 44382 49038 44434
rect 51762 44382 51774 44434
rect 51826 44382 51838 44434
rect 52882 44382 52894 44434
rect 52946 44382 52958 44434
rect 53442 44382 53454 44434
rect 53506 44382 53518 44434
rect 55346 44382 55358 44434
rect 55410 44382 55422 44434
rect 56354 44382 56366 44434
rect 56418 44382 56430 44434
rect 38446 44370 38498 44382
rect 42926 44370 42978 44382
rect 3726 44322 3778 44334
rect 3726 44258 3778 44270
rect 3950 44322 4002 44334
rect 3950 44258 4002 44270
rect 4286 44322 4338 44334
rect 6190 44322 6242 44334
rect 8094 44322 8146 44334
rect 4834 44270 4846 44322
rect 4898 44270 4910 44322
rect 5282 44270 5294 44322
rect 5346 44270 5358 44322
rect 6626 44270 6638 44322
rect 6690 44270 6702 44322
rect 7522 44270 7534 44322
rect 7586 44270 7598 44322
rect 4286 44258 4338 44270
rect 6190 44258 6242 44270
rect 8094 44258 8146 44270
rect 11342 44322 11394 44334
rect 30494 44322 30546 44334
rect 14354 44270 14366 44322
rect 14418 44270 14430 44322
rect 17826 44270 17838 44322
rect 17890 44270 17902 44322
rect 22194 44270 22206 44322
rect 22258 44270 22270 44322
rect 27234 44270 27246 44322
rect 27298 44270 27310 44322
rect 27682 44270 27694 44322
rect 27746 44270 27758 44322
rect 28466 44270 28478 44322
rect 28530 44270 28542 44322
rect 28914 44270 28926 44322
rect 28978 44270 28990 44322
rect 29922 44270 29934 44322
rect 29986 44270 29998 44322
rect 11342 44258 11394 44270
rect 30494 44258 30546 44270
rect 31614 44322 31666 44334
rect 31614 44258 31666 44270
rect 31838 44322 31890 44334
rect 37102 44322 37154 44334
rect 34066 44270 34078 44322
rect 34130 44270 34142 44322
rect 34850 44270 34862 44322
rect 34914 44270 34926 44322
rect 31838 44258 31890 44270
rect 37102 44258 37154 44270
rect 38894 44322 38946 44334
rect 38894 44258 38946 44270
rect 39342 44322 39394 44334
rect 50990 44322 51042 44334
rect 54350 44322 54402 44334
rect 40674 44270 40686 44322
rect 40738 44270 40750 44322
rect 45826 44270 45838 44322
rect 45890 44270 45902 44322
rect 51426 44270 51438 44322
rect 51490 44270 51502 44322
rect 39342 44258 39394 44270
rect 50990 44258 51042 44270
rect 54350 44258 54402 44270
rect 54574 44322 54626 44334
rect 54574 44258 54626 44270
rect 55022 44322 55074 44334
rect 56130 44270 56142 44322
rect 56194 44270 56206 44322
rect 55022 44258 55074 44270
rect 4062 44210 4114 44222
rect 26910 44210 26962 44222
rect 1474 44158 1486 44210
rect 1538 44158 1550 44210
rect 9090 44158 9102 44210
rect 9154 44158 9166 44210
rect 12226 44158 12238 44210
rect 12290 44158 12302 44210
rect 20066 44158 20078 44210
rect 20130 44158 20142 44210
rect 24882 44158 24894 44210
rect 24946 44158 24958 44210
rect 4062 44146 4114 44158
rect 3054 44098 3106 44110
rect 3054 44034 3106 44046
rect 8206 44098 8258 44110
rect 8206 44034 8258 44046
rect 10670 44098 10722 44110
rect 11106 44102 11118 44154
rect 11170 44102 11182 44154
rect 26910 44146 26962 44158
rect 38110 44210 38162 44222
rect 38110 44146 38162 44158
rect 39118 44210 39170 44222
rect 54126 44210 54178 44222
rect 43474 44158 43486 44210
rect 43538 44158 43550 44210
rect 48514 44158 48526 44210
rect 48578 44158 48590 44210
rect 39118 44146 39170 44158
rect 54126 44146 54178 44158
rect 54462 44210 54514 44222
rect 54462 44146 54514 44158
rect 13806 44098 13858 44110
rect 11666 44046 11678 44098
rect 11730 44046 11742 44098
rect 10670 44034 10722 44046
rect 13806 44034 13858 44046
rect 16046 44098 16098 44110
rect 16046 44034 16098 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 30606 44098 30658 44110
rect 30606 44034 30658 44046
rect 32510 44098 32562 44110
rect 32510 44034 32562 44046
rect 36430 44098 36482 44110
rect 36430 44034 36482 44046
rect 36878 44098 36930 44110
rect 36878 44034 36930 44046
rect 37998 44098 38050 44110
rect 37998 44034 38050 44046
rect 42814 44098 42866 44110
rect 42814 44034 42866 44046
rect 45054 44098 45106 44110
rect 45054 44034 45106 44046
rect 47406 44098 47458 44110
rect 47406 44034 47458 44046
rect 52334 44098 52386 44110
rect 52334 44034 52386 44046
rect 52670 44098 52722 44110
rect 52670 44034 52722 44046
rect 53902 44098 53954 44110
rect 53902 44034 53954 44046
rect 672 43930 56784 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 43806 43930
rect 43858 43878 43910 43930
rect 43962 43878 44014 43930
rect 44066 43878 56784 43930
rect 672 43844 56784 43878
rect 45054 43762 45106 43774
rect 45054 43698 45106 43710
rect 3166 43650 3218 43662
rect 3166 43586 3218 43598
rect 5182 43650 5234 43662
rect 5182 43586 5234 43598
rect 10782 43650 10834 43662
rect 10782 43586 10834 43598
rect 11342 43650 11394 43662
rect 11342 43586 11394 43598
rect 12238 43650 12290 43662
rect 12238 43586 12290 43598
rect 15598 43650 15650 43662
rect 15598 43586 15650 43598
rect 16382 43650 16434 43662
rect 16382 43586 16434 43598
rect 16830 43650 16882 43662
rect 34750 43650 34802 43662
rect 41694 43650 41746 43662
rect 28690 43598 28702 43650
rect 28754 43598 28766 43650
rect 33170 43598 33182 43650
rect 33234 43598 33246 43650
rect 39666 43598 39678 43650
rect 39730 43598 39742 43650
rect 41234 43598 41246 43650
rect 41298 43598 41310 43650
rect 16830 43586 16882 43598
rect 34750 43586 34802 43598
rect 41694 43586 41746 43598
rect 43374 43650 43426 43662
rect 43374 43586 43426 43598
rect 43598 43650 43650 43662
rect 48178 43598 48190 43650
rect 48242 43598 48254 43650
rect 43598 43586 43650 43598
rect 4062 43538 4114 43550
rect 5518 43538 5570 43550
rect 11790 43538 11842 43550
rect 15374 43538 15426 43550
rect 1474 43486 1486 43538
rect 1538 43486 1550 43538
rect 3602 43486 3614 43538
rect 3666 43486 3678 43538
rect 4274 43486 4286 43538
rect 4338 43486 4350 43538
rect 6178 43486 6190 43538
rect 6242 43486 6254 43538
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 9090 43486 9102 43538
rect 9154 43486 9166 43538
rect 13234 43486 13246 43538
rect 13298 43486 13310 43538
rect 4062 43474 4114 43486
rect 5518 43474 5570 43486
rect 11790 43474 11842 43486
rect 15374 43474 15426 43486
rect 15822 43538 15874 43550
rect 35534 43538 35586 43550
rect 44494 43538 44546 43550
rect 45166 43538 45218 43550
rect 17154 43486 17166 43538
rect 17218 43486 17230 43538
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 19058 43486 19070 43538
rect 19122 43486 19134 43538
rect 19842 43486 19854 43538
rect 19906 43486 19918 43538
rect 22194 43486 22206 43538
rect 22258 43486 22270 43538
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 24994 43486 25006 43538
rect 25058 43486 25070 43538
rect 26338 43486 26350 43538
rect 26402 43486 26414 43538
rect 27234 43486 27246 43538
rect 27298 43486 27310 43538
rect 32498 43486 32510 43538
rect 32562 43486 32574 43538
rect 35186 43486 35198 43538
rect 35250 43486 35262 43538
rect 37314 43486 37326 43538
rect 37378 43486 37390 43538
rect 42242 43486 42254 43538
rect 42306 43486 42318 43538
rect 44818 43486 44830 43538
rect 44882 43486 44894 43538
rect 15822 43474 15874 43486
rect 35534 43474 35586 43486
rect 44494 43474 44546 43486
rect 45166 43474 45218 43486
rect 49198 43538 49250 43550
rect 49198 43474 49250 43486
rect 50542 43538 50594 43550
rect 50542 43474 50594 43486
rect 50766 43538 50818 43550
rect 50766 43474 50818 43486
rect 52110 43538 52162 43550
rect 52110 43474 52162 43486
rect 52558 43538 52610 43550
rect 52558 43474 52610 43486
rect 52782 43538 52834 43550
rect 54114 43486 54126 43538
rect 54178 43486 54190 43538
rect 52782 43474 52834 43486
rect 11230 43426 11282 43438
rect 6290 43374 6302 43426
rect 6354 43374 6366 43426
rect 7410 43374 7422 43426
rect 7474 43374 7486 43426
rect 11230 43362 11282 43374
rect 11566 43426 11618 43438
rect 16046 43426 16098 43438
rect 13682 43374 13694 43426
rect 13746 43374 13758 43426
rect 11566 43362 11618 43374
rect 16046 43362 16098 43374
rect 16494 43426 16546 43438
rect 16494 43362 16546 43374
rect 18286 43426 18338 43438
rect 18286 43362 18338 43374
rect 24222 43426 24274 43438
rect 24222 43362 24274 43374
rect 25678 43426 25730 43438
rect 35646 43426 35698 43438
rect 39342 43426 39394 43438
rect 32050 43374 32062 43426
rect 32114 43374 32126 43426
rect 33506 43374 33518 43426
rect 33570 43374 33582 43426
rect 36754 43374 36766 43426
rect 36818 43374 36830 43426
rect 25678 43362 25730 43374
rect 35646 43362 35698 43374
rect 39342 43362 39394 43374
rect 39678 43426 39730 43438
rect 40462 43426 40514 43438
rect 39778 43374 39790 43426
rect 39842 43374 39854 43426
rect 39678 43362 39730 43374
rect 40462 43362 40514 43374
rect 40798 43426 40850 43438
rect 41918 43426 41970 43438
rect 40898 43374 40910 43426
rect 40962 43374 40974 43426
rect 40798 43362 40850 43374
rect 41918 43362 41970 43374
rect 43150 43426 43202 43438
rect 43150 43362 43202 43374
rect 44158 43426 44210 43438
rect 44158 43362 44210 43374
rect 45502 43426 45554 43438
rect 51102 43426 51154 43438
rect 47842 43374 47854 43426
rect 47906 43374 47918 43426
rect 49410 43374 49422 43426
rect 49474 43374 49486 43426
rect 49746 43374 49758 43426
rect 49810 43374 49822 43426
rect 45502 43362 45554 43374
rect 51102 43362 51154 43374
rect 51326 43426 51378 43438
rect 51326 43362 51378 43374
rect 51998 43426 52050 43438
rect 51998 43362 52050 43374
rect 52334 43426 52386 43438
rect 55806 43426 55858 43438
rect 54562 43374 54574 43426
rect 54626 43374 54638 43426
rect 52334 43362 52386 43374
rect 55806 43362 55858 43374
rect 56366 43426 56418 43438
rect 56366 43362 56418 43374
rect 3838 43314 3890 43326
rect 2034 43262 2046 43314
rect 2098 43262 2110 43314
rect 3838 43250 3890 43262
rect 3950 43314 4002 43326
rect 3950 43250 4002 43262
rect 8542 43314 8594 43326
rect 12126 43314 12178 43326
rect 9650 43262 9662 43314
rect 9714 43262 9726 43314
rect 8542 43250 8594 43262
rect 12126 43250 12178 43262
rect 14926 43314 14978 43326
rect 23774 43314 23826 43326
rect 30270 43314 30322 43326
rect 17826 43262 17838 43314
rect 17890 43262 17902 43314
rect 22642 43262 22654 43314
rect 22706 43262 22718 43314
rect 25218 43262 25230 43314
rect 25282 43262 25294 43314
rect 29138 43262 29150 43314
rect 29202 43262 29214 43314
rect 14926 43250 14978 43262
rect 23774 43250 23826 43262
rect 30270 43250 30322 43262
rect 30830 43314 30882 43326
rect 30830 43250 30882 43262
rect 35758 43314 35810 43326
rect 35758 43250 35810 43262
rect 36430 43314 36482 43326
rect 38894 43314 38946 43326
rect 37762 43262 37774 43314
rect 37826 43262 37838 43314
rect 36430 43250 36482 43262
rect 38894 43250 38946 43262
rect 39566 43314 39618 43326
rect 39566 43250 39618 43262
rect 40686 43314 40738 43326
rect 40686 43250 40738 43262
rect 41582 43314 41634 43326
rect 41582 43250 41634 43262
rect 41806 43314 41858 43326
rect 41806 43250 41858 43262
rect 42926 43314 42978 43326
rect 42926 43250 42978 43262
rect 43038 43314 43090 43326
rect 43038 43250 43090 43262
rect 44270 43314 44322 43326
rect 44270 43250 44322 43262
rect 45390 43314 45442 43326
rect 45390 43250 45442 43262
rect 45838 43314 45890 43326
rect 46622 43314 46674 43326
rect 46162 43262 46174 43314
rect 46226 43262 46238 43314
rect 45838 43250 45890 43262
rect 46622 43250 46674 43262
rect 48862 43314 48914 43326
rect 48862 43250 48914 43262
rect 50430 43314 50482 43326
rect 53566 43314 53618 43326
rect 53218 43262 53230 43314
rect 53282 43262 53294 43314
rect 50430 43250 50482 43262
rect 53566 43250 53618 43262
rect 56254 43314 56306 43326
rect 56254 43250 56306 43262
rect 672 43146 56784 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 44466 43146
rect 44518 43094 44570 43146
rect 44622 43094 44674 43146
rect 44726 43094 56784 43146
rect 672 43060 56784 43094
rect 8206 42978 8258 42990
rect 1810 42926 1822 42978
rect 1874 42926 1886 42978
rect 4386 42926 4398 42978
rect 4450 42926 4462 42978
rect 8206 42914 8258 42926
rect 10446 42978 10498 42990
rect 36430 42978 36482 42990
rect 45054 42978 45106 42990
rect 12674 42926 12686 42978
rect 12738 42926 12750 42978
rect 27458 42926 27470 42978
rect 27522 42926 27534 42978
rect 35298 42926 35310 42978
rect 35362 42926 35374 42978
rect 37538 42926 37550 42978
rect 37602 42926 37614 42978
rect 39106 42926 39118 42978
rect 39170 42926 39182 42978
rect 43922 42926 43934 42978
rect 43986 42926 43998 42978
rect 10446 42914 10498 42926
rect 36430 42914 36482 42926
rect 45054 42914 45106 42926
rect 46286 42978 46338 42990
rect 55234 42926 55246 42978
rect 55298 42926 55310 42978
rect 46286 42914 46338 42926
rect 4846 42866 4898 42878
rect 9550 42866 9602 42878
rect 7186 42814 7198 42866
rect 7250 42814 7262 42866
rect 7522 42814 7534 42866
rect 7586 42814 7598 42866
rect 4846 42802 4898 42814
rect 9550 42802 9602 42814
rect 9774 42866 9826 42878
rect 19742 42866 19794 42878
rect 27918 42866 27970 42878
rect 47406 42866 47458 42878
rect 53678 42866 53730 42878
rect 10994 42814 11006 42866
rect 11058 42814 11070 42866
rect 11442 42814 11454 42866
rect 11506 42814 11518 42866
rect 14914 42814 14926 42866
rect 14978 42814 14990 42866
rect 18050 42814 18062 42866
rect 18114 42814 18126 42866
rect 20738 42814 20750 42866
rect 20802 42814 20814 42866
rect 30706 42814 30718 42866
rect 30770 42814 30782 42866
rect 33618 42814 33630 42866
rect 33682 42814 33694 42866
rect 41234 42814 41246 42866
rect 41298 42814 41310 42866
rect 45714 42814 45726 42866
rect 45778 42814 45790 42866
rect 49970 42814 49982 42866
rect 50034 42814 50046 42866
rect 53890 42814 53902 42866
rect 53954 42814 53966 42866
rect 56354 42814 56366 42866
rect 56418 42814 56430 42866
rect 9774 42802 9826 42814
rect 19742 42802 19794 42814
rect 27918 42802 27970 42814
rect 47406 42802 47458 42814
rect 53678 42802 53730 42814
rect 7870 42754 7922 42766
rect 3714 42702 3726 42754
rect 3778 42702 3790 42754
rect 4274 42702 4286 42754
rect 4338 42702 4350 42754
rect 5394 42702 5406 42754
rect 5458 42702 5470 42754
rect 6402 42702 6414 42754
rect 6466 42702 6478 42754
rect 7870 42690 7922 42702
rect 8990 42754 9042 42766
rect 21422 42754 21474 42766
rect 38670 42754 38722 42766
rect 11554 42702 11566 42754
rect 11618 42702 11630 42754
rect 14354 42702 14366 42754
rect 14418 42702 14430 42754
rect 17602 42702 17614 42754
rect 17666 42702 17678 42754
rect 20066 42702 20078 42754
rect 20130 42702 20142 42754
rect 20514 42702 20526 42754
rect 20578 42702 20590 42754
rect 21746 42702 21758 42754
rect 21810 42702 21822 42754
rect 22754 42702 22766 42754
rect 22818 42702 22830 42754
rect 26786 42702 26798 42754
rect 26850 42702 26862 42754
rect 27234 42702 27246 42754
rect 27298 42702 27310 42754
rect 28690 42702 28702 42754
rect 28754 42702 28766 42754
rect 29474 42702 29486 42754
rect 29538 42702 29550 42754
rect 30818 42702 30830 42754
rect 30882 42702 30894 42754
rect 34850 42702 34862 42754
rect 34914 42702 34926 42754
rect 37090 42702 37102 42754
rect 37154 42702 37166 42754
rect 8990 42690 9042 42702
rect 21422 42690 21474 42702
rect 38670 42690 38722 42702
rect 39454 42754 39506 42766
rect 45502 42754 45554 42766
rect 43362 42702 43374 42754
rect 43426 42702 43438 42754
rect 39454 42690 39506 42702
rect 45502 42690 45554 42702
rect 45950 42754 46002 42766
rect 46846 42754 46898 42766
rect 46050 42702 46062 42754
rect 46114 42702 46126 42754
rect 46610 42702 46622 42754
rect 46674 42702 46686 42754
rect 45950 42690 46002 42702
rect 46846 42690 46898 42702
rect 47070 42754 47122 42766
rect 47070 42690 47122 42702
rect 47294 42754 47346 42766
rect 54126 42754 54178 42766
rect 52098 42702 52110 42754
rect 52162 42702 52174 42754
rect 47294 42690 47346 42702
rect 54126 42690 54178 42702
rect 54350 42754 54402 42766
rect 54910 42754 54962 42766
rect 54350 42690 54402 42702
rect 54574 42698 54626 42710
rect 3390 42642 3442 42654
rect 16046 42642 16098 42654
rect 26462 42642 26514 42654
rect 39678 42642 39730 42654
rect 42814 42642 42866 42654
rect 1362 42590 1374 42642
rect 1426 42590 1438 42642
rect 12226 42590 12238 42642
rect 12290 42590 12302 42642
rect 17714 42590 17726 42642
rect 17778 42590 17790 42642
rect 34066 42590 34078 42642
rect 34130 42590 34142 42642
rect 40786 42590 40798 42642
rect 40850 42590 40862 42642
rect 3390 42578 3442 42590
rect 16046 42578 16098 42590
rect 26462 42578 26514 42590
rect 39678 42578 39730 42590
rect 42814 42578 42866 42590
rect 54462 42642 54514 42654
rect 54910 42690 54962 42702
rect 56030 42754 56082 42766
rect 56030 42690 56082 42702
rect 54574 42634 54626 42646
rect 54462 42578 54514 42590
rect 2942 42530 2994 42542
rect 2942 42466 2994 42478
rect 9214 42530 9266 42542
rect 9214 42466 9266 42478
rect 9662 42530 9714 42542
rect 9662 42466 9714 42478
rect 10782 42530 10834 42542
rect 10782 42466 10834 42478
rect 13806 42530 13858 42542
rect 13806 42466 13858 42478
rect 19294 42530 19346 42542
rect 19294 42466 19346 42478
rect 31390 42530 31442 42542
rect 31390 42466 31442 42478
rect 31726 42530 31778 42542
rect 31726 42466 31778 42478
rect 32510 42530 32562 42542
rect 32510 42466 32562 42478
rect 42366 42530 42418 42542
rect 42366 42466 42418 42478
rect 42926 42530 42978 42542
rect 42926 42466 42978 42478
rect 672 42362 56784 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 43806 42362
rect 43858 42310 43910 42362
rect 43962 42310 44014 42362
rect 44066 42310 56784 42362
rect 672 42276 56784 42310
rect 5854 42194 5906 42206
rect 5854 42130 5906 42142
rect 6190 42194 6242 42206
rect 6190 42130 6242 42142
rect 8990 42194 9042 42206
rect 8990 42130 9042 42142
rect 36766 42194 36818 42206
rect 36766 42130 36818 42142
rect 43262 42194 43314 42206
rect 43262 42130 43314 42142
rect 43598 42194 43650 42206
rect 43598 42130 43650 42142
rect 50430 42194 50482 42206
rect 50430 42130 50482 42142
rect 54014 42194 54066 42206
rect 54014 42130 54066 42142
rect 54574 42194 54626 42206
rect 54574 42130 54626 42142
rect 30606 42082 30658 42094
rect 38110 42082 38162 42094
rect 42254 42082 42306 42094
rect 6850 42030 6862 42082
rect 6914 42030 6926 42082
rect 9202 42030 9214 42082
rect 9266 42030 9278 42082
rect 35746 42030 35758 42082
rect 35810 42030 35822 42082
rect 39218 42030 39230 42082
rect 39282 42030 39294 42082
rect 51202 42030 51214 42082
rect 51266 42030 51278 42082
rect 56130 42030 56142 42082
rect 56194 42030 56206 42082
rect 30606 42018 30658 42030
rect 38110 42018 38162 42030
rect 42254 42018 42306 42030
rect 3278 41970 3330 41982
rect 1250 41918 1262 41970
rect 1314 41918 1326 41970
rect 3278 41906 3330 41918
rect 3614 41970 3666 41982
rect 3614 41906 3666 41918
rect 3726 41970 3778 41982
rect 3726 41906 3778 41918
rect 4062 41970 4114 41982
rect 4062 41906 4114 41918
rect 4286 41970 4338 41982
rect 12126 41970 12178 41982
rect 9314 41918 9326 41970
rect 9378 41918 9390 41970
rect 10434 41918 10446 41970
rect 10498 41918 10510 41970
rect 4286 41906 4338 41918
rect 12126 41906 12178 41918
rect 12798 41970 12850 41982
rect 12798 41906 12850 41918
rect 12910 41970 12962 41982
rect 14814 41970 14866 41982
rect 16830 41970 16882 41982
rect 18286 41970 18338 41982
rect 21646 41970 21698 41982
rect 32286 41970 32338 41982
rect 34974 41970 35026 41982
rect 38222 41970 38274 41982
rect 13346 41918 13358 41970
rect 13410 41918 13422 41970
rect 14242 41918 14254 41970
rect 14306 41918 14318 41970
rect 15698 41918 15710 41970
rect 15762 41918 15774 41970
rect 16146 41918 16158 41970
rect 16210 41918 16222 41970
rect 17154 41918 17166 41970
rect 17218 41918 17230 41970
rect 17602 41918 17614 41970
rect 17666 41918 17678 41970
rect 19058 41918 19070 41970
rect 19122 41918 19134 41970
rect 19954 41918 19966 41970
rect 20018 41918 20030 41970
rect 21970 41918 21982 41970
rect 22034 41918 22046 41970
rect 22530 41918 22542 41970
rect 22594 41918 22606 41970
rect 23650 41918 23662 41970
rect 23714 41918 23726 41970
rect 24770 41918 24782 41970
rect 24834 41918 24846 41970
rect 25442 41918 25454 41970
rect 25506 41918 25518 41970
rect 31042 41918 31054 41970
rect 31106 41918 31118 41970
rect 31490 41918 31502 41970
rect 31554 41918 31566 41970
rect 32610 41918 32622 41970
rect 32674 41918 32686 41970
rect 33618 41918 33630 41970
rect 33682 41918 33694 41970
rect 35410 41918 35422 41970
rect 35474 41918 35486 41970
rect 35634 41918 35646 41970
rect 35698 41918 35710 41970
rect 38546 41918 38558 41970
rect 38610 41918 38622 41970
rect 45938 41918 45950 41970
rect 46002 41918 46014 41970
rect 48066 41918 48078 41970
rect 48130 41918 48142 41970
rect 48738 41918 48750 41970
rect 48802 41918 48814 41970
rect 52434 41918 52446 41970
rect 52498 41918 52510 41970
rect 12910 41906 12962 41918
rect 14814 41906 14866 41918
rect 16830 41906 16882 41918
rect 18286 41906 18338 41918
rect 21646 41906 21698 41918
rect 32286 41906 32338 41918
rect 34974 41906 35026 41918
rect 38222 41906 38274 41918
rect 3390 41858 3442 41870
rect 16494 41858 16546 41870
rect 1586 41806 1598 41858
rect 1650 41806 1662 41858
rect 5282 41806 5294 41858
rect 5346 41806 5358 41858
rect 5618 41806 5630 41858
rect 5682 41806 5694 41858
rect 9986 41806 9998 41858
rect 10050 41806 10062 41858
rect 10882 41806 10894 41858
rect 10946 41806 10958 41858
rect 15474 41806 15486 41858
rect 15538 41806 15550 41858
rect 3390 41794 3442 41806
rect 16494 41794 16546 41806
rect 23102 41858 23154 41870
rect 34414 41858 34466 41870
rect 31602 41806 31614 41858
rect 31666 41806 31678 41858
rect 23102 41794 23154 41806
rect 34414 41794 34466 41806
rect 34526 41858 34578 41870
rect 34526 41794 34578 41806
rect 35198 41858 35250 41870
rect 42590 41858 42642 41870
rect 36978 41806 36990 41858
rect 37042 41806 37054 41858
rect 37426 41806 37438 41858
rect 37490 41806 37502 41858
rect 41570 41806 41582 41858
rect 41634 41806 41646 41858
rect 41906 41806 41918 41858
rect 41970 41806 41982 41858
rect 35198 41794 35250 41806
rect 42590 41794 42642 41806
rect 43038 41858 43090 41870
rect 43038 41794 43090 41806
rect 51438 41858 51490 41870
rect 51438 41794 51490 41806
rect 2830 41746 2882 41758
rect 2830 41682 2882 41694
rect 4062 41746 4114 41758
rect 8430 41746 8482 41758
rect 7298 41694 7310 41746
rect 7362 41694 7374 41746
rect 4062 41682 4114 41694
rect 8430 41682 8482 41694
rect 9662 41746 9714 41758
rect 27022 41746 27074 41758
rect 10994 41694 11006 41746
rect 11058 41694 11070 41746
rect 17826 41694 17838 41746
rect 17890 41694 17902 41746
rect 22642 41694 22654 41746
rect 22706 41694 22718 41746
rect 25890 41694 25902 41746
rect 25954 41694 25966 41746
rect 9662 41682 9714 41694
rect 27022 41682 27074 41694
rect 34750 41746 34802 41758
rect 34750 41682 34802 41694
rect 36430 41746 36482 41758
rect 36430 41682 36482 41694
rect 37998 41746 38050 41758
rect 40798 41746 40850 41758
rect 39666 41694 39678 41746
rect 39730 41694 39742 41746
rect 37998 41682 38050 41694
rect 40798 41682 40850 41694
rect 44270 41746 44322 41758
rect 46510 41746 46562 41758
rect 51214 41746 51266 41758
rect 45378 41694 45390 41746
rect 45442 41694 45454 41746
rect 47618 41694 47630 41746
rect 47682 41694 47694 41746
rect 49298 41694 49310 41746
rect 49362 41694 49374 41746
rect 52882 41694 52894 41746
rect 52946 41694 52958 41746
rect 55682 41694 55694 41746
rect 55746 41694 55758 41746
rect 44270 41682 44322 41694
rect 46510 41682 46562 41694
rect 51214 41682 51266 41694
rect 672 41578 56784 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 44466 41578
rect 44518 41526 44570 41578
rect 44622 41526 44674 41578
rect 44726 41526 56784 41578
rect 672 41492 56784 41526
rect 12798 41410 12850 41422
rect 20190 41410 20242 41422
rect 37102 41410 37154 41422
rect 2258 41358 2270 41410
rect 2322 41358 2334 41410
rect 7074 41358 7086 41410
rect 7138 41358 7150 41410
rect 8082 41358 8094 41410
rect 8146 41358 8158 41410
rect 12450 41358 12462 41410
rect 12514 41358 12526 41410
rect 13122 41358 13134 41410
rect 13186 41358 13198 41410
rect 26338 41358 26350 41410
rect 26402 41358 26414 41410
rect 28914 41358 28926 41410
rect 28978 41358 28990 41410
rect 33394 41358 33406 41410
rect 33458 41358 33470 41410
rect 12798 41346 12850 41358
rect 20190 41346 20242 41358
rect 37102 41346 37154 41358
rect 37326 41410 37378 41422
rect 42590 41410 42642 41422
rect 38434 41358 38446 41410
rect 38498 41358 38510 41410
rect 40898 41358 40910 41410
rect 40962 41358 40974 41410
rect 37326 41346 37378 41358
rect 42590 41346 42642 41358
rect 43262 41410 43314 41422
rect 43262 41346 43314 41358
rect 43822 41410 43874 41422
rect 43822 41346 43874 41358
rect 46286 41410 46338 41422
rect 46286 41346 46338 41358
rect 48190 41410 48242 41422
rect 48190 41346 48242 41358
rect 48302 41410 48354 41422
rect 48302 41346 48354 41358
rect 48526 41410 48578 41422
rect 49970 41358 49982 41410
rect 50034 41358 50046 41410
rect 56242 41358 56254 41410
rect 56306 41358 56318 41410
rect 48526 41346 48578 41358
rect 10334 41298 10386 41310
rect 16046 41298 16098 41310
rect 20638 41298 20690 41310
rect 22094 41298 22146 41310
rect 48078 41298 48130 41310
rect 4498 41246 4510 41298
rect 4562 41246 4574 41298
rect 9874 41246 9886 41298
rect 9938 41246 9950 41298
rect 14802 41246 14814 41298
rect 14866 41246 14878 41298
rect 17378 41246 17390 41298
rect 17442 41246 17454 41298
rect 17938 41246 17950 41298
rect 18002 41246 18014 41298
rect 18946 41246 18958 41298
rect 19010 41246 19022 41298
rect 21634 41246 21646 41298
rect 21698 41246 21710 41298
rect 26226 41246 26238 41298
rect 26290 41246 26302 41298
rect 35634 41246 35646 41298
rect 35698 41246 35710 41298
rect 44930 41246 44942 41298
rect 44994 41246 45006 41298
rect 47170 41246 47182 41298
rect 47234 41246 47246 41298
rect 50194 41246 50206 41298
rect 50258 41246 50270 41298
rect 51314 41246 51326 41298
rect 51378 41246 51390 41298
rect 53554 41246 53566 41298
rect 53618 41246 53630 41298
rect 10334 41234 10386 41246
rect 16046 41234 16098 41246
rect 20638 41234 20690 41246
rect 22094 41234 22146 41246
rect 48078 41234 48130 41246
rect 7758 41186 7810 41198
rect 29598 41186 29650 41198
rect 37438 41186 37490 41198
rect 42478 41186 42530 41198
rect 2706 41134 2718 41186
rect 2770 41134 2782 41186
rect 3826 41134 3838 41186
rect 3890 41134 3902 41186
rect 4274 41134 4286 41186
rect 4338 41134 4350 41186
rect 5058 41134 5070 41186
rect 5122 41134 5134 41186
rect 5506 41134 5518 41186
rect 5570 41134 5582 41186
rect 6514 41134 6526 41186
rect 6578 41134 6590 41186
rect 7298 41134 7310 41186
rect 7362 41134 7374 41186
rect 9314 41134 9326 41186
rect 9378 41134 9390 41186
rect 9762 41134 9774 41186
rect 9826 41134 9838 41186
rect 10434 41134 10446 41186
rect 10498 41134 10510 41186
rect 11106 41134 11118 41186
rect 11170 41134 11182 41186
rect 12002 41134 12014 41186
rect 12066 41134 12078 41186
rect 13346 41134 13358 41186
rect 13410 41134 13422 41186
rect 14354 41134 14366 41186
rect 14418 41134 14430 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 20962 41134 20974 41186
rect 21026 41134 21038 41186
rect 21522 41134 21534 41186
rect 21586 41134 21598 41186
rect 22642 41134 22654 41186
rect 22706 41134 22718 41186
rect 23650 41134 23662 41186
rect 23714 41134 23726 41186
rect 25778 41134 25790 41186
rect 25842 41134 25854 41186
rect 28354 41134 28366 41186
rect 28418 41134 28430 41186
rect 28690 41134 28702 41186
rect 28754 41134 28766 41186
rect 30034 41134 30046 41186
rect 30098 41134 30110 41186
rect 30930 41134 30942 41186
rect 30994 41134 31006 41186
rect 32946 41134 32958 41186
rect 33010 41134 33022 41186
rect 35074 41134 35086 41186
rect 35138 41134 35150 41186
rect 37874 41134 37886 41186
rect 37938 41134 37950 41186
rect 40338 41134 40350 41186
rect 40402 41134 40414 41186
rect 7758 41122 7810 41134
rect 29598 41122 29650 41134
rect 37438 41122 37490 41134
rect 42478 41122 42530 41134
rect 42814 41186 42866 41198
rect 46622 41186 46674 41198
rect 50430 41186 50482 41198
rect 55358 41186 55410 41198
rect 43026 41134 43038 41186
rect 43090 41134 43102 41186
rect 45378 41134 45390 41186
rect 45442 41134 45454 41186
rect 47394 41134 47406 41186
rect 47458 41134 47470 41186
rect 49298 41134 49310 41186
rect 49362 41134 49374 41186
rect 49634 41134 49646 41186
rect 49698 41134 49710 41186
rect 50866 41134 50878 41186
rect 50930 41134 50942 41186
rect 42814 41122 42866 41134
rect 46622 41122 46674 41134
rect 50430 41122 50482 41134
rect 55358 41122 55410 41134
rect 55918 41186 55970 41198
rect 55918 41122 55970 41134
rect 3502 41074 3554 41086
rect 3502 41010 3554 41022
rect 8878 41074 8930 41086
rect 8878 41010 8930 41022
rect 27918 41074 27970 41086
rect 49982 41074 50034 41086
rect 49186 41022 49198 41074
rect 49250 41022 49262 41074
rect 27918 41010 27970 41022
rect 49982 41010 50034 41022
rect 52558 41074 52610 41086
rect 53218 41022 53230 41074
rect 53282 41022 53294 41074
rect 52558 41010 52610 41022
rect 1150 40962 1202 40974
rect 1150 40898 1202 40910
rect 16830 40962 16882 40974
rect 16830 40898 16882 40910
rect 17166 40962 17218 40974
rect 17166 40898 17218 40910
rect 27470 40962 27522 40974
rect 27470 40898 27522 40910
rect 34526 40962 34578 40974
rect 34526 40898 34578 40910
rect 36766 40962 36818 40974
rect 36766 40898 36818 40910
rect 39566 40962 39618 40974
rect 39566 40898 39618 40910
rect 42030 40962 42082 40974
rect 42030 40898 42082 40910
rect 43374 40962 43426 40974
rect 43374 40898 43426 40910
rect 48974 40962 49026 40974
rect 48974 40898 49026 40910
rect 54798 40962 54850 40974
rect 54798 40898 54850 40910
rect 55246 40962 55298 40974
rect 55246 40898 55298 40910
rect 672 40794 56784 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 43806 40794
rect 43858 40742 43910 40794
rect 43962 40742 44014 40794
rect 44066 40742 56784 40794
rect 672 40708 56784 40742
rect 30494 40626 30546 40638
rect 30494 40562 30546 40574
rect 42926 40626 42978 40638
rect 42926 40562 42978 40574
rect 8318 40514 8370 40526
rect 21982 40514 22034 40526
rect 30942 40514 30994 40526
rect 5394 40462 5406 40514
rect 5458 40462 5470 40514
rect 6290 40462 6302 40514
rect 6354 40462 6366 40514
rect 18386 40462 18398 40514
rect 18450 40462 18462 40514
rect 28914 40462 28926 40514
rect 28978 40462 28990 40514
rect 8318 40450 8370 40462
rect 21982 40450 22034 40462
rect 30942 40450 30994 40462
rect 42814 40514 42866 40526
rect 51214 40514 51266 40526
rect 46610 40462 46622 40514
rect 46674 40462 46686 40514
rect 52210 40462 52222 40514
rect 52274 40462 52286 40514
rect 55906 40462 55918 40514
rect 55970 40462 55982 40514
rect 42814 40450 42866 40462
rect 51214 40450 51266 40462
rect 2606 40402 2658 40414
rect 5518 40402 5570 40414
rect 9774 40402 9826 40414
rect 12238 40402 12290 40414
rect 19966 40402 20018 40414
rect 23438 40402 23490 40414
rect 32398 40402 32450 40414
rect 36318 40402 36370 40414
rect 1586 40350 1598 40402
rect 1650 40350 1662 40402
rect 1922 40350 1934 40402
rect 1986 40350 1998 40402
rect 3154 40350 3166 40402
rect 3218 40350 3230 40402
rect 4162 40350 4174 40402
rect 4226 40350 4238 40402
rect 4946 40350 4958 40402
rect 5010 40350 5022 40402
rect 8754 40350 8766 40402
rect 8818 40350 8830 40402
rect 9090 40350 9102 40402
rect 9154 40350 9166 40402
rect 10322 40350 10334 40402
rect 10386 40350 10398 40402
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 13906 40350 13918 40402
rect 13970 40350 13982 40402
rect 14466 40350 14478 40402
rect 14530 40350 14542 40402
rect 15138 40350 15150 40402
rect 15202 40350 15214 40402
rect 15586 40350 15598 40402
rect 15650 40350 15662 40402
rect 16706 40350 16718 40402
rect 16770 40350 16782 40402
rect 22306 40350 22318 40402
rect 22370 40350 22382 40402
rect 22754 40350 22766 40402
rect 22818 40350 22830 40402
rect 24098 40350 24110 40402
rect 24162 40350 24174 40402
rect 24994 40350 25006 40402
rect 25058 40350 25070 40402
rect 26226 40350 26238 40402
rect 26290 40350 26302 40402
rect 31266 40350 31278 40402
rect 31330 40350 31342 40402
rect 31714 40350 31726 40402
rect 31778 40350 31790 40402
rect 32946 40350 32958 40402
rect 33010 40350 33022 40402
rect 33954 40350 33966 40402
rect 34018 40350 34030 40402
rect 35074 40350 35086 40402
rect 35138 40350 35150 40402
rect 2606 40338 2658 40350
rect 5518 40338 5570 40350
rect 9774 40338 9826 40350
rect 12238 40338 12290 40350
rect 19966 40338 20018 40350
rect 23438 40338 23490 40350
rect 32398 40338 32450 40350
rect 36318 40338 36370 40350
rect 36654 40402 36706 40414
rect 38782 40402 38834 40414
rect 37202 40350 37214 40402
rect 37266 40350 37278 40402
rect 39554 40350 39566 40402
rect 39618 40350 39630 40402
rect 36654 40338 36706 40350
rect 38782 40338 38834 40350
rect 40114 40344 40126 40396
rect 40178 40344 40190 40396
rect 40786 40350 40798 40402
rect 40850 40350 40862 40402
rect 41234 40350 41246 40402
rect 41298 40350 41310 40402
rect 42354 40350 42366 40402
rect 42418 40350 42430 40402
rect 43362 40350 43374 40402
rect 43426 40350 43438 40402
rect 44370 40350 44382 40402
rect 44434 40350 44446 40402
rect 48850 40350 48862 40402
rect 48914 40350 48926 40402
rect 1150 40290 1202 40302
rect 1150 40226 1202 40238
rect 5182 40290 5234 40302
rect 13582 40290 13634 40302
rect 35422 40290 35474 40302
rect 9314 40238 9326 40290
rect 9378 40238 9390 40290
rect 11890 40238 11902 40290
rect 11954 40238 11966 40290
rect 12786 40238 12798 40290
rect 12850 40238 12862 40290
rect 14578 40238 14590 40290
rect 14642 40238 14654 40290
rect 18834 40238 18846 40290
rect 18898 40238 18910 40290
rect 22978 40238 22990 40290
rect 23042 40238 23054 40290
rect 29362 40238 29374 40290
rect 29426 40238 29438 40290
rect 31938 40238 31950 40290
rect 32002 40238 32014 40290
rect 5182 40226 5234 40238
rect 13582 40226 13634 40238
rect 35422 40226 35474 40238
rect 35758 40290 35810 40302
rect 35758 40226 35810 40238
rect 36430 40290 36482 40302
rect 39230 40290 39282 40302
rect 51326 40290 51378 40302
rect 37538 40238 37550 40290
rect 37602 40238 37614 40290
rect 40226 40238 40238 40290
rect 40290 40238 40302 40290
rect 49298 40238 49310 40290
rect 49362 40238 49374 40290
rect 36430 40226 36482 40238
rect 39230 40226 39282 40238
rect 51326 40226 51378 40238
rect 5406 40178 5458 40190
rect 7870 40178 7922 40190
rect 2146 40126 2158 40178
rect 2210 40126 2222 40178
rect 6738 40126 6750 40178
rect 6802 40126 6814 40178
rect 5406 40114 5458 40126
rect 7870 40114 7922 40126
rect 13134 40178 13186 40190
rect 27806 40178 27858 40190
rect 26674 40126 26686 40178
rect 26738 40126 26750 40178
rect 13134 40114 13186 40126
rect 27806 40114 27858 40126
rect 35534 40178 35586 40190
rect 35534 40114 35586 40126
rect 35646 40178 35698 40190
rect 45950 40178 46002 40190
rect 48190 40178 48242 40190
rect 43586 40126 43598 40178
rect 43650 40126 43662 40178
rect 44818 40126 44830 40178
rect 44882 40126 44894 40178
rect 47058 40126 47070 40178
rect 47122 40126 47134 40178
rect 35646 40114 35698 40126
rect 45950 40114 46002 40126
rect 48190 40114 48242 40126
rect 50430 40178 50482 40190
rect 50430 40114 50482 40126
rect 50878 40178 50930 40190
rect 50878 40114 50930 40126
rect 51102 40178 51154 40190
rect 53790 40178 53842 40190
rect 52658 40126 52670 40178
rect 52722 40126 52734 40178
rect 51102 40114 51154 40126
rect 53790 40114 53842 40126
rect 54350 40178 54402 40190
rect 55458 40126 55470 40178
rect 55522 40126 55534 40178
rect 54350 40114 54402 40126
rect 672 40010 56784 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 44466 40010
rect 44518 39958 44570 40010
rect 44622 39958 44674 40010
rect 44726 39958 56784 40010
rect 672 39924 56784 39958
rect 1038 39842 1090 39854
rect 1710 39842 1762 39854
rect 2718 39842 2770 39854
rect 6862 39842 6914 39854
rect 1362 39790 1374 39842
rect 1426 39790 1438 39842
rect 2034 39790 2046 39842
rect 2098 39790 2110 39842
rect 3938 39790 3950 39842
rect 4002 39790 4014 39842
rect 6514 39790 6526 39842
rect 6578 39790 6590 39842
rect 1038 39778 1090 39790
rect 1710 39778 1762 39790
rect 2718 39778 2770 39790
rect 6862 39778 6914 39790
rect 7310 39842 7362 39854
rect 16158 39842 16210 39854
rect 13458 39790 13470 39842
rect 13522 39790 13534 39842
rect 7310 39778 7362 39790
rect 16158 39778 16210 39790
rect 20078 39842 20130 39854
rect 36430 39842 36482 39854
rect 21522 39790 21534 39842
rect 21586 39790 21598 39842
rect 27458 39790 27470 39842
rect 27522 39790 27534 39842
rect 33618 39790 33630 39842
rect 33682 39790 33694 39842
rect 20078 39778 20130 39790
rect 36430 39778 36482 39790
rect 39566 39842 39618 39854
rect 39566 39778 39618 39790
rect 39790 39842 39842 39854
rect 48414 39842 48466 39854
rect 53566 39842 53618 39854
rect 41234 39790 41246 39842
rect 41298 39790 41310 39842
rect 45042 39790 45054 39842
rect 45106 39790 45118 39842
rect 47506 39790 47518 39842
rect 47570 39790 47582 39842
rect 49298 39790 49310 39842
rect 49362 39790 49374 39842
rect 39790 39778 39842 39790
rect 48414 39778 48466 39790
rect 53566 39778 53618 39790
rect 54574 39842 54626 39854
rect 56242 39790 56254 39842
rect 56306 39790 56318 39842
rect 54574 39778 54626 39790
rect 2382 39730 2434 39742
rect 2382 39666 2434 39678
rect 2494 39730 2546 39742
rect 2494 39666 2546 39678
rect 7198 39730 7250 39742
rect 7198 39666 7250 39678
rect 8878 39730 8930 39742
rect 39454 39730 39506 39742
rect 9874 39678 9886 39730
rect 9938 39678 9950 39730
rect 18834 39678 18846 39730
rect 18898 39678 18910 39730
rect 30146 39678 30158 39730
rect 30210 39678 30222 39730
rect 35186 39678 35198 39730
rect 35250 39678 35262 39730
rect 37762 39678 37774 39730
rect 37826 39678 37838 39730
rect 8878 39666 8930 39678
rect 39454 39666 39506 39678
rect 40238 39730 40290 39742
rect 40238 39666 40290 39678
rect 48190 39730 48242 39742
rect 51538 39678 51550 39730
rect 51602 39678 51614 39730
rect 48190 39666 48242 39678
rect 4622 39618 4674 39630
rect 7870 39618 7922 39630
rect 3266 39566 3278 39618
rect 3330 39566 3342 39618
rect 3714 39566 3726 39618
rect 3778 39566 3790 39618
rect 4946 39566 4958 39618
rect 5010 39566 5022 39618
rect 6066 39566 6078 39618
rect 6130 39566 6142 39618
rect 4622 39554 4674 39566
rect 7870 39554 7922 39566
rect 7982 39618 8034 39630
rect 7982 39554 8034 39566
rect 8430 39618 8482 39630
rect 41918 39618 41970 39630
rect 46174 39618 46226 39630
rect 9202 39566 9214 39618
rect 9266 39566 9278 39618
rect 9762 39566 9774 39618
rect 9826 39566 9838 39618
rect 10434 39566 10446 39618
rect 10498 39566 10510 39618
rect 10882 39566 10894 39618
rect 10946 39566 10958 39618
rect 11890 39566 11902 39618
rect 11954 39566 11966 39618
rect 12898 39566 12910 39618
rect 12962 39566 12974 39618
rect 18498 39566 18510 39618
rect 18562 39566 18574 39618
rect 20850 39566 20862 39618
rect 20914 39566 20926 39618
rect 21410 39566 21422 39618
rect 21474 39566 21486 39618
rect 22082 39566 22094 39618
rect 22146 39566 22158 39618
rect 22530 39566 22542 39618
rect 22594 39566 22606 39618
rect 23538 39566 23550 39618
rect 23602 39566 23614 39618
rect 26898 39566 26910 39618
rect 26962 39566 26974 39618
rect 27234 39566 27246 39618
rect 27298 39566 27310 39618
rect 28018 39566 28030 39618
rect 28082 39566 28094 39618
rect 28690 39566 28702 39618
rect 28754 39566 28766 39618
rect 29474 39566 29486 39618
rect 29538 39566 29550 39618
rect 30370 39566 30382 39618
rect 30434 39566 30446 39618
rect 34066 39566 34078 39618
rect 34130 39566 34142 39618
rect 34850 39566 34862 39618
rect 34914 39566 34926 39618
rect 37314 39566 37326 39618
rect 37378 39566 37390 39618
rect 40562 39566 40574 39618
rect 40626 39566 40638 39618
rect 41010 39566 41022 39618
rect 41074 39566 41086 39618
rect 42242 39566 42254 39618
rect 42306 39566 42318 39618
rect 43250 39566 43262 39618
rect 43314 39566 43326 39618
rect 45490 39566 45502 39618
rect 45554 39566 45566 39618
rect 8430 39554 8482 39566
rect 41918 39554 41970 39566
rect 46174 39554 46226 39566
rect 46398 39618 46450 39630
rect 46398 39554 46450 39566
rect 47182 39618 47234 39630
rect 47182 39554 47234 39566
rect 48078 39618 48130 39630
rect 53678 39618 53730 39630
rect 48850 39566 48862 39618
rect 48914 39566 48926 39618
rect 50978 39566 50990 39618
rect 51042 39566 51054 39618
rect 48078 39554 48130 39566
rect 53678 39554 53730 39566
rect 53790 39618 53842 39630
rect 53790 39554 53842 39566
rect 54350 39618 54402 39630
rect 54350 39554 54402 39566
rect 54798 39618 54850 39630
rect 54798 39554 54850 39566
rect 55022 39618 55074 39630
rect 56018 39566 56030 39618
rect 56082 39566 56094 39618
rect 55022 39554 55074 39566
rect 2942 39506 2994 39518
rect 2942 39442 2994 39454
rect 8206 39506 8258 39518
rect 8206 39442 8258 39454
rect 16046 39506 16098 39518
rect 16046 39442 16098 39454
rect 20526 39506 20578 39518
rect 20526 39442 20578 39454
rect 26462 39506 26514 39518
rect 26462 39442 26514 39454
rect 53342 39506 53394 39518
rect 53342 39442 53394 39454
rect 54462 39506 54514 39518
rect 54462 39442 54514 39454
rect 7310 39394 7362 39406
rect 7310 39330 7362 39342
rect 14590 39394 14642 39406
rect 14590 39330 14642 39342
rect 30942 39394 30994 39406
rect 30942 39330 30994 39342
rect 31278 39394 31330 39406
rect 31278 39330 31330 39342
rect 32510 39394 32562 39406
rect 32510 39330 32562 39342
rect 39006 39394 39058 39406
rect 39006 39330 39058 39342
rect 43934 39394 43986 39406
rect 50430 39394 50482 39406
rect 46722 39342 46734 39394
rect 46786 39342 46798 39394
rect 43934 39330 43986 39342
rect 50430 39330 50482 39342
rect 52670 39394 52722 39406
rect 52670 39330 52722 39342
rect 53118 39394 53170 39406
rect 53118 39330 53170 39342
rect 672 39226 56784 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 43806 39226
rect 43858 39174 43910 39226
rect 43962 39174 44014 39226
rect 44066 39174 56784 39226
rect 672 39140 56784 39174
rect 11790 39058 11842 39070
rect 11790 38994 11842 39006
rect 30382 39058 30434 39070
rect 30382 38994 30434 39006
rect 35646 39058 35698 39070
rect 35646 38994 35698 39006
rect 43486 39058 43538 39070
rect 43486 38994 43538 39006
rect 48190 39058 48242 39070
rect 48190 38994 48242 39006
rect 51998 39058 52050 39070
rect 51998 38994 52050 39006
rect 53342 39058 53394 39070
rect 53342 38994 53394 39006
rect 11902 38946 11954 38958
rect 1250 38894 1262 38946
rect 1314 38894 1326 38946
rect 11902 38882 11954 38894
rect 14366 38946 14418 38958
rect 35758 38946 35810 38958
rect 21298 38894 21310 38946
rect 21362 38894 21374 38946
rect 23538 38894 23550 38946
rect 23602 38894 23614 38946
rect 31378 38894 31390 38946
rect 31442 38894 31454 38946
rect 35074 38894 35086 38946
rect 35138 38894 35150 38946
rect 14366 38882 14418 38894
rect 35758 38882 35810 38894
rect 36766 38946 36818 38958
rect 50766 38946 50818 38958
rect 39666 38894 39678 38946
rect 39730 38894 39742 38946
rect 44370 38894 44382 38946
rect 44434 38894 44446 38946
rect 46610 38894 46622 38946
rect 46674 38894 46686 38946
rect 36766 38882 36818 38894
rect 50766 38882 50818 38894
rect 52222 38946 52274 38958
rect 52222 38882 52274 38894
rect 53118 38946 53170 38958
rect 53118 38882 53170 38894
rect 53678 38946 53730 38958
rect 53678 38882 53730 38894
rect 55694 38946 55746 38958
rect 55694 38882 55746 38894
rect 3278 38834 3330 38846
rect 3278 38770 3330 38782
rect 3838 38834 3890 38846
rect 3838 38770 3890 38782
rect 4174 38834 4226 38846
rect 4174 38770 4226 38782
rect 4398 38834 4450 38846
rect 4398 38770 4450 38782
rect 5294 38834 5346 38846
rect 8206 38834 8258 38846
rect 9662 38834 9714 38846
rect 12686 38834 12738 38846
rect 6066 38782 6078 38834
rect 6130 38782 6142 38834
rect 8642 38782 8654 38834
rect 8706 38782 8718 38834
rect 9090 38782 9102 38834
rect 9154 38782 9166 38834
rect 10322 38782 10334 38834
rect 10386 38782 10398 38834
rect 11330 38782 11342 38834
rect 11394 38782 11406 38834
rect 5294 38770 5346 38782
rect 8206 38770 8258 38782
rect 9662 38770 9714 38782
rect 12686 38770 12738 38782
rect 13022 38834 13074 38846
rect 15822 38834 15874 38846
rect 36206 38834 36258 38846
rect 14802 38782 14814 38834
rect 14866 38782 14878 38834
rect 15250 38782 15262 38834
rect 15314 38782 15326 38834
rect 16594 38782 16606 38834
rect 16658 38782 16670 38834
rect 17490 38782 17502 38834
rect 17554 38782 17566 38834
rect 18274 38782 18286 38834
rect 18338 38782 18350 38834
rect 26226 38782 26238 38834
rect 26290 38782 26302 38834
rect 28690 38782 28702 38834
rect 28754 38782 28766 38834
rect 13022 38770 13074 38782
rect 15822 38770 15874 38782
rect 36206 38770 36258 38782
rect 36654 38834 36706 38846
rect 36654 38770 36706 38782
rect 36878 38834 36930 38846
rect 49086 38834 49138 38846
rect 37314 38782 37326 38834
rect 37378 38782 37390 38834
rect 41906 38782 41918 38834
rect 41970 38782 41982 38834
rect 36878 38770 36930 38782
rect 49086 38770 49138 38782
rect 50542 38834 50594 38846
rect 50542 38770 50594 38782
rect 51214 38834 51266 38846
rect 51214 38770 51266 38782
rect 52446 38834 52498 38846
rect 52446 38770 52498 38782
rect 52670 38834 52722 38846
rect 52670 38770 52722 38782
rect 54014 38834 54066 38846
rect 54014 38770 54066 38782
rect 55582 38834 55634 38846
rect 55582 38770 55634 38782
rect 55806 38834 55858 38846
rect 55806 38770 55858 38782
rect 3390 38722 3442 38734
rect 55246 38722 55298 38734
rect 1698 38670 1710 38722
rect 1762 38670 1774 38722
rect 4946 38670 4958 38722
rect 5010 38670 5022 38722
rect 6626 38670 6638 38722
rect 6690 38670 6702 38722
rect 9202 38670 9214 38722
rect 9266 38670 9278 38722
rect 18834 38670 18846 38722
rect 18898 38670 18910 38722
rect 21634 38670 21646 38722
rect 21698 38670 21710 38722
rect 23986 38670 23998 38722
rect 24050 38670 24062 38722
rect 26674 38670 26686 38722
rect 26738 38670 26750 38722
rect 29250 38670 29262 38722
rect 29314 38670 29326 38722
rect 34626 38670 34638 38722
rect 34690 38670 34702 38722
rect 37874 38670 37886 38722
rect 37938 38670 37950 38722
rect 40002 38670 40014 38722
rect 40066 38670 40078 38722
rect 42354 38670 42366 38722
rect 42418 38670 42430 38722
rect 44706 38670 44718 38722
rect 44770 38670 44782 38722
rect 46946 38670 46958 38722
rect 47010 38670 47022 38722
rect 49410 38670 49422 38722
rect 49474 38670 49486 38722
rect 49858 38670 49870 38722
rect 49922 38670 49934 38722
rect 54338 38670 54350 38722
rect 54402 38670 54414 38722
rect 54898 38670 54910 38722
rect 54962 38670 54974 38722
rect 3390 38658 3442 38670
rect 55246 38658 55298 38670
rect 2830 38610 2882 38622
rect 2830 38546 2882 38558
rect 3614 38610 3666 38622
rect 3614 38546 3666 38558
rect 4062 38610 4114 38622
rect 4062 38546 4114 38558
rect 7758 38610 7810 38622
rect 7758 38546 7810 38558
rect 12910 38610 12962 38622
rect 19966 38610 20018 38622
rect 15362 38558 15374 38610
rect 15426 38558 15438 38610
rect 12910 38546 12962 38558
rect 19966 38546 20018 38558
rect 22878 38610 22930 38622
rect 22878 38546 22930 38558
rect 25118 38610 25170 38622
rect 25118 38546 25170 38558
rect 27806 38610 27858 38622
rect 32958 38610 33010 38622
rect 31826 38558 31838 38610
rect 31890 38558 31902 38610
rect 27806 38546 27858 38558
rect 32958 38546 33010 38558
rect 33518 38610 33570 38622
rect 33518 38546 33570 38558
rect 39006 38610 39058 38622
rect 39006 38546 39058 38558
rect 41246 38610 41298 38622
rect 41246 38546 41298 38558
rect 45950 38610 46002 38622
rect 45950 38546 46002 38558
rect 48750 38610 48802 38622
rect 48750 38546 48802 38558
rect 50990 38610 51042 38622
rect 50990 38546 51042 38558
rect 51102 38610 51154 38622
rect 51102 38546 51154 38558
rect 52558 38610 52610 38622
rect 52558 38546 52610 38558
rect 54686 38610 54738 38622
rect 54686 38546 54738 38558
rect 56030 38610 56082 38622
rect 56030 38546 56082 38558
rect 672 38442 56784 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 44466 38442
rect 44518 38390 44570 38442
rect 44622 38390 44674 38442
rect 44726 38390 56784 38442
rect 672 38356 56784 38390
rect 7086 38274 7138 38286
rect 7086 38210 7138 38222
rect 7310 38274 7362 38286
rect 7310 38210 7362 38222
rect 9550 38274 9602 38286
rect 9550 38210 9602 38222
rect 12126 38274 12178 38286
rect 22766 38274 22818 38286
rect 48190 38274 48242 38286
rect 13234 38222 13246 38274
rect 13298 38222 13310 38274
rect 26450 38222 26462 38274
rect 26514 38222 26526 38274
rect 29250 38222 29262 38274
rect 29314 38222 29326 38274
rect 33618 38222 33630 38274
rect 33682 38222 33694 38274
rect 41458 38222 41470 38274
rect 41522 38222 41534 38274
rect 44930 38222 44942 38274
rect 44994 38222 45006 38274
rect 12126 38210 12178 38222
rect 22766 38210 22818 38222
rect 48190 38210 48242 38222
rect 50430 38274 50482 38286
rect 50430 38210 50482 38222
rect 7422 38162 7474 38174
rect 1586 38110 1598 38162
rect 1650 38110 1662 38162
rect 4610 38110 4622 38162
rect 4674 38110 4686 38162
rect 7422 38098 7474 38110
rect 7758 38162 7810 38174
rect 7758 38098 7810 38110
rect 8318 38162 8370 38174
rect 8318 38098 8370 38110
rect 8878 38162 8930 38174
rect 8878 38098 8930 38110
rect 8990 38162 9042 38174
rect 18846 38162 18898 38174
rect 20302 38162 20354 38174
rect 29710 38162 29762 38174
rect 10994 38110 11006 38162
rect 11058 38110 11070 38162
rect 15138 38110 15150 38162
rect 15202 38110 15214 38162
rect 19842 38110 19854 38162
rect 19906 38110 19918 38162
rect 23874 38110 23886 38162
rect 23938 38110 23950 38162
rect 8990 38098 9042 38110
rect 18846 38098 18898 38110
rect 20302 38098 20354 38110
rect 29710 38098 29762 38110
rect 34078 38162 34130 38174
rect 47294 38162 47346 38174
rect 37538 38110 37550 38162
rect 37602 38110 37614 38162
rect 34078 38098 34130 38110
rect 47294 38098 47346 38110
rect 48078 38162 48130 38174
rect 49298 38110 49310 38162
rect 49362 38110 49374 38162
rect 51762 38110 51774 38162
rect 51826 38110 51838 38162
rect 54114 38110 54126 38162
rect 54178 38110 54190 38162
rect 56354 38110 56366 38162
rect 56418 38110 56430 38162
rect 48078 38098 48130 38110
rect 3614 38050 3666 38062
rect 8094 38050 8146 38062
rect 1250 37998 1262 38050
rect 1314 37998 1326 38050
rect 3938 37998 3950 38050
rect 4002 37998 4014 38050
rect 4498 37998 4510 38050
rect 4562 37998 4574 38050
rect 5170 37998 5182 38050
rect 5234 37998 5246 38050
rect 5618 37998 5630 38050
rect 5682 37998 5694 38050
rect 6626 37998 6638 38050
rect 6690 37998 6702 38050
rect 3614 37986 3666 37998
rect 8094 37986 8146 37998
rect 8206 38050 8258 38062
rect 9774 38050 9826 38062
rect 9314 37998 9326 38050
rect 9378 37998 9390 38050
rect 8206 37986 8258 37998
rect 9774 37986 9826 37998
rect 9886 38050 9938 38062
rect 15710 38050 15762 38062
rect 29934 38050 29986 38062
rect 44270 38050 44322 38062
rect 56030 38050 56082 38062
rect 10546 37998 10558 38050
rect 10610 37998 10622 38050
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 19282 37998 19294 38050
rect 19346 37998 19358 38050
rect 19618 37998 19630 38050
rect 19682 37998 19694 38050
rect 21074 37998 21086 38050
rect 21138 37998 21150 38050
rect 21858 37998 21870 38050
rect 21922 37998 21934 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 26002 37998 26014 38050
rect 26066 37998 26078 38050
rect 28690 37998 28702 38050
rect 28754 37998 28766 38050
rect 29026 37998 29038 38050
rect 29090 37998 29102 38050
rect 30482 37998 30494 38050
rect 30546 37998 30558 38050
rect 31266 37998 31278 38050
rect 31330 37998 31342 38050
rect 32946 37998 32958 38050
rect 33010 37998 33022 38050
rect 33394 37998 33406 38050
rect 33458 37998 33470 38050
rect 34626 37998 34638 38050
rect 34690 37998 34702 38050
rect 35634 37998 35646 38050
rect 35698 37998 35710 38050
rect 37874 37998 37886 38050
rect 37938 37998 37950 38050
rect 42802 37998 42814 38050
rect 42866 37998 42878 38050
rect 43698 37998 43710 38050
rect 43762 37998 43774 38050
rect 45042 37998 45054 38050
rect 45106 37998 45118 38050
rect 45602 37998 45614 38050
rect 45666 37998 45678 38050
rect 53554 37998 53566 38050
rect 53618 37998 53630 38050
rect 9886 37986 9938 37998
rect 15710 37986 15762 37998
rect 29934 37986 29986 37998
rect 44270 37986 44322 37998
rect 56030 37986 56082 37998
rect 9662 37938 9714 37950
rect 28254 37938 28306 37950
rect 12786 37886 12798 37938
rect 12850 37886 12862 37938
rect 9662 37874 9714 37886
rect 28254 37874 28306 37886
rect 32622 37938 32674 37950
rect 42478 37938 42530 37950
rect 41906 37886 41918 37938
rect 41970 37886 41982 37938
rect 32622 37874 32674 37886
rect 42478 37874 42530 37886
rect 45950 37938 46002 37950
rect 45950 37874 46002 37886
rect 46734 37938 46786 37950
rect 47282 37886 47294 37938
rect 47346 37886 47358 37938
rect 48850 37886 48862 37938
rect 48914 37886 48926 37938
rect 51426 37886 51438 37938
rect 51490 37886 51502 37938
rect 46734 37874 46786 37886
rect 2830 37826 2882 37838
rect 2830 37762 2882 37774
rect 14366 37826 14418 37838
rect 14366 37762 14418 37774
rect 16046 37826 16098 37838
rect 16046 37762 16098 37774
rect 23102 37826 23154 37838
rect 23102 37762 23154 37774
rect 27582 37826 27634 37838
rect 27582 37762 27634 37774
rect 36318 37826 36370 37838
rect 36318 37762 36370 37774
rect 40350 37826 40402 37838
rect 40350 37762 40402 37774
rect 46958 37826 47010 37838
rect 46958 37762 47010 37774
rect 47518 37826 47570 37838
rect 47518 37762 47570 37774
rect 48190 37826 48242 37838
rect 48190 37762 48242 37774
rect 53006 37826 53058 37838
rect 53006 37762 53058 37774
rect 55246 37826 55298 37838
rect 55246 37762 55298 37774
rect 672 37658 56784 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 43806 37658
rect 43858 37606 43910 37658
rect 43962 37606 44014 37658
rect 44066 37606 56784 37658
rect 672 37572 56784 37606
rect 19966 37490 20018 37502
rect 19966 37426 20018 37438
rect 50654 37490 50706 37502
rect 50654 37426 50706 37438
rect 28478 37378 28530 37390
rect 8082 37326 8094 37378
rect 8146 37326 8158 37378
rect 46274 37326 46286 37378
rect 46338 37326 46350 37378
rect 48402 37326 48414 37378
rect 48466 37326 48478 37378
rect 49074 37326 49086 37378
rect 49138 37326 49150 37378
rect 52434 37326 52446 37378
rect 52498 37326 52510 37378
rect 28478 37314 28530 37326
rect 2942 37266 2994 37278
rect 15934 37266 15986 37278
rect 25678 37266 25730 37278
rect 29934 37266 29986 37278
rect 1362 37214 1374 37266
rect 1426 37214 1438 37266
rect 2146 37214 2158 37266
rect 2210 37214 2222 37266
rect 3490 37214 3502 37266
rect 3554 37214 3566 37266
rect 3938 37214 3950 37266
rect 4002 37214 4014 37266
rect 5058 37214 5070 37266
rect 5122 37214 5134 37266
rect 5842 37214 5854 37266
rect 5906 37214 5918 37266
rect 10322 37214 10334 37266
rect 10386 37214 10398 37266
rect 14914 37214 14926 37266
rect 14978 37214 14990 37266
rect 15362 37214 15374 37266
rect 15426 37214 15438 37266
rect 16482 37214 16494 37266
rect 16546 37214 16558 37266
rect 17602 37214 17614 37266
rect 17666 37214 17678 37266
rect 18274 37214 18286 37266
rect 18338 37214 18350 37266
rect 22194 37214 22206 37266
rect 22258 37214 22270 37266
rect 24546 37214 24558 37266
rect 24610 37214 24622 37266
rect 24994 37214 25006 37266
rect 25058 37214 25070 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 27234 37214 27246 37266
rect 27298 37214 27310 37266
rect 28802 37214 28814 37266
rect 28866 37214 28878 37266
rect 29362 37214 29374 37266
rect 29426 37214 29438 37266
rect 30482 37214 30494 37266
rect 30546 37214 30558 37266
rect 31390 37261 31442 37273
rect 34190 37266 34242 37278
rect 43262 37266 43314 37278
rect 51102 37266 51154 37278
rect 2942 37202 2994 37214
rect 15934 37202 15986 37214
rect 25678 37202 25730 37214
rect 29934 37202 29986 37214
rect 32834 37214 32846 37266
rect 32898 37214 32910 37266
rect 33394 37214 33406 37266
rect 33458 37214 33470 37266
rect 34626 37214 34638 37266
rect 34690 37214 34702 37266
rect 35634 37214 35646 37266
rect 35698 37214 35710 37266
rect 36754 37214 36766 37266
rect 36818 37214 36830 37266
rect 39106 37214 39118 37266
rect 39170 37214 39182 37266
rect 39666 37214 39678 37266
rect 39730 37214 39742 37266
rect 40338 37214 40350 37266
rect 40402 37214 40414 37266
rect 40898 37214 40910 37266
rect 40962 37214 40974 37266
rect 41906 37214 41918 37266
rect 41970 37214 41982 37266
rect 45602 37214 45614 37266
rect 45666 37214 45678 37266
rect 54562 37214 54574 37266
rect 54626 37214 54638 37266
rect 31390 37197 31442 37209
rect 34190 37202 34242 37214
rect 43262 37202 43314 37214
rect 51102 37202 51154 37214
rect 4398 37154 4450 37166
rect 14478 37154 14530 37166
rect 24222 37154 24274 37166
rect 32510 37154 32562 37166
rect 38782 37154 38834 37166
rect 42702 37154 42754 37166
rect 44158 37154 44210 37166
rect 44718 37154 44770 37166
rect 3378 37102 3390 37154
rect 3442 37102 3454 37154
rect 5282 37102 5294 37154
rect 5346 37102 5358 37154
rect 6178 37102 6190 37154
rect 6242 37102 6254 37154
rect 8418 37102 8430 37154
rect 8482 37102 8494 37154
rect 10770 37102 10782 37154
rect 10834 37102 10846 37154
rect 18834 37102 18846 37154
rect 18898 37102 18910 37154
rect 22530 37102 22542 37154
rect 22594 37102 22606 37154
rect 25218 37102 25230 37154
rect 25282 37102 25294 37154
rect 29474 37102 29486 37154
rect 29538 37102 29550 37154
rect 33506 37102 33518 37154
rect 33570 37102 33582 37154
rect 37202 37102 37214 37154
rect 37266 37102 37278 37154
rect 39778 37102 39790 37154
rect 39842 37102 39854 37154
rect 43586 37102 43598 37154
rect 43650 37102 43662 37154
rect 44482 37102 44494 37154
rect 44546 37102 44558 37154
rect 4398 37090 4450 37102
rect 14478 37090 14530 37102
rect 24222 37090 24274 37102
rect 32510 37090 32562 37102
rect 38782 37090 38834 37102
rect 42702 37090 42754 37102
rect 44158 37090 44210 37102
rect 44718 37090 44770 37102
rect 7422 37042 7474 37054
rect 7422 36978 7474 36990
rect 9662 37042 9714 37054
rect 9662 36978 9714 36990
rect 11902 37042 11954 37054
rect 23774 37042 23826 37054
rect 15474 36990 15486 37042
rect 15538 36990 15550 37042
rect 11902 36978 11954 36990
rect 23774 36978 23826 36990
rect 38334 37042 38386 37054
rect 38334 36978 38386 36990
rect 42814 37042 42866 37054
rect 42814 36978 42866 36990
rect 43038 37042 43090 37054
rect 54014 37042 54066 37054
rect 56254 37042 56306 37054
rect 49522 36990 49534 37042
rect 49586 36990 49598 37042
rect 51426 36990 51438 37042
rect 51490 36990 51502 37042
rect 52882 36990 52894 37042
rect 52946 36990 52958 37042
rect 55122 36990 55134 37042
rect 55186 36990 55198 37042
rect 43038 36978 43090 36990
rect 54014 36978 54066 36990
rect 56254 36978 56306 36990
rect 672 36874 56784 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 44466 36874
rect 44518 36822 44570 36874
rect 44622 36822 44674 36874
rect 44726 36822 56784 36874
rect 672 36788 56784 36822
rect 6862 36706 6914 36718
rect 7534 36706 7586 36718
rect 7186 36654 7198 36706
rect 7250 36654 7262 36706
rect 6862 36642 6914 36654
rect 7534 36642 7586 36654
rect 9214 36706 9266 36718
rect 9214 36642 9266 36654
rect 9438 36706 9490 36718
rect 9438 36642 9490 36654
rect 9662 36706 9714 36718
rect 9662 36642 9714 36654
rect 16046 36706 16098 36718
rect 47070 36706 47122 36718
rect 17378 36654 17390 36706
rect 17442 36654 17454 36706
rect 25554 36654 25566 36706
rect 25618 36654 25630 36706
rect 36194 36654 36206 36706
rect 36258 36654 36270 36706
rect 42130 36654 42142 36706
rect 42194 36654 42206 36706
rect 16046 36642 16098 36654
rect 47070 36642 47122 36654
rect 54126 36706 54178 36718
rect 54126 36642 54178 36654
rect 54238 36706 54290 36718
rect 54786 36654 54798 36706
rect 54850 36654 54862 36706
rect 54238 36642 54290 36654
rect 3782 36594 3834 36606
rect 8318 36594 8370 36606
rect 9774 36594 9826 36606
rect 18958 36594 19010 36606
rect 20414 36594 20466 36606
rect 1586 36542 1598 36594
rect 1650 36542 1662 36594
rect 4274 36542 4286 36594
rect 4338 36542 4350 36594
rect 7858 36542 7870 36594
rect 7922 36542 7934 36594
rect 8866 36542 8878 36594
rect 8930 36542 8942 36594
rect 11106 36542 11118 36594
rect 11170 36542 11182 36594
rect 14914 36542 14926 36594
rect 14978 36542 14990 36594
rect 19954 36542 19966 36594
rect 20018 36542 20030 36594
rect 3782 36530 3834 36542
rect 8318 36530 8370 36542
rect 9774 36530 9826 36542
rect 18958 36530 19010 36542
rect 20414 36530 20466 36542
rect 24558 36594 24610 36606
rect 24558 36530 24610 36542
rect 26014 36594 26066 36606
rect 35198 36594 35250 36606
rect 30146 36542 30158 36594
rect 30210 36542 30222 36594
rect 33506 36542 33518 36594
rect 33570 36542 33582 36594
rect 26014 36530 26066 36542
rect 35198 36530 35250 36542
rect 36654 36594 36706 36606
rect 36654 36530 36706 36542
rect 42590 36594 42642 36606
rect 47294 36594 47346 36606
rect 45266 36542 45278 36594
rect 45330 36542 45342 36594
rect 42590 36530 42642 36542
rect 47294 36530 47346 36542
rect 55918 36594 55970 36606
rect 55918 36530 55970 36542
rect 56142 36594 56194 36606
rect 56142 36530 56194 36542
rect 2830 36482 2882 36494
rect 4734 36482 4786 36494
rect 34750 36482 34802 36494
rect 46958 36482 47010 36494
rect 1250 36430 1262 36482
rect 1314 36430 1326 36482
rect 4050 36430 4062 36482
rect 4114 36430 4126 36482
rect 5506 36430 5518 36482
rect 5570 36430 5582 36482
rect 6290 36430 6302 36482
rect 6354 36430 6366 36482
rect 10434 36430 10446 36482
rect 10498 36430 10510 36482
rect 10994 36430 11006 36482
rect 11058 36430 11070 36482
rect 11666 36430 11678 36482
rect 11730 36430 11742 36482
rect 12114 36430 12126 36482
rect 12178 36430 12190 36482
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 13122 36430 13134 36482
rect 13186 36430 13198 36482
rect 14466 36430 14478 36482
rect 14530 36430 14542 36482
rect 19394 36430 19406 36482
rect 19458 36430 19470 36482
rect 19730 36430 19742 36482
rect 19794 36430 19806 36482
rect 20962 36430 20974 36482
rect 21026 36430 21038 36482
rect 22082 36430 22094 36482
rect 22146 36430 22158 36482
rect 24994 36430 25006 36482
rect 25058 36430 25070 36482
rect 25442 36430 25454 36482
rect 25506 36430 25518 36482
rect 26786 36430 26798 36482
rect 26850 36430 26862 36482
rect 27570 36430 27582 36482
rect 27634 36430 27646 36482
rect 33170 36430 33182 36482
rect 33234 36430 33246 36482
rect 35522 36430 35534 36482
rect 35586 36430 35598 36482
rect 35970 36430 35982 36482
rect 36034 36430 36046 36482
rect 37426 36430 37438 36482
rect 37490 36430 37502 36482
rect 38210 36430 38222 36482
rect 38274 36430 38286 36482
rect 41570 36430 41582 36482
rect 41634 36430 41646 36482
rect 41906 36430 41918 36482
rect 41970 36430 41982 36482
rect 43138 36430 43150 36482
rect 43202 36430 43214 36482
rect 44146 36430 44158 36482
rect 44210 36430 44222 36482
rect 2830 36418 2882 36430
rect 4734 36418 4786 36430
rect 34750 36418 34802 36430
rect 46958 36418 47010 36430
rect 47518 36482 47570 36494
rect 53678 36482 53730 36494
rect 49522 36430 49534 36482
rect 49586 36430 49598 36482
rect 47518 36418 47570 36430
rect 53678 36418 53730 36430
rect 53902 36482 53954 36494
rect 53902 36418 53954 36430
rect 54350 36482 54402 36494
rect 54350 36418 54402 36430
rect 3278 36370 3330 36382
rect 3278 36306 3330 36318
rect 8206 36370 8258 36382
rect 8206 36306 8258 36318
rect 10110 36370 10162 36382
rect 41134 36370 41186 36382
rect 55358 36370 55410 36382
rect 16930 36318 16942 36370
rect 16994 36318 17006 36370
rect 29810 36318 29822 36370
rect 29874 36318 29886 36370
rect 44930 36318 44942 36370
rect 44994 36318 45006 36370
rect 52210 36318 52222 36370
rect 52274 36318 52286 36370
rect 10110 36306 10162 36318
rect 41134 36306 41186 36318
rect 55358 36306 55410 36318
rect 18510 36258 18562 36270
rect 18510 36194 18562 36206
rect 31390 36258 31442 36270
rect 31390 36194 31442 36206
rect 46510 36258 46562 36270
rect 46510 36194 46562 36206
rect 55134 36258 55186 36270
rect 55134 36194 55186 36206
rect 56254 36258 56306 36270
rect 56254 36194 56306 36206
rect 672 36090 56784 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 43806 36090
rect 43858 36038 43910 36090
rect 43962 36038 44014 36090
rect 44066 36038 56784 36090
rect 672 36004 56784 36038
rect 23326 35922 23378 35934
rect 23326 35858 23378 35870
rect 44270 35922 44322 35934
rect 44270 35858 44322 35870
rect 48190 35922 48242 35934
rect 48190 35858 48242 35870
rect 55358 35922 55410 35934
rect 55358 35858 55410 35870
rect 4398 35810 4450 35822
rect 4398 35746 4450 35758
rect 4958 35810 5010 35822
rect 30606 35810 30658 35822
rect 21746 35758 21758 35810
rect 21810 35758 21822 35810
rect 4958 35746 5010 35758
rect 30606 35746 30658 35758
rect 38894 35810 38946 35822
rect 53230 35810 53282 35822
rect 48850 35758 48862 35810
rect 48914 35758 48926 35810
rect 52546 35758 52558 35810
rect 52610 35758 52622 35810
rect 38894 35746 38946 35758
rect 53230 35746 53282 35758
rect 54238 35810 54290 35822
rect 54238 35746 54290 35758
rect 54798 35810 54850 35822
rect 54798 35746 54850 35758
rect 55806 35810 55858 35822
rect 55806 35746 55858 35758
rect 1486 35693 1538 35705
rect 10446 35698 10498 35710
rect 20078 35698 20130 35710
rect 32510 35698 32562 35710
rect 40574 35698 40626 35710
rect 43374 35698 43426 35710
rect 52110 35698 52162 35710
rect 2370 35646 2382 35698
rect 2434 35646 2446 35698
rect 2818 35646 2830 35698
rect 2882 35646 2894 35698
rect 3602 35646 3614 35698
rect 3666 35646 3678 35698
rect 3938 35646 3950 35698
rect 4002 35646 4014 35698
rect 5282 35646 5294 35698
rect 5346 35646 5358 35698
rect 5730 35646 5742 35698
rect 5794 35646 5806 35698
rect 6962 35646 6974 35698
rect 7026 35646 7038 35698
rect 7970 35646 7982 35698
rect 8034 35646 8046 35698
rect 9314 35646 9326 35698
rect 9378 35646 9390 35698
rect 9762 35646 9774 35698
rect 9826 35646 9838 35698
rect 11218 35646 11230 35698
rect 11282 35646 11294 35698
rect 12114 35646 12126 35698
rect 12178 35646 12190 35698
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 23986 35646 23998 35698
rect 24050 35646 24062 35698
rect 26114 35646 26126 35698
rect 26178 35646 26190 35698
rect 28690 35646 28702 35698
rect 28754 35646 28766 35698
rect 31042 35646 31054 35698
rect 31106 35646 31118 35698
rect 32162 35646 32174 35698
rect 32226 35646 32238 35698
rect 33282 35646 33294 35698
rect 33346 35646 33358 35698
rect 33730 35646 33742 35698
rect 33794 35646 33806 35698
rect 37986 35646 37998 35698
rect 38050 35646 38062 35698
rect 39218 35646 39230 35698
rect 39282 35646 39294 35698
rect 39778 35646 39790 35698
rect 39842 35646 39854 35698
rect 40898 35646 40910 35698
rect 40962 35646 40974 35698
rect 42018 35646 42030 35698
rect 42082 35646 42094 35698
rect 45826 35646 45838 35698
rect 45890 35646 45902 35698
rect 46610 35646 46622 35698
rect 46674 35646 46686 35698
rect 1486 35629 1538 35641
rect 10446 35634 10498 35646
rect 20078 35634 20130 35646
rect 32510 35634 32562 35646
rect 40574 35634 40626 35646
rect 43374 35634 43426 35646
rect 52110 35634 52162 35646
rect 52334 35698 52386 35710
rect 52334 35634 52386 35646
rect 52670 35698 52722 35710
rect 52670 35634 52722 35646
rect 53454 35698 53506 35710
rect 53454 35634 53506 35646
rect 54126 35698 54178 35710
rect 54126 35634 54178 35646
rect 54910 35698 54962 35710
rect 54910 35634 54962 35646
rect 55134 35698 55186 35710
rect 55134 35634 55186 35646
rect 55694 35698 55746 35710
rect 55694 35634 55746 35646
rect 6414 35586 6466 35598
rect 6414 35522 6466 35534
rect 8990 35586 9042 35598
rect 19518 35586 19570 35598
rect 9986 35534 9998 35586
rect 10050 35534 10062 35586
rect 14354 35534 14366 35586
rect 14418 35534 14430 35586
rect 8990 35522 9042 35534
rect 19518 35522 19570 35534
rect 19742 35586 19794 35598
rect 34190 35586 34242 35598
rect 42926 35586 42978 35598
rect 22082 35534 22094 35586
rect 22146 35534 22158 35586
rect 26674 35534 26686 35586
rect 26738 35534 26750 35586
rect 33170 35534 33182 35586
rect 33234 35534 33246 35586
rect 37538 35534 37550 35586
rect 37602 35534 37614 35586
rect 19742 35522 19794 35534
rect 34190 35522 34242 35534
rect 42926 35522 42978 35534
rect 43486 35586 43538 35598
rect 43486 35522 43538 35534
rect 43710 35586 43762 35598
rect 50878 35586 50930 35598
rect 45378 35534 45390 35586
rect 45442 35534 45454 35586
rect 46946 35534 46958 35586
rect 47010 35534 47022 35586
rect 49186 35534 49198 35586
rect 49250 35534 49262 35586
rect 43710 35522 43762 35534
rect 50878 35522 50930 35534
rect 51214 35586 51266 35598
rect 51214 35522 51266 35534
rect 51438 35586 51490 35598
rect 51438 35522 51490 35534
rect 52894 35586 52946 35598
rect 52894 35522 52946 35534
rect 15486 35474 15538 35486
rect 3378 35422 3390 35474
rect 3442 35422 3454 35474
rect 5954 35422 5966 35474
rect 6018 35422 6030 35474
rect 15486 35410 15538 35422
rect 19854 35474 19906 35486
rect 25566 35474 25618 35486
rect 24434 35422 24446 35474
rect 24498 35422 24510 35474
rect 19854 35410 19906 35422
rect 25566 35410 25618 35422
rect 27806 35474 27858 35486
rect 30270 35474 30322 35486
rect 29138 35422 29150 35474
rect 29202 35422 29214 35474
rect 27806 35410 27858 35422
rect 30270 35410 30322 35422
rect 36430 35474 36482 35486
rect 43038 35474 43090 35486
rect 39890 35422 39902 35474
rect 39954 35422 39966 35474
rect 36430 35410 36482 35422
rect 43038 35410 43090 35422
rect 50430 35474 50482 35486
rect 50430 35410 50482 35422
rect 50990 35474 51042 35486
rect 54686 35474 54738 35486
rect 53778 35422 53790 35474
rect 53842 35422 53854 35474
rect 50990 35410 51042 35422
rect 54686 35410 54738 35422
rect 55918 35474 55970 35486
rect 55918 35410 55970 35422
rect 56142 35474 56194 35486
rect 56142 35410 56194 35422
rect 672 35306 56784 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 44466 35306
rect 44518 35254 44570 35306
rect 44622 35254 44674 35306
rect 44726 35254 56784 35306
rect 672 35220 56784 35254
rect 19630 35138 19682 35150
rect 19630 35074 19682 35086
rect 32510 35138 32562 35150
rect 44830 35138 44882 35150
rect 33618 35086 33630 35138
rect 33682 35086 33694 35138
rect 35634 35086 35646 35138
rect 35698 35086 35710 35138
rect 32510 35074 32562 35086
rect 44830 35074 44882 35086
rect 47182 35138 47234 35150
rect 47182 35074 47234 35086
rect 54798 35138 54850 35150
rect 54798 35074 54850 35086
rect 55246 35138 55298 35150
rect 55246 35074 55298 35086
rect 2830 35026 2882 35038
rect 1586 34974 1598 35026
rect 1650 34974 1662 35026
rect 2830 34962 2882 34974
rect 3390 35026 3442 35038
rect 7982 35026 8034 35038
rect 5282 34974 5294 35026
rect 5346 34974 5358 35026
rect 3390 34962 3442 34974
rect 7982 34962 8034 34974
rect 8094 35026 8146 35038
rect 19070 35026 19122 35038
rect 10994 34974 11006 35026
rect 11058 34974 11070 35026
rect 14802 34974 14814 35026
rect 14866 34974 14878 35026
rect 17266 34974 17278 35026
rect 17330 34974 17342 35026
rect 8094 34962 8146 34974
rect 19070 34962 19122 34974
rect 19182 35026 19234 35038
rect 22206 35026 22258 35038
rect 28702 35026 28754 35038
rect 47406 35026 47458 35038
rect 54686 35026 54738 35038
rect 21746 34974 21758 35026
rect 21810 34974 21822 35026
rect 25666 34974 25678 35026
rect 25730 34974 25742 35026
rect 28242 34974 28254 35026
rect 28306 34974 28318 35026
rect 41570 34974 41582 35026
rect 41634 34974 41646 35026
rect 43138 34974 43150 35026
rect 43202 34974 43214 35026
rect 45938 34974 45950 35026
rect 46002 34974 46014 35026
rect 49970 34974 49982 35026
rect 50034 34974 50046 35026
rect 51314 34974 51326 35026
rect 51378 34974 51390 35026
rect 19182 34962 19234 34974
rect 22206 34962 22258 34974
rect 28702 34962 28754 34974
rect 47406 34962 47458 34974
rect 54686 34962 54738 34974
rect 56142 35026 56194 35038
rect 56142 34962 56194 34974
rect 3502 34914 3554 34926
rect 3502 34850 3554 34862
rect 3614 34914 3666 34926
rect 3614 34850 3666 34862
rect 3726 34914 3778 34926
rect 7758 34914 7810 34926
rect 11678 34914 11730 34926
rect 19742 34914 19794 34926
rect 3938 34862 3950 34914
rect 4002 34862 4014 34914
rect 4610 34862 4622 34914
rect 4674 34862 4686 34914
rect 5058 34862 5070 34914
rect 5122 34862 5134 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 6290 34862 6302 34914
rect 6354 34862 6366 34914
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 10322 34862 10334 34914
rect 10386 34862 10398 34914
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 12002 34862 12014 34914
rect 12066 34862 12078 34914
rect 13010 34862 13022 34914
rect 13074 34862 13086 34914
rect 15362 34862 15374 34914
rect 15426 34862 15438 34914
rect 3726 34850 3778 34862
rect 7758 34850 7810 34862
rect 11678 34850 11730 34862
rect 19742 34850 19794 34862
rect 19966 34914 20018 34926
rect 36318 34914 36370 34926
rect 46958 34914 47010 34926
rect 54574 34914 54626 34926
rect 20178 34862 20190 34914
rect 20242 34862 20254 34914
rect 21074 34862 21086 34914
rect 21138 34862 21150 34914
rect 21634 34862 21646 34914
rect 21698 34862 21710 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 23874 34862 23886 34914
rect 23938 34862 23950 34914
rect 25218 34862 25230 34914
rect 25282 34862 25294 34914
rect 27682 34862 27694 34914
rect 27746 34862 27758 34914
rect 28018 34862 28030 34914
rect 28082 34862 28094 34914
rect 29474 34862 29486 34914
rect 29538 34862 29550 34914
rect 30370 34862 30382 34914
rect 30434 34862 30446 34914
rect 35074 34862 35086 34914
rect 35138 34862 35150 34914
rect 35410 34862 35422 34914
rect 35474 34862 35486 34914
rect 36866 34862 36878 34914
rect 36930 34862 36942 34914
rect 37762 34862 37774 34914
rect 37826 34862 37838 34914
rect 42018 34862 42030 34914
rect 42082 34862 42094 34914
rect 46386 34862 46398 34914
rect 46450 34862 46462 34914
rect 52210 34862 52222 34914
rect 52274 34862 52286 34914
rect 19966 34850 20018 34862
rect 36318 34850 36370 34862
rect 46958 34850 47010 34862
rect 54574 34850 54626 34862
rect 4286 34802 4338 34814
rect 1250 34750 1262 34802
rect 1314 34750 1326 34802
rect 4286 34738 4338 34750
rect 9998 34802 10050 34814
rect 19854 34802 19906 34814
rect 16930 34750 16942 34802
rect 16994 34750 17006 34802
rect 9998 34738 10050 34750
rect 19854 34738 19906 34750
rect 20750 34802 20802 34814
rect 20750 34738 20802 34750
rect 27246 34802 27298 34814
rect 34638 34802 34690 34814
rect 47070 34802 47122 34814
rect 34066 34750 34078 34802
rect 34130 34750 34142 34802
rect 42690 34750 42702 34802
rect 42754 34750 42766 34802
rect 27246 34738 27298 34750
rect 34638 34738 34690 34750
rect 47070 34738 47122 34750
rect 54350 34802 54402 34814
rect 54350 34738 54402 34750
rect 55358 34802 55410 34814
rect 56130 34750 56142 34802
rect 56194 34750 56206 34802
rect 55358 34738 55410 34750
rect 13694 34690 13746 34702
rect 13694 34626 13746 34638
rect 18510 34690 18562 34702
rect 18510 34626 18562 34638
rect 19070 34690 19122 34702
rect 19070 34626 19122 34638
rect 26798 34690 26850 34702
rect 26798 34626 26850 34638
rect 40350 34690 40402 34702
rect 40350 34626 40402 34638
rect 44270 34690 44322 34702
rect 44270 34626 44322 34638
rect 54126 34690 54178 34702
rect 54126 34626 54178 34638
rect 55918 34690 55970 34702
rect 55918 34626 55970 34638
rect 672 34522 56784 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 43806 34522
rect 43858 34470 43910 34522
rect 43962 34470 44014 34522
rect 44066 34470 56784 34522
rect 672 34436 56784 34470
rect 19070 34354 19122 34366
rect 19070 34290 19122 34302
rect 35198 34354 35250 34366
rect 35198 34290 35250 34302
rect 45614 34354 45666 34366
rect 45614 34290 45666 34302
rect 50318 34354 50370 34366
rect 50318 34290 50370 34302
rect 54686 34354 54738 34366
rect 54686 34290 54738 34302
rect 5070 34242 5122 34254
rect 14030 34242 14082 34254
rect 10546 34190 10558 34242
rect 10610 34190 10622 34242
rect 5070 34178 5122 34190
rect 14030 34178 14082 34190
rect 29822 34242 29874 34254
rect 37326 34242 37378 34254
rect 50878 34242 50930 34254
rect 33618 34190 33630 34242
rect 33682 34190 33694 34242
rect 46274 34190 46286 34242
rect 46338 34190 46350 34242
rect 48290 34190 48302 34242
rect 48354 34190 48366 34242
rect 29822 34178 29874 34190
rect 37326 34178 37378 34190
rect 50878 34178 50930 34190
rect 52558 34242 52610 34254
rect 52558 34178 52610 34190
rect 55694 34242 55746 34254
rect 55694 34178 55746 34190
rect 3838 34130 3890 34142
rect 1250 34078 1262 34130
rect 1314 34078 1326 34130
rect 3838 34066 3890 34078
rect 3950 34130 4002 34142
rect 3950 34066 4002 34078
rect 4174 34130 4226 34142
rect 4174 34066 4226 34078
rect 4846 34130 4898 34142
rect 15486 34130 15538 34142
rect 18622 34130 18674 34142
rect 6066 34078 6078 34130
rect 6130 34078 6142 34130
rect 9874 34078 9886 34130
rect 9938 34078 9950 34130
rect 14466 34078 14478 34130
rect 14530 34078 14542 34130
rect 14802 34078 14814 34130
rect 14866 34078 14878 34130
rect 16146 34078 16158 34130
rect 16210 34078 16222 34130
rect 17042 34078 17054 34130
rect 17106 34078 17118 34130
rect 4846 34066 4898 34078
rect 15486 34066 15538 34078
rect 18622 34066 18674 34078
rect 19630 34130 19682 34142
rect 19630 34066 19682 34078
rect 20078 34130 20130 34142
rect 20078 34066 20130 34078
rect 20526 34130 20578 34142
rect 20526 34066 20578 34078
rect 20862 34130 20914 34142
rect 26014 34130 26066 34142
rect 31278 34130 31330 34142
rect 36766 34130 36818 34142
rect 39566 34130 39618 34142
rect 45278 34130 45330 34142
rect 22418 34078 22430 34130
rect 22482 34078 22494 34130
rect 24882 34078 24894 34130
rect 24946 34078 24958 34130
rect 25330 34078 25342 34130
rect 25394 34078 25406 34130
rect 26674 34078 26686 34130
rect 26738 34078 26750 34130
rect 27570 34078 27582 34130
rect 27634 34078 27646 34130
rect 30258 34078 30270 34130
rect 30322 34078 30334 34130
rect 30594 34078 30606 34130
rect 30658 34078 30670 34130
rect 32050 34078 32062 34130
rect 32114 34078 32126 34130
rect 32834 34078 32846 34130
rect 32898 34078 32910 34130
rect 38098 34078 38110 34130
rect 38162 34078 38174 34130
rect 38994 34078 39006 34130
rect 39058 34078 39070 34130
rect 40338 34078 40350 34130
rect 40402 34078 40414 34130
rect 40786 34078 40798 34130
rect 40850 34078 40862 34130
rect 43362 34078 43374 34130
rect 43426 34078 43438 34130
rect 44818 34078 44830 34130
rect 44882 34078 44894 34130
rect 20862 34066 20914 34078
rect 26014 34066 26066 34078
rect 31278 34066 31330 34078
rect 36766 34066 36818 34078
rect 39566 34066 39618 34078
rect 45278 34066 45330 34078
rect 46062 34130 46114 34142
rect 46062 34066 46114 34078
rect 47854 34130 47906 34142
rect 47854 34066 47906 34078
rect 50542 34130 50594 34142
rect 50542 34066 50594 34078
rect 52222 34130 52274 34142
rect 55358 34130 55410 34142
rect 53106 34078 53118 34130
rect 53170 34078 53182 34130
rect 52222 34066 52274 34078
rect 55358 34066 55410 34078
rect 55918 34130 55970 34142
rect 55918 34066 55970 34078
rect 3278 34018 3330 34030
rect 3278 33954 3330 33966
rect 4398 34018 4450 34030
rect 4398 33954 4450 33966
rect 5294 34018 5346 34030
rect 5294 33954 5346 33966
rect 5518 34018 5570 34030
rect 18510 34018 18562 34030
rect 6514 33966 6526 34018
rect 6578 33966 6590 34018
rect 15026 33966 15038 34018
rect 15090 33966 15102 34018
rect 5518 33954 5570 33966
rect 18510 33954 18562 33966
rect 18958 34018 19010 34030
rect 18958 33954 19010 33966
rect 19406 34018 19458 34030
rect 19406 33954 19458 33966
rect 20750 34018 20802 34030
rect 20750 33954 20802 33966
rect 24558 34018 24610 34030
rect 37438 34018 37490 34030
rect 41246 34018 41298 34030
rect 46286 34018 46338 34030
rect 25554 33966 25566 34018
rect 25618 33966 25630 34018
rect 30818 33966 30830 34018
rect 30882 33966 30894 34018
rect 34066 33966 34078 34018
rect 34130 33966 34142 34018
rect 40226 33966 40238 34018
rect 40290 33966 40302 34018
rect 42802 33966 42814 34018
rect 42866 33966 42878 34018
rect 44706 33966 44718 34018
rect 44770 33966 44782 34018
rect 24558 33954 24610 33966
rect 37438 33954 37490 33966
rect 41246 33954 41298 33966
rect 46286 33954 46338 33966
rect 46398 34018 46450 34030
rect 47182 34018 47234 34030
rect 46610 33966 46622 34018
rect 46674 33966 46686 34018
rect 46398 33954 46450 33966
rect 47182 33954 47234 33966
rect 47294 34018 47346 34030
rect 50766 34018 50818 34030
rect 48626 33966 48638 34018
rect 48690 33966 48702 34018
rect 47294 33954 47346 33966
rect 50766 33954 50818 33966
rect 50990 34018 51042 34030
rect 50990 33954 51042 33966
rect 51998 34018 52050 34030
rect 53554 33966 53566 34018
rect 53618 33966 53630 34018
rect 51998 33954 52050 33966
rect 2830 33906 2882 33918
rect 1698 33854 1710 33906
rect 1762 33854 1774 33906
rect 2830 33842 2882 33854
rect 3390 33906 3442 33918
rect 3390 33842 3442 33854
rect 3614 33906 3666 33918
rect 3614 33842 3666 33854
rect 7646 33906 7698 33918
rect 7646 33842 7698 33854
rect 8206 33906 8258 33918
rect 12126 33906 12178 33918
rect 9314 33854 9326 33906
rect 9378 33854 9390 33906
rect 10994 33854 11006 33906
rect 11058 33854 11070 33906
rect 8206 33842 8258 33854
rect 12126 33842 12178 33854
rect 19854 33906 19906 33918
rect 24110 33906 24162 33918
rect 22978 33854 22990 33906
rect 23042 33854 23054 33906
rect 19854 33842 19906 33854
rect 24110 33842 24162 33854
rect 37214 33906 37266 33918
rect 37214 33842 37266 33854
rect 41694 33906 41746 33918
rect 41694 33842 41746 33854
rect 47406 33906 47458 33918
rect 47406 33842 47458 33854
rect 49870 33906 49922 33918
rect 49870 33842 49922 33854
rect 55246 33906 55298 33918
rect 55246 33842 55298 33854
rect 55470 33906 55522 33918
rect 55470 33842 55522 33854
rect 672 33738 56784 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 44466 33738
rect 44518 33686 44570 33738
rect 44622 33686 44674 33738
rect 44726 33686 56784 33738
rect 672 33652 56784 33686
rect 2494 33570 2546 33582
rect 1362 33518 1374 33570
rect 1426 33518 1438 33570
rect 2494 33506 2546 33518
rect 2718 33570 2770 33582
rect 6526 33570 6578 33582
rect 18510 33570 18562 33582
rect 39566 33570 39618 33582
rect 55022 33570 55074 33582
rect 3938 33518 3950 33570
rect 4002 33518 4014 33570
rect 13906 33518 13918 33570
rect 13970 33518 13982 33570
rect 20514 33518 20526 33570
rect 20578 33518 20590 33570
rect 33058 33518 33070 33570
rect 33122 33518 33134 33570
rect 38434 33518 38446 33570
rect 38498 33518 38510 33570
rect 40898 33518 40910 33570
rect 40962 33518 40974 33570
rect 53890 33518 53902 33570
rect 53954 33518 53966 33570
rect 2718 33506 2770 33518
rect 6526 33506 6578 33518
rect 18510 33506 18562 33518
rect 39566 33506 39618 33518
rect 55022 33506 55074 33518
rect 2382 33458 2434 33470
rect 2034 33406 2046 33458
rect 2098 33406 2110 33458
rect 2382 33394 2434 33406
rect 6638 33458 6690 33470
rect 14366 33458 14418 33470
rect 19518 33458 19570 33470
rect 8082 33406 8094 33458
rect 8146 33406 8158 33458
rect 9874 33406 9886 33458
rect 9938 33406 9950 33458
rect 17378 33406 17390 33458
rect 17442 33406 17454 33458
rect 6638 33394 6690 33406
rect 14366 33394 14418 33406
rect 19518 33394 19570 33406
rect 20974 33458 21026 33470
rect 28030 33458 28082 33470
rect 52670 33458 52722 33470
rect 27570 33406 27582 33458
rect 27634 33406 27646 33458
rect 32946 33406 32958 33458
rect 33010 33406 33022 33458
rect 35858 33406 35870 33458
rect 35922 33406 35934 33458
rect 40786 33406 40798 33458
rect 40850 33406 40862 33458
rect 44594 33406 44606 33458
rect 44658 33406 44670 33458
rect 47506 33406 47518 33458
rect 47570 33406 47582 33458
rect 48738 33406 48750 33458
rect 48802 33406 48814 33458
rect 20974 33394 21026 33406
rect 28030 33394 28082 33406
rect 52670 33394 52722 33406
rect 56030 33458 56082 33470
rect 56354 33406 56366 33458
rect 56418 33406 56430 33458
rect 56030 33394 56082 33406
rect 4398 33346 4450 33358
rect 7086 33346 7138 33358
rect 1138 33294 1150 33346
rect 1202 33294 1214 33346
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 3378 33294 3390 33346
rect 3442 33294 3454 33346
rect 3714 33294 3726 33346
rect 3778 33294 3790 33346
rect 5058 33294 5070 33346
rect 5122 33294 5134 33346
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 4398 33282 4450 33294
rect 7086 33282 7138 33294
rect 7422 33346 7474 33358
rect 10334 33346 10386 33358
rect 36990 33346 37042 33358
rect 45278 33346 45330 33358
rect 47182 33346 47234 33358
rect 8194 33294 8206 33346
rect 8258 33294 8270 33346
rect 9202 33294 9214 33346
rect 9266 33294 9278 33346
rect 9762 33294 9774 33346
rect 9826 33294 9838 33346
rect 10882 33294 10894 33346
rect 10946 33294 10958 33346
rect 12002 33294 12014 33346
rect 12066 33294 12078 33346
rect 13234 33294 13246 33346
rect 13298 33294 13310 33346
rect 13794 33294 13806 33346
rect 13858 33294 13870 33346
rect 14914 33294 14926 33346
rect 14978 33294 14990 33346
rect 16034 33294 16046 33346
rect 16098 33294 16110 33346
rect 19954 33294 19966 33346
rect 20018 33294 20030 33346
rect 7422 33282 7474 33294
rect 10334 33282 10386 33294
rect 20402 33282 20414 33334
rect 20466 33282 20478 33334
rect 21746 33294 21758 33346
rect 21810 33294 21822 33346
rect 22642 33294 22654 33346
rect 22706 33294 22718 33346
rect 27010 33294 27022 33346
rect 27074 33294 27086 33346
rect 27346 33294 27358 33346
rect 27410 33294 27422 33346
rect 28578 33294 28590 33346
rect 28642 33294 28654 33346
rect 29698 33294 29710 33346
rect 29762 33294 29774 33346
rect 32498 33294 32510 33346
rect 32562 33294 32574 33346
rect 35410 33294 35422 33346
rect 35474 33294 35486 33346
rect 37986 33294 37998 33346
rect 38050 33294 38062 33346
rect 44034 33294 44046 33346
rect 44098 33294 44110 33346
rect 44370 33294 44382 33346
rect 44434 33294 44446 33346
rect 45602 33294 45614 33346
rect 45666 33294 45678 33346
rect 46610 33294 46622 33346
rect 46674 33294 46686 33346
rect 36990 33282 37042 33294
rect 45278 33282 45330 33294
rect 47182 33282 47234 33294
rect 50654 33346 50706 33358
rect 50654 33282 50706 33294
rect 51326 33346 51378 33358
rect 51326 33282 51378 33294
rect 51550 33346 51602 33358
rect 52222 33346 52274 33358
rect 51874 33294 51886 33346
rect 51938 33294 51950 33346
rect 51550 33282 51602 33294
rect 52222 33282 52274 33294
rect 52446 33346 52498 33358
rect 52446 33282 52498 33294
rect 2942 33234 2994 33246
rect 2942 33170 2994 33182
rect 8878 33234 8930 33246
rect 8878 33170 8930 33182
rect 12910 33234 12962 33246
rect 26574 33234 26626 33246
rect 43598 33234 43650 33246
rect 50430 33234 50482 33246
rect 16930 33182 16942 33234
rect 16994 33182 17006 33234
rect 40450 33182 40462 33234
rect 40514 33182 40526 33234
rect 48402 33182 48414 33234
rect 48466 33182 48478 33234
rect 12910 33170 12962 33182
rect 26574 33170 26626 33182
rect 43598 33170 43650 33182
rect 50430 33170 50482 33182
rect 51438 33234 51490 33246
rect 51438 33170 51490 33182
rect 52334 33234 52386 33246
rect 53442 33182 53454 33234
rect 53506 33182 53518 33234
rect 52334 33170 52386 33182
rect 34190 33122 34242 33134
rect 34190 33058 34242 33070
rect 42030 33122 42082 33134
rect 42030 33058 42082 33070
rect 49982 33122 50034 33134
rect 50978 33070 50990 33122
rect 51042 33070 51054 33122
rect 49982 33058 50034 33070
rect 672 32954 56784 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 43806 32954
rect 43858 32902 43910 32954
rect 43962 32902 44014 32954
rect 44066 32902 56784 32954
rect 672 32868 56784 32902
rect 7982 32786 8034 32798
rect 7982 32722 8034 32734
rect 45950 32786 46002 32798
rect 45950 32722 46002 32734
rect 50094 32786 50146 32798
rect 50094 32722 50146 32734
rect 8430 32674 8482 32686
rect 1250 32622 1262 32674
rect 1314 32622 1326 32674
rect 4162 32622 4174 32674
rect 4226 32622 4238 32674
rect 8430 32610 8482 32622
rect 15486 32674 15538 32686
rect 26126 32674 26178 32686
rect 20850 32622 20862 32674
rect 20914 32622 20926 32674
rect 15486 32610 15538 32622
rect 26126 32610 26178 32622
rect 28814 32674 28866 32686
rect 40350 32674 40402 32686
rect 37986 32622 37998 32674
rect 38050 32622 38062 32674
rect 44370 32622 44382 32674
rect 44434 32622 44446 32674
rect 28814 32610 28866 32622
rect 40350 32610 40402 32622
rect 3838 32562 3890 32574
rect 9886 32562 9938 32574
rect 15038 32562 15090 32574
rect 24446 32562 24498 32574
rect 38558 32562 38610 32574
rect 41806 32562 41858 32574
rect 48638 32562 48690 32574
rect 6402 32510 6414 32562
rect 6466 32510 6478 32562
rect 8754 32510 8766 32562
rect 8818 32510 8830 32562
rect 9202 32510 9214 32562
rect 9266 32510 9278 32562
rect 10658 32510 10670 32562
rect 10722 32510 10734 32562
rect 11442 32510 11454 32562
rect 11506 32510 11518 32562
rect 13458 32510 13470 32562
rect 13522 32510 13534 32562
rect 15810 32510 15822 32562
rect 15874 32510 15886 32562
rect 16258 32510 16270 32562
rect 16322 32510 16334 32562
rect 17490 32510 17502 32562
rect 17554 32510 17566 32562
rect 18498 32510 18510 32562
rect 18562 32510 18574 32562
rect 23090 32510 23102 32562
rect 23154 32510 23166 32562
rect 23874 32510 23886 32562
rect 23938 32510 23950 32562
rect 24098 32510 24110 32562
rect 24162 32510 24174 32562
rect 25330 32510 25342 32562
rect 25394 32510 25406 32562
rect 25666 32510 25678 32562
rect 25730 32510 25742 32562
rect 29922 32510 29934 32562
rect 29986 32510 29998 32562
rect 32274 32510 32286 32562
rect 32338 32510 32350 32562
rect 33058 32510 33070 32562
rect 33122 32510 33134 32562
rect 34402 32510 34414 32562
rect 34466 32510 34478 32562
rect 34850 32510 34862 32562
rect 34914 32510 34926 32562
rect 39218 32510 39230 32562
rect 39282 32510 39294 32562
rect 40674 32510 40686 32562
rect 40738 32510 40750 32562
rect 41122 32510 41134 32562
rect 41186 32510 41198 32562
rect 42466 32510 42478 32562
rect 42530 32510 42542 32562
rect 43474 32510 43486 32562
rect 43538 32510 43550 32562
rect 46610 32510 46622 32562
rect 46674 32510 46686 32562
rect 3838 32498 3890 32510
rect 9886 32498 9938 32510
rect 15038 32498 15090 32510
rect 24446 32498 24498 32510
rect 38558 32498 38610 32510
rect 41806 32498 41858 32510
rect 48638 32498 48690 32510
rect 48974 32562 49026 32574
rect 48974 32498 49026 32510
rect 50878 32562 50930 32574
rect 50878 32498 50930 32510
rect 51102 32562 51154 32574
rect 51102 32498 51154 32510
rect 51998 32562 52050 32574
rect 51998 32498 52050 32510
rect 52670 32562 52722 32574
rect 52670 32498 52722 32510
rect 52894 32562 52946 32574
rect 52894 32498 52946 32510
rect 54574 32562 54626 32574
rect 54574 32498 54626 32510
rect 54798 32562 54850 32574
rect 54798 32498 54850 32510
rect 3278 32450 3330 32462
rect 1698 32398 1710 32450
rect 1762 32398 1774 32450
rect 3278 32386 3330 32398
rect 3390 32450 3442 32462
rect 5854 32450 5906 32462
rect 16942 32450 16994 32462
rect 29262 32450 29314 32462
rect 33854 32450 33906 32462
rect 35310 32450 35362 32462
rect 4946 32398 4958 32450
rect 5010 32398 5022 32450
rect 6738 32398 6750 32450
rect 6802 32398 6814 32450
rect 9426 32398 9438 32450
rect 9490 32398 9502 32450
rect 21298 32398 21310 32450
rect 21362 32398 21374 32450
rect 30482 32398 30494 32450
rect 30546 32398 30558 32450
rect 34290 32398 34302 32450
rect 34354 32398 34366 32450
rect 3390 32386 3442 32398
rect 5854 32386 5906 32398
rect 16942 32386 16994 32398
rect 29262 32386 29314 32398
rect 33854 32386 33906 32398
rect 35310 32386 35362 32398
rect 38782 32450 38834 32462
rect 38782 32386 38834 32398
rect 38894 32450 38946 32462
rect 48750 32450 48802 32462
rect 53342 32450 53394 32462
rect 55694 32450 55746 32462
rect 46946 32398 46958 32450
rect 47010 32398 47022 32450
rect 49298 32398 49310 32450
rect 49362 32398 49374 32450
rect 49858 32398 49870 32450
rect 49922 32398 49934 32450
rect 53778 32398 53790 32450
rect 53842 32398 53854 32450
rect 56018 32398 56030 32450
rect 56082 32398 56094 32450
rect 38894 32386 38946 32398
rect 48750 32386 48802 32398
rect 53342 32386 53394 32398
rect 55694 32386 55746 32398
rect 2830 32338 2882 32350
rect 2830 32274 2882 32286
rect 3950 32338 4002 32350
rect 3950 32274 4002 32286
rect 4174 32338 4226 32350
rect 4174 32274 4226 32286
rect 4286 32338 4338 32350
rect 4286 32274 4338 32286
rect 5294 32338 5346 32350
rect 5294 32274 5346 32286
rect 5518 32338 5570 32350
rect 5518 32274 5570 32286
rect 5742 32338 5794 32350
rect 22430 32338 22482 32350
rect 28926 32338 28978 32350
rect 13906 32286 13918 32338
rect 13970 32286 13982 32338
rect 16482 32286 16494 32338
rect 16546 32286 16558 32338
rect 25106 32286 25118 32338
rect 25170 32286 25182 32338
rect 5742 32274 5794 32286
rect 22430 32274 22482 32286
rect 28926 32274 28978 32286
rect 29374 32338 29426 32350
rect 29374 32274 29426 32286
rect 29598 32338 29650 32350
rect 29598 32274 29650 32286
rect 31614 32338 31666 32350
rect 31614 32274 31666 32286
rect 36430 32338 36482 32350
rect 38670 32338 38722 32350
rect 48190 32338 48242 32350
rect 37538 32286 37550 32338
rect 37602 32286 37614 32338
rect 41346 32286 41358 32338
rect 41410 32286 41422 32338
rect 44818 32286 44830 32338
rect 44882 32286 44894 32338
rect 36430 32274 36482 32286
rect 38670 32274 38722 32286
rect 48190 32274 48242 32286
rect 50430 32338 50482 32350
rect 53118 32338 53170 32350
rect 51426 32286 51438 32338
rect 51490 32286 51502 32338
rect 52322 32286 52334 32338
rect 52386 32286 52398 32338
rect 50430 32274 50482 32286
rect 53118 32274 53170 32286
rect 53230 32338 53282 32350
rect 53230 32274 53282 32286
rect 54126 32338 54178 32350
rect 54126 32274 54178 32286
rect 55022 32338 55074 32350
rect 55022 32274 55074 32286
rect 55134 32338 55186 32350
rect 55134 32274 55186 32286
rect 55246 32338 55298 32350
rect 55246 32274 55298 32286
rect 672 32170 56784 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 44466 32170
rect 44518 32118 44570 32170
rect 44622 32118 44674 32170
rect 44726 32118 56784 32170
rect 672 32084 56784 32118
rect 2830 32002 2882 32014
rect 2830 31938 2882 31950
rect 34190 32002 34242 32014
rect 34190 31938 34242 31950
rect 50206 32002 50258 32014
rect 50206 31938 50258 31950
rect 52894 32002 52946 32014
rect 52894 31938 52946 31950
rect 7534 31890 7586 31902
rect 1586 31838 1598 31890
rect 1650 31838 1662 31890
rect 3602 31838 3614 31890
rect 3666 31838 3678 31890
rect 4946 31838 4958 31890
rect 5010 31838 5022 31890
rect 7534 31826 7586 31838
rect 7646 31890 7698 31902
rect 7646 31826 7698 31838
rect 8206 31890 8258 31902
rect 10334 31890 10386 31902
rect 16046 31890 16098 31902
rect 34750 31890 34802 31902
rect 9874 31838 9886 31890
rect 9938 31838 9950 31890
rect 14914 31838 14926 31890
rect 14978 31838 14990 31890
rect 20402 31838 20414 31890
rect 20466 31838 20478 31890
rect 22642 31838 22654 31890
rect 22706 31838 22718 31890
rect 25218 31838 25230 31890
rect 25282 31838 25294 31890
rect 25554 31838 25566 31890
rect 25618 31838 25630 31890
rect 27458 31838 27470 31890
rect 27522 31838 27534 31890
rect 33058 31838 33070 31890
rect 33122 31838 33134 31890
rect 8206 31826 8258 31838
rect 10334 31826 10386 31838
rect 16046 31826 16098 31838
rect 34750 31826 34802 31838
rect 34974 31890 35026 31902
rect 34974 31826 35026 31838
rect 35422 31890 35474 31902
rect 35422 31826 35474 31838
rect 35534 31890 35586 31902
rect 41246 31890 41298 31902
rect 47182 31890 47234 31902
rect 37314 31838 37326 31890
rect 37378 31838 37390 31890
rect 42242 31838 42254 31890
rect 42306 31838 42318 31890
rect 45378 31838 45390 31890
rect 45442 31838 45454 31890
rect 35534 31826 35586 31838
rect 41246 31826 41298 31838
rect 47182 31826 47234 31838
rect 47406 31890 47458 31902
rect 47406 31826 47458 31838
rect 48190 31890 48242 31902
rect 50654 31890 50706 31902
rect 55246 31890 55298 31902
rect 49410 31838 49422 31890
rect 49474 31838 49486 31890
rect 51762 31838 51774 31890
rect 51826 31838 51838 31890
rect 54114 31838 54126 31890
rect 54178 31838 54190 31890
rect 56354 31838 56366 31890
rect 56418 31838 56430 31890
rect 48190 31826 48242 31838
rect 50654 31826 50706 31838
rect 55246 31826 55298 31838
rect 5406 31778 5458 31790
rect 7870 31778 7922 31790
rect 1250 31726 1262 31778
rect 1314 31726 1326 31778
rect 3378 31726 3390 31778
rect 3442 31726 3454 31778
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 4834 31726 4846 31778
rect 4898 31726 4910 31778
rect 6178 31726 6190 31778
rect 6242 31726 6254 31778
rect 7074 31726 7086 31778
rect 7138 31726 7150 31778
rect 5406 31714 5458 31726
rect 7870 31714 7922 31726
rect 8318 31778 8370 31790
rect 19966 31778 20018 31790
rect 23886 31778 23938 31790
rect 9202 31726 9214 31778
rect 9266 31726 9278 31778
rect 9762 31726 9774 31778
rect 9826 31726 9838 31778
rect 10882 31726 10894 31778
rect 10946 31726 10958 31778
rect 11890 31726 11902 31778
rect 11954 31726 11966 31778
rect 18274 31726 18286 31778
rect 18338 31726 18350 31778
rect 19394 31726 19406 31778
rect 19458 31726 19470 31778
rect 20626 31726 20638 31778
rect 20690 31726 20702 31778
rect 20962 31726 20974 31778
rect 21026 31726 21038 31778
rect 8318 31714 8370 31726
rect 19966 31714 20018 31726
rect 23886 31714 23938 31726
rect 25006 31778 25058 31790
rect 27918 31778 27970 31790
rect 34638 31778 34690 31790
rect 26898 31726 26910 31778
rect 26962 31726 26974 31778
rect 27346 31726 27358 31778
rect 27410 31726 27422 31778
rect 28578 31726 28590 31778
rect 28642 31726 28654 31778
rect 29586 31726 29598 31778
rect 29650 31726 29662 31778
rect 32498 31726 32510 31778
rect 32562 31726 32574 31778
rect 25006 31714 25058 31726
rect 27918 31714 27970 31726
rect 34638 31714 34690 31726
rect 35198 31778 35250 31790
rect 35198 31714 35250 31726
rect 35310 31778 35362 31790
rect 48078 31778 48130 31790
rect 35858 31726 35870 31778
rect 35922 31726 35934 31778
rect 36754 31726 36766 31778
rect 36818 31726 36830 31778
rect 37090 31726 37102 31778
rect 37154 31726 37166 31778
rect 37874 31726 37886 31778
rect 37938 31726 37950 31778
rect 38434 31726 38446 31778
rect 38498 31726 38510 31778
rect 39330 31726 39342 31778
rect 39394 31726 39406 31778
rect 41682 31726 41694 31778
rect 41746 31726 41758 31778
rect 42018 31726 42030 31778
rect 42082 31726 42094 31778
rect 42802 31726 42814 31778
rect 42866 31726 42878 31778
rect 43250 31726 43262 31778
rect 43314 31726 43326 31778
rect 44258 31726 44270 31778
rect 44322 31726 44334 31778
rect 45042 31726 45054 31778
rect 45106 31726 45118 31778
rect 35310 31714 35362 31726
rect 48078 31714 48130 31726
rect 48414 31778 48466 31790
rect 48414 31714 48466 31726
rect 48526 31778 48578 31790
rect 48526 31714 48578 31726
rect 49086 31778 49138 31790
rect 50094 31778 50146 31790
rect 49746 31726 49758 31778
rect 49810 31726 49822 31778
rect 49086 31714 49138 31726
rect 50094 31714 50146 31726
rect 50430 31778 50482 31790
rect 50430 31714 50482 31726
rect 56030 31778 56082 31790
rect 56030 31714 56082 31726
rect 3950 31666 4002 31678
rect 3950 31602 4002 31614
rect 8878 31666 8930 31678
rect 21422 31666 21474 31678
rect 24670 31666 24722 31678
rect 14466 31614 14478 31666
rect 14530 31614 14542 31666
rect 22306 31614 22318 31666
rect 22370 31614 22382 31666
rect 8878 31602 8930 31614
rect 21422 31602 21474 31614
rect 24670 31602 24722 31614
rect 26462 31666 26514 31678
rect 26462 31602 26514 31614
rect 36318 31666 36370 31678
rect 51314 31614 51326 31666
rect 51378 31614 51390 31666
rect 53666 31614 53678 31666
rect 53730 31614 53742 31666
rect 36318 31602 36370 31614
rect 8206 31554 8258 31566
rect 8206 31490 8258 31502
rect 46622 31554 46674 31566
rect 46622 31490 46674 31502
rect 47070 31554 47122 31566
rect 47070 31490 47122 31502
rect 50206 31554 50258 31566
rect 50206 31490 50258 31502
rect 672 31386 56784 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 43806 31386
rect 43858 31334 43910 31386
rect 43962 31334 44014 31386
rect 44066 31334 56784 31386
rect 672 31300 56784 31334
rect 22430 31218 22482 31230
rect 22430 31154 22482 31166
rect 42814 31218 42866 31230
rect 42814 31154 42866 31166
rect 48526 31218 48578 31230
rect 48526 31154 48578 31166
rect 51326 31218 51378 31230
rect 51326 31154 51378 31166
rect 53790 31218 53842 31230
rect 53790 31154 53842 31166
rect 56030 31218 56082 31230
rect 56030 31154 56082 31166
rect 5070 31106 5122 31118
rect 8206 31106 8258 31118
rect 6178 31054 6190 31106
rect 6242 31054 6254 31106
rect 5070 31042 5122 31054
rect 8206 31042 8258 31054
rect 16830 31106 16882 31118
rect 26126 31106 26178 31118
rect 20850 31054 20862 31106
rect 20914 31054 20926 31106
rect 16830 31042 16882 31054
rect 26126 31042 26178 31054
rect 28926 31106 28978 31118
rect 43486 31106 43538 31118
rect 29922 31054 29934 31106
rect 29986 31054 29998 31106
rect 36530 31054 36542 31106
rect 36594 31054 36606 31106
rect 38770 31054 38782 31106
rect 38834 31054 38846 31106
rect 47506 31054 47518 31106
rect 47570 31054 47582 31106
rect 28926 31042 28978 31054
rect 43486 31042 43538 31054
rect 4958 30994 5010 31006
rect 1362 30942 1374 30994
rect 1426 30942 1438 30994
rect 2370 30942 2382 30994
rect 2434 30942 2446 30994
rect 3602 30942 3614 30994
rect 3666 30942 3678 30994
rect 3938 30942 3950 30994
rect 4002 30942 4014 30994
rect 4958 30930 5010 30942
rect 5182 30994 5234 31006
rect 9886 30994 9938 31006
rect 18510 30994 18562 31006
rect 27470 30994 27522 31006
rect 35870 30994 35922 31006
rect 48414 30994 48466 31006
rect 51214 30994 51266 31006
rect 8530 30942 8542 30994
rect 8594 30942 8606 30994
rect 8978 30942 8990 30994
rect 9042 30942 9054 30994
rect 10322 30942 10334 30994
rect 10386 30942 10398 30994
rect 11330 30942 11342 30994
rect 11394 30942 11406 30994
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 13906 30942 13918 30994
rect 13970 30942 13982 30994
rect 15138 30942 15150 30994
rect 15202 30942 15214 30994
rect 16258 30942 16270 30994
rect 16322 30942 16334 30994
rect 17154 30942 17166 30994
rect 17218 30942 17230 30994
rect 17602 30942 17614 30994
rect 17666 30942 17678 30994
rect 18834 30942 18846 30994
rect 18898 30942 18910 30994
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 23090 30942 23102 30994
rect 23154 30942 23166 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 24098 30942 24110 30994
rect 24162 30942 24174 30994
rect 24546 30942 24558 30994
rect 24610 30942 24622 30994
rect 25218 30942 25230 30994
rect 25282 30942 25294 30994
rect 25666 30942 25678 30994
rect 25730 30942 25742 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 32386 30942 32398 30994
rect 32450 30942 32462 30994
rect 32722 30942 32734 30994
rect 32786 30942 32798 30994
rect 34066 30942 34078 30994
rect 34130 30942 34142 30994
rect 34962 30942 34974 30994
rect 35026 30942 35038 30994
rect 41122 30942 41134 30994
rect 41186 30942 41198 30994
rect 45154 30942 45166 30994
rect 45218 30942 45230 30994
rect 47842 30942 47854 30994
rect 47906 30942 47918 30994
rect 49186 30942 49198 30994
rect 49250 30942 49262 30994
rect 52210 30942 52222 30994
rect 52274 30942 52286 30994
rect 54338 30942 54350 30994
rect 54402 30942 54414 30994
rect 5182 30930 5234 30942
rect 9886 30930 9938 30942
rect 18510 30930 18562 30942
rect 27470 30930 27522 30942
rect 35870 30930 35922 30942
rect 48414 30930 48466 30942
rect 51214 30930 51266 30942
rect 2942 30882 2994 30894
rect 2942 30818 2994 30830
rect 4398 30882 4450 30894
rect 4398 30818 4450 30830
rect 5518 30882 5570 30894
rect 5518 30818 5570 30830
rect 13134 30882 13186 30894
rect 14590 30882 14642 30894
rect 31950 30882 32002 30894
rect 14130 30830 14142 30882
rect 14194 30830 14206 30882
rect 17826 30830 17838 30882
rect 17890 30830 17902 30882
rect 21186 30830 21198 30882
rect 21250 30830 21262 30882
rect 25106 30830 25118 30882
rect 25170 30830 25182 30882
rect 26674 30830 26686 30882
rect 26738 30830 26750 30882
rect 30370 30830 30382 30882
rect 30434 30830 30446 30882
rect 13134 30818 13186 30830
rect 14590 30818 14642 30830
rect 31950 30818 32002 30830
rect 33406 30882 33458 30894
rect 33406 30818 33458 30830
rect 35534 30882 35586 30894
rect 35534 30818 35586 30830
rect 35646 30882 35698 30894
rect 44382 30882 44434 30894
rect 39106 30830 39118 30882
rect 39170 30830 39182 30882
rect 41570 30830 41582 30882
rect 41634 30830 41646 30882
rect 35646 30818 35698 30830
rect 44382 30818 44434 30830
rect 44494 30882 44546 30894
rect 44494 30818 44546 30830
rect 44718 30882 44770 30894
rect 44718 30818 44770 30830
rect 47406 30882 47458 30894
rect 47406 30818 47458 30830
rect 47518 30882 47570 30894
rect 47518 30818 47570 30830
rect 48526 30882 48578 30894
rect 52658 30830 52670 30882
rect 52722 30830 52734 30882
rect 48526 30818 48578 30830
rect 7758 30770 7810 30782
rect 27806 30770 27858 30782
rect 3378 30718 3390 30770
rect 3442 30718 3454 30770
rect 6626 30718 6638 30770
rect 6690 30718 6702 30770
rect 9202 30718 9214 30770
rect 9266 30718 9278 30770
rect 21298 30718 21310 30770
rect 21362 30718 21374 30770
rect 7758 30706 7810 30718
rect 27806 30706 27858 30718
rect 28814 30770 28866 30782
rect 28814 30706 28866 30718
rect 29038 30770 29090 30782
rect 29038 30706 29090 30718
rect 29262 30770 29314 30782
rect 29262 30706 29314 30718
rect 31502 30770 31554 30782
rect 38110 30770 38162 30782
rect 32946 30718 32958 30770
rect 33010 30718 33022 30770
rect 36978 30718 36990 30770
rect 37042 30718 37054 30770
rect 31502 30706 31554 30718
rect 38110 30706 38162 30718
rect 40350 30770 40402 30782
rect 40350 30706 40402 30718
rect 43598 30770 43650 30782
rect 46734 30770 46786 30782
rect 45602 30718 45614 30770
rect 45666 30718 45678 30770
rect 43598 30706 43650 30718
rect 46734 30706 46786 30718
rect 47182 30770 47234 30782
rect 50766 30770 50818 30782
rect 49634 30718 49646 30770
rect 49698 30718 49710 30770
rect 47182 30706 47234 30718
rect 50766 30706 50818 30718
rect 51326 30770 51378 30782
rect 54898 30718 54910 30770
rect 54962 30718 54974 30770
rect 51326 30706 51378 30718
rect 672 30602 56784 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 44466 30602
rect 44518 30550 44570 30602
rect 44622 30550 44674 30602
rect 44726 30550 56784 30602
rect 672 30516 56784 30550
rect 2830 30434 2882 30446
rect 2830 30370 2882 30382
rect 9326 30434 9378 30446
rect 9326 30370 9378 30382
rect 9550 30434 9602 30446
rect 9550 30370 9602 30382
rect 13806 30434 13858 30446
rect 19070 30434 19122 30446
rect 14914 30382 14926 30434
rect 14978 30382 14990 30434
rect 17938 30382 17950 30434
rect 18002 30382 18014 30434
rect 13806 30370 13858 30382
rect 19070 30370 19122 30382
rect 27246 30434 27298 30446
rect 27246 30370 27298 30382
rect 29934 30434 29986 30446
rect 29934 30370 29986 30382
rect 30046 30434 30098 30446
rect 30046 30370 30098 30382
rect 30158 30434 30210 30446
rect 38446 30434 38498 30446
rect 36642 30382 36654 30434
rect 36706 30382 36718 30434
rect 30158 30370 30210 30382
rect 38446 30370 38498 30382
rect 38670 30434 38722 30446
rect 52222 30434 52274 30446
rect 38670 30370 38722 30382
rect 39342 30378 39394 30390
rect 50082 30382 50094 30434
rect 50146 30382 50158 30434
rect 16830 30322 16882 30334
rect 1586 30270 1598 30322
rect 1650 30270 1662 30322
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 12674 30270 12686 30322
rect 12738 30270 12750 30322
rect 16830 30258 16882 30270
rect 16942 30322 16994 30334
rect 38222 30322 38274 30334
rect 20514 30270 20526 30322
rect 20578 30270 20590 30322
rect 26002 30270 26014 30322
rect 26066 30270 26078 30322
rect 28354 30270 28366 30322
rect 28418 30270 28430 30322
rect 30482 30270 30494 30322
rect 30546 30270 30558 30322
rect 33394 30270 33406 30322
rect 33458 30270 33470 30322
rect 16942 30258 16994 30270
rect 38222 30258 38274 30270
rect 39230 30322 39282 30334
rect 52222 30370 52274 30382
rect 52334 30434 52386 30446
rect 52334 30370 52386 30382
rect 56142 30434 56194 30446
rect 56142 30370 56194 30382
rect 39342 30314 39394 30326
rect 47406 30322 47458 30334
rect 41234 30270 41246 30322
rect 41298 30270 41310 30322
rect 45042 30270 45054 30322
rect 45106 30270 45118 30322
rect 47170 30270 47182 30322
rect 47234 30270 47246 30322
rect 39230 30258 39282 30270
rect 47406 30258 47458 30270
rect 48974 30322 49026 30334
rect 48974 30258 49026 30270
rect 51214 30322 51266 30334
rect 51214 30258 51266 30270
rect 52110 30322 52162 30334
rect 55918 30322 55970 30334
rect 53666 30270 53678 30322
rect 53730 30270 53742 30322
rect 52110 30258 52162 30270
rect 55918 30258 55970 30270
rect 5294 30210 5346 30222
rect 7758 30210 7810 30222
rect 9438 30210 9490 30222
rect 10110 30210 10162 30222
rect 1250 30158 1262 30210
rect 1314 30158 1326 30210
rect 4050 30158 4062 30210
rect 4114 30158 4126 30210
rect 4498 30158 4510 30210
rect 4562 30158 4574 30210
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 6626 30158 6638 30210
rect 6690 30158 6702 30210
rect 9090 30158 9102 30210
rect 9154 30158 9166 30210
rect 9762 30158 9774 30210
rect 9826 30158 9838 30210
rect 5294 30146 5346 30158
rect 7758 30146 7810 30158
rect 9438 30146 9490 30158
rect 10110 30146 10162 30158
rect 10222 30210 10274 30222
rect 10222 30146 10274 30158
rect 10334 30210 10386 30222
rect 10334 30146 10386 30158
rect 10558 30210 10610 30222
rect 16046 30210 16098 30222
rect 20974 30210 21026 30222
rect 29486 30210 29538 30222
rect 31502 30210 31554 30222
rect 40238 30210 40290 30222
rect 41918 30210 41970 30222
rect 46174 30210 46226 30222
rect 46958 30210 47010 30222
rect 12226 30158 12238 30210
rect 12290 30158 12302 30210
rect 14466 30158 14478 30210
rect 14530 30158 14542 30210
rect 17378 30158 17390 30210
rect 17442 30158 17454 30210
rect 19954 30158 19966 30210
rect 20018 30158 20030 30210
rect 20402 30158 20414 30210
rect 20466 30158 20478 30210
rect 21522 30158 21534 30210
rect 21586 30158 21598 30210
rect 22642 30158 22654 30210
rect 22706 30158 22718 30210
rect 30370 30158 30382 30210
rect 30434 30158 30446 30210
rect 32722 30158 32734 30210
rect 32786 30158 32798 30210
rect 33170 30158 33182 30210
rect 33234 30158 33246 30210
rect 33954 30158 33966 30210
rect 34018 30158 34030 30210
rect 34514 30158 34526 30210
rect 34578 30158 34590 30210
rect 35522 30158 35534 30210
rect 35586 30158 35598 30210
rect 40562 30158 40574 30210
rect 40626 30158 40638 30210
rect 41010 30158 41022 30210
rect 41074 30158 41086 30210
rect 42354 30158 42366 30210
rect 42418 30158 42430 30210
rect 43250 30158 43262 30210
rect 43314 30158 43326 30210
rect 44482 30158 44494 30210
rect 44546 30158 44558 30210
rect 46722 30158 46734 30210
rect 46786 30158 46798 30210
rect 10558 30146 10610 30158
rect 16046 30146 16098 30158
rect 20974 30146 21026 30158
rect 29486 30146 29538 30158
rect 31502 30146 31554 30158
rect 40238 30146 40290 30158
rect 41918 30146 41970 30158
rect 46174 30146 46226 30158
rect 46958 30146 47010 30158
rect 47294 30210 47346 30222
rect 47294 30146 47346 30158
rect 48302 30210 48354 30222
rect 51662 30210 51714 30222
rect 49522 30158 49534 30210
rect 49586 30158 49598 30210
rect 48302 30146 48354 30158
rect 51662 30146 51714 30158
rect 51886 30210 51938 30222
rect 51886 30146 51938 30158
rect 54910 30210 54962 30222
rect 54910 30146 54962 30158
rect 3614 30098 3666 30110
rect 3614 30034 3666 30046
rect 8206 30098 8258 30110
rect 8206 30034 8258 30046
rect 19518 30098 19570 30110
rect 31278 30098 31330 30110
rect 25666 30046 25678 30098
rect 25730 30046 25742 30098
rect 27906 30046 27918 30098
rect 27970 30046 27982 30098
rect 19518 30034 19570 30046
rect 31278 30034 31330 30046
rect 32398 30098 32450 30110
rect 38334 30098 38386 30110
rect 56030 30098 56082 30110
rect 36194 30046 36206 30098
rect 36258 30046 36270 30098
rect 53330 30046 53342 30098
rect 53394 30046 53406 30098
rect 32398 30034 32450 30046
rect 38334 30034 38386 30046
rect 56030 30034 56082 30046
rect 7870 29986 7922 29998
rect 7870 29922 7922 29934
rect 8318 29986 8370 29998
rect 8318 29922 8370 29934
rect 16830 29986 16882 29998
rect 37774 29986 37826 29998
rect 31826 29934 31838 29986
rect 31890 29934 31902 29986
rect 16830 29922 16882 29934
rect 37774 29922 37826 29934
rect 39230 29986 39282 29998
rect 39230 29922 39282 29934
rect 48190 29986 48242 29998
rect 48190 29922 48242 29934
rect 48526 29986 48578 29998
rect 48526 29922 48578 29934
rect 48638 29986 48690 29998
rect 48638 29922 48690 29934
rect 49086 29986 49138 29998
rect 49086 29922 49138 29934
rect 672 29818 56784 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 43806 29818
rect 43858 29766 43910 29818
rect 43962 29766 44014 29818
rect 44066 29766 56784 29818
rect 672 29732 56784 29766
rect 5854 29650 5906 29662
rect 5854 29586 5906 29598
rect 6302 29650 6354 29662
rect 6302 29586 6354 29598
rect 8990 29650 9042 29662
rect 8990 29586 9042 29598
rect 12910 29650 12962 29662
rect 12910 29586 12962 29598
rect 23326 29650 23378 29662
rect 23326 29586 23378 29598
rect 27806 29650 27858 29662
rect 27806 29586 27858 29598
rect 34750 29650 34802 29662
rect 34750 29586 34802 29598
rect 36430 29650 36482 29662
rect 36430 29586 36482 29598
rect 42142 29650 42194 29662
rect 42142 29586 42194 29598
rect 53230 29650 53282 29662
rect 53230 29586 53282 29598
rect 55470 29650 55522 29662
rect 55470 29586 55522 29598
rect 4174 29538 4226 29550
rect 1250 29486 1262 29538
rect 1314 29486 1326 29538
rect 4174 29474 4226 29486
rect 6414 29538 6466 29550
rect 6414 29474 6466 29486
rect 20078 29538 20130 29550
rect 33966 29538 34018 29550
rect 21746 29486 21758 29538
rect 21810 29486 21822 29538
rect 23986 29486 23998 29538
rect 24050 29486 24062 29538
rect 26226 29486 26238 29538
rect 26290 29486 26302 29538
rect 20078 29474 20130 29486
rect 33966 29474 34018 29486
rect 46846 29538 46898 29550
rect 52546 29486 52558 29538
rect 52610 29486 52622 29538
rect 46846 29474 46898 29486
rect 2830 29426 2882 29438
rect 2830 29362 2882 29374
rect 3838 29426 3890 29438
rect 3838 29362 3890 29374
rect 4062 29426 4114 29438
rect 4062 29362 4114 29374
rect 4398 29426 4450 29438
rect 4398 29362 4450 29374
rect 5182 29426 5234 29438
rect 5182 29362 5234 29374
rect 5406 29426 5458 29438
rect 5406 29362 5458 29374
rect 5966 29426 6018 29438
rect 9326 29426 9378 29438
rect 7410 29374 7422 29426
rect 7474 29374 7486 29426
rect 5966 29362 6018 29374
rect 9326 29362 9378 29374
rect 9662 29426 9714 29438
rect 9662 29362 9714 29374
rect 9886 29426 9938 29438
rect 9886 29362 9938 29374
rect 11678 29426 11730 29438
rect 14466 29374 14478 29426
rect 14530 29374 14542 29426
rect 17166 29421 17218 29433
rect 20862 29426 20914 29438
rect 11678 29362 11730 29374
rect 17826 29374 17838 29426
rect 17890 29374 17902 29426
rect 18498 29374 18510 29426
rect 18562 29374 18574 29426
rect 19170 29374 19182 29426
rect 19234 29374 19246 29426
rect 19618 29374 19630 29426
rect 19682 29374 19694 29426
rect 17166 29357 17218 29369
rect 20862 29362 20914 29374
rect 21086 29426 21138 29438
rect 32510 29426 32562 29438
rect 35646 29426 35698 29438
rect 46622 29426 46674 29438
rect 50318 29426 50370 29438
rect 28690 29374 28702 29426
rect 28754 29374 28766 29426
rect 30818 29374 30830 29426
rect 30882 29374 30894 29426
rect 31826 29374 31838 29426
rect 31890 29374 31902 29426
rect 33058 29374 33070 29426
rect 33122 29374 33134 29426
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 34850 29374 34862 29426
rect 34914 29374 34926 29426
rect 37202 29374 37214 29426
rect 37266 29374 37278 29426
rect 37650 29374 37662 29426
rect 37714 29374 37726 29426
rect 38322 29374 38334 29426
rect 38386 29374 38398 29426
rect 38770 29374 38782 29426
rect 38834 29374 38846 29426
rect 39778 29374 39790 29426
rect 39842 29374 39854 29426
rect 40450 29374 40462 29426
rect 40514 29374 40526 29426
rect 45826 29374 45838 29426
rect 45890 29374 45902 29426
rect 47506 29374 47518 29426
rect 47570 29374 47582 29426
rect 49522 29374 49534 29426
rect 49586 29374 49598 29426
rect 21086 29362 21138 29374
rect 32510 29362 32562 29374
rect 35646 29362 35698 29374
rect 46622 29362 46674 29374
rect 50318 29362 50370 29374
rect 50766 29426 50818 29438
rect 50766 29362 50818 29374
rect 50990 29426 51042 29438
rect 52782 29426 52834 29438
rect 52098 29374 52110 29426
rect 52162 29374 52174 29426
rect 50990 29362 51042 29374
rect 52782 29362 52834 29374
rect 53342 29426 53394 29438
rect 53890 29374 53902 29426
rect 53954 29374 53966 29426
rect 53342 29362 53394 29374
rect 3278 29314 3330 29326
rect 1586 29262 1598 29314
rect 1650 29262 1662 29314
rect 3278 29250 3330 29262
rect 4958 29314 5010 29326
rect 11230 29314 11282 29326
rect 7746 29262 7758 29314
rect 7810 29262 7822 29314
rect 4958 29250 5010 29262
rect 11230 29250 11282 29262
rect 11902 29314 11954 29326
rect 11902 29250 11954 29262
rect 12238 29314 12290 29326
rect 16382 29314 16434 29326
rect 20638 29314 20690 29326
rect 34302 29314 34354 29326
rect 35534 29314 35586 29326
rect 14130 29262 14142 29314
rect 14194 29262 14206 29314
rect 19058 29262 19070 29314
rect 19122 29262 19134 29314
rect 22082 29262 22094 29314
rect 22146 29262 22158 29314
rect 24434 29262 24446 29314
rect 24498 29262 24510 29314
rect 26562 29262 26574 29314
rect 26626 29262 26638 29314
rect 32946 29262 32958 29314
rect 33010 29262 33022 29314
rect 34514 29262 34526 29314
rect 34578 29262 34590 29314
rect 12238 29250 12290 29262
rect 16382 29250 16434 29262
rect 20638 29250 20690 29262
rect 34302 29250 34354 29262
rect 35534 29250 35586 29262
rect 36318 29314 36370 29326
rect 36318 29250 36370 29262
rect 36766 29314 36818 29326
rect 46398 29314 46450 29326
rect 37762 29262 37774 29314
rect 37826 29262 37838 29314
rect 45490 29262 45502 29314
rect 45554 29262 45566 29314
rect 36766 29250 36818 29262
rect 46398 29250 46450 29262
rect 46958 29314 47010 29326
rect 46958 29250 47010 29262
rect 49870 29314 49922 29326
rect 49870 29250 49922 29262
rect 50206 29314 50258 29326
rect 50206 29250 50258 29262
rect 52446 29314 52498 29326
rect 54226 29262 54238 29314
rect 54290 29262 54302 29314
rect 52446 29250 52498 29262
rect 3390 29202 3442 29214
rect 3390 29138 3442 29150
rect 5070 29202 5122 29214
rect 5070 29138 5122 29150
rect 9550 29202 9602 29214
rect 9550 29138 9602 29150
rect 11342 29202 11394 29214
rect 11342 29138 11394 29150
rect 12126 29202 12178 29214
rect 12126 29138 12178 29150
rect 16494 29202 16546 29214
rect 16494 29138 16546 29150
rect 20750 29202 20802 29214
rect 20750 29138 20802 29150
rect 25566 29202 25618 29214
rect 30270 29202 30322 29214
rect 29138 29150 29150 29202
rect 29202 29150 29214 29202
rect 25566 29138 25618 29150
rect 30270 29138 30322 29150
rect 35086 29202 35138 29214
rect 35086 29138 35138 29150
rect 35310 29202 35362 29214
rect 44270 29202 44322 29214
rect 49086 29202 49138 29214
rect 41010 29150 41022 29202
rect 41074 29150 41086 29202
rect 47954 29150 47966 29202
rect 48018 29150 48030 29202
rect 35310 29138 35362 29150
rect 44270 29138 44322 29150
rect 49086 29138 49138 29150
rect 49758 29202 49810 29214
rect 49758 29138 49810 29150
rect 51102 29202 51154 29214
rect 51102 29138 51154 29150
rect 52558 29202 52610 29214
rect 52558 29138 52610 29150
rect 53230 29202 53282 29214
rect 53230 29138 53282 29150
rect 55918 29202 55970 29214
rect 56242 29150 56254 29202
rect 56306 29150 56318 29202
rect 55918 29138 55970 29150
rect 672 29034 56784 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 44466 29034
rect 44518 28982 44570 29034
rect 44622 28982 44674 29034
rect 44726 28982 56784 29034
rect 672 28948 56784 28982
rect 2830 28866 2882 28878
rect 2830 28802 2882 28814
rect 11902 28866 11954 28878
rect 11902 28802 11954 28814
rect 18510 28866 18562 28878
rect 18510 28802 18562 28814
rect 19070 28866 19122 28878
rect 19070 28802 19122 28814
rect 19182 28866 19234 28878
rect 19182 28802 19234 28814
rect 19406 28866 19458 28878
rect 19406 28802 19458 28814
rect 19854 28866 19906 28878
rect 19854 28802 19906 28814
rect 20078 28866 20130 28878
rect 31726 28866 31778 28878
rect 26450 28814 26462 28866
rect 26514 28814 26526 28866
rect 29026 28814 29038 28866
rect 29090 28814 29102 28866
rect 20078 28802 20130 28814
rect 31726 28802 31778 28814
rect 38334 28866 38386 28878
rect 38334 28802 38386 28814
rect 38782 28866 38834 28878
rect 46286 28866 46338 28878
rect 40898 28814 40910 28866
rect 40962 28814 40974 28866
rect 38782 28802 38834 28814
rect 46286 28802 46338 28814
rect 46398 28866 46450 28878
rect 46398 28802 46450 28814
rect 46510 28866 46562 28878
rect 46510 28802 46562 28814
rect 46734 28866 46786 28878
rect 53342 28866 53394 28878
rect 51090 28814 51102 28866
rect 51154 28814 51166 28866
rect 46734 28802 46786 28814
rect 53342 28802 53394 28814
rect 55022 28866 55074 28878
rect 55022 28802 55074 28814
rect 55918 28866 55970 28878
rect 56242 28814 56254 28866
rect 56306 28814 56318 28866
rect 55918 28802 55970 28814
rect 3502 28754 3554 28766
rect 9326 28754 9378 28766
rect 20190 28754 20242 28766
rect 1586 28702 1598 28754
rect 1650 28702 1662 28754
rect 4946 28702 4958 28754
rect 5010 28702 5022 28754
rect 7522 28702 7534 28754
rect 7586 28702 7598 28754
rect 10770 28702 10782 28754
rect 10834 28702 10846 28754
rect 13570 28702 13582 28754
rect 13634 28702 13646 28754
rect 17378 28702 17390 28754
rect 17442 28702 17454 28754
rect 3502 28690 3554 28702
rect 9326 28690 9378 28702
rect 20190 28690 20242 28702
rect 20638 28754 20690 28766
rect 27582 28754 27634 28766
rect 21634 28702 21646 28754
rect 21698 28702 21710 28754
rect 20638 28690 20690 28702
rect 27582 28690 27634 28702
rect 28030 28754 28082 28766
rect 28030 28690 28082 28702
rect 31614 28754 31666 28766
rect 31614 28690 31666 28702
rect 32398 28754 32450 28766
rect 36094 28754 36146 28766
rect 47406 28754 47458 28766
rect 33394 28702 33406 28754
rect 33458 28702 33470 28754
rect 37202 28702 37214 28754
rect 37266 28702 37278 28754
rect 43698 28702 43710 28754
rect 43762 28702 43774 28754
rect 32398 28690 32450 28702
rect 36094 28690 36146 28702
rect 47406 28690 47458 28702
rect 47630 28754 47682 28766
rect 49298 28702 49310 28754
rect 49362 28702 49374 28754
rect 50082 28702 50094 28754
rect 50146 28702 50158 28754
rect 47630 28690 47682 28702
rect 3278 28642 3330 28654
rect 3278 28578 3330 28590
rect 3614 28642 3666 28654
rect 3614 28578 3666 28590
rect 3950 28642 4002 28654
rect 5406 28642 5458 28654
rect 8206 28642 8258 28654
rect 4386 28590 4398 28642
rect 4450 28590 4462 28642
rect 4834 28590 4846 28642
rect 4898 28590 4910 28642
rect 6066 28590 6078 28642
rect 6130 28590 6142 28642
rect 7074 28590 7086 28642
rect 7138 28590 7150 28642
rect 7746 28590 7758 28642
rect 7810 28590 7822 28642
rect 3950 28578 4002 28590
rect 5406 28578 5458 28590
rect 8206 28578 8258 28590
rect 8878 28642 8930 28654
rect 8878 28578 8930 28590
rect 9102 28642 9154 28654
rect 9102 28578 9154 28590
rect 12574 28642 12626 28654
rect 14254 28642 14306 28654
rect 22094 28642 22146 28654
rect 29710 28642 29762 28654
rect 34078 28642 34130 28654
rect 35982 28642 36034 28654
rect 13010 28590 13022 28642
rect 13074 28590 13086 28642
rect 13346 28590 13358 28642
rect 13410 28590 13422 28642
rect 14578 28590 14590 28642
rect 14642 28590 14654 28642
rect 15586 28590 15598 28642
rect 15650 28590 15662 28642
rect 16930 28590 16942 28642
rect 16994 28590 17006 28642
rect 19618 28590 19630 28642
rect 19682 28590 19694 28642
rect 20962 28590 20974 28642
rect 21026 28590 21038 28642
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 22642 28590 22654 28642
rect 22706 28590 22718 28642
rect 23650 28590 23662 28642
rect 23714 28590 23726 28642
rect 28354 28590 28366 28642
rect 28418 28590 28430 28642
rect 28914 28590 28926 28642
rect 28978 28590 28990 28642
rect 30034 28590 30046 28642
rect 30098 28590 30110 28642
rect 31042 28590 31054 28642
rect 31106 28590 31118 28642
rect 32722 28590 32734 28642
rect 32786 28590 32798 28642
rect 33170 28590 33182 28642
rect 33234 28590 33246 28642
rect 34402 28590 34414 28642
rect 34466 28590 34478 28642
rect 35522 28590 35534 28642
rect 35586 28590 35598 28642
rect 12574 28578 12626 28590
rect 14254 28578 14306 28590
rect 22094 28578 22146 28590
rect 29710 28578 29762 28590
rect 34078 28578 34130 28590
rect 35982 28578 36034 28590
rect 36318 28642 36370 28654
rect 39006 28642 39058 28654
rect 36642 28590 36654 28642
rect 36706 28590 36718 28642
rect 36318 28578 36370 28590
rect 39006 28578 39058 28590
rect 39454 28642 39506 28654
rect 47294 28642 47346 28654
rect 40450 28590 40462 28642
rect 40514 28590 40526 28642
rect 43138 28590 43150 28642
rect 43202 28590 43214 28642
rect 43474 28590 43486 28642
rect 43538 28590 43550 28642
rect 44258 28590 44270 28642
rect 44322 28590 44334 28642
rect 44706 28590 44718 28642
rect 44770 28590 44782 28642
rect 45714 28590 45726 28642
rect 45778 28590 45790 28642
rect 39454 28578 39506 28590
rect 47294 28578 47346 28590
rect 48190 28642 48242 28654
rect 49758 28642 49810 28654
rect 48962 28590 48974 28642
rect 49026 28590 49038 28642
rect 48190 28578 48242 28590
rect 49758 28578 49810 28590
rect 52894 28642 52946 28654
rect 52894 28578 52946 28590
rect 53118 28642 53170 28654
rect 53118 28578 53170 28590
rect 53902 28642 53954 28654
rect 53902 28578 53954 28590
rect 54126 28642 54178 28654
rect 54126 28578 54178 28590
rect 54350 28642 54402 28654
rect 54350 28578 54402 28590
rect 8990 28530 9042 28542
rect 19294 28530 19346 28542
rect 38894 28530 38946 28542
rect 1250 28478 1262 28530
rect 1314 28478 1326 28530
rect 10322 28478 10334 28530
rect 10386 28478 10398 28530
rect 26002 28478 26014 28530
rect 26066 28478 26078 28530
rect 8990 28466 9042 28478
rect 19294 28466 19346 28478
rect 38894 28466 38946 28478
rect 42702 28530 42754 28542
rect 53230 28530 53282 28542
rect 50642 28478 50654 28530
rect 50706 28478 50718 28530
rect 42702 28466 42754 28478
rect 53230 28466 53282 28478
rect 54014 28530 54066 28542
rect 54014 28466 54066 28478
rect 8318 28418 8370 28430
rect 8318 28354 8370 28366
rect 31726 28418 31778 28430
rect 31726 28354 31778 28366
rect 42030 28418 42082 28430
rect 42030 28354 42082 28366
rect 48526 28418 48578 28430
rect 48526 28354 48578 28366
rect 52222 28418 52274 28430
rect 52222 28354 52274 28366
rect 52670 28418 52722 28430
rect 52670 28354 52722 28366
rect 54574 28418 54626 28430
rect 54574 28354 54626 28366
rect 54910 28418 54962 28430
rect 54910 28354 54962 28366
rect 55246 28418 55298 28430
rect 55246 28354 55298 28366
rect 672 28250 56784 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 43806 28250
rect 43858 28198 43910 28250
rect 43962 28198 44014 28250
rect 44066 28198 56784 28250
rect 672 28164 56784 28198
rect 11454 28082 11506 28094
rect 11454 28018 11506 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 32510 28082 32562 28094
rect 32510 28018 32562 28030
rect 33070 28082 33122 28094
rect 33070 28018 33122 28030
rect 38110 28082 38162 28094
rect 38110 28018 38162 28030
rect 43374 28082 43426 28094
rect 43374 28018 43426 28030
rect 44606 28082 44658 28094
rect 44606 28018 44658 28030
rect 51998 28082 52050 28094
rect 51998 28018 52050 28030
rect 53342 28082 53394 28094
rect 53342 28018 53394 28030
rect 53902 28082 53954 28094
rect 53902 28018 53954 28030
rect 4398 27970 4450 27982
rect 13694 27970 13746 27982
rect 39790 27970 39842 27982
rect 9314 27918 9326 27970
rect 9378 27918 9390 27970
rect 9874 27918 9886 27970
rect 9938 27918 9950 27970
rect 17490 27918 17502 27970
rect 17554 27918 17566 27970
rect 21858 27918 21870 27970
rect 21922 27918 21934 27970
rect 38882 27918 38894 27970
rect 38946 27918 38958 27970
rect 4398 27906 4450 27918
rect 13694 27906 13746 27918
rect 39790 27906 39842 27918
rect 44494 27970 44546 27982
rect 46386 27918 46398 27970
rect 46450 27918 46462 27970
rect 52210 27918 52222 27970
rect 52274 27918 52286 27970
rect 44494 27906 44546 27918
rect 12798 27858 12850 27870
rect 1362 27806 1374 27858
rect 1426 27806 1438 27858
rect 2370 27806 2382 27858
rect 2434 27806 2446 27858
rect 3490 27806 3502 27858
rect 3554 27806 3566 27858
rect 3938 27806 3950 27858
rect 4002 27806 4014 27858
rect 5282 27806 5294 27858
rect 5346 27806 5358 27858
rect 5842 27806 5854 27858
rect 5906 27806 5918 27858
rect 7186 27806 7198 27858
rect 7250 27806 7262 27858
rect 7970 27806 7982 27858
rect 8034 27806 8046 27858
rect 9202 27806 9214 27858
rect 9266 27806 9278 27858
rect 12798 27794 12850 27806
rect 13358 27858 13410 27870
rect 19070 27858 19122 27870
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 14578 27806 14590 27858
rect 14642 27806 14654 27858
rect 15698 27806 15710 27858
rect 15762 27806 15774 27858
rect 16706 27806 16718 27858
rect 16770 27806 16782 27858
rect 13358 27794 13410 27806
rect 19070 27794 19122 27806
rect 19630 27858 19682 27870
rect 19630 27794 19682 27806
rect 19742 27858 19794 27870
rect 19742 27794 19794 27806
rect 20078 27858 20130 27870
rect 20078 27794 20130 27806
rect 20638 27858 20690 27870
rect 20638 27794 20690 27806
rect 23438 27858 23490 27870
rect 25566 27858 25618 27870
rect 35198 27858 35250 27870
rect 24210 27806 24222 27858
rect 24274 27806 24286 27858
rect 24770 27806 24782 27858
rect 24834 27806 24846 27858
rect 25890 27806 25902 27858
rect 25954 27806 25966 27858
rect 27010 27806 27022 27858
rect 27074 27806 27086 27858
rect 27682 27806 27694 27858
rect 27746 27806 27758 27858
rect 30146 27806 30158 27858
rect 30210 27806 30222 27858
rect 30818 27806 30830 27858
rect 30882 27806 30894 27858
rect 34626 27806 34638 27858
rect 34690 27806 34702 27858
rect 23438 27794 23490 27806
rect 25566 27794 25618 27806
rect 35198 27794 35250 27806
rect 35758 27858 35810 27870
rect 38558 27858 38610 27870
rect 39678 27858 39730 27870
rect 36530 27806 36542 27858
rect 36594 27806 36606 27858
rect 39218 27806 39230 27858
rect 39282 27806 39294 27858
rect 35758 27794 35810 27806
rect 38558 27794 38610 27806
rect 39678 27794 39730 27806
rect 40014 27858 40066 27870
rect 40014 27794 40066 27806
rect 40126 27858 40178 27870
rect 40126 27794 40178 27806
rect 40910 27858 40962 27870
rect 44942 27858 44994 27870
rect 41794 27806 41806 27858
rect 41858 27806 41870 27858
rect 40910 27794 40962 27806
rect 44942 27794 44994 27806
rect 45054 27858 45106 27870
rect 45054 27794 45106 27806
rect 45502 27858 45554 27870
rect 52110 27858 52162 27870
rect 50306 27806 50318 27858
rect 50370 27806 50382 27858
rect 45502 27794 45554 27806
rect 52110 27794 52162 27806
rect 52558 27858 52610 27870
rect 52558 27794 52610 27806
rect 52782 27858 52834 27870
rect 55570 27806 55582 27858
rect 55634 27806 55646 27858
rect 52782 27794 52834 27806
rect 2942 27746 2994 27758
rect 4958 27746 5010 27758
rect 3378 27694 3390 27746
rect 3442 27694 3454 27746
rect 2942 27682 2994 27694
rect 4958 27682 5010 27694
rect 6414 27746 6466 27758
rect 6414 27682 6466 27694
rect 8542 27746 8594 27758
rect 8542 27682 8594 27694
rect 8878 27746 8930 27758
rect 12126 27746 12178 27758
rect 10210 27694 10222 27746
rect 10274 27694 10286 27746
rect 8878 27682 8930 27694
rect 12126 27682 12178 27694
rect 12238 27746 12290 27758
rect 12238 27682 12290 27694
rect 13022 27746 13074 27758
rect 15150 27746 15202 27758
rect 14690 27694 14702 27746
rect 14754 27694 14766 27746
rect 13022 27682 13074 27694
rect 15150 27682 15202 27694
rect 21310 27746 21362 27758
rect 21310 27682 21362 27694
rect 23886 27746 23938 27758
rect 35422 27746 35474 27758
rect 38894 27746 38946 27758
rect 45278 27746 45330 27758
rect 53342 27746 53394 27758
rect 24882 27694 24894 27746
rect 24946 27694 24958 27746
rect 27906 27694 27918 27746
rect 27970 27694 27982 27746
rect 31378 27694 31390 27746
rect 31442 27694 31454 27746
rect 34178 27694 34190 27746
rect 34242 27694 34254 27746
rect 36978 27694 36990 27746
rect 37042 27694 37054 27746
rect 42130 27694 42142 27746
rect 42194 27694 42206 27746
rect 48066 27694 48078 27746
rect 48130 27694 48142 27746
rect 23886 27682 23938 27694
rect 35422 27682 35474 27694
rect 38894 27682 38946 27694
rect 45278 27682 45330 27694
rect 53342 27682 53394 27694
rect 53454 27746 53506 27758
rect 55010 27694 55022 27746
rect 55074 27694 55086 27746
rect 56354 27694 56366 27746
rect 56418 27694 56430 27746
rect 53454 27682 53506 27694
rect 8766 27634 8818 27646
rect 5954 27582 5966 27634
rect 6018 27582 6030 27634
rect 8766 27570 8818 27582
rect 11902 27634 11954 27646
rect 11902 27570 11954 27582
rect 13246 27634 13298 27646
rect 19854 27634 19906 27646
rect 17938 27582 17950 27634
rect 18002 27582 18014 27634
rect 13246 27570 13298 27582
rect 19854 27570 19906 27582
rect 20974 27634 21026 27646
rect 20974 27570 21026 27582
rect 21198 27634 21250 27646
rect 35646 27634 35698 27646
rect 22306 27582 22318 27634
rect 22370 27582 22382 27634
rect 30370 27582 30382 27634
rect 30434 27582 30446 27634
rect 21198 27570 21250 27582
rect 35646 27570 35698 27582
rect 38782 27634 38834 27646
rect 38782 27570 38834 27582
rect 40686 27634 40738 27646
rect 40686 27570 40738 27582
rect 40798 27634 40850 27646
rect 40798 27570 40850 27582
rect 41134 27634 41186 27646
rect 41134 27570 41186 27582
rect 56030 27634 56082 27646
rect 56030 27570 56082 27582
rect 672 27466 56784 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 44466 27466
rect 44518 27414 44570 27466
rect 44622 27414 44674 27466
rect 44726 27414 56784 27466
rect 672 27380 56784 27414
rect 2830 27298 2882 27310
rect 1698 27246 1710 27298
rect 1762 27246 1774 27298
rect 2830 27234 2882 27246
rect 3502 27298 3554 27310
rect 3502 27234 3554 27246
rect 7758 27298 7810 27310
rect 7758 27234 7810 27246
rect 7870 27298 7922 27310
rect 12014 27298 12066 27310
rect 20302 27298 20354 27310
rect 31838 27298 31890 27310
rect 38670 27298 38722 27310
rect 10098 27246 10110 27298
rect 10162 27246 10174 27298
rect 13906 27246 13918 27298
rect 13970 27246 13982 27298
rect 19170 27246 19182 27298
rect 19234 27246 19246 27298
rect 27570 27246 27582 27298
rect 27634 27246 27646 27298
rect 37538 27246 37550 27298
rect 37602 27246 37614 27298
rect 7870 27234 7922 27246
rect 12014 27234 12066 27246
rect 20302 27234 20354 27246
rect 31838 27234 31890 27246
rect 38670 27234 38722 27246
rect 41694 27298 41746 27310
rect 47294 27298 47346 27310
rect 54910 27298 54962 27310
rect 45490 27246 45502 27298
rect 45554 27246 45566 27298
rect 53778 27246 53790 27298
rect 53842 27246 53854 27298
rect 41694 27234 41746 27246
rect 47294 27234 47346 27246
rect 54910 27234 54962 27246
rect 55022 27298 55074 27310
rect 55022 27234 55074 27246
rect 56142 27298 56194 27310
rect 56142 27234 56194 27246
rect 3614 27186 3666 27198
rect 3614 27122 3666 27134
rect 3950 27186 4002 27198
rect 5406 27186 5458 27198
rect 4946 27134 4958 27186
rect 5010 27134 5022 27186
rect 3950 27122 4002 27134
rect 5406 27122 5458 27134
rect 7982 27186 8034 27198
rect 7982 27122 8034 27134
rect 11902 27186 11954 27198
rect 11902 27122 11954 27134
rect 12462 27186 12514 27198
rect 12462 27122 12514 27134
rect 12910 27186 12962 27198
rect 12910 27122 12962 27134
rect 14366 27186 14418 27198
rect 22206 27186 22258 27198
rect 21746 27134 21758 27186
rect 21810 27134 21822 27186
rect 14366 27122 14418 27134
rect 22206 27122 22258 27134
rect 26574 27186 26626 27198
rect 26574 27122 26626 27134
rect 31726 27186 31778 27198
rect 40910 27186 40962 27198
rect 33730 27134 33742 27186
rect 33794 27134 33806 27186
rect 35186 27134 35198 27186
rect 35250 27134 35262 27186
rect 31726 27122 31778 27134
rect 40910 27122 40962 27134
rect 41806 27186 41858 27198
rect 41806 27122 41858 27134
rect 42254 27186 42306 27198
rect 47406 27186 47458 27198
rect 52670 27186 52722 27198
rect 43250 27134 43262 27186
rect 43314 27134 43326 27186
rect 49410 27134 49422 27186
rect 49474 27134 49486 27186
rect 50866 27134 50878 27186
rect 50930 27134 50942 27186
rect 42254 27122 42306 27134
rect 47406 27122 47458 27134
rect 52670 27122 52722 27134
rect 8430 27074 8482 27086
rect 12350 27074 12402 27086
rect 1138 27022 1150 27074
rect 1202 27022 1214 27074
rect 4386 27022 4398 27074
rect 4450 27022 4462 27074
rect 4722 27022 4734 27074
rect 4786 27022 4798 27074
rect 6066 27022 6078 27074
rect 6130 27022 6142 27074
rect 6962 27022 6974 27074
rect 7026 27022 7038 27074
rect 10658 27022 10670 27074
rect 10722 27022 10734 27074
rect 8430 27010 8482 27022
rect 12350 27010 12402 27022
rect 12686 27074 12738 27086
rect 20750 27074 20802 27086
rect 22430 27074 22482 27086
rect 28030 27074 28082 27086
rect 39118 27074 39170 27086
rect 13234 27022 13246 27074
rect 13298 27022 13310 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 15026 27022 15038 27074
rect 15090 27022 15102 27074
rect 16034 27022 16046 27074
rect 16098 27022 16110 27074
rect 18722 27022 18734 27074
rect 18786 27022 18798 27074
rect 21074 27022 21086 27074
rect 21138 27022 21150 27074
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 22754 27022 22766 27074
rect 22818 27022 22830 27074
rect 23762 27022 23774 27074
rect 23826 27022 23838 27074
rect 26898 27022 26910 27074
rect 26962 27022 26974 27074
rect 12686 27010 12738 27022
rect 20750 27010 20802 27022
rect 22430 27010 22482 27022
rect 27346 27010 27358 27062
rect 27410 27010 27422 27062
rect 28578 27022 28590 27074
rect 28642 27022 28654 27074
rect 29586 27022 29598 27074
rect 29650 27022 29662 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 37090 27022 37102 27074
rect 37154 27022 37166 27074
rect 28030 27010 28082 27022
rect 39118 27010 39170 27022
rect 40238 27074 40290 27086
rect 40238 27010 40290 27022
rect 40574 27074 40626 27086
rect 40574 27010 40626 27022
rect 41134 27074 41186 27086
rect 41134 27010 41186 27022
rect 41582 27074 41634 27086
rect 42802 27022 42814 27074
rect 42866 27022 42878 27074
rect 45042 27022 45054 27074
rect 45106 27022 45118 27074
rect 49858 27022 49870 27074
rect 49922 27022 49934 27074
rect 50418 27022 50430 27074
rect 50482 27022 50494 27074
rect 41582 27010 41634 27022
rect 31278 26962 31330 26974
rect 31278 26898 31330 26910
rect 31390 26962 31442 26974
rect 39342 26962 39394 26974
rect 34066 26910 34078 26962
rect 34130 26910 34142 26962
rect 31390 26898 31442 26910
rect 39342 26898 39394 26910
rect 40462 26962 40514 26974
rect 40462 26898 40514 26910
rect 48190 26962 48242 26974
rect 55918 26962 55970 26974
rect 54226 26910 54238 26962
rect 54290 26910 54302 26962
rect 56130 26910 56142 26962
rect 56194 26910 56206 26962
rect 48190 26898 48242 26910
rect 55918 26898 55970 26910
rect 3502 26850 3554 26862
rect 3502 26786 3554 26798
rect 8990 26850 9042 26862
rect 8990 26786 9042 26798
rect 32510 26850 32562 26862
rect 32510 26786 32562 26798
rect 36430 26850 36482 26862
rect 42142 26850 42194 26862
rect 39666 26798 39678 26850
rect 39730 26798 39742 26850
rect 36430 26786 36482 26798
rect 42142 26786 42194 26798
rect 44382 26850 44434 26862
rect 44382 26786 44434 26798
rect 46622 26850 46674 26862
rect 46622 26786 46674 26798
rect 47182 26850 47234 26862
rect 47182 26786 47234 26798
rect 52110 26850 52162 26862
rect 52110 26786 52162 26798
rect 54798 26850 54850 26862
rect 54798 26786 54850 26798
rect 672 26682 56784 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 43806 26682
rect 43858 26630 43910 26682
rect 43962 26630 44014 26682
rect 44066 26630 56784 26682
rect 672 26596 56784 26630
rect 2830 26514 2882 26526
rect 2830 26450 2882 26462
rect 9214 26514 9266 26526
rect 9214 26450 9266 26462
rect 9774 26514 9826 26526
rect 9774 26450 9826 26462
rect 10334 26514 10386 26526
rect 10334 26450 10386 26462
rect 35758 26514 35810 26526
rect 35758 26450 35810 26462
rect 43150 26514 43202 26526
rect 51998 26514 52050 26526
rect 49746 26462 49758 26514
rect 49810 26462 49822 26514
rect 43150 26450 43202 26462
rect 51998 26450 52050 26462
rect 55246 26514 55298 26526
rect 55246 26450 55298 26462
rect 3278 26402 3330 26414
rect 17278 26402 17330 26414
rect 21310 26402 21362 26414
rect 28702 26402 28754 26414
rect 6626 26350 6638 26402
rect 6690 26350 6702 26402
rect 7634 26350 7646 26402
rect 7698 26350 7710 26402
rect 18386 26350 18398 26402
rect 18450 26350 18462 26402
rect 26226 26350 26238 26402
rect 26290 26350 26302 26402
rect 3278 26338 3330 26350
rect 17278 26338 17330 26350
rect 21310 26338 21362 26350
rect 28702 26338 28754 26350
rect 35646 26402 35698 26414
rect 49198 26402 49250 26414
rect 37874 26350 37886 26402
rect 37938 26350 37950 26402
rect 46610 26350 46622 26402
rect 46674 26350 46686 26402
rect 48738 26350 48750 26402
rect 48802 26350 48814 26402
rect 35646 26338 35698 26350
rect 49198 26338 49250 26350
rect 49422 26402 49474 26414
rect 49422 26338 49474 26350
rect 52558 26402 52610 26414
rect 52558 26338 52610 26350
rect 3950 26290 4002 26302
rect 1250 26238 1262 26290
rect 1314 26238 1326 26290
rect 3950 26226 4002 26238
rect 4174 26290 4226 26302
rect 9662 26290 9714 26302
rect 13022 26290 13074 26302
rect 4386 26238 4398 26290
rect 4450 26238 4462 26290
rect 12786 26238 12798 26290
rect 12850 26238 12862 26290
rect 4174 26226 4226 26238
rect 9662 26226 9714 26238
rect 13022 26226 13074 26238
rect 13246 26290 13298 26302
rect 16830 26290 16882 26302
rect 13458 26238 13470 26290
rect 13522 26238 13534 26290
rect 13246 26226 13298 26238
rect 16830 26226 16882 26238
rect 17054 26290 17106 26302
rect 17054 26226 17106 26238
rect 20974 26290 21026 26302
rect 27806 26290 27858 26302
rect 30382 26290 30434 26302
rect 40126 26290 40178 26302
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 22194 26238 22206 26290
rect 22258 26238 22270 26290
rect 23314 26238 23326 26290
rect 23378 26238 23390 26290
rect 24322 26238 24334 26290
rect 24386 26238 24398 26290
rect 26114 26238 26126 26290
rect 26178 26238 26190 26290
rect 29026 26238 29038 26290
rect 29090 26238 29102 26290
rect 29586 26238 29598 26290
rect 29650 26238 29662 26290
rect 30930 26238 30942 26290
rect 30994 26238 31006 26290
rect 31826 26238 31838 26290
rect 31890 26238 31902 26290
rect 32386 26238 32398 26290
rect 32450 26238 32462 26290
rect 34514 26238 34526 26290
rect 34578 26238 34590 26290
rect 20974 26226 21026 26238
rect 27806 26226 27858 26238
rect 30382 26226 30434 26238
rect 40126 26226 40178 26238
rect 40798 26290 40850 26302
rect 40798 26226 40850 26238
rect 41470 26290 41522 26302
rect 41470 26226 41522 26238
rect 42926 26290 42978 26302
rect 42926 26226 42978 26238
rect 43262 26290 43314 26302
rect 43262 26226 43314 26238
rect 45614 26290 45666 26302
rect 50542 26290 50594 26302
rect 52222 26290 52274 26302
rect 45938 26238 45950 26290
rect 46002 26238 46014 26290
rect 51202 26238 51214 26290
rect 51266 26238 51278 26290
rect 45614 26226 45666 26238
rect 50542 26226 50594 26238
rect 52222 26226 52274 26238
rect 52446 26290 52498 26302
rect 52446 26226 52498 26238
rect 52670 26290 52722 26302
rect 53554 26238 53566 26290
rect 53618 26238 53630 26290
rect 56130 26238 56142 26290
rect 56194 26238 56206 26290
rect 52670 26226 52722 26238
rect 9774 26178 9826 26190
rect 6290 26126 6302 26178
rect 6354 26126 6366 26178
rect 8082 26126 8094 26178
rect 8146 26126 8158 26178
rect 9774 26114 9826 26126
rect 10222 26178 10274 26190
rect 10222 26114 10274 26126
rect 10334 26178 10386 26190
rect 10334 26114 10386 26126
rect 17614 26178 17666 26190
rect 20862 26178 20914 26190
rect 18834 26126 18846 26178
rect 18898 26126 18910 26178
rect 17614 26114 17666 26126
rect 20862 26114 20914 26126
rect 22766 26178 22818 26190
rect 22766 26114 22818 26126
rect 25006 26178 25058 26190
rect 34974 26178 35026 26190
rect 26562 26126 26574 26178
rect 26626 26126 26638 26178
rect 29698 26126 29710 26178
rect 29762 26126 29774 26178
rect 25006 26114 25058 26126
rect 34974 26114 35026 26126
rect 36542 26178 36594 26190
rect 36542 26114 36594 26126
rect 36654 26178 36706 26190
rect 40574 26178 40626 26190
rect 36754 26126 36766 26178
rect 36818 26126 36830 26178
rect 38322 26126 38334 26178
rect 38386 26126 38398 26178
rect 36654 26114 36706 26126
rect 40574 26114 40626 26126
rect 41246 26178 41298 26190
rect 41246 26114 41298 26126
rect 41358 26178 41410 26190
rect 42254 26178 42306 26190
rect 41906 26126 41918 26178
rect 41970 26126 41982 26178
rect 41358 26114 41410 26126
rect 42254 26114 42306 26126
rect 42478 26178 42530 26190
rect 42478 26114 42530 26126
rect 43374 26178 43426 26190
rect 43374 26114 43426 26126
rect 45278 26178 45330 26190
rect 45278 26114 45330 26126
rect 45390 26178 45442 26190
rect 51314 26126 51326 26178
rect 51378 26126 51390 26178
rect 54002 26126 54014 26178
rect 54066 26126 54078 26178
rect 55906 26126 55918 26178
rect 55970 26126 55982 26178
rect 45390 26114 45442 26126
rect 3390 26066 3442 26078
rect 1698 26014 1710 26066
rect 1762 26014 1774 26066
rect 3390 26002 3442 26014
rect 3838 26066 3890 26078
rect 3838 26002 3890 26014
rect 4062 26066 4114 26078
rect 4062 26002 4114 26014
rect 5070 26066 5122 26078
rect 13134 26066 13186 26078
rect 6178 26014 6190 26066
rect 6242 26014 6254 26066
rect 5070 26002 5122 26014
rect 13134 26002 13186 26014
rect 17502 26066 17554 26078
rect 17502 26002 17554 26014
rect 17726 26066 17778 26078
rect 17726 26002 17778 26014
rect 19966 26066 20018 26078
rect 19966 26002 20018 26014
rect 20638 26066 20690 26078
rect 24894 26066 24946 26078
rect 34078 26066 34130 26078
rect 22306 26014 22318 26066
rect 22370 26014 22382 26066
rect 32946 26014 32958 26066
rect 33010 26014 33022 26066
rect 20638 26002 20690 26014
rect 24894 26002 24946 26014
rect 34078 26002 34130 26014
rect 35086 26066 35138 26078
rect 35086 26002 35138 26014
rect 35198 26066 35250 26078
rect 35198 26002 35250 26014
rect 35310 26066 35362 26078
rect 35310 26002 35362 26014
rect 36318 26066 36370 26078
rect 36318 26002 36370 26014
rect 36430 26066 36482 26078
rect 36430 26002 36482 26014
rect 39454 26066 39506 26078
rect 39454 26002 39506 26014
rect 40462 26066 40514 26078
rect 40462 26002 40514 26014
rect 42702 26066 42754 26078
rect 42702 26002 42754 26014
rect 50206 26066 50258 26078
rect 50206 26002 50258 26014
rect 672 25898 56784 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 44466 25898
rect 44518 25846 44570 25898
rect 44622 25846 44674 25898
rect 44726 25846 56784 25898
rect 672 25812 56784 25846
rect 2942 25730 2994 25742
rect 1810 25678 1822 25730
rect 1874 25678 1886 25730
rect 2942 25666 2994 25678
rect 4398 25730 4450 25742
rect 4398 25666 4450 25678
rect 10782 25730 10834 25742
rect 24782 25730 24834 25742
rect 27694 25730 27746 25742
rect 30382 25730 30434 25742
rect 12226 25678 12238 25730
rect 12290 25678 12302 25730
rect 26562 25678 26574 25730
rect 26626 25678 26638 25730
rect 29250 25678 29262 25730
rect 29314 25678 29326 25730
rect 10782 25666 10834 25678
rect 4062 25618 4114 25630
rect 6974 25618 7026 25630
rect 5842 25566 5854 25618
rect 5906 25566 5918 25618
rect 4062 25554 4114 25566
rect 6974 25554 7026 25566
rect 7646 25618 7698 25630
rect 7646 25554 7698 25566
rect 7758 25618 7810 25630
rect 11230 25618 11282 25630
rect 21634 25622 21646 25674
rect 21698 25622 21710 25674
rect 24782 25666 24834 25678
rect 27694 25666 27746 25678
rect 30382 25666 30434 25678
rect 36542 25730 36594 25742
rect 40686 25730 40738 25742
rect 39666 25678 39678 25730
rect 39730 25678 39742 25730
rect 36542 25666 36594 25678
rect 40686 25666 40738 25678
rect 41918 25730 41970 25742
rect 41918 25666 41970 25678
rect 42030 25730 42082 25742
rect 48190 25730 48242 25742
rect 52110 25730 52162 25742
rect 47282 25678 47294 25730
rect 47346 25678 47358 25730
rect 49298 25678 49310 25730
rect 49362 25678 49374 25730
rect 42030 25666 42082 25678
rect 48190 25666 48242 25678
rect 52110 25666 52162 25678
rect 52670 25730 52722 25742
rect 52670 25666 52722 25678
rect 31614 25618 31666 25630
rect 7858 25566 7870 25618
rect 7922 25566 7934 25618
rect 9650 25566 9662 25618
rect 9714 25566 9726 25618
rect 17714 25566 17726 25618
rect 17778 25566 17790 25618
rect 7758 25554 7810 25566
rect 11230 25554 11282 25566
rect 31614 25554 31666 25566
rect 31726 25618 31778 25630
rect 40798 25618 40850 25630
rect 42702 25618 42754 25630
rect 33618 25566 33630 25618
rect 33682 25566 33694 25618
rect 34850 25566 34862 25618
rect 34914 25566 34926 25618
rect 37538 25566 37550 25618
rect 37602 25566 37614 25618
rect 41010 25566 41022 25618
rect 41074 25566 41086 25618
rect 31726 25554 31778 25566
rect 40798 25554 40850 25566
rect 42702 25554 42754 25566
rect 43150 25618 43202 25630
rect 44146 25566 44158 25618
rect 44210 25566 44222 25618
rect 50978 25566 50990 25618
rect 51042 25566 51054 25618
rect 52994 25566 53006 25618
rect 53058 25566 53070 25618
rect 53890 25566 53902 25618
rect 53954 25566 53966 25618
rect 56242 25566 56254 25618
rect 56306 25566 56318 25618
rect 43150 25554 43202 25566
rect 4398 25506 4450 25518
rect 1250 25454 1262 25506
rect 1314 25454 1326 25506
rect 4398 25442 4450 25454
rect 4734 25506 4786 25518
rect 4734 25442 4786 25454
rect 7422 25506 7474 25518
rect 12910 25506 12962 25518
rect 18174 25506 18226 25518
rect 20638 25506 20690 25518
rect 22318 25506 22370 25518
rect 25006 25506 25058 25518
rect 39118 25506 39170 25518
rect 11666 25454 11678 25506
rect 11730 25454 11742 25506
rect 12002 25454 12014 25506
rect 12066 25454 12078 25506
rect 13234 25454 13246 25506
rect 13298 25454 13310 25506
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 17042 25454 17054 25506
rect 17106 25454 17118 25506
rect 17602 25454 17614 25506
rect 17666 25454 17678 25506
rect 18722 25454 18734 25506
rect 18786 25454 18798 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 20962 25454 20974 25506
rect 21026 25454 21038 25506
rect 7422 25442 7474 25454
rect 12910 25442 12962 25454
rect 18174 25442 18226 25454
rect 20638 25442 20690 25454
rect 21410 25442 21422 25494
rect 21474 25442 21486 25494
rect 22642 25454 22654 25506
rect 22706 25454 22718 25506
rect 23650 25454 23662 25506
rect 23714 25454 23726 25506
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 26114 25454 26126 25506
rect 26178 25454 26190 25506
rect 28802 25454 28814 25506
rect 28866 25454 28878 25506
rect 33730 25454 33742 25506
rect 33794 25454 33806 25506
rect 34402 25454 34414 25506
rect 34466 25454 34478 25506
rect 36978 25454 36990 25506
rect 37042 25454 37054 25506
rect 22318 25442 22370 25454
rect 25006 25442 25058 25454
rect 39118 25442 39170 25454
rect 40462 25506 40514 25518
rect 41470 25506 41522 25518
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 40462 25442 40514 25454
rect 41470 25442 41522 25454
rect 42142 25506 42194 25518
rect 44606 25506 44658 25518
rect 46734 25506 46786 25518
rect 55918 25506 55970 25518
rect 43586 25454 43598 25506
rect 43650 25454 43662 25506
rect 44034 25454 44046 25506
rect 44098 25454 44110 25506
rect 45378 25454 45390 25506
rect 45442 25454 45454 25506
rect 46162 25454 46174 25506
rect 46226 25454 46238 25506
rect 50530 25454 50542 25506
rect 50594 25454 50606 25506
rect 42142 25442 42194 25454
rect 44606 25442 44658 25454
rect 46734 25442 46786 25454
rect 55918 25442 55970 25454
rect 7534 25394 7586 25406
rect 16718 25394 16770 25406
rect 5394 25342 5406 25394
rect 5458 25342 5470 25394
rect 9202 25342 9214 25394
rect 9266 25342 9278 25394
rect 7534 25330 7586 25342
rect 16718 25330 16770 25342
rect 24894 25394 24946 25406
rect 24894 25330 24946 25342
rect 36430 25394 36482 25406
rect 41234 25342 41246 25394
rect 41298 25342 41310 25394
rect 42690 25342 42702 25394
rect 42754 25342 42766 25394
rect 49746 25342 49758 25394
rect 49810 25342 49822 25394
rect 53554 25342 53566 25394
rect 53618 25342 53630 25394
rect 36430 25330 36482 25342
rect 31726 25282 31778 25294
rect 31726 25218 31778 25230
rect 32622 25282 32674 25294
rect 32622 25218 32674 25230
rect 32958 25282 33010 25294
rect 32958 25218 33010 25230
rect 35982 25282 36034 25294
rect 35982 25218 36034 25230
rect 38670 25282 38722 25294
rect 38670 25218 38722 25230
rect 39342 25282 39394 25294
rect 39342 25218 39394 25230
rect 42478 25282 42530 25294
rect 42478 25218 42530 25230
rect 46958 25282 47010 25294
rect 46958 25218 47010 25230
rect 55134 25282 55186 25294
rect 55134 25218 55186 25230
rect 672 25114 56784 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 43806 25114
rect 43858 25062 43910 25114
rect 43962 25062 44014 25114
rect 44066 25062 56784 25114
rect 672 25028 56784 25062
rect 5070 24946 5122 24958
rect 5070 24882 5122 24894
rect 5518 24946 5570 24958
rect 5518 24882 5570 24894
rect 25566 24946 25618 24958
rect 25566 24882 25618 24894
rect 41246 24946 41298 24958
rect 41246 24882 41298 24894
rect 44270 24946 44322 24958
rect 44270 24882 44322 24894
rect 48974 24946 49026 24958
rect 48974 24882 49026 24894
rect 52446 24946 52498 24958
rect 52446 24882 52498 24894
rect 6414 24834 6466 24846
rect 6414 24770 6466 24782
rect 6862 24834 6914 24846
rect 6862 24770 6914 24782
rect 21086 24834 21138 24846
rect 23986 24782 23998 24834
rect 24050 24782 24062 24834
rect 26226 24782 26238 24834
rect 26290 24782 26302 24834
rect 34066 24782 34078 24834
rect 34130 24782 34142 24834
rect 36530 24782 36542 24834
rect 36594 24782 36606 24834
rect 39666 24782 39678 24834
rect 39730 24782 39742 24834
rect 41906 24782 41918 24834
rect 41970 24782 41982 24834
rect 47394 24782 47406 24834
rect 47458 24782 47470 24834
rect 51090 24782 51102 24834
rect 51154 24782 51166 24834
rect 21086 24770 21138 24782
rect 2830 24722 2882 24734
rect 6302 24722 6354 24734
rect 21310 24722 21362 24734
rect 32734 24722 32786 24734
rect 1474 24670 1486 24722
rect 1538 24670 1550 24722
rect 1922 24670 1934 24722
rect 1986 24670 1998 24722
rect 3266 24670 3278 24722
rect 3330 24670 3342 24722
rect 4162 24670 4174 24722
rect 4226 24670 4238 24722
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 7634 24670 7646 24722
rect 7698 24670 7710 24722
rect 8418 24670 8430 24722
rect 8482 24670 8494 24722
rect 9090 24670 9102 24722
rect 9154 24670 9166 24722
rect 9986 24670 9998 24722
rect 10050 24670 10062 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 17042 24670 17054 24722
rect 17106 24670 17118 24722
rect 17378 24670 17390 24722
rect 17442 24670 17454 24722
rect 18162 24670 18174 24722
rect 18226 24670 18238 24722
rect 18834 24670 18846 24722
rect 18898 24670 18910 24722
rect 19618 24670 19630 24722
rect 19682 24670 19694 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 28802 24670 28814 24722
rect 28866 24670 28878 24722
rect 29250 24670 29262 24722
rect 29314 24670 29326 24722
rect 30706 24670 30718 24722
rect 30770 24670 30782 24722
rect 31490 24670 31502 24722
rect 31554 24670 31566 24722
rect 2830 24658 2882 24670
rect 6302 24658 6354 24670
rect 21310 24658 21362 24670
rect 32734 24658 32786 24670
rect 32958 24722 33010 24734
rect 39230 24722 39282 24734
rect 33282 24670 33294 24722
rect 33346 24670 33358 24722
rect 42018 24670 42030 24722
rect 42082 24670 42094 24722
rect 45826 24670 45838 24722
rect 45890 24670 45902 24722
rect 53890 24670 53902 24722
rect 53954 24670 53966 24722
rect 56130 24670 56142 24722
rect 56194 24670 56206 24722
rect 32958 24658 33010 24670
rect 39230 24658 39282 24670
rect 1150 24610 1202 24622
rect 4958 24610 5010 24622
rect 2146 24558 2158 24610
rect 2210 24558 2222 24610
rect 1150 24546 1202 24558
rect 4958 24546 5010 24558
rect 5406 24610 5458 24622
rect 5406 24546 5458 24558
rect 5518 24610 5570 24622
rect 5518 24546 5570 24558
rect 6078 24610 6130 24622
rect 6078 24546 6130 24558
rect 16606 24610 16658 24622
rect 16606 24546 16658 24558
rect 20638 24610 20690 24622
rect 20638 24546 20690 24558
rect 20862 24610 20914 24622
rect 27806 24610 27858 24622
rect 24434 24558 24446 24610
rect 24498 24558 24510 24610
rect 20862 24546 20914 24558
rect 27806 24546 27858 24558
rect 28478 24610 28530 24622
rect 28478 24546 28530 24558
rect 29934 24610 29986 24622
rect 38894 24610 38946 24622
rect 34402 24558 34414 24610
rect 34466 24558 34478 24610
rect 29934 24546 29986 24558
rect 38894 24546 38946 24558
rect 39006 24610 39058 24622
rect 39006 24546 39058 24558
rect 41694 24610 41746 24622
rect 47842 24558 47854 24610
rect 47906 24558 47918 24610
rect 50642 24558 50654 24610
rect 50706 24558 50718 24610
rect 52770 24558 52782 24610
rect 52834 24558 52846 24610
rect 53218 24558 53230 24610
rect 53282 24558 53294 24610
rect 54226 24558 54238 24610
rect 54290 24558 54302 24610
rect 56354 24558 56366 24610
rect 56418 24558 56430 24610
rect 41694 24546 41746 24558
rect 6526 24498 6578 24510
rect 15710 24498 15762 24510
rect 23326 24498 23378 24510
rect 32846 24498 32898 24510
rect 7858 24446 7870 24498
rect 7922 24446 7934 24498
rect 14578 24446 14590 24498
rect 14642 24446 14654 24498
rect 17602 24446 17614 24498
rect 17666 24446 17678 24498
rect 22194 24446 22206 24498
rect 22258 24446 22270 24498
rect 26674 24446 26686 24498
rect 26738 24446 26750 24498
rect 29474 24446 29486 24498
rect 29538 24446 29550 24498
rect 6526 24434 6578 24446
rect 15710 24434 15762 24446
rect 23326 24434 23378 24446
rect 32846 24434 32898 24446
rect 35646 24498 35698 24510
rect 38110 24498 38162 24510
rect 46510 24498 46562 24510
rect 49534 24498 49586 24510
rect 36978 24446 36990 24498
rect 37042 24446 37054 24498
rect 40114 24446 40126 24498
rect 40178 24446 40190 24498
rect 45378 24446 45390 24498
rect 45442 24446 45454 24498
rect 46834 24446 46846 24498
rect 46898 24446 46910 24498
rect 35646 24434 35698 24446
rect 38110 24434 38162 24446
rect 46510 24434 46562 24446
rect 49534 24434 49586 24446
rect 52110 24498 52162 24510
rect 52110 24434 52162 24446
rect 55470 24498 55522 24510
rect 55470 24434 55522 24446
rect 672 24330 56784 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 44466 24330
rect 44518 24278 44570 24330
rect 44622 24278 44674 24330
rect 44726 24278 56784 24330
rect 672 24244 56784 24278
rect 8990 24162 9042 24174
rect 3714 24110 3726 24162
rect 3778 24110 3790 24162
rect 6066 24110 6078 24162
rect 6130 24110 6142 24162
rect 8990 24098 9042 24110
rect 12910 24162 12962 24174
rect 12910 24098 12962 24110
rect 20862 24162 20914 24174
rect 20862 24098 20914 24110
rect 21646 24162 21698 24174
rect 32510 24162 32562 24174
rect 53678 24162 53730 24174
rect 22754 24110 22766 24162
rect 22818 24110 22830 24162
rect 30258 24110 30270 24162
rect 30322 24110 30334 24162
rect 33618 24110 33630 24162
rect 33682 24110 33694 24162
rect 41458 24110 41470 24162
rect 41522 24110 41534 24162
rect 52546 24110 52558 24162
rect 52610 24110 52622 24162
rect 21646 24098 21698 24110
rect 32510 24098 32562 24110
rect 53678 24098 53730 24110
rect 55918 24162 55970 24174
rect 55918 24098 55970 24110
rect 5070 24050 5122 24062
rect 16718 24050 16770 24062
rect 20750 24050 20802 24062
rect 9538 23998 9550 24050
rect 9602 23998 9614 24050
rect 9874 23998 9886 24050
rect 9938 23998 9950 24050
rect 11666 23998 11678 24050
rect 11730 23998 11742 24050
rect 14690 23998 14702 24050
rect 14754 23998 14766 24050
rect 17714 23998 17726 24050
rect 17778 23998 17790 24050
rect 5070 23986 5122 23998
rect 16718 23986 16770 23998
rect 20750 23986 20802 23998
rect 21422 24050 21474 24062
rect 21422 23986 21474 23998
rect 21758 24050 21810 24062
rect 26562 23998 26574 24050
rect 26626 23998 26638 24050
rect 34850 23998 34862 24050
rect 34914 23998 34926 24050
rect 37426 23998 37438 24050
rect 37490 23998 37502 24050
rect 43138 23998 43150 24050
rect 43202 23998 43214 24050
rect 45266 23998 45278 24050
rect 45330 23998 45342 24050
rect 48850 23998 48862 24050
rect 48914 23998 48926 24050
rect 54226 23998 54238 24050
rect 54290 23998 54302 24050
rect 54562 23998 54574 24050
rect 54626 23998 54638 24050
rect 56242 23998 56254 24050
rect 56306 23998 56318 24050
rect 21758 23986 21810 23998
rect 3054 23938 3106 23950
rect 6750 23938 6802 23950
rect 9326 23938 9378 23950
rect 18174 23938 18226 23950
rect 21310 23938 21362 23950
rect 23886 23938 23938 23950
rect 1698 23886 1710 23938
rect 1762 23886 1774 23938
rect 2594 23886 2606 23938
rect 2658 23886 2670 23938
rect 3826 23886 3838 23938
rect 3890 23886 3902 23938
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 5394 23886 5406 23938
rect 5458 23886 5470 23938
rect 5954 23886 5966 23938
rect 6018 23886 6030 23938
rect 7074 23886 7086 23938
rect 7138 23886 7150 23938
rect 8082 23886 8094 23938
rect 8146 23886 8158 23938
rect 11330 23886 11342 23938
rect 11394 23886 11406 23938
rect 14242 23886 14254 23938
rect 14306 23886 14318 23938
rect 17042 23886 17054 23938
rect 17106 23886 17118 23938
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 18834 23886 18846 23938
rect 18898 23886 18910 23938
rect 19730 23886 19742 23938
rect 19794 23886 19806 23938
rect 22194 23886 22206 23938
rect 22258 23886 22270 23938
rect 25890 23892 25902 23944
rect 25954 23892 25966 23944
rect 27022 23938 27074 23950
rect 35646 23938 35698 23950
rect 38110 23938 38162 23950
rect 54014 23938 54066 23950
rect 26338 23886 26350 23938
rect 26402 23886 26414 23938
rect 27682 23886 27694 23938
rect 27746 23886 27758 23938
rect 28690 23886 28702 23938
rect 28754 23886 28766 23938
rect 29698 23886 29710 23938
rect 29762 23886 29774 23938
rect 35074 23886 35086 23938
rect 35138 23886 35150 23938
rect 36754 23886 36766 23938
rect 36818 23886 36830 23938
rect 37202 23886 37214 23938
rect 37266 23886 37278 23938
rect 38434 23886 38446 23938
rect 38498 23886 38510 23938
rect 39554 23886 39566 23938
rect 39618 23886 39630 23938
rect 44930 23886 44942 23938
rect 44994 23886 45006 23938
rect 48066 23886 48078 23938
rect 48130 23886 48142 23938
rect 52994 23886 53006 23938
rect 53058 23886 53070 23938
rect 3054 23874 3106 23886
rect 6750 23874 6802 23886
rect 9326 23874 9378 23886
rect 18174 23874 18226 23886
rect 21310 23874 21362 23886
rect 23886 23874 23938 23886
rect 27022 23874 27074 23886
rect 35646 23874 35698 23886
rect 38110 23874 38162 23886
rect 54014 23874 54066 23886
rect 4734 23826 4786 23838
rect 25566 23826 25618 23838
rect 36430 23826 36482 23838
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 34066 23774 34078 23826
rect 34130 23774 34142 23826
rect 41906 23774 41918 23826
rect 41970 23774 41982 23826
rect 42690 23774 42702 23826
rect 42754 23774 42766 23826
rect 50978 23774 50990 23826
rect 51042 23774 51054 23826
rect 4734 23762 4786 23774
rect 25566 23762 25618 23774
rect 36430 23762 36482 23774
rect 15934 23714 15986 23726
rect 15934 23650 15986 23662
rect 31390 23714 31442 23726
rect 31390 23650 31442 23662
rect 35982 23714 36034 23726
rect 35982 23650 36034 23662
rect 40350 23714 40402 23726
rect 40350 23650 40402 23662
rect 44270 23714 44322 23726
rect 44270 23650 44322 23662
rect 46510 23714 46562 23726
rect 46510 23650 46562 23662
rect 51438 23714 51490 23726
rect 51438 23650 51490 23662
rect 672 23546 56784 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 43806 23546
rect 43858 23494 43910 23546
rect 43962 23494 44014 23546
rect 44066 23494 56784 23546
rect 672 23460 56784 23494
rect 2942 23378 2994 23390
rect 2942 23314 2994 23326
rect 6750 23378 6802 23390
rect 6750 23314 6802 23326
rect 19406 23378 19458 23390
rect 19406 23314 19458 23326
rect 51214 23378 51266 23390
rect 51214 23314 51266 23326
rect 54574 23378 54626 23390
rect 54574 23314 54626 23326
rect 4062 23266 4114 23278
rect 15374 23266 15426 23278
rect 35646 23266 35698 23278
rect 14466 23214 14478 23266
rect 14530 23214 14542 23266
rect 21522 23214 21534 23266
rect 21586 23214 21598 23266
rect 4062 23202 4114 23214
rect 15374 23202 15426 23214
rect 35646 23202 35698 23214
rect 36318 23266 36370 23278
rect 53790 23266 53842 23278
rect 49634 23214 49646 23266
rect 49698 23214 49710 23266
rect 52210 23214 52222 23266
rect 52274 23214 52286 23266
rect 36318 23202 36370 23214
rect 53790 23202 53842 23214
rect 55134 23266 55186 23278
rect 55134 23202 55186 23214
rect 8990 23154 9042 23166
rect 17278 23154 17330 23166
rect 23102 23154 23154 23166
rect 25006 23154 25058 23166
rect 30606 23154 30658 23166
rect 32622 23154 32674 23166
rect 35758 23154 35810 23166
rect 36990 23154 37042 23166
rect 1250 23102 1262 23154
rect 1314 23102 1326 23154
rect 5170 23102 5182 23154
rect 5234 23102 5246 23154
rect 7858 23102 7870 23154
rect 7922 23102 7934 23154
rect 8306 23102 8318 23154
rect 8370 23102 8382 23154
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 10658 23102 10670 23154
rect 10722 23102 10734 23154
rect 16258 23102 16270 23154
rect 16322 23102 16334 23154
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 18946 23102 18958 23154
rect 19010 23102 19022 23154
rect 23874 23102 23886 23154
rect 23938 23102 23950 23154
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 25666 23102 25678 23154
rect 25730 23102 25742 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 29026 23102 29038 23154
rect 29090 23102 29102 23154
rect 31154 23102 31166 23154
rect 31218 23102 31230 23154
rect 32050 23102 32062 23154
rect 32114 23102 32126 23154
rect 33394 23102 33406 23154
rect 33458 23102 33470 23154
rect 33842 23102 33854 23154
rect 33906 23102 33918 23154
rect 35186 23102 35198 23154
rect 35250 23102 35262 23154
rect 36642 23102 36654 23154
rect 36706 23102 36718 23154
rect 8990 23090 9042 23102
rect 17278 23090 17330 23102
rect 23102 23090 23154 23102
rect 25006 23090 25058 23102
rect 30606 23090 30658 23102
rect 32622 23090 32674 23102
rect 35758 23090 35810 23102
rect 36990 23090 37042 23102
rect 37214 23154 37266 23166
rect 37214 23090 37266 23102
rect 37662 23154 37714 23166
rect 39902 23154 39954 23166
rect 47070 23154 47122 23166
rect 54798 23154 54850 23166
rect 38658 23102 38670 23154
rect 38722 23102 38734 23154
rect 38994 23102 39006 23154
rect 39058 23102 39070 23154
rect 40226 23102 40238 23154
rect 40290 23102 40302 23154
rect 41346 23102 41358 23154
rect 41410 23102 41422 23154
rect 45714 23102 45726 23154
rect 45778 23102 45790 23154
rect 46498 23102 46510 23154
rect 46562 23102 46574 23154
rect 47842 23102 47854 23154
rect 47906 23102 47918 23154
rect 48290 23102 48302 23154
rect 48354 23102 48366 23154
rect 37662 23090 37714 23102
rect 39902 23090 39954 23102
rect 47070 23090 47122 23102
rect 54798 23090 54850 23102
rect 55022 23154 55074 23166
rect 55022 23090 55074 23102
rect 55246 23154 55298 23166
rect 55246 23090 55298 23102
rect 55918 23154 55970 23166
rect 55918 23090 55970 23102
rect 7534 23042 7586 23054
rect 15486 23042 15538 23054
rect 5506 22990 5518 23042
rect 5570 22990 5582 23042
rect 8530 22990 8542 23042
rect 8594 22990 8606 23042
rect 14130 22990 14142 23042
rect 14194 22990 14206 23042
rect 7534 22978 7586 22990
rect 15486 22978 15538 22990
rect 15822 23042 15874 23054
rect 23550 23042 23602 23054
rect 34302 23042 34354 23054
rect 21858 22990 21870 23042
rect 21922 22990 21934 23042
rect 29474 22990 29486 23042
rect 29538 22990 29550 23042
rect 15822 22978 15874 22990
rect 23550 22978 23602 22990
rect 34302 22978 34354 22990
rect 35534 23042 35586 23054
rect 35534 22978 35586 22990
rect 38222 23042 38274 23054
rect 38222 22978 38274 22990
rect 48750 23042 48802 23054
rect 52658 22990 52670 23042
rect 52722 22990 52734 23042
rect 56242 22990 56254 23042
rect 56306 22990 56318 23042
rect 48750 22978 48802 22990
rect 3726 22930 3778 22942
rect 1810 22878 1822 22930
rect 1874 22878 1886 22930
rect 3378 22878 3390 22930
rect 3442 22878 3454 22930
rect 3726 22866 3778 22878
rect 4174 22930 4226 22942
rect 4174 22866 4226 22878
rect 12910 22930 12962 22942
rect 12910 22866 12962 22878
rect 15262 22930 15314 22942
rect 19518 22930 19570 22942
rect 16818 22878 16830 22930
rect 16882 22878 16894 22930
rect 15262 22866 15314 22878
rect 19518 22866 19570 22878
rect 19630 22930 19682 22942
rect 36430 22930 36482 22942
rect 24546 22878 24558 22930
rect 24610 22878 24622 22930
rect 33282 22878 33294 22930
rect 33346 22878 33358 22930
rect 19630 22866 19682 22878
rect 36430 22866 36482 22878
rect 37102 22930 37154 22942
rect 39218 22878 39230 22930
rect 39282 22878 39294 22930
rect 47730 22878 47742 22930
rect 47794 22878 47806 22930
rect 50082 22878 50094 22930
rect 50146 22878 50158 22930
rect 37102 22866 37154 22878
rect 672 22762 56784 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 44466 22762
rect 44518 22710 44570 22762
rect 44622 22710 44674 22762
rect 44726 22710 56784 22762
rect 672 22676 56784 22710
rect 16046 22594 16098 22606
rect 10210 22542 10222 22594
rect 10274 22542 10286 22594
rect 16046 22530 16098 22542
rect 17278 22594 17330 22606
rect 17278 22530 17330 22542
rect 17390 22594 17442 22606
rect 27694 22594 27746 22606
rect 18386 22542 18398 22594
rect 18450 22542 18462 22594
rect 20962 22542 20974 22594
rect 21026 22542 21038 22594
rect 47182 22594 47234 22606
rect 17390 22530 17442 22542
rect 27694 22530 27746 22542
rect 41470 22538 41522 22550
rect 11790 22482 11842 22494
rect 13246 22482 13298 22494
rect 1362 22430 1374 22482
rect 1426 22430 1438 22482
rect 3714 22430 3726 22482
rect 3778 22430 3790 22482
rect 6962 22430 6974 22482
rect 7026 22430 7038 22482
rect 12786 22430 12798 22482
rect 12850 22430 12862 22482
rect 11790 22418 11842 22430
rect 13246 22418 13298 22430
rect 16158 22482 16210 22494
rect 16158 22418 16210 22430
rect 16942 22482 16994 22494
rect 16942 22418 16994 22430
rect 19966 22482 20018 22494
rect 28142 22482 28194 22494
rect 32846 22482 32898 22494
rect 40462 22482 40514 22494
rect 26562 22430 26574 22482
rect 26626 22430 26638 22482
rect 29138 22430 29150 22482
rect 29202 22430 29214 22482
rect 33842 22430 33854 22482
rect 33906 22430 33918 22482
rect 37090 22430 37102 22482
rect 37154 22430 37166 22482
rect 19966 22418 20018 22430
rect 28142 22418 28194 22430
rect 32846 22418 32898 22430
rect 40462 22418 40514 22430
rect 40798 22482 40850 22494
rect 40798 22418 40850 22430
rect 41022 22482 41074 22494
rect 49298 22542 49310 22594
rect 49362 22542 49374 22594
rect 51314 22542 51326 22594
rect 51378 22542 51390 22594
rect 54114 22542 54126 22594
rect 54178 22542 54190 22594
rect 56242 22542 56254 22594
rect 56306 22542 56318 22594
rect 47182 22530 47234 22542
rect 41470 22474 41522 22486
rect 41582 22482 41634 22494
rect 46062 22482 46114 22494
rect 48190 22482 48242 22494
rect 41022 22418 41074 22430
rect 43138 22430 43150 22482
rect 43202 22430 43214 22482
rect 46834 22430 46846 22482
rect 46898 22430 46910 22482
rect 47506 22430 47518 22482
rect 47570 22430 47582 22482
rect 41582 22418 41634 22430
rect 46062 22418 46114 22430
rect 48190 22418 48242 22430
rect 53006 22482 53058 22494
rect 53006 22418 53058 22430
rect 1934 22370 1986 22382
rect 4174 22370 4226 22382
rect 11342 22370 11394 22382
rect 17166 22370 17218 22382
rect 1138 22318 1150 22370
rect 1202 22318 1214 22370
rect 3042 22318 3054 22370
rect 3106 22318 3118 22370
rect 3602 22318 3614 22370
rect 3666 22318 3678 22370
rect 4946 22318 4958 22370
rect 5010 22318 5022 22370
rect 5842 22318 5854 22370
rect 5906 22318 5918 22370
rect 9762 22318 9774 22370
rect 9826 22318 9838 22370
rect 12114 22318 12126 22370
rect 12178 22318 12190 22370
rect 12562 22318 12574 22370
rect 12626 22318 12638 22370
rect 13794 22318 13806 22370
rect 13858 22318 13870 22370
rect 14802 22318 14814 22370
rect 14866 22318 14878 22370
rect 15810 22318 15822 22370
rect 15874 22318 15886 22370
rect 1934 22306 1986 22318
rect 4174 22306 4226 22318
rect 11342 22306 11394 22318
rect 17166 22306 17218 22318
rect 19518 22370 19570 22382
rect 21422 22370 21474 22382
rect 29822 22370 29874 22382
rect 34526 22370 34578 22382
rect 43822 22370 43874 22382
rect 45950 22370 46002 22382
rect 53118 22370 53170 22382
rect 20290 22318 20302 22370
rect 20354 22318 20366 22370
rect 20738 22318 20750 22370
rect 20802 22318 20814 22370
rect 21970 22318 21982 22370
rect 22034 22318 22046 22370
rect 22978 22318 22990 22370
rect 23042 22318 23054 22370
rect 26114 22318 26126 22370
rect 26178 22318 26190 22370
rect 28578 22318 28590 22370
rect 28642 22318 28654 22370
rect 28914 22318 28926 22370
rect 28978 22318 28990 22370
rect 30370 22318 30382 22370
rect 30434 22318 30446 22370
rect 31154 22318 31166 22370
rect 31218 22318 31230 22370
rect 33170 22318 33182 22370
rect 33234 22318 33246 22370
rect 33618 22318 33630 22370
rect 33682 22318 33694 22370
rect 34850 22318 34862 22370
rect 34914 22318 34926 22370
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 36530 22318 36542 22370
rect 36594 22318 36606 22370
rect 42578 22318 42590 22370
rect 42642 22318 42654 22370
rect 42914 22318 42926 22370
rect 42978 22318 42990 22370
rect 44146 22318 44158 22370
rect 44210 22318 44222 22370
rect 45154 22318 45166 22370
rect 45218 22318 45230 22370
rect 46610 22318 46622 22370
rect 46674 22318 46686 22370
rect 50754 22318 50766 22370
rect 50818 22318 50830 22370
rect 53554 22318 53566 22370
rect 53618 22318 53630 22370
rect 56018 22318 56030 22370
rect 56082 22318 56094 22370
rect 19518 22306 19570 22318
rect 21422 22306 21474 22318
rect 29822 22306 29874 22318
rect 34526 22306 34578 22318
rect 43822 22306 43874 22318
rect 45950 22306 46002 22318
rect 53118 22306 53170 22318
rect 2718 22258 2770 22270
rect 40910 22258 40962 22270
rect 6514 22206 6526 22258
rect 6578 22206 6590 22258
rect 17938 22206 17950 22258
rect 18002 22206 18014 22258
rect 2718 22194 2770 22206
rect 40910 22194 40962 22206
rect 42142 22258 42194 22270
rect 49746 22206 49758 22258
rect 49810 22206 49822 22258
rect 53666 22206 53678 22258
rect 53730 22206 53742 22258
rect 42142 22194 42194 22206
rect 2270 22146 2322 22158
rect 2270 22082 2322 22094
rect 8094 22146 8146 22158
rect 8094 22082 8146 22094
rect 38222 22146 38274 22158
rect 38222 22082 38274 22094
rect 40350 22146 40402 22158
rect 40350 22082 40402 22094
rect 41582 22146 41634 22158
rect 41582 22082 41634 22094
rect 46062 22146 46114 22158
rect 46062 22082 46114 22094
rect 52446 22146 52498 22158
rect 52446 22082 52498 22094
rect 53006 22146 53058 22158
rect 53006 22082 53058 22094
rect 55246 22146 55298 22158
rect 55246 22082 55298 22094
rect 672 21978 56784 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 43806 21978
rect 43858 21926 43910 21978
rect 43962 21926 44014 21978
rect 44066 21926 56784 21978
rect 672 21892 56784 21926
rect 12126 21810 12178 21822
rect 12126 21746 12178 21758
rect 19966 21810 20018 21822
rect 19966 21746 20018 21758
rect 22430 21810 22482 21822
rect 22430 21746 22482 21758
rect 27022 21810 27074 21822
rect 27022 21746 27074 21758
rect 32510 21810 32562 21822
rect 32510 21746 32562 21758
rect 34638 21810 34690 21822
rect 42926 21810 42978 21822
rect 40562 21758 40574 21810
rect 40626 21758 40638 21810
rect 34638 21746 34690 21758
rect 42926 21746 42978 21758
rect 47070 21810 47122 21822
rect 47070 21746 47122 21758
rect 4286 21698 4338 21710
rect 28478 21698 28530 21710
rect 2706 21646 2718 21698
rect 2770 21646 2782 21698
rect 10546 21646 10558 21698
rect 10610 21646 10622 21698
rect 4286 21634 4338 21646
rect 28478 21634 28530 21646
rect 32398 21698 32450 21710
rect 55694 21698 55746 21710
rect 41346 21646 41358 21698
rect 41410 21646 41422 21698
rect 32398 21634 32450 21646
rect 55694 21634 55746 21646
rect 8206 21586 8258 21598
rect 7186 21534 7198 21586
rect 7250 21534 7262 21586
rect 7522 21534 7534 21586
rect 7586 21534 7598 21586
rect 8206 21522 8258 21534
rect 8430 21586 8482 21598
rect 17278 21586 17330 21598
rect 24782 21586 24834 21598
rect 29934 21586 29986 21598
rect 38110 21586 38162 21598
rect 39566 21586 39618 21598
rect 8754 21534 8766 21586
rect 8818 21534 8830 21586
rect 9762 21534 9774 21586
rect 9826 21534 9838 21586
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 13682 21534 13694 21586
rect 13746 21534 13758 21586
rect 14802 21534 14814 21586
rect 14866 21534 14878 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 16818 21534 16830 21586
rect 16882 21534 16894 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 20738 21534 20750 21586
rect 20802 21534 20814 21586
rect 23090 21534 23102 21586
rect 23154 21534 23166 21586
rect 25442 21534 25454 21586
rect 25506 21534 25518 21586
rect 28802 21534 28814 21586
rect 28866 21534 28878 21586
rect 29250 21534 29262 21586
rect 29314 21534 29326 21586
rect 30706 21534 30718 21586
rect 30770 21534 30782 21586
rect 31602 21534 31614 21586
rect 31666 21534 31678 21586
rect 32946 21534 32958 21586
rect 33010 21534 33022 21586
rect 36418 21534 36430 21586
rect 36482 21534 36494 21586
rect 37314 21534 37326 21586
rect 37378 21534 37390 21586
rect 38658 21534 38670 21586
rect 38722 21534 38734 21586
rect 39218 21534 39230 21586
rect 39282 21534 39294 21586
rect 8430 21522 8482 21534
rect 17278 21522 17330 21534
rect 24782 21522 24834 21534
rect 29934 21522 29986 21534
rect 38110 21522 38162 21534
rect 39566 21522 39618 21534
rect 40014 21586 40066 21598
rect 51214 21586 51266 21598
rect 40562 21534 40574 21586
rect 40626 21534 40638 21586
rect 45378 21534 45390 21586
rect 45442 21534 45454 21586
rect 49186 21534 49198 21586
rect 49250 21534 49262 21586
rect 49970 21534 49982 21586
rect 50034 21534 50046 21586
rect 40014 21522 40066 21534
rect 51214 21522 51266 21534
rect 51550 21586 51602 21598
rect 51550 21522 51602 21534
rect 53006 21586 53058 21598
rect 55470 21586 55522 21598
rect 53442 21534 53454 21586
rect 53506 21534 53518 21586
rect 53006 21522 53058 21534
rect 55470 21522 55522 21534
rect 55918 21586 55970 21598
rect 55918 21522 55970 21534
rect 1374 21474 1426 21486
rect 6750 21474 6802 21486
rect 12798 21474 12850 21486
rect 14254 21474 14306 21486
rect 50766 21474 50818 21486
rect 1698 21422 1710 21474
rect 1762 21422 1774 21474
rect 7746 21422 7758 21474
rect 7810 21422 7822 21474
rect 10882 21422 10894 21474
rect 10946 21422 10958 21474
rect 13794 21422 13806 21474
rect 13858 21422 13870 21474
rect 16482 21422 16494 21474
rect 16546 21422 16558 21474
rect 21186 21422 21198 21474
rect 21250 21422 21262 21474
rect 23538 21422 23550 21474
rect 23602 21422 23614 21474
rect 33506 21422 33518 21474
rect 33570 21422 33582 21474
rect 40226 21422 40238 21474
rect 40290 21422 40302 21474
rect 48738 21422 48750 21474
rect 48802 21422 48814 21474
rect 1374 21410 1426 21422
rect 6750 21410 6802 21422
rect 12798 21410 12850 21422
rect 14254 21410 14306 21422
rect 50766 21410 50818 21422
rect 51326 21474 51378 21486
rect 53778 21422 53790 21474
rect 53842 21422 53854 21474
rect 51326 21410 51378 21422
rect 2046 21362 2098 21374
rect 5294 21362 5346 21374
rect 1026 21310 1038 21362
rect 1090 21310 1102 21362
rect 3154 21310 3166 21362
rect 3218 21310 3230 21362
rect 4946 21310 4958 21362
rect 5010 21310 5022 21362
rect 2046 21298 2098 21310
rect 5294 21298 5346 21310
rect 17614 21362 17666 21374
rect 40798 21362 40850 21374
rect 47630 21362 47682 21374
rect 52334 21362 52386 21374
rect 18834 21310 18846 21362
rect 18898 21310 18910 21362
rect 25890 21310 25902 21362
rect 25954 21310 25966 21362
rect 29474 21310 29486 21362
rect 29538 21310 29550 21362
rect 38546 21310 38558 21362
rect 38610 21310 38622 21362
rect 41794 21310 41806 21362
rect 41858 21310 41870 21362
rect 45938 21310 45950 21362
rect 46002 21310 46014 21362
rect 49746 21310 49758 21362
rect 49810 21310 49822 21362
rect 50418 21310 50430 21362
rect 50482 21310 50494 21362
rect 17614 21298 17666 21310
rect 40798 21298 40850 21310
rect 47630 21298 47682 21310
rect 52334 21298 52386 21310
rect 52446 21362 52498 21374
rect 52446 21298 52498 21310
rect 52558 21362 52610 21374
rect 52558 21298 52610 21310
rect 55022 21362 55074 21374
rect 55022 21298 55074 21310
rect 56030 21362 56082 21374
rect 56030 21298 56082 21310
rect 56142 21362 56194 21374
rect 56142 21298 56194 21310
rect 672 21194 56784 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 44466 21194
rect 44518 21142 44570 21194
rect 44622 21142 44674 21194
rect 44726 21142 56784 21194
rect 672 21108 56784 21142
rect 2830 21026 2882 21038
rect 13806 21026 13858 21038
rect 21646 21026 21698 21038
rect 29934 21026 29986 21038
rect 37774 21026 37826 21038
rect 1698 20974 1710 21026
rect 1762 20974 1774 21026
rect 4274 20974 4286 21026
rect 4338 20974 4350 21026
rect 20514 20974 20526 21026
rect 20578 20974 20590 21026
rect 22754 20974 22766 21026
rect 22818 20974 22830 21026
rect 33394 20974 33406 21026
rect 33458 20974 33470 21026
rect 36642 20974 36654 21026
rect 36706 20974 36718 21026
rect 2830 20962 2882 20974
rect 13806 20962 13858 20974
rect 21646 20962 21698 20974
rect 29934 20962 29986 20974
rect 37774 20962 37826 20974
rect 41246 21026 41298 21038
rect 41246 20962 41298 20974
rect 41358 21026 41410 21038
rect 41358 20962 41410 20974
rect 41470 21026 41522 21038
rect 47518 21026 47570 21038
rect 55246 21026 55298 21038
rect 44146 20974 44158 21026
rect 44210 20974 44222 21026
rect 47170 20974 47182 21026
rect 47234 20974 47246 21026
rect 49186 20974 49198 21026
rect 49250 20974 49262 21026
rect 50194 20974 50206 21026
rect 50258 20974 50270 21026
rect 54114 20974 54126 21026
rect 54178 20974 54190 21026
rect 41470 20962 41522 20974
rect 47518 20962 47570 20974
rect 55246 20962 55298 20974
rect 56030 21026 56082 21038
rect 56354 20974 56366 21026
rect 56418 20974 56430 21026
rect 56030 20962 56082 20974
rect 3278 20914 3330 20926
rect 3278 20850 3330 20862
rect 4734 20914 4786 20926
rect 10670 20914 10722 20926
rect 9426 20862 9438 20914
rect 9490 20862 9502 20914
rect 4734 20850 4786 20862
rect 10670 20850 10722 20862
rect 11342 20914 11394 20926
rect 11342 20850 11394 20862
rect 11566 20914 11618 20926
rect 16046 20914 16098 20926
rect 12674 20862 12686 20914
rect 12738 20862 12750 20914
rect 14802 20862 14814 20914
rect 14866 20862 14878 20914
rect 11566 20850 11618 20862
rect 16046 20850 16098 20862
rect 17166 20914 17218 20926
rect 39118 20914 39170 20926
rect 18162 20862 18174 20914
rect 18226 20862 18238 20914
rect 25554 20862 25566 20914
rect 25618 20862 25630 20914
rect 28690 20862 28702 20914
rect 28754 20862 28766 20914
rect 30594 20862 30606 20914
rect 30658 20862 30670 20914
rect 17166 20850 17218 20862
rect 39118 20850 39170 20862
rect 39230 20914 39282 20926
rect 39230 20850 39282 20862
rect 40350 20914 40402 20926
rect 40350 20850 40402 20862
rect 40686 20914 40738 20926
rect 40686 20850 40738 20862
rect 43038 20914 43090 20926
rect 46846 20914 46898 20926
rect 46498 20862 46510 20914
rect 46562 20862 46574 20914
rect 43038 20850 43090 20862
rect 46846 20850 46898 20862
rect 52334 20914 52386 20926
rect 52334 20850 52386 20862
rect 52782 20914 52834 20926
rect 52782 20850 52834 20862
rect 11118 20802 11170 20814
rect 23886 20802 23938 20814
rect 31278 20802 31330 20814
rect 1250 20750 1262 20802
rect 1314 20750 1326 20802
rect 3602 20750 3614 20802
rect 3666 20750 3678 20802
rect 4162 20750 4174 20802
rect 4226 20750 4238 20802
rect 5506 20750 5518 20802
rect 5570 20750 5582 20802
rect 6290 20750 6302 20802
rect 6354 20750 6366 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 17826 20750 17838 20802
rect 17890 20750 17902 20802
rect 19954 20750 19966 20802
rect 20018 20750 20030 20802
rect 24882 20750 24894 20802
rect 24946 20750 24958 20802
rect 25330 20750 25342 20802
rect 25394 20750 25406 20802
rect 26114 20750 26126 20802
rect 26178 20750 26190 20802
rect 26562 20750 26574 20802
rect 26626 20750 26638 20802
rect 27570 20750 27582 20802
rect 27634 20750 27646 20802
rect 30482 20750 30494 20802
rect 30546 20750 30558 20802
rect 11118 20738 11170 20750
rect 23886 20738 23938 20750
rect 31278 20738 31330 20750
rect 32398 20802 32450 20814
rect 33854 20802 33906 20814
rect 38894 20802 38946 20814
rect 40574 20802 40626 20814
rect 32722 20750 32734 20802
rect 32786 20750 32798 20802
rect 33282 20750 33294 20802
rect 33346 20750 33358 20802
rect 34402 20750 34414 20802
rect 34466 20750 34478 20802
rect 35410 20750 35422 20802
rect 35474 20750 35486 20802
rect 39666 20750 39678 20802
rect 39730 20750 39742 20802
rect 32398 20738 32450 20750
rect 33854 20738 33906 20750
rect 38894 20738 38946 20750
rect 40574 20738 40626 20750
rect 40798 20802 40850 20814
rect 42366 20802 42418 20814
rect 41570 20750 41582 20802
rect 41634 20750 41646 20802
rect 40798 20738 40850 20750
rect 42366 20738 42418 20750
rect 42814 20802 42866 20814
rect 48862 20802 48914 20814
rect 43586 20750 43598 20802
rect 43650 20750 43662 20802
rect 52546 20750 52558 20802
rect 52610 20750 52622 20802
rect 53666 20750 53678 20802
rect 53730 20750 53742 20802
rect 42814 20738 42866 20750
rect 48862 20738 48914 20750
rect 11230 20690 11282 20702
rect 17278 20690 17330 20702
rect 24558 20690 24610 20702
rect 42590 20690 42642 20702
rect 9090 20638 9102 20690
rect 9154 20638 9166 20690
rect 14466 20638 14478 20690
rect 14530 20638 14542 20690
rect 22306 20638 22318 20690
rect 22370 20638 22382 20690
rect 28354 20638 28366 20690
rect 28418 20638 28430 20690
rect 36194 20638 36206 20690
rect 36258 20638 36270 20690
rect 39218 20638 39230 20690
rect 39282 20638 39294 20690
rect 11230 20626 11282 20638
rect 17278 20626 17330 20638
rect 24558 20626 24610 20638
rect 42590 20626 42642 20638
rect 48638 20690 48690 20702
rect 49746 20638 49758 20690
rect 49810 20638 49822 20690
rect 52882 20638 52894 20690
rect 52946 20638 52958 20690
rect 48638 20626 48690 20638
rect 19406 20578 19458 20590
rect 19406 20514 19458 20526
rect 31614 20578 31666 20590
rect 31614 20514 31666 20526
rect 41918 20578 41970 20590
rect 41918 20514 41970 20526
rect 42142 20578 42194 20590
rect 42142 20514 42194 20526
rect 45278 20578 45330 20590
rect 45278 20514 45330 20526
rect 51326 20578 51378 20590
rect 51326 20514 51378 20526
rect 51886 20578 51938 20590
rect 51886 20514 51938 20526
rect 51998 20578 52050 20590
rect 51998 20514 52050 20526
rect 672 20410 56784 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 43806 20410
rect 43858 20358 43910 20410
rect 43962 20358 44014 20410
rect 44066 20358 56784 20410
rect 672 20324 56784 20358
rect 32622 20242 32674 20254
rect 32622 20178 32674 20190
rect 33182 20242 33234 20254
rect 33182 20178 33234 20190
rect 38670 20242 38722 20254
rect 38670 20178 38722 20190
rect 51326 20242 51378 20254
rect 51326 20178 51378 20190
rect 52894 20242 52946 20254
rect 52894 20178 52946 20190
rect 4958 20130 5010 20142
rect 18510 20130 18562 20142
rect 22654 20130 22706 20142
rect 41470 20130 41522 20142
rect 2706 20078 2718 20130
rect 2770 20078 2782 20130
rect 11554 20078 11566 20130
rect 11618 20078 11630 20130
rect 21074 20078 21086 20130
rect 21138 20078 21150 20130
rect 34738 20078 34750 20130
rect 34802 20078 34814 20130
rect 4958 20066 5010 20078
rect 18510 20066 18562 20078
rect 22654 20066 22706 20078
rect 41470 20066 41522 20078
rect 53230 20130 53282 20142
rect 53230 20066 53282 20078
rect 3614 20018 3666 20030
rect 14814 20018 14866 20030
rect 16830 20018 16882 20030
rect 24782 20018 24834 20030
rect 41358 20018 41410 20030
rect 5394 19966 5406 20018
rect 5458 19966 5470 20018
rect 5730 19966 5742 20018
rect 5794 19966 5806 20018
rect 6514 19966 6526 20018
rect 6578 19966 6590 20018
rect 7186 19966 7198 20018
rect 7250 19966 7262 20018
rect 7970 19966 7982 20018
rect 8034 19966 8046 20018
rect 8754 19966 8766 20018
rect 8818 19966 8830 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 15362 19966 15374 20018
rect 15426 19966 15438 20018
rect 16482 19966 16494 20018
rect 16546 19966 16558 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 18050 19966 18062 20018
rect 18114 19966 18126 20018
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 23986 19966 23998 20018
rect 24050 19966 24062 20018
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 26226 19966 26238 20018
rect 26290 19966 26302 20018
rect 28690 19966 28702 20018
rect 28754 19966 28766 20018
rect 31042 19966 31054 20018
rect 31106 19966 31118 20018
rect 37090 19966 37102 20018
rect 37154 19966 37166 20018
rect 39330 19966 39342 20018
rect 39394 19966 39406 20018
rect 3614 19954 3666 19966
rect 14814 19954 14866 19966
rect 16830 19954 16882 19966
rect 24782 19954 24834 19966
rect 41358 19954 41410 19966
rect 42702 20018 42754 20030
rect 46734 20018 46786 20030
rect 45378 19966 45390 20018
rect 45442 19966 45454 20018
rect 45826 19966 45838 20018
rect 45890 19966 45902 20018
rect 47058 19966 47070 20018
rect 47122 19966 47134 20018
rect 48066 19966 48078 20018
rect 48130 19966 48142 20018
rect 48738 19966 48750 20018
rect 48802 19966 48814 20018
rect 49746 19966 49758 20018
rect 49810 19966 49822 20018
rect 53890 19966 53902 20018
rect 53954 19966 53966 20018
rect 42702 19954 42754 19966
rect 46734 19954 46786 19966
rect 10782 19906 10834 19918
rect 2370 19854 2382 19906
rect 2434 19854 2446 19906
rect 3266 19854 3278 19906
rect 3330 19854 3342 19906
rect 3938 19854 3950 19906
rect 4002 19854 4014 19906
rect 9202 19854 9214 19906
rect 9266 19854 9278 19906
rect 10782 19842 10834 19854
rect 11118 19906 11170 19918
rect 11790 19906 11842 19918
rect 11330 19854 11342 19906
rect 11394 19854 11406 19906
rect 11118 19842 11170 19854
rect 11790 19842 11842 19854
rect 12126 19906 12178 19918
rect 23102 19906 23154 19918
rect 30270 19906 30322 19918
rect 45054 19906 45106 19918
rect 13570 19854 13582 19906
rect 13634 19854 13646 19906
rect 17490 19854 17502 19906
rect 17554 19854 17566 19906
rect 21410 19854 21422 19906
rect 21474 19854 21486 19906
rect 29138 19854 29150 19906
rect 29202 19854 29214 19906
rect 37538 19854 37550 19906
rect 37602 19854 37614 19906
rect 42130 19854 42142 19906
rect 42194 19854 42206 19906
rect 42354 19854 42366 19906
rect 42418 19854 42430 19906
rect 48962 19854 48974 19906
rect 49026 19854 49038 19906
rect 50082 19854 50094 19906
rect 50146 19854 50158 19906
rect 52098 19854 52110 19906
rect 52162 19854 52174 19906
rect 52658 19854 52670 19906
rect 52722 19854 52734 19906
rect 56242 19854 56254 19906
rect 56306 19854 56318 19906
rect 12126 19842 12178 19854
rect 23102 19842 23154 19854
rect 30270 19842 30322 19854
rect 45054 19842 45106 19854
rect 1150 19794 1202 19806
rect 1150 19730 1202 19742
rect 4286 19794 4338 19806
rect 10334 19794 10386 19806
rect 5954 19742 5966 19794
rect 6018 19742 6030 19794
rect 4286 19730 4338 19742
rect 10334 19730 10386 19742
rect 11006 19794 11058 19806
rect 11006 19730 11058 19742
rect 12014 19794 12066 19806
rect 40910 19794 40962 19806
rect 24098 19742 24110 19794
rect 24162 19742 24174 19794
rect 31490 19742 31502 19794
rect 31554 19742 31566 19794
rect 34290 19742 34302 19794
rect 34354 19742 34366 19794
rect 39778 19742 39790 19794
rect 39842 19742 39854 19794
rect 12014 19730 12066 19742
rect 40910 19730 40962 19742
rect 43038 19794 43090 19806
rect 55470 19794 55522 19806
rect 46050 19742 46062 19794
rect 46114 19742 46126 19794
rect 54338 19742 54350 19794
rect 54402 19742 54414 19794
rect 43038 19730 43090 19742
rect 55470 19730 55522 19742
rect 55918 19794 55970 19806
rect 55918 19730 55970 19742
rect 672 19626 56784 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 44466 19626
rect 44518 19574 44570 19626
rect 44622 19574 44674 19626
rect 44726 19574 56784 19626
rect 672 19540 56784 19574
rect 9214 19458 9266 19470
rect 9214 19394 9266 19406
rect 9326 19458 9378 19470
rect 9326 19394 9378 19406
rect 13358 19458 13410 19470
rect 16046 19458 16098 19470
rect 39566 19458 39618 19470
rect 14914 19406 14926 19458
rect 14978 19406 14990 19458
rect 20290 19406 20302 19458
rect 20354 19406 20366 19458
rect 25330 19406 25342 19458
rect 25394 19406 25406 19458
rect 27906 19406 27918 19458
rect 27970 19406 27982 19458
rect 33058 19406 33070 19458
rect 33122 19406 33134 19458
rect 37538 19406 37550 19458
rect 37602 19406 37614 19458
rect 13358 19394 13410 19406
rect 16046 19394 16098 19406
rect 39566 19394 39618 19406
rect 42142 19458 42194 19470
rect 42142 19394 42194 19406
rect 42814 19458 42866 19470
rect 42814 19394 42866 19406
rect 48414 19458 48466 19470
rect 54126 19458 54178 19470
rect 49186 19406 49198 19458
rect 49250 19406 49262 19458
rect 52434 19406 52446 19458
rect 52498 19406 52510 19458
rect 48414 19394 48466 19406
rect 54126 19394 54178 19406
rect 55022 19458 55074 19470
rect 55022 19394 55074 19406
rect 56030 19458 56082 19470
rect 56354 19406 56366 19458
rect 56418 19406 56430 19458
rect 56030 19394 56082 19406
rect 1486 19346 1538 19358
rect 5070 19346 5122 19358
rect 9774 19346 9826 19358
rect 13470 19346 13522 19358
rect 20750 19346 20802 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 6066 19294 6078 19346
rect 6130 19294 6142 19346
rect 10770 19294 10782 19346
rect 10834 19294 10846 19346
rect 18050 19294 18062 19346
rect 18114 19294 18126 19346
rect 1486 19282 1538 19294
rect 5070 19282 5122 19294
rect 9774 19282 9826 19294
rect 13470 19282 13522 19294
rect 20750 19282 20802 19294
rect 26910 19346 26962 19358
rect 26910 19282 26962 19294
rect 30718 19346 30770 19358
rect 30718 19282 30770 19294
rect 30830 19346 30882 19358
rect 30830 19282 30882 19294
rect 31054 19346 31106 19358
rect 44270 19346 44322 19358
rect 53566 19346 53618 19358
rect 35186 19294 35198 19346
rect 35250 19294 35262 19346
rect 41010 19294 41022 19346
rect 41074 19294 41086 19346
rect 45266 19294 45278 19346
rect 45330 19294 45342 19346
rect 48066 19294 48078 19346
rect 48130 19294 48142 19346
rect 50194 19294 50206 19346
rect 50258 19294 50270 19346
rect 31054 19282 31106 19294
rect 44270 19282 44322 19294
rect 53566 19282 53618 19294
rect 54238 19346 54290 19358
rect 54238 19282 54290 19294
rect 55246 19346 55298 19358
rect 55246 19282 55298 19294
rect 3166 19234 3218 19246
rect 6526 19234 6578 19246
rect 9438 19234 9490 19246
rect 11230 19234 11282 19246
rect 16830 19234 16882 19246
rect 26462 19234 26514 19246
rect 28366 19234 28418 19246
rect 31166 19234 31218 19246
rect 1922 19182 1934 19234
rect 1986 19182 1998 19234
rect 2370 19182 2382 19234
rect 2434 19182 2446 19234
rect 3602 19182 3614 19234
rect 3666 19182 3678 19234
rect 4610 19182 4622 19234
rect 4674 19182 4686 19234
rect 5394 19182 5406 19234
rect 5458 19182 5470 19234
rect 5842 19182 5854 19234
rect 5906 19182 5918 19234
rect 7074 19182 7086 19234
rect 7138 19182 7150 19234
rect 8194 19182 8206 19234
rect 8258 19182 8270 19234
rect 8866 19182 8878 19234
rect 8930 19182 8942 19234
rect 10210 19182 10222 19234
rect 10274 19182 10286 19234
rect 3166 19170 3218 19182
rect 6526 19170 6578 19182
rect 9438 19170 9490 19182
rect 10546 19170 10558 19222
rect 10610 19170 10622 19222
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 12002 19182 12014 19234
rect 12066 19182 12078 19234
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 18386 19182 18398 19234
rect 18450 19182 18462 19234
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 21298 19182 21310 19234
rect 21362 19182 21374 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22306 19182 22318 19234
rect 22370 19182 22382 19234
rect 27234 19182 27246 19234
rect 27298 19182 27310 19234
rect 27682 19182 27694 19234
rect 27746 19182 27758 19234
rect 28914 19182 28926 19234
rect 28978 19182 28990 19234
rect 29922 19182 29934 19234
rect 29986 19182 29998 19234
rect 11230 19170 11282 19182
rect 16830 19170 16882 19182
rect 26462 19170 26514 19182
rect 28366 19170 28418 19182
rect 31166 19170 31218 19182
rect 31614 19234 31666 19246
rect 31614 19170 31666 19182
rect 31838 19234 31890 19246
rect 42590 19234 42642 19246
rect 54014 19234 54066 19246
rect 55358 19234 55410 19246
rect 36978 19182 36990 19234
rect 37042 19182 37054 19234
rect 43026 19182 43038 19234
rect 43090 19182 43102 19234
rect 43250 19182 43262 19234
rect 43314 19182 43326 19234
rect 44594 19182 44606 19234
rect 44658 19182 44670 19234
rect 45154 19182 45166 19234
rect 45218 19182 45230 19234
rect 45826 19182 45838 19234
rect 45890 19182 45902 19234
rect 46386 19182 46398 19234
rect 46450 19182 46462 19234
rect 47394 19182 47406 19234
rect 47458 19182 47470 19234
rect 48962 19182 48974 19234
rect 49026 19182 49038 19234
rect 51874 19182 51886 19234
rect 51938 19182 51950 19234
rect 54450 19182 54462 19234
rect 54514 19182 54526 19234
rect 54674 19182 54686 19234
rect 54738 19182 54750 19234
rect 31838 19170 31890 19182
rect 42590 19170 42642 19182
rect 54014 19170 54066 19182
rect 55358 19170 55410 19182
rect 19294 19122 19346 19134
rect 31726 19122 31778 19134
rect 24882 19070 24894 19122
rect 24946 19070 24958 19122
rect 32610 19070 32622 19122
rect 32674 19070 32686 19122
rect 34850 19070 34862 19122
rect 34914 19070 34926 19122
rect 40562 19070 40574 19122
rect 40626 19070 40638 19122
rect 42914 19070 42926 19122
rect 42978 19070 42990 19122
rect 49746 19070 49758 19122
rect 49810 19070 49822 19122
rect 19294 19058 19346 19070
rect 31726 19058 31778 19070
rect 34190 19010 34242 19022
rect 34190 18946 34242 18958
rect 36430 19010 36482 19022
rect 36430 18946 36482 18958
rect 38670 19010 38722 19022
rect 38670 18946 38722 18958
rect 39342 19010 39394 19022
rect 39342 18946 39394 18958
rect 39678 19010 39730 19022
rect 39678 18946 39730 18958
rect 51326 19010 51378 19022
rect 51326 18946 51378 18958
rect 672 18842 56784 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 43806 18842
rect 43858 18790 43910 18842
rect 43962 18790 44014 18842
rect 44066 18790 56784 18842
rect 672 18756 56784 18790
rect 24670 18674 24722 18686
rect 24670 18610 24722 18622
rect 27806 18674 27858 18686
rect 43262 18674 43314 18686
rect 40562 18622 40574 18674
rect 40626 18622 40638 18674
rect 27806 18610 27858 18622
rect 43262 18610 43314 18622
rect 44270 18674 44322 18686
rect 44270 18610 44322 18622
rect 53006 18674 53058 18686
rect 53006 18610 53058 18622
rect 41022 18562 41074 18574
rect 51214 18562 51266 18574
rect 20850 18510 20862 18562
rect 20914 18510 20926 18562
rect 23090 18510 23102 18562
rect 23154 18510 23166 18562
rect 28690 18510 28702 18562
rect 28754 18510 28766 18562
rect 34290 18510 34302 18562
rect 34354 18510 34366 18562
rect 45826 18510 45838 18562
rect 45890 18510 45902 18562
rect 49074 18510 49086 18562
rect 49138 18510 49150 18562
rect 52098 18510 52110 18562
rect 52162 18510 52174 18562
rect 41022 18498 41074 18510
rect 51214 18498 51266 18510
rect 2046 18450 2098 18462
rect 4286 18450 4338 18462
rect 6526 18450 6578 18462
rect 10670 18450 10722 18462
rect 14590 18450 14642 18462
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 5394 18398 5406 18450
rect 5458 18398 5470 18450
rect 5842 18398 5854 18450
rect 5906 18398 5918 18450
rect 7298 18398 7310 18450
rect 7362 18398 7374 18450
rect 8194 18398 8206 18450
rect 8258 18398 8270 18450
rect 9314 18398 9326 18450
rect 9378 18398 9390 18450
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 10994 18398 11006 18450
rect 11058 18398 11070 18450
rect 12114 18398 12126 18450
rect 12178 18398 12190 18450
rect 13010 18398 13022 18450
rect 13074 18398 13086 18450
rect 2046 18386 2098 18398
rect 4286 18386 4338 18398
rect 6526 18386 6578 18398
rect 10670 18386 10722 18398
rect 14590 18386 14642 18398
rect 15038 18450 15090 18462
rect 16718 18450 16770 18462
rect 22430 18450 22482 18462
rect 30270 18450 30322 18462
rect 32510 18450 32562 18462
rect 33966 18450 34018 18462
rect 35086 18450 35138 18462
rect 37998 18450 38050 18462
rect 49646 18450 49698 18462
rect 51326 18450 51378 18462
rect 52894 18450 52946 18462
rect 56254 18450 56306 18462
rect 15474 18398 15486 18450
rect 15538 18398 15550 18450
rect 15810 18398 15822 18450
rect 15874 18398 15886 18450
rect 17154 18398 17166 18450
rect 17218 18398 17230 18450
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 26226 18398 26238 18450
rect 26290 18398 26302 18450
rect 30818 18398 30830 18450
rect 30882 18398 30894 18450
rect 31714 18398 31726 18450
rect 31778 18398 31790 18450
rect 33058 18398 33070 18450
rect 33122 18398 33134 18450
rect 33506 18398 33518 18450
rect 33570 18398 33582 18450
rect 34402 18398 34414 18450
rect 34466 18398 34478 18450
rect 34626 18398 34638 18450
rect 34690 18398 34702 18450
rect 36642 18398 36654 18450
rect 36706 18398 36718 18450
rect 37090 18398 37102 18450
rect 37154 18398 37166 18450
rect 38546 18398 38558 18450
rect 38610 18398 38622 18450
rect 39330 18398 39342 18450
rect 39394 18398 39406 18450
rect 40562 18398 40574 18450
rect 40626 18398 40638 18450
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 41570 18398 41582 18450
rect 41634 18398 41646 18450
rect 45938 18398 45950 18450
rect 46002 18398 46014 18450
rect 46946 18398 46958 18450
rect 47010 18398 47022 18450
rect 50306 18398 50318 18450
rect 50370 18398 50382 18450
rect 51986 18398 51998 18450
rect 52050 18398 52062 18450
rect 54114 18398 54126 18450
rect 54178 18398 54190 18450
rect 15038 18386 15090 18398
rect 16718 18386 16770 18398
rect 22430 18386 22482 18398
rect 30270 18386 30322 18398
rect 32510 18386 32562 18398
rect 33966 18386 34018 18398
rect 35086 18386 35138 18398
rect 37998 18386 38050 18398
rect 49646 18386 49698 18398
rect 51326 18386 51378 18398
rect 52894 18386 52946 18398
rect 56254 18386 56306 18398
rect 5070 18338 5122 18350
rect 8990 18338 9042 18350
rect 34862 18338 34914 18350
rect 1026 18286 1038 18338
rect 1090 18286 1102 18338
rect 3154 18286 3166 18338
rect 3218 18286 3230 18338
rect 6066 18286 6078 18338
rect 6130 18286 6142 18338
rect 9986 18286 9998 18338
rect 10050 18286 10062 18338
rect 13346 18286 13358 18338
rect 13410 18286 13422 18338
rect 16034 18286 16046 18338
rect 16098 18286 16110 18338
rect 26674 18286 26686 18338
rect 26738 18286 26750 18338
rect 29026 18286 29038 18338
rect 29090 18286 29102 18338
rect 5070 18274 5122 18286
rect 8990 18274 9042 18286
rect 34862 18274 34914 18286
rect 35422 18338 35474 18350
rect 35422 18274 35474 18286
rect 35534 18338 35586 18350
rect 35534 18274 35586 18286
rect 36318 18338 36370 18350
rect 41134 18338 41186 18350
rect 49982 18338 50034 18350
rect 37314 18286 37326 18338
rect 37378 18286 37390 18338
rect 46722 18286 46734 18338
rect 46786 18286 46798 18338
rect 48738 18286 48750 18338
rect 48802 18286 48814 18338
rect 36318 18274 36370 18286
rect 41134 18274 41186 18286
rect 49982 18274 50034 18286
rect 50878 18338 50930 18350
rect 52558 18338 52610 18350
rect 52322 18286 52334 18338
rect 52386 18286 52398 18338
rect 50878 18274 50930 18286
rect 52558 18274 52610 18286
rect 56366 18338 56418 18350
rect 56366 18274 56418 18286
rect 1374 18226 1426 18238
rect 47518 18226 47570 18238
rect 1698 18174 1710 18226
rect 1762 18174 1774 18226
rect 21298 18174 21310 18226
rect 21362 18174 21374 18226
rect 23538 18174 23550 18226
rect 23602 18174 23614 18226
rect 32946 18174 32958 18226
rect 33010 18174 33022 18226
rect 42130 18174 42142 18226
rect 42194 18174 42206 18226
rect 45378 18174 45390 18226
rect 45442 18174 45454 18226
rect 1374 18162 1426 18174
rect 47518 18162 47570 18174
rect 49758 18226 49810 18238
rect 49758 18162 49810 18174
rect 49870 18226 49922 18238
rect 49870 18162 49922 18174
rect 51102 18226 51154 18238
rect 53678 18226 53730 18238
rect 55806 18226 55858 18238
rect 53330 18174 53342 18226
rect 53394 18174 53406 18226
rect 54674 18174 54686 18226
rect 54738 18174 54750 18226
rect 51102 18162 51154 18174
rect 53678 18162 53730 18174
rect 55806 18162 55858 18174
rect 672 18058 56784 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 44466 18058
rect 44518 18006 44570 18058
rect 44622 18006 44674 18058
rect 44726 18006 56784 18058
rect 672 17972 56784 18006
rect 11230 17890 11282 17902
rect 3378 17838 3390 17890
rect 3442 17838 3454 17890
rect 5730 17838 5742 17890
rect 5794 17838 5806 17890
rect 11230 17826 11282 17838
rect 11454 17890 11506 17902
rect 31726 17890 31778 17902
rect 34974 17890 35026 17902
rect 12674 17838 12686 17890
rect 12738 17838 12750 17890
rect 14914 17838 14926 17890
rect 14978 17838 14990 17890
rect 20178 17838 20190 17890
rect 20242 17838 20254 17890
rect 33058 17838 33070 17890
rect 33122 17838 33134 17890
rect 11454 17826 11506 17838
rect 31726 17826 31778 17838
rect 34974 17826 35026 17838
rect 35086 17890 35138 17902
rect 43710 17890 43762 17902
rect 37314 17838 37326 17890
rect 37378 17838 37390 17890
rect 35086 17826 35138 17838
rect 43710 17826 43762 17838
rect 43934 17890 43986 17902
rect 43934 17826 43986 17838
rect 46622 17890 46674 17902
rect 46622 17826 46674 17838
rect 47182 17890 47234 17902
rect 53678 17890 53730 17902
rect 51986 17838 51998 17890
rect 52050 17838 52062 17890
rect 56354 17838 56366 17890
rect 56418 17838 56430 17890
rect 47182 17826 47234 17838
rect 53678 17826 53730 17838
rect 6190 17778 6242 17790
rect 16942 17778 16994 17790
rect 9538 17726 9550 17778
rect 9602 17726 9614 17778
rect 6190 17714 6242 17726
rect 16942 17714 16994 17726
rect 17054 17778 17106 17790
rect 36318 17778 36370 17790
rect 47070 17778 47122 17790
rect 17154 17726 17166 17778
rect 17218 17726 17230 17778
rect 25890 17726 25902 17778
rect 25954 17726 25966 17778
rect 29026 17726 29038 17778
rect 29090 17726 29102 17778
rect 41234 17726 41246 17778
rect 41298 17726 41310 17778
rect 45490 17726 45502 17778
rect 45554 17726 45566 17778
rect 17054 17714 17106 17726
rect 36318 17714 36370 17726
rect 47070 17714 47122 17726
rect 54910 17778 54962 17790
rect 54910 17714 54962 17726
rect 2942 17666 2994 17678
rect 11118 17666 11170 17678
rect 16046 17666 16098 17678
rect 1362 17614 1374 17666
rect 1426 17614 1438 17666
rect 2146 17614 2158 17666
rect 2210 17614 2222 17666
rect 3602 17614 3614 17666
rect 3666 17614 3678 17666
rect 3938 17614 3950 17666
rect 4002 17614 4014 17666
rect 5058 17614 5070 17666
rect 5122 17614 5134 17666
rect 5506 17614 5518 17666
rect 5570 17614 5582 17666
rect 6962 17614 6974 17666
rect 7026 17614 7038 17666
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 9090 17614 9102 17666
rect 9154 17614 9166 17666
rect 12226 17614 12238 17666
rect 12290 17614 12302 17666
rect 14466 17614 14478 17666
rect 14530 17614 14542 17666
rect 2942 17602 2994 17614
rect 11118 17602 11170 17614
rect 16046 17602 16098 17614
rect 16718 17666 16770 17678
rect 19518 17666 19570 17678
rect 29710 17666 29762 17678
rect 31614 17666 31666 17678
rect 18050 17614 18062 17666
rect 18114 17614 18126 17666
rect 18946 17614 18958 17666
rect 19010 17614 19022 17666
rect 20402 17614 20414 17666
rect 20466 17614 20478 17666
rect 20738 17614 20750 17666
rect 20802 17614 20814 17666
rect 26226 17614 26238 17666
rect 26290 17614 26302 17666
rect 28354 17614 28366 17666
rect 28418 17614 28430 17666
rect 28914 17614 28926 17666
rect 28978 17614 28990 17666
rect 30146 17614 30158 17666
rect 30210 17614 30222 17666
rect 31042 17614 31054 17666
rect 31106 17614 31118 17666
rect 16718 17602 16770 17614
rect 19518 17602 19570 17614
rect 29710 17602 29762 17614
rect 31614 17602 31666 17614
rect 34526 17666 34578 17678
rect 34526 17602 34578 17614
rect 35198 17666 35250 17678
rect 37998 17666 38050 17678
rect 41918 17666 41970 17678
rect 44046 17666 44098 17678
rect 47406 17666 47458 17678
rect 54238 17666 54290 17678
rect 36642 17614 36654 17666
rect 36706 17614 36718 17666
rect 37090 17614 37102 17666
rect 37154 17614 37166 17666
rect 38546 17614 38558 17666
rect 38610 17614 38622 17666
rect 39330 17614 39342 17666
rect 39394 17614 39406 17666
rect 40562 17614 40574 17666
rect 40626 17614 40638 17666
rect 41010 17614 41022 17666
rect 41074 17614 41086 17666
rect 42242 17614 42254 17666
rect 42306 17614 42318 17666
rect 43250 17614 43262 17666
rect 43314 17614 43326 17666
rect 45042 17614 45054 17666
rect 45106 17614 45118 17666
rect 48178 17614 48190 17666
rect 48242 17614 48254 17666
rect 35198 17602 35250 17614
rect 37998 17602 38050 17614
rect 41918 17602 41970 17614
rect 44046 17602 44098 17614
rect 47406 17602 47458 17614
rect 54238 17602 54290 17614
rect 55022 17666 55074 17678
rect 55346 17614 55358 17666
rect 55410 17614 55422 17666
rect 56130 17614 56142 17666
rect 56194 17614 56206 17666
rect 55022 17602 55074 17614
rect 4398 17554 4450 17566
rect 4398 17490 4450 17502
rect 4734 17554 4786 17566
rect 21198 17554 21250 17566
rect 16930 17502 16942 17554
rect 16994 17502 17006 17554
rect 4734 17490 4786 17502
rect 21198 17490 21250 17502
rect 28030 17554 28082 17566
rect 40238 17554 40290 17566
rect 53566 17554 53618 17566
rect 32610 17502 32622 17554
rect 32674 17502 32686 17554
rect 48850 17502 48862 17554
rect 48914 17502 48926 17554
rect 50978 17502 50990 17554
rect 51042 17502 51054 17554
rect 51538 17502 51550 17554
rect 51602 17502 51614 17554
rect 28030 17490 28082 17502
rect 40238 17490 40290 17502
rect 53566 17490 53618 17502
rect 54014 17554 54066 17566
rect 54014 17490 54066 17502
rect 10670 17442 10722 17454
rect 10670 17378 10722 17390
rect 13806 17442 13858 17454
rect 13806 17378 13858 17390
rect 24670 17442 24722 17454
rect 24670 17378 24722 17390
rect 31726 17442 31778 17454
rect 31726 17378 31778 17390
rect 34190 17442 34242 17454
rect 34190 17378 34242 17390
rect 53118 17442 53170 17454
rect 53118 17378 53170 17390
rect 54350 17442 54402 17454
rect 54786 17390 54798 17442
rect 54850 17390 54862 17442
rect 54350 17378 54402 17390
rect 672 17274 56784 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 43806 17274
rect 43858 17222 43910 17274
rect 43962 17222 44014 17274
rect 44066 17222 56784 17274
rect 672 17188 56784 17222
rect 3390 17106 3442 17118
rect 3390 17042 3442 17054
rect 8542 17106 8594 17118
rect 8542 17042 8594 17054
rect 14926 17106 14978 17118
rect 14926 17042 14978 17054
rect 15486 17106 15538 17118
rect 15486 17042 15538 17054
rect 17726 17106 17778 17118
rect 17726 17042 17778 17054
rect 19966 17106 20018 17118
rect 19966 17042 20018 17054
rect 30270 17106 30322 17118
rect 30270 17042 30322 17054
rect 38110 17106 38162 17118
rect 38110 17042 38162 17054
rect 40350 17106 40402 17118
rect 40350 17042 40402 17054
rect 42590 17106 42642 17118
rect 42590 17042 42642 17054
rect 50318 17106 50370 17118
rect 53566 17106 53618 17118
rect 51314 17054 51326 17106
rect 51378 17054 51390 17106
rect 50318 17042 50370 17054
rect 53566 17042 53618 17054
rect 5406 16994 5458 17006
rect 8990 16994 9042 17006
rect 23774 16994 23826 17006
rect 43486 16994 43538 17006
rect 1810 16942 1822 16994
rect 1874 16942 1886 16994
rect 6962 16942 6974 16994
rect 7026 16942 7038 16994
rect 13346 16942 13358 16994
rect 13410 16942 13422 16994
rect 16146 16942 16158 16994
rect 16210 16942 16222 16994
rect 18386 16942 18398 16994
rect 18450 16942 18462 16994
rect 21746 16942 21758 16994
rect 21810 16942 21822 16994
rect 28690 16942 28702 16994
rect 28754 16942 28766 16994
rect 32834 16942 32846 16994
rect 32898 16942 32910 16994
rect 48178 16942 48190 16994
rect 48242 16942 48254 16994
rect 52322 16942 52334 16994
rect 52386 16942 52398 16994
rect 55122 16942 55134 16994
rect 55186 16942 55198 16994
rect 5406 16930 5458 16942
rect 8990 16930 9042 16942
rect 23774 16930 23826 16942
rect 43486 16930 43538 16942
rect 3726 16882 3778 16894
rect 3726 16818 3778 16830
rect 4286 16882 4338 16894
rect 4286 16818 4338 16830
rect 5966 16882 6018 16894
rect 15374 16882 15426 16894
rect 9314 16830 9326 16882
rect 9378 16830 9390 16882
rect 9762 16830 9774 16882
rect 9826 16830 9838 16882
rect 10546 16830 10558 16882
rect 10610 16830 10622 16882
rect 11218 16830 11230 16882
rect 11282 16830 11294 16882
rect 12002 16830 12014 16882
rect 12066 16830 12078 16882
rect 5966 16818 6018 16830
rect 15374 16818 15426 16830
rect 23326 16882 23378 16894
rect 25230 16882 25282 16894
rect 42926 16882 42978 16894
rect 24098 16830 24110 16882
rect 24162 16830 24174 16882
rect 24546 16830 24558 16882
rect 24610 16830 24622 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 26786 16830 26798 16882
rect 26850 16830 26862 16882
rect 32946 16830 32958 16882
rect 33010 16830 33022 16882
rect 33282 16830 33294 16882
rect 33346 16830 33358 16882
rect 33842 16830 33854 16882
rect 33906 16830 33918 16882
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 38770 16830 38782 16882
rect 38834 16830 38846 16882
rect 40898 16830 40910 16882
rect 40962 16830 40974 16882
rect 23326 16818 23378 16830
rect 25230 16818 25282 16830
rect 42926 16818 42978 16830
rect 43374 16882 43426 16894
rect 46286 16882 46338 16894
rect 45938 16830 45950 16882
rect 46002 16830 46014 16882
rect 43374 16818 43426 16830
rect 46286 16818 46338 16830
rect 46958 16882 47010 16894
rect 46958 16818 47010 16830
rect 47630 16882 47682 16894
rect 47630 16818 47682 16830
rect 50206 16882 50258 16894
rect 50206 16818 50258 16830
rect 50766 16882 50818 16894
rect 50766 16818 50818 16830
rect 50990 16882 51042 16894
rect 55694 16882 55746 16894
rect 52434 16830 52446 16882
rect 52498 16830 52510 16882
rect 50990 16818 51042 16830
rect 55694 16818 55746 16830
rect 32510 16770 32562 16782
rect 2258 16718 2270 16770
rect 2322 16718 2334 16770
rect 5618 16718 5630 16770
rect 5682 16718 5694 16770
rect 9986 16718 9998 16770
rect 10050 16718 10062 16770
rect 13794 16718 13806 16770
rect 13858 16718 13870 16770
rect 16482 16718 16494 16770
rect 16546 16718 16558 16770
rect 18834 16718 18846 16770
rect 18898 16718 18910 16770
rect 22194 16718 22206 16770
rect 22258 16718 22270 16770
rect 24770 16718 24782 16770
rect 24834 16718 24846 16770
rect 32510 16706 32562 16718
rect 32734 16770 32786 16782
rect 43598 16770 43650 16782
rect 47294 16770 47346 16782
rect 49758 16770 49810 16782
rect 36978 16718 36990 16770
rect 37042 16718 37054 16770
rect 45378 16718 45390 16770
rect 45442 16718 45454 16770
rect 48626 16718 48638 16770
rect 48690 16718 48702 16770
rect 32734 16706 32786 16718
rect 43598 16706 43650 16718
rect 47294 16706 47346 16718
rect 49758 16706 49810 16718
rect 52782 16770 52834 16782
rect 52782 16706 52834 16718
rect 52894 16770 52946 16782
rect 52894 16706 52946 16718
rect 53118 16770 53170 16782
rect 54674 16718 54686 16770
rect 54738 16718 54750 16770
rect 53118 16706 53170 16718
rect 4174 16658 4226 16670
rect 4174 16594 4226 16606
rect 4398 16658 4450 16670
rect 15486 16658 15538 16670
rect 35422 16658 35474 16670
rect 44270 16658 44322 16670
rect 7410 16606 7422 16658
rect 7474 16606 7486 16658
rect 29138 16606 29150 16658
rect 29202 16606 29214 16658
rect 34290 16606 34302 16658
rect 34354 16606 34366 16658
rect 39218 16606 39230 16658
rect 39282 16606 39294 16658
rect 41458 16606 41470 16658
rect 41522 16606 41534 16658
rect 4398 16594 4450 16606
rect 15486 16594 15538 16606
rect 35422 16594 35474 16606
rect 44270 16594 44322 16606
rect 46622 16658 46674 16670
rect 46622 16594 46674 16606
rect 46846 16658 46898 16670
rect 46846 16594 46898 16606
rect 47406 16658 47458 16670
rect 47406 16594 47458 16606
rect 50318 16658 50370 16670
rect 56018 16606 56030 16658
rect 56082 16606 56094 16658
rect 50318 16594 50370 16606
rect 672 16490 56784 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 44466 16490
rect 44518 16438 44570 16490
rect 44622 16438 44674 16490
rect 44726 16438 56784 16490
rect 672 16404 56784 16438
rect 2830 16322 2882 16334
rect 6862 16322 6914 16334
rect 7422 16322 7474 16334
rect 4274 16270 4286 16322
rect 4338 16270 4350 16322
rect 7074 16270 7086 16322
rect 7138 16270 7150 16322
rect 2830 16258 2882 16270
rect 6862 16258 6914 16270
rect 7422 16258 7474 16270
rect 7758 16322 7810 16334
rect 7758 16258 7810 16270
rect 8990 16322 9042 16334
rect 13022 16322 13074 16334
rect 10322 16270 10334 16322
rect 10386 16270 10398 16322
rect 8990 16258 9042 16270
rect 13022 16258 13074 16270
rect 13582 16322 13634 16334
rect 28366 16322 28418 16334
rect 36654 16322 36706 16334
rect 40574 16322 40626 16334
rect 21186 16270 21198 16322
rect 21250 16270 21262 16322
rect 30594 16270 30606 16322
rect 30658 16270 30670 16322
rect 35522 16270 35534 16322
rect 35586 16270 35598 16322
rect 38322 16270 38334 16322
rect 38386 16270 38398 16322
rect 13582 16258 13634 16270
rect 28366 16258 28418 16270
rect 36654 16258 36706 16270
rect 40574 16258 40626 16270
rect 42702 16322 42754 16334
rect 42702 16258 42754 16270
rect 46398 16322 46450 16334
rect 46398 16258 46450 16270
rect 48862 16322 48914 16334
rect 48862 16258 48914 16270
rect 49198 16322 49250 16334
rect 49198 16258 49250 16270
rect 49310 16322 49362 16334
rect 49310 16258 49362 16270
rect 49646 16322 49698 16334
rect 54798 16322 54850 16334
rect 53442 16270 53454 16322
rect 53506 16270 53518 16322
rect 49646 16258 49698 16270
rect 54798 16258 54850 16270
rect 56030 16322 56082 16334
rect 56354 16270 56366 16322
rect 56418 16270 56430 16322
rect 56030 16258 56082 16270
rect 8878 16210 8930 16222
rect 1586 16158 1598 16210
rect 1650 16158 1662 16210
rect 8082 16158 8094 16210
rect 8146 16158 8158 16210
rect 8878 16146 8930 16158
rect 10782 16210 10834 16222
rect 16046 16210 16098 16222
rect 20190 16210 20242 16222
rect 45390 16210 45442 16222
rect 14802 16158 14814 16210
rect 14866 16158 14878 16210
rect 18498 16158 18510 16210
rect 18562 16158 18574 16210
rect 27234 16158 27246 16210
rect 27298 16158 27310 16210
rect 32946 16158 32958 16210
rect 33010 16158 33022 16210
rect 41458 16158 41470 16210
rect 41522 16158 41534 16210
rect 44370 16158 44382 16210
rect 44434 16158 44446 16210
rect 10782 16146 10834 16158
rect 16046 16146 16098 16158
rect 20190 16146 20242 16158
rect 45390 16146 45442 16158
rect 45502 16210 45554 16222
rect 45502 16146 45554 16158
rect 47182 16210 47234 16222
rect 47182 16146 47234 16158
rect 47406 16210 47458 16222
rect 47406 16146 47458 16158
rect 49422 16210 49474 16222
rect 49422 16146 49474 16158
rect 51550 16210 51602 16222
rect 51550 16146 51602 16158
rect 4958 16098 5010 16110
rect 13358 16098 13410 16110
rect 1250 16046 1262 16098
rect 1314 16046 1326 16098
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 4050 16046 4062 16098
rect 4114 16046 4126 16098
rect 5506 16046 5518 16098
rect 5570 16046 5582 16098
rect 6290 16046 6302 16098
rect 6354 16046 6366 16098
rect 9650 16046 9662 16098
rect 9714 16046 9726 16098
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 11330 16046 11342 16098
rect 11394 16046 11406 16098
rect 12450 16046 12462 16098
rect 12514 16046 12526 16098
rect 4958 16034 5010 16046
rect 13358 16034 13410 16046
rect 14030 16098 14082 16110
rect 19742 16098 19794 16110
rect 21870 16098 21922 16110
rect 45614 16098 45666 16110
rect 14354 16046 14366 16098
rect 14418 16046 14430 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 20962 16046 20974 16098
rect 21026 16046 21038 16098
rect 22418 16046 22430 16098
rect 22482 16046 22494 16098
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 26674 16046 26686 16098
rect 26738 16046 26750 16098
rect 30034 16046 30046 16098
rect 30098 16046 30110 16098
rect 32610 16046 32622 16098
rect 32674 16046 32686 16098
rect 34962 16046 34974 16098
rect 35026 16046 35038 16098
rect 38882 16046 38894 16098
rect 38946 16046 38958 16098
rect 41010 16046 41022 16098
rect 41074 16046 41086 16098
rect 44818 16046 44830 16098
rect 44882 16046 44894 16098
rect 14030 16034 14082 16046
rect 19742 16034 19794 16046
rect 21870 16034 21922 16046
rect 45614 16034 45666 16046
rect 46062 16098 46114 16110
rect 46062 16034 46114 16046
rect 46174 16098 46226 16110
rect 46174 16034 46226 16046
rect 46622 16098 46674 16110
rect 46622 16034 46674 16046
rect 46734 16098 46786 16110
rect 46734 16034 46786 16046
rect 48190 16098 48242 16110
rect 48190 16034 48242 16046
rect 48638 16098 48690 16110
rect 48638 16034 48690 16046
rect 51438 16098 51490 16110
rect 51438 16034 51490 16046
rect 51998 16098 52050 16110
rect 51998 16034 52050 16046
rect 52334 16098 52386 16110
rect 52334 16034 52386 16046
rect 54574 16098 54626 16110
rect 54574 16034 54626 16046
rect 54686 16098 54738 16110
rect 55246 16098 55298 16110
rect 54898 16046 54910 16098
rect 54962 16046 54974 16098
rect 54686 16034 54738 16046
rect 55246 16034 55298 16046
rect 3278 15986 3330 15998
rect 3278 15922 3330 15934
rect 9326 15986 9378 15998
rect 9326 15922 9378 15934
rect 12910 15986 12962 15998
rect 12910 15922 12962 15934
rect 13470 15986 13522 15998
rect 37214 15986 37266 15998
rect 18162 15934 18174 15986
rect 18226 15934 18238 15986
rect 13470 15922 13522 15934
rect 37214 15922 37266 15934
rect 40462 15986 40514 15998
rect 40462 15922 40514 15934
rect 48750 15986 48802 15998
rect 48750 15922 48802 15934
rect 50094 15986 50146 15998
rect 50094 15922 50146 15934
rect 50206 15986 50258 15998
rect 50206 15922 50258 15934
rect 50542 15986 50594 15998
rect 53890 15934 53902 15986
rect 53954 15934 53966 15986
rect 50542 15922 50594 15934
rect 31726 15874 31778 15886
rect 31726 15810 31778 15822
rect 34190 15874 34242 15886
rect 34190 15810 34242 15822
rect 43262 15874 43314 15886
rect 43262 15810 43314 15822
rect 47518 15874 47570 15886
rect 47518 15810 47570 15822
rect 50766 15874 50818 15886
rect 50766 15810 50818 15822
rect 50878 15874 50930 15886
rect 51874 15822 51886 15874
rect 51938 15822 51950 15874
rect 50878 15810 50930 15822
rect 672 15706 56784 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 43806 15706
rect 43858 15654 43910 15706
rect 43962 15654 44014 15706
rect 44066 15654 56784 15706
rect 672 15620 56784 15654
rect 1150 15538 1202 15550
rect 1150 15474 1202 15486
rect 22430 15538 22482 15550
rect 22430 15474 22482 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 46286 15538 46338 15550
rect 46286 15474 46338 15486
rect 48302 15538 48354 15550
rect 48302 15474 48354 15486
rect 52110 15538 52162 15550
rect 52110 15474 52162 15486
rect 56142 15538 56194 15550
rect 56142 15474 56194 15486
rect 3726 15426 3778 15438
rect 2706 15374 2718 15426
rect 2770 15374 2782 15426
rect 3726 15362 3778 15374
rect 5742 15426 5794 15438
rect 31950 15426 32002 15438
rect 10546 15374 10558 15426
rect 10610 15374 10622 15426
rect 5742 15362 5794 15374
rect 31950 15362 32002 15374
rect 37550 15426 37602 15438
rect 42802 15374 42814 15426
rect 42866 15374 42878 15426
rect 53666 15374 53678 15426
rect 53730 15374 53742 15426
rect 54562 15374 54574 15426
rect 54626 15374 54638 15426
rect 37550 15362 37602 15374
rect 3278 15314 3330 15326
rect 3278 15250 3330 15262
rect 3502 15314 3554 15326
rect 3502 15250 3554 15262
rect 4174 15314 4226 15326
rect 4174 15250 4226 15262
rect 4958 15314 5010 15326
rect 18510 15314 18562 15326
rect 33630 15314 33682 15326
rect 46846 15314 46898 15326
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 6626 15262 6638 15314
rect 6690 15262 6702 15314
rect 7970 15262 7982 15314
rect 8034 15262 8046 15314
rect 8866 15262 8878 15314
rect 8930 15262 8942 15314
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 13570 15262 13582 15314
rect 13634 15262 13646 15314
rect 14354 15262 14366 15314
rect 14418 15262 14430 15314
rect 14802 15262 14814 15314
rect 14866 15262 14878 15314
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 17154 15262 17166 15314
rect 17218 15262 17230 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 20738 15262 20750 15314
rect 20802 15262 20814 15314
rect 24434 15262 24446 15314
rect 24498 15262 24510 15314
rect 32274 15262 32286 15314
rect 32338 15262 32350 15314
rect 32722 15262 32734 15314
rect 32786 15262 32798 15314
rect 34178 15262 34190 15314
rect 34242 15262 34254 15314
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 37874 15262 37886 15314
rect 37938 15262 37950 15314
rect 38434 15262 38446 15314
rect 38498 15262 38510 15314
rect 39106 15262 39118 15314
rect 39170 15262 39182 15314
rect 39554 15262 39566 15314
rect 39618 15262 39630 15314
rect 40674 15262 40686 15314
rect 40738 15262 40750 15314
rect 44706 15262 44718 15314
rect 44770 15262 44782 15314
rect 4958 15250 5010 15262
rect 18510 15250 18562 15262
rect 33630 15250 33682 15262
rect 46846 15250 46898 15262
rect 47182 15314 47234 15326
rect 47182 15250 47234 15262
rect 47406 15314 47458 15326
rect 47406 15250 47458 15262
rect 47742 15314 47794 15326
rect 51438 15314 51490 15326
rect 49970 15262 49982 15314
rect 50034 15262 50046 15314
rect 50642 15262 50654 15314
rect 50706 15262 50718 15314
rect 47742 15250 47794 15262
rect 51438 15250 51490 15262
rect 3950 15202 4002 15214
rect 7198 15202 7250 15214
rect 9662 15202 9714 15214
rect 12126 15202 12178 15214
rect 2370 15150 2382 15202
rect 2434 15150 2446 15202
rect 5282 15150 5294 15202
rect 5346 15150 5358 15202
rect 9314 15150 9326 15202
rect 9378 15150 9390 15202
rect 10882 15150 10894 15202
rect 10946 15150 10958 15202
rect 3950 15138 4002 15150
rect 7198 15138 7250 15150
rect 9662 15138 9714 15150
rect 12126 15138 12178 15150
rect 12798 15202 12850 15214
rect 16830 15202 16882 15214
rect 43374 15202 43426 15214
rect 13794 15150 13806 15202
rect 13858 15150 13870 15202
rect 17826 15150 17838 15202
rect 17890 15150 17902 15202
rect 21298 15150 21310 15202
rect 21362 15150 21374 15202
rect 24882 15150 24894 15202
rect 24946 15150 24958 15202
rect 38546 15150 38558 15202
rect 38610 15150 38622 15202
rect 42354 15150 42366 15202
rect 42418 15150 42430 15202
rect 12798 15138 12850 15150
rect 16830 15138 16882 15150
rect 43374 15138 43426 15150
rect 43486 15202 43538 15214
rect 46958 15202 47010 15214
rect 45154 15150 45166 15202
rect 45218 15150 45230 15202
rect 43486 15138 43538 15150
rect 46958 15138 47010 15150
rect 47518 15202 47570 15214
rect 49410 15150 49422 15202
rect 49474 15150 49486 15202
rect 50418 15150 50430 15202
rect 50482 15150 50494 15202
rect 51090 15150 51102 15202
rect 51154 15150 51166 15202
rect 53330 15150 53342 15202
rect 53394 15150 53406 15202
rect 54898 15150 54910 15202
rect 54962 15150 54974 15202
rect 47518 15138 47570 15150
rect 4062 15090 4114 15102
rect 26126 15090 26178 15102
rect 41246 15090 41298 15102
rect 6738 15038 6750 15090
rect 6802 15038 6814 15090
rect 32946 15038 32958 15090
rect 33010 15038 33022 15090
rect 4062 15026 4114 15038
rect 26126 15026 26178 15038
rect 41246 15026 41298 15038
rect 672 14922 56784 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 44466 14922
rect 44518 14870 44570 14922
rect 44622 14870 44674 14922
rect 44726 14870 56784 14922
rect 672 14836 56784 14870
rect 2382 14754 2434 14766
rect 2382 14690 2434 14702
rect 4622 14754 4674 14766
rect 18622 14754 18674 14766
rect 44942 14754 44994 14766
rect 8866 14702 8878 14754
rect 8930 14702 8942 14754
rect 17490 14702 17502 14754
rect 17554 14702 17566 14754
rect 29586 14702 29598 14754
rect 29650 14702 29662 14754
rect 35970 14702 35982 14754
rect 36034 14702 36046 14754
rect 42018 14702 42030 14754
rect 42082 14702 42094 14754
rect 4622 14690 4674 14702
rect 18622 14690 18674 14702
rect 44942 14690 44994 14702
rect 45166 14754 45218 14766
rect 45166 14690 45218 14702
rect 49870 14754 49922 14766
rect 53342 14754 53394 14766
rect 50866 14702 50878 14754
rect 50930 14702 50942 14754
rect 52546 14702 52558 14754
rect 52610 14702 52622 14754
rect 49870 14690 49922 14702
rect 53342 14690 53394 14702
rect 56030 14754 56082 14766
rect 56354 14702 56366 14754
rect 56418 14702 56430 14754
rect 56030 14690 56082 14702
rect 1598 14642 1650 14654
rect 1598 14578 1650 14590
rect 1822 14642 1874 14654
rect 1822 14578 1874 14590
rect 2494 14642 2546 14654
rect 9886 14642 9938 14654
rect 19070 14642 19122 14654
rect 24670 14642 24722 14654
rect 26126 14642 26178 14654
rect 3490 14590 3502 14642
rect 3554 14590 3566 14642
rect 6066 14590 6078 14642
rect 6130 14590 6142 14642
rect 10882 14590 10894 14642
rect 10946 14590 10958 14642
rect 14802 14590 14814 14642
rect 14866 14590 14878 14642
rect 20066 14590 20078 14642
rect 20130 14590 20142 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 2494 14578 2546 14590
rect 9886 14578 9938 14590
rect 19070 14578 19122 14590
rect 24670 14578 24722 14590
rect 26126 14578 26178 14590
rect 41022 14642 41074 14654
rect 48638 14642 48690 14654
rect 46162 14590 46174 14642
rect 46226 14590 46238 14642
rect 41022 14578 41074 14590
rect 48638 14578 48690 14590
rect 48750 14642 48802 14654
rect 48750 14578 48802 14590
rect 48974 14642 49026 14654
rect 49522 14590 49534 14642
rect 49586 14590 49598 14642
rect 54450 14590 54462 14642
rect 54514 14590 54526 14642
rect 48974 14578 49026 14590
rect 1150 14530 1202 14542
rect 11342 14530 11394 14542
rect 20750 14530 20802 14542
rect 30270 14530 30322 14542
rect 36654 14530 36706 14542
rect 42702 14530 42754 14542
rect 44830 14530 44882 14542
rect 52894 14530 52946 14542
rect 2146 14478 2158 14530
rect 2210 14478 2222 14530
rect 3042 14478 3054 14530
rect 3106 14478 3118 14530
rect 5394 14478 5406 14530
rect 5458 14478 5470 14530
rect 5842 14478 5854 14530
rect 5906 14478 5918 14530
rect 6626 14478 6638 14530
rect 6690 14478 6702 14530
rect 7298 14478 7310 14530
rect 7362 14478 7374 14530
rect 8082 14478 8094 14530
rect 8146 14478 8158 14530
rect 9090 14478 9102 14530
rect 9154 14478 9166 14530
rect 10322 14478 10334 14530
rect 10386 14478 10398 14530
rect 10658 14478 10670 14530
rect 10722 14478 10734 14530
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 12114 14478 12126 14530
rect 12178 14478 12190 14530
rect 12898 14478 12910 14530
rect 12962 14478 12974 14530
rect 14466 14478 14478 14530
rect 14530 14478 14542 14530
rect 17042 14478 17054 14530
rect 17106 14478 17118 14530
rect 19506 14478 19518 14530
rect 19570 14478 19582 14530
rect 19954 14478 19966 14530
rect 20018 14478 20030 14530
rect 21074 14478 21086 14530
rect 21138 14478 21150 14530
rect 21298 14478 21310 14530
rect 21362 14478 21374 14530
rect 22082 14478 22094 14530
rect 22146 14478 22158 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 25554 14478 25566 14530
rect 25618 14478 25630 14530
rect 26786 14478 26798 14530
rect 26850 14478 26862 14530
rect 27794 14478 27806 14530
rect 27858 14478 27870 14530
rect 28914 14478 28926 14530
rect 28978 14478 28990 14530
rect 29474 14478 29486 14530
rect 29538 14478 29550 14530
rect 30594 14478 30606 14530
rect 30658 14478 30670 14530
rect 31602 14478 31614 14530
rect 31666 14478 31678 14530
rect 35410 14478 35422 14530
rect 35474 14478 35486 14530
rect 35858 14478 35870 14530
rect 35922 14478 35934 14530
rect 36978 14478 36990 14530
rect 37042 14478 37054 14530
rect 37986 14478 37998 14530
rect 38050 14478 38062 14530
rect 41346 14478 41358 14530
rect 41410 14478 41422 14530
rect 41794 14478 41806 14530
rect 41858 14478 41870 14530
rect 43026 14478 43038 14530
rect 43090 14478 43102 14530
rect 44034 14478 44046 14530
rect 44098 14478 44110 14530
rect 45714 14478 45726 14530
rect 45778 14478 45790 14530
rect 54898 14478 54910 14530
rect 54962 14478 54974 14530
rect 1150 14466 1202 14478
rect 11342 14466 11394 14478
rect 20750 14466 20802 14478
rect 30270 14466 30322 14478
rect 36654 14466 36706 14478
rect 42702 14466 42754 14478
rect 44830 14466 44882 14478
rect 52894 14466 52946 14478
rect 1038 14418 1090 14430
rect 5070 14418 5122 14430
rect 1474 14366 1486 14418
rect 1538 14366 1550 14418
rect 1038 14354 1090 14366
rect 5070 14354 5122 14366
rect 28590 14418 28642 14430
rect 28590 14354 28642 14366
rect 34974 14418 35026 14430
rect 34974 14354 35026 14366
rect 48414 14418 48466 14430
rect 50418 14366 50430 14418
rect 50482 14366 50494 14418
rect 48414 14354 48466 14366
rect 16046 14306 16098 14318
rect 16046 14242 16098 14254
rect 47294 14306 47346 14318
rect 47294 14242 47346 14254
rect 48190 14306 48242 14318
rect 48190 14242 48242 14254
rect 51998 14306 52050 14318
rect 51998 14242 52050 14254
rect 672 14138 56784 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 43806 14138
rect 43858 14086 43910 14138
rect 43962 14086 44014 14138
rect 44066 14086 56784 14138
rect 672 14052 56784 14086
rect 4958 13970 5010 13982
rect 4958 13906 5010 13918
rect 12126 13970 12178 13982
rect 12126 13906 12178 13918
rect 13246 13970 13298 13982
rect 13246 13906 13298 13918
rect 13582 13970 13634 13982
rect 13582 13906 13634 13918
rect 19070 13970 19122 13982
rect 19070 13906 19122 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 30494 13970 30546 13982
rect 30494 13906 30546 13918
rect 39118 13970 39170 13982
rect 39118 13906 39170 13918
rect 43486 13970 43538 13982
rect 43486 13906 43538 13918
rect 48526 13970 48578 13982
rect 48526 13906 48578 13918
rect 55582 13970 55634 13982
rect 55582 13906 55634 13918
rect 1710 13858 1762 13870
rect 5966 13858 6018 13870
rect 14814 13858 14866 13870
rect 2146 13806 2158 13858
rect 2210 13806 2222 13858
rect 10546 13806 10558 13858
rect 10610 13806 10622 13858
rect 1710 13794 1762 13806
rect 5966 13794 6018 13806
rect 14814 13794 14866 13806
rect 18622 13858 18674 13870
rect 20638 13858 20690 13870
rect 32286 13858 32338 13870
rect 44158 13858 44210 13870
rect 19842 13806 19854 13858
rect 19906 13806 19918 13858
rect 28914 13806 28926 13858
rect 28978 13806 28990 13858
rect 37538 13806 37550 13858
rect 37602 13806 37614 13858
rect 18622 13794 18674 13806
rect 20638 13794 20690 13806
rect 32286 13794 32338 13806
rect 44158 13794 44210 13806
rect 52894 13858 52946 13870
rect 52894 13794 52946 13806
rect 55694 13858 55746 13870
rect 55694 13794 55746 13806
rect 7422 13746 7474 13758
rect 16270 13746 16322 13758
rect 19294 13746 19346 13758
rect 33966 13746 34018 13758
rect 47966 13746 48018 13758
rect 51102 13746 51154 13758
rect 6290 13694 6302 13746
rect 6354 13694 6366 13746
rect 6850 13694 6862 13746
rect 6914 13694 6926 13746
rect 7970 13694 7982 13746
rect 8034 13694 8046 13746
rect 8194 13694 8206 13746
rect 8258 13694 8270 13746
rect 8978 13694 8990 13746
rect 9042 13694 9054 13746
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 15250 13694 15262 13746
rect 15314 13694 15326 13746
rect 15586 13694 15598 13746
rect 15650 13694 15662 13746
rect 16818 13694 16830 13746
rect 16882 13694 16894 13746
rect 17826 13694 17838 13746
rect 17890 13694 17902 13746
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 20962 13694 20974 13746
rect 21026 13694 21038 13746
rect 21410 13694 21422 13746
rect 21474 13694 21486 13746
rect 22754 13694 22766 13746
rect 22818 13694 22830 13746
rect 23650 13694 23662 13746
rect 23714 13694 23726 13746
rect 25890 13694 25902 13746
rect 25954 13694 25966 13746
rect 32722 13694 32734 13746
rect 32786 13694 32798 13746
rect 33058 13694 33070 13746
rect 33122 13694 33134 13746
rect 34402 13694 34414 13746
rect 34466 13694 34478 13746
rect 35298 13694 35310 13746
rect 35362 13694 35374 13746
rect 39778 13694 39790 13746
rect 39842 13694 39854 13746
rect 44482 13694 44494 13746
rect 44546 13694 44558 13746
rect 44930 13694 44942 13746
rect 44994 13694 45006 13746
rect 46162 13694 46174 13746
rect 46226 13694 46238 13746
rect 47170 13694 47182 13746
rect 47234 13694 47246 13746
rect 50082 13694 50094 13746
rect 50146 13694 50158 13746
rect 7422 13682 7474 13694
rect 16270 13682 16322 13694
rect 19294 13682 19346 13694
rect 33966 13682 34018 13694
rect 47966 13682 48018 13694
rect 51102 13682 51154 13694
rect 52334 13746 52386 13758
rect 55010 13694 55022 13746
rect 55074 13694 55086 13746
rect 56130 13694 56142 13746
rect 56194 13694 56206 13746
rect 52334 13682 52386 13694
rect 5070 13634 5122 13646
rect 1026 13582 1038 13634
rect 1090 13582 1102 13634
rect 5070 13570 5122 13582
rect 5294 13634 5346 13646
rect 18734 13634 18786 13646
rect 9538 13582 9550 13634
rect 9602 13582 9614 13634
rect 10994 13582 11006 13634
rect 11058 13582 11070 13634
rect 13906 13582 13918 13634
rect 13970 13582 13982 13634
rect 14354 13582 14366 13634
rect 14418 13582 14430 13634
rect 15810 13582 15822 13634
rect 15874 13582 15886 13634
rect 5294 13570 5346 13582
rect 18734 13570 18786 13582
rect 22094 13634 22146 13646
rect 43598 13634 43650 13646
rect 29250 13582 29262 13634
rect 29314 13582 29326 13634
rect 33282 13582 33294 13634
rect 33346 13582 33358 13634
rect 37986 13582 37998 13634
rect 38050 13582 38062 13634
rect 40226 13582 40238 13634
rect 40290 13582 40302 13634
rect 22094 13570 22146 13582
rect 43598 13570 43650 13582
rect 45614 13634 45666 13646
rect 45614 13570 45666 13582
rect 50878 13634 50930 13646
rect 50878 13570 50930 13582
rect 51998 13634 52050 13646
rect 51998 13570 52050 13582
rect 52558 13634 52610 13646
rect 52558 13570 52610 13582
rect 53006 13634 53058 13646
rect 54562 13582 54574 13634
rect 54626 13582 54638 13634
rect 56354 13582 56366 13634
rect 56418 13582 56430 13634
rect 53006 13570 53058 13582
rect 1374 13522 1426 13534
rect 3726 13522 3778 13534
rect 18510 13522 18562 13534
rect 2594 13470 2606 13522
rect 2658 13470 2670 13522
rect 6962 13470 6974 13522
rect 7026 13470 7038 13522
rect 1374 13458 1426 13470
rect 3726 13458 3778 13470
rect 18510 13458 18562 13470
rect 19742 13522 19794 13534
rect 19742 13458 19794 13470
rect 19966 13522 20018 13534
rect 41358 13522 41410 13534
rect 48078 13522 48130 13534
rect 52110 13522 52162 13534
rect 21634 13470 21646 13522
rect 21698 13470 21710 13522
rect 25442 13470 25454 13522
rect 25506 13470 25518 13522
rect 45154 13470 45166 13522
rect 45218 13470 45230 13522
rect 49634 13470 49646 13522
rect 49698 13470 49710 13522
rect 51426 13470 51438 13522
rect 51490 13470 51502 13522
rect 19966 13458 20018 13470
rect 41358 13458 41410 13470
rect 48078 13458 48130 13470
rect 52110 13458 52162 13470
rect 53454 13522 53506 13534
rect 53454 13458 53506 13470
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 1150 13186 1202 13198
rect 15486 13186 15538 13198
rect 23102 13186 23154 13198
rect 28814 13186 28866 13198
rect 2258 13134 2270 13186
rect 2322 13134 2334 13186
rect 4498 13134 4510 13186
rect 4562 13134 4574 13186
rect 7970 13134 7982 13186
rect 8034 13134 8046 13186
rect 17826 13134 17838 13186
rect 17890 13134 17902 13186
rect 25778 13134 25790 13186
rect 25842 13134 25854 13186
rect 1150 13122 1202 13134
rect 15486 13122 15538 13134
rect 23102 13122 23154 13134
rect 28814 13122 28866 13134
rect 34190 13186 34242 13198
rect 36654 13186 36706 13198
rect 45614 13186 45666 13198
rect 35522 13134 35534 13186
rect 35586 13134 35598 13186
rect 37762 13134 37774 13186
rect 37826 13134 37838 13186
rect 41234 13134 41246 13186
rect 41298 13134 41310 13186
rect 34190 13122 34242 13134
rect 36654 13122 36706 13134
rect 45614 13122 45666 13134
rect 46622 13186 46674 13198
rect 46622 13122 46674 13134
rect 46958 13186 47010 13198
rect 46958 13122 47010 13134
rect 47182 13186 47234 13198
rect 47182 13122 47234 13134
rect 47406 13186 47458 13198
rect 47406 13122 47458 13134
rect 48862 13186 48914 13198
rect 48862 13122 48914 13134
rect 52110 13186 52162 13198
rect 52110 13122 52162 13134
rect 52446 13186 52498 13198
rect 52446 13122 52498 13134
rect 53006 13186 53058 13198
rect 53006 13122 53058 13134
rect 53230 13186 53282 13198
rect 54674 13134 54686 13186
rect 54738 13134 54750 13186
rect 56242 13134 56254 13186
rect 56306 13134 56318 13186
rect 53230 13122 53282 13134
rect 3502 13074 3554 13086
rect 3502 13010 3554 13022
rect 8990 13074 9042 13086
rect 8990 13010 9042 13022
rect 9550 13074 9602 13086
rect 16046 13074 16098 13086
rect 22990 13074 23042 13086
rect 11106 13022 11118 13074
rect 11170 13022 11182 13074
rect 14242 13022 14254 13074
rect 14306 13022 14318 13074
rect 20402 13022 20414 13074
rect 20466 13022 20478 13074
rect 9550 13010 9602 13022
rect 16046 13010 16098 13022
rect 22990 13010 23042 13022
rect 23214 13074 23266 13086
rect 46062 13074 46114 13086
rect 27682 13022 27694 13074
rect 27746 13022 27758 13074
rect 33058 13022 33070 13074
rect 33122 13022 33134 13074
rect 44482 13022 44494 13074
rect 44546 13022 44558 13074
rect 23214 13010 23266 13022
rect 46062 13010 46114 13022
rect 46174 13074 46226 13086
rect 51886 13074 51938 13086
rect 50194 13022 50206 13074
rect 50258 13022 50270 13074
rect 46174 13010 46226 13022
rect 51886 13010 51938 13022
rect 52894 13074 52946 13086
rect 52894 13010 52946 13022
rect 6974 12962 7026 12974
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 3826 12910 3838 12962
rect 3890 12910 3902 12962
rect 4386 12910 4398 12962
rect 4450 12910 4462 12962
rect 5058 12910 5070 12962
rect 5122 12910 5134 12962
rect 5730 12910 5742 12962
rect 5794 12910 5806 12962
rect 6626 12910 6638 12962
rect 6690 12910 6702 12962
rect 6974 12898 7026 12910
rect 7422 12962 7474 12974
rect 7422 12898 7474 12910
rect 7534 12962 7586 12974
rect 7534 12898 7586 12910
rect 7646 12962 7698 12974
rect 9102 12962 9154 12974
rect 15822 12962 15874 12974
rect 8194 12910 8206 12962
rect 8258 12910 8270 12962
rect 10546 12910 10558 12962
rect 10610 12910 10622 12962
rect 10882 12910 10894 12962
rect 10946 12910 10958 12962
rect 11666 12910 11678 12962
rect 11730 12910 11742 12962
rect 12338 12910 12350 12962
rect 12402 12910 12414 12962
rect 13122 12910 13134 12962
rect 13186 12910 13198 12962
rect 13906 12910 13918 12962
rect 13970 12910 13982 12962
rect 7646 12898 7698 12910
rect 9102 12898 9154 12910
rect 15822 12898 15874 12910
rect 16158 12962 16210 12974
rect 20862 12962 20914 12974
rect 17266 12910 17278 12962
rect 17330 12910 17342 12962
rect 19730 12910 19742 12962
rect 19794 12910 19806 12962
rect 20178 12910 20190 12962
rect 20242 12910 20254 12962
rect 16158 12898 16210 12910
rect 20862 12898 20914 12910
rect 21086 12962 21138 12974
rect 41694 12962 41746 12974
rect 46510 12962 46562 12974
rect 48750 12962 48802 12974
rect 21522 12910 21534 12962
rect 21586 12910 21598 12962
rect 22530 12910 22542 12962
rect 22594 12910 22606 12962
rect 32610 12910 32622 12962
rect 32674 12910 32686 12962
rect 34962 12910 34974 12962
rect 35026 12910 35038 12962
rect 37314 12910 37326 12962
rect 37378 12910 37390 12962
rect 40674 12910 40686 12962
rect 40738 12910 40750 12962
rect 41010 12910 41022 12962
rect 41074 12910 41086 12962
rect 42242 12910 42254 12962
rect 42306 12910 42318 12962
rect 43362 12910 43374 12962
rect 43426 12910 43438 12962
rect 44034 12910 44046 12962
rect 44098 12910 44110 12962
rect 48626 12910 48638 12962
rect 48690 12910 48702 12962
rect 21086 12898 21138 12910
rect 41694 12898 41746 12910
rect 46510 12898 46562 12910
rect 48750 12898 48802 12910
rect 48974 12962 49026 12974
rect 48974 12898 49026 12910
rect 52334 12962 52386 12974
rect 52334 12898 52386 12910
rect 55918 12962 55970 12974
rect 55918 12898 55970 12910
rect 10110 12850 10162 12862
rect 10110 12786 10162 12798
rect 16718 12850 16770 12862
rect 16718 12786 16770 12798
rect 18958 12850 19010 12862
rect 18958 12786 19010 12798
rect 19406 12850 19458 12862
rect 40238 12850 40290 12862
rect 26226 12798 26238 12850
rect 26290 12798 26302 12850
rect 27234 12798 27246 12850
rect 27298 12798 27310 12850
rect 19406 12786 19458 12798
rect 40238 12786 40290 12798
rect 47070 12850 47122 12862
rect 49858 12798 49870 12850
rect 49922 12798 49934 12850
rect 52434 12798 52446 12850
rect 52498 12798 52510 12850
rect 55122 12798 55134 12850
rect 55186 12798 55198 12850
rect 47070 12786 47122 12798
rect 8990 12738 9042 12750
rect 8990 12674 9042 12686
rect 9438 12738 9490 12750
rect 9438 12674 9490 12686
rect 9774 12738 9826 12750
rect 9774 12674 9826 12686
rect 16830 12738 16882 12750
rect 16830 12674 16882 12686
rect 24670 12738 24722 12750
rect 24670 12674 24722 12686
rect 38894 12738 38946 12750
rect 38894 12674 38946 12686
rect 48078 12738 48130 12750
rect 48078 12674 48130 12686
rect 48302 12738 48354 12750
rect 48302 12674 48354 12686
rect 51438 12738 51490 12750
rect 51438 12674 51490 12686
rect 53566 12738 53618 12750
rect 53566 12674 53618 12686
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 19070 12402 19122 12414
rect 19070 12338 19122 12350
rect 20638 12402 20690 12414
rect 20638 12338 20690 12350
rect 32734 12402 32786 12414
rect 32734 12338 32786 12350
rect 41694 12402 41746 12414
rect 41694 12338 41746 12350
rect 50990 12402 51042 12414
rect 50990 12338 51042 12350
rect 52110 12402 52162 12414
rect 52110 12338 52162 12350
rect 1150 12290 1202 12302
rect 1150 12226 1202 12238
rect 4958 12290 5010 12302
rect 4958 12226 5010 12238
rect 5406 12290 5458 12302
rect 5406 12226 5458 12238
rect 8990 12290 9042 12302
rect 19966 12290 20018 12302
rect 13346 12238 13358 12290
rect 13410 12238 13422 12290
rect 8990 12226 9042 12238
rect 19966 12226 20018 12238
rect 20750 12290 20802 12302
rect 48302 12290 48354 12302
rect 30146 12238 30158 12290
rect 30210 12238 30222 12290
rect 31154 12238 31166 12290
rect 31218 12238 31230 12290
rect 20750 12226 20802 12238
rect 48302 12226 48354 12238
rect 7086 12178 7138 12190
rect 19854 12178 19906 12190
rect 1474 12126 1486 12178
rect 1538 12126 1550 12178
rect 1922 12126 1934 12178
rect 1986 12126 1998 12178
rect 3266 12126 3278 12178
rect 3330 12126 3342 12178
rect 4162 12126 4174 12178
rect 4226 12126 4238 12178
rect 5730 12126 5742 12178
rect 5794 12126 5806 12178
rect 6290 12126 6302 12178
rect 6354 12126 6366 12178
rect 7410 12126 7422 12178
rect 7474 12126 7486 12178
rect 8530 12126 8542 12178
rect 8594 12126 8606 12178
rect 9314 12126 9326 12178
rect 9378 12126 9390 12178
rect 9874 12126 9886 12178
rect 9938 12126 9950 12178
rect 10546 12126 10558 12178
rect 10610 12126 10622 12178
rect 11218 12126 11230 12178
rect 11282 12126 11294 12178
rect 12002 12126 12014 12178
rect 12066 12126 12078 12178
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 16146 12126 16158 12178
rect 16210 12126 16222 12178
rect 17490 12126 17502 12178
rect 17554 12126 17566 12178
rect 18386 12126 18398 12178
rect 18450 12126 18462 12178
rect 7086 12114 7138 12126
rect 19854 12114 19906 12126
rect 20078 12178 20130 12190
rect 23102 12178 23154 12190
rect 25006 12178 25058 12190
rect 47294 12178 47346 12190
rect 20962 12126 20974 12178
rect 21026 12126 21038 12178
rect 21410 12126 21422 12178
rect 21474 12126 21486 12178
rect 23874 12126 23886 12178
rect 23938 12126 23950 12178
rect 24434 12126 24446 12178
rect 24498 12126 24510 12178
rect 25554 12126 25566 12178
rect 25618 12126 25630 12178
rect 26562 12126 26574 12178
rect 26626 12126 26638 12178
rect 33954 12126 33966 12178
rect 34018 12126 34030 12178
rect 38210 12126 38222 12178
rect 38274 12126 38286 12178
rect 39218 12126 39230 12178
rect 39282 12126 39294 12178
rect 40338 12126 40350 12178
rect 40402 12126 40414 12178
rect 40786 12126 40798 12178
rect 40850 12126 40862 12178
rect 43250 12126 43262 12178
rect 43314 12126 43326 12178
rect 20078 12114 20130 12126
rect 23102 12114 23154 12126
rect 25006 12114 25058 12126
rect 47294 12114 47346 12126
rect 47966 12178 48018 12190
rect 47966 12114 48018 12126
rect 49758 12178 49810 12190
rect 49758 12114 49810 12126
rect 52446 12178 52498 12190
rect 56030 12178 56082 12190
rect 54002 12126 54014 12178
rect 54066 12126 54078 12178
rect 52446 12114 52498 12126
rect 56030 12114 56082 12126
rect 2606 12066 2658 12078
rect 2146 12014 2158 12066
rect 2210 12014 2222 12066
rect 2606 12002 2658 12014
rect 6862 12066 6914 12078
rect 6862 12002 6914 12014
rect 15374 12066 15426 12078
rect 16830 12066 16882 12078
rect 16370 12014 16382 12066
rect 16434 12014 16446 12066
rect 15374 12002 15426 12014
rect 16830 12002 16882 12014
rect 19182 12066 19234 12078
rect 23550 12066 23602 12078
rect 36766 12066 36818 12078
rect 21970 12014 21982 12066
rect 22034 12014 22046 12066
rect 29810 12014 29822 12066
rect 29874 12014 29886 12066
rect 31602 12014 31614 12066
rect 31666 12014 31678 12066
rect 34514 12014 34526 12066
rect 34578 12014 34590 12066
rect 19182 12002 19234 12014
rect 23550 12002 23602 12014
rect 36766 12002 36818 12014
rect 39790 12066 39842 12078
rect 39790 12002 39842 12014
rect 41246 12066 41298 12078
rect 41246 12002 41298 12014
rect 47518 12066 47570 12078
rect 47518 12002 47570 12014
rect 47742 12066 47794 12078
rect 47742 12002 47794 12014
rect 48638 12066 48690 12078
rect 49410 12014 49422 12066
rect 49474 12014 49486 12066
rect 50306 12014 50318 12066
rect 50370 12014 50382 12066
rect 50642 12014 50654 12066
rect 50706 12014 50718 12066
rect 52658 12014 52670 12066
rect 52722 12014 52734 12066
rect 52994 12014 53006 12066
rect 53058 12014 53070 12066
rect 54450 12014 54462 12066
rect 54514 12014 54526 12066
rect 56354 12014 56366 12066
rect 56418 12014 56430 12066
rect 48638 12002 48690 12014
rect 5070 11954 5122 11966
rect 14926 11954 14978 11966
rect 6402 11902 6414 11954
rect 6466 11902 6478 11954
rect 9986 11902 9998 11954
rect 10050 11902 10062 11954
rect 13794 11902 13806 11954
rect 13858 11902 13870 11954
rect 5070 11890 5122 11902
rect 14926 11890 14978 11902
rect 19630 11954 19682 11966
rect 28590 11954 28642 11966
rect 24546 11902 24558 11954
rect 24610 11902 24622 11954
rect 19630 11890 19682 11902
rect 28590 11890 28642 11902
rect 35646 11954 35698 11966
rect 35646 11890 35698 11902
rect 36318 11954 36370 11966
rect 36318 11890 36370 11902
rect 36430 11954 36482 11966
rect 36430 11890 36482 11902
rect 36542 11954 36594 11966
rect 48190 11954 48242 11966
rect 40226 11902 40238 11954
rect 40290 11902 40302 11954
rect 42802 11902 42814 11954
rect 42866 11902 42878 11954
rect 36542 11890 36594 11902
rect 48190 11890 48242 11902
rect 48414 11954 48466 11966
rect 48414 11890 48466 11902
rect 51326 11954 51378 11966
rect 51326 11890 51378 11902
rect 55582 11954 55634 11966
rect 55582 11890 55634 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 2830 11618 2882 11630
rect 2830 11554 2882 11566
rect 3390 11618 3442 11630
rect 8206 11618 8258 11630
rect 48190 11618 48242 11630
rect 51886 11618 51938 11630
rect 4498 11566 4510 11618
rect 4562 11566 4574 11618
rect 20178 11566 20190 11618
rect 20242 11566 20254 11618
rect 36530 11566 36542 11618
rect 36594 11566 36606 11618
rect 43026 11566 43038 11618
rect 43090 11566 43102 11618
rect 50754 11566 50766 11618
rect 50818 11566 50830 11618
rect 3390 11554 3442 11566
rect 8206 11554 8258 11566
rect 48190 11554 48242 11566
rect 51886 11554 51938 11566
rect 52446 11618 52498 11630
rect 52446 11554 52498 11566
rect 55022 11618 55074 11630
rect 56354 11566 56366 11618
rect 56418 11566 56430 11618
rect 55022 11554 55074 11566
rect 5854 11506 5906 11518
rect 10222 11506 10274 11518
rect 28702 11506 28754 11518
rect 1586 11454 1598 11506
rect 1650 11454 1662 11506
rect 6962 11454 6974 11506
rect 7026 11454 7038 11506
rect 11218 11454 11230 11506
rect 11282 11454 11294 11506
rect 14802 11454 14814 11506
rect 14866 11454 14878 11506
rect 17602 11454 17614 11506
rect 17666 11454 17678 11506
rect 25554 11454 25566 11506
rect 25618 11454 25630 11506
rect 28242 11454 28254 11506
rect 28306 11454 28318 11506
rect 5854 11442 5906 11454
rect 10222 11442 10274 11454
rect 28702 11442 28754 11454
rect 36094 11506 36146 11518
rect 36094 11442 36146 11454
rect 37550 11506 37602 11518
rect 42030 11506 42082 11518
rect 47406 11506 47458 11518
rect 38434 11454 38446 11506
rect 38498 11454 38510 11506
rect 38994 11454 39006 11506
rect 39058 11454 39070 11506
rect 46274 11454 46286 11506
rect 46338 11454 46350 11506
rect 48738 11454 48750 11506
rect 48802 11454 48814 11506
rect 49074 11454 49086 11506
rect 49138 11454 49150 11506
rect 53666 11454 53678 11506
rect 53730 11454 53742 11506
rect 55346 11454 55358 11506
rect 55410 11454 55422 11506
rect 37550 11442 37602 11454
rect 42030 11442 42082 11454
rect 47406 11442 47458 11454
rect 5406 11394 5458 11406
rect 1250 11342 1262 11394
rect 1314 11342 1326 11394
rect 4946 11342 4958 11394
rect 5010 11342 5022 11394
rect 5406 11330 5458 11342
rect 5630 11394 5682 11406
rect 5630 11330 5682 11342
rect 5966 11394 6018 11406
rect 8878 11394 8930 11406
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 5966 11330 6018 11342
rect 8878 11330 8930 11342
rect 9550 11394 9602 11406
rect 9550 11330 9602 11342
rect 9774 11394 9826 11406
rect 11902 11394 11954 11406
rect 18734 11394 18786 11406
rect 20862 11394 20914 11406
rect 26798 11394 26850 11406
rect 35870 11394 35922 11406
rect 43486 11394 43538 11406
rect 48526 11394 48578 11406
rect 56030 11394 56082 11406
rect 10546 11342 10558 11394
rect 10610 11342 10622 11394
rect 11106 11342 11118 11394
rect 11170 11342 11182 11394
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 13234 11342 13246 11394
rect 13298 11342 13310 11394
rect 14354 11342 14366 11394
rect 14418 11342 14430 11394
rect 19506 11342 19518 11394
rect 19570 11342 19582 11394
rect 19954 11342 19966 11394
rect 20018 11342 20030 11394
rect 21186 11342 21198 11394
rect 21250 11342 21262 11394
rect 22194 11342 22206 11394
rect 22258 11342 22270 11394
rect 25218 11342 25230 11394
rect 25282 11342 25294 11394
rect 27570 11342 27582 11394
rect 27634 11342 27646 11394
rect 28018 11342 28030 11394
rect 28082 11342 28094 11394
rect 29474 11342 29486 11394
rect 29538 11342 29550 11394
rect 30258 11342 30270 11394
rect 30322 11342 30334 11394
rect 34402 11342 34414 11394
rect 34466 11342 34478 11394
rect 35298 11342 35310 11394
rect 35362 11342 35374 11394
rect 35522 11342 35534 11394
rect 35586 11342 35598 11394
rect 36642 11342 36654 11394
rect 36706 11342 36718 11394
rect 37090 11342 37102 11394
rect 37154 11342 37166 11394
rect 42466 11342 42478 11394
rect 42530 11342 42542 11394
rect 42802 11342 42814 11394
rect 42866 11342 42878 11394
rect 44146 11342 44158 11394
rect 44210 11342 44222 11394
rect 45042 11342 45054 11394
rect 45106 11342 45118 11394
rect 45714 11342 45726 11394
rect 45778 11342 45790 11394
rect 54002 11342 54014 11394
rect 54066 11342 54078 11394
rect 9774 11330 9826 11342
rect 11902 11330 11954 11342
rect 18734 11330 18786 11342
rect 20862 11330 20914 11342
rect 26798 11330 26850 11342
rect 35870 11330 35922 11342
rect 43486 11330 43538 11342
rect 48526 11330 48578 11342
rect 56030 11330 56082 11342
rect 9326 11282 9378 11294
rect 13806 11282 13858 11294
rect 19182 11282 19234 11294
rect 9650 11230 9662 11282
rect 9714 11230 9726 11282
rect 17154 11230 17166 11282
rect 17218 11230 17230 11282
rect 9326 11218 9378 11230
rect 13806 11218 13858 11230
rect 19182 11218 19234 11230
rect 27246 11282 27298 11294
rect 50306 11230 50318 11282
rect 50370 11230 50382 11282
rect 27246 11218 27298 11230
rect 9102 11170 9154 11182
rect 9102 11106 9154 11118
rect 13918 11170 13970 11182
rect 13918 11106 13970 11118
rect 16046 11170 16098 11182
rect 16046 11106 16098 11118
rect 39230 11170 39282 11182
rect 39230 11106 39282 11118
rect 39566 11170 39618 11182
rect 39566 11106 39618 11118
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 10894 10834 10946 10846
rect 10894 10770 10946 10782
rect 22542 10834 22594 10846
rect 22542 10770 22594 10782
rect 36654 10834 36706 10846
rect 36654 10770 36706 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 43150 10834 43202 10846
rect 43150 10770 43202 10782
rect 52334 10834 52386 10846
rect 52334 10770 52386 10782
rect 52670 10834 52722 10846
rect 52670 10770 52722 10782
rect 4398 10722 4450 10734
rect 4398 10658 4450 10670
rect 11454 10722 11506 10734
rect 11454 10658 11506 10670
rect 16382 10722 16434 10734
rect 29262 10722 29314 10734
rect 20962 10670 20974 10722
rect 21026 10670 21038 10722
rect 16382 10658 16434 10670
rect 29262 10658 29314 10670
rect 35646 10722 35698 10734
rect 44270 10722 44322 10734
rect 38210 10670 38222 10722
rect 38274 10670 38286 10722
rect 35646 10658 35698 10670
rect 44270 10658 44322 10670
rect 49534 10722 49586 10734
rect 49534 10658 49586 10670
rect 52782 10722 52834 10734
rect 52782 10658 52834 10670
rect 2942 10610 2994 10622
rect 5518 10610 5570 10622
rect 7198 10610 7250 10622
rect 11342 10610 11394 10622
rect 1362 10558 1374 10610
rect 1426 10558 1438 10610
rect 2146 10558 2158 10610
rect 2210 10558 2222 10610
rect 3602 10558 3614 10610
rect 3666 10558 3678 10610
rect 4050 10558 4062 10610
rect 4114 10558 4126 10610
rect 5954 10558 5966 10610
rect 6018 10558 6030 10610
rect 6290 10558 6302 10610
rect 6354 10558 6366 10610
rect 7634 10558 7646 10610
rect 7698 10558 7710 10610
rect 8530 10558 8542 10610
rect 8594 10558 8606 10610
rect 9202 10558 9214 10610
rect 9266 10558 9278 10610
rect 2942 10546 2994 10558
rect 5518 10546 5570 10558
rect 7198 10546 7250 10558
rect 11342 10546 11394 10558
rect 11566 10610 11618 10622
rect 14590 10610 14642 10622
rect 12898 10558 12910 10610
rect 12962 10558 12974 10610
rect 14018 10558 14030 10610
rect 14082 10558 14094 10610
rect 15250 10558 15262 10610
rect 15314 10558 15326 10610
rect 15698 10558 15710 10610
rect 15762 10558 15774 10610
rect 16706 10558 16718 10610
rect 16770 10558 16782 10610
rect 17266 10570 17278 10622
rect 17330 10570 17342 10622
rect 17838 10610 17890 10622
rect 24446 10610 24498 10622
rect 30942 10610 30994 10622
rect 35758 10610 35810 10622
rect 36766 10610 36818 10622
rect 44158 10610 44210 10622
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 19394 10558 19406 10610
rect 19458 10558 19470 10610
rect 23314 10558 23326 10610
rect 23378 10558 23390 10610
rect 23762 10558 23774 10610
rect 23826 10558 23838 10610
rect 24994 10558 25006 10610
rect 25058 10558 25070 10610
rect 26002 10558 26014 10610
rect 26066 10558 26078 10610
rect 29586 10558 29598 10610
rect 29650 10558 29662 10610
rect 30146 10558 30158 10610
rect 30210 10558 30222 10610
rect 31266 10558 31278 10610
rect 31330 10558 31342 10610
rect 32274 10558 32286 10610
rect 32338 10558 32350 10610
rect 32946 10558 32958 10610
rect 33010 10558 33022 10610
rect 36306 10558 36318 10610
rect 36370 10558 36382 10610
rect 41570 10558 41582 10610
rect 41634 10558 41646 10610
rect 11566 10546 11618 10558
rect 14590 10546 14642 10558
rect 17838 10546 17890 10558
rect 24446 10546 24498 10558
rect 30942 10546 30994 10558
rect 35758 10546 35810 10558
rect 36766 10546 36818 10558
rect 44158 10546 44210 10558
rect 47742 10610 47794 10622
rect 47742 10546 47794 10558
rect 48414 10610 48466 10622
rect 48414 10546 48466 10558
rect 48750 10610 48802 10622
rect 48750 10546 48802 10558
rect 48974 10610 49026 10622
rect 50990 10610 51042 10622
rect 56030 10610 56082 10622
rect 49298 10558 49310 10610
rect 49362 10558 49374 10610
rect 50418 10558 50430 10610
rect 50482 10558 50494 10610
rect 51986 10558 51998 10610
rect 52050 10558 52062 10610
rect 53442 10558 53454 10610
rect 53506 10558 53518 10610
rect 48974 10546 49026 10558
rect 50990 10546 51042 10558
rect 56030 10546 56082 10558
rect 4958 10498 5010 10510
rect 4958 10434 5010 10446
rect 6974 10498 7026 10510
rect 6974 10434 7026 10446
rect 16046 10498 16098 10510
rect 16046 10434 16098 10446
rect 22990 10498 23042 10510
rect 22990 10434 23042 10446
rect 37102 10498 37154 10510
rect 44382 10498 44434 10510
rect 38658 10446 38670 10498
rect 38722 10446 38734 10498
rect 42018 10446 42030 10498
rect 42082 10446 42094 10498
rect 37102 10434 37154 10446
rect 44382 10434 44434 10446
rect 47966 10498 48018 10510
rect 47966 10434 48018 10446
rect 48078 10498 48130 10510
rect 48078 10434 48130 10446
rect 48526 10498 48578 10510
rect 50194 10446 50206 10498
rect 50258 10446 50270 10498
rect 50642 10446 50654 10498
rect 50706 10446 50718 10498
rect 53778 10446 53790 10498
rect 53842 10446 53854 10498
rect 56354 10446 56366 10498
rect 56418 10446 56430 10498
rect 48526 10434 48578 10446
rect 5070 10386 5122 10398
rect 3378 10334 3390 10386
rect 3442 10334 3454 10386
rect 5070 10322 5122 10334
rect 5294 10386 5346 10398
rect 11790 10386 11842 10398
rect 34638 10386 34690 10398
rect 44606 10386 44658 10398
rect 6514 10334 6526 10386
rect 6578 10334 6590 10386
rect 9762 10334 9774 10386
rect 9826 10334 9838 10386
rect 15026 10334 15038 10386
rect 15090 10334 15102 10386
rect 17378 10334 17390 10386
rect 17442 10334 17454 10386
rect 21410 10334 21422 10386
rect 21474 10334 21486 10386
rect 23986 10334 23998 10386
rect 24050 10334 24062 10386
rect 30258 10334 30270 10386
rect 30322 10334 30334 10386
rect 33506 10334 33518 10386
rect 33570 10334 33582 10386
rect 36642 10334 36654 10386
rect 36706 10334 36718 10386
rect 5294 10322 5346 10334
rect 11790 10322 11842 10334
rect 34638 10322 34690 10334
rect 44606 10322 44658 10334
rect 49422 10386 49474 10398
rect 49422 10322 49474 10334
rect 49646 10386 49698 10398
rect 49646 10322 49698 10334
rect 51326 10386 51378 10398
rect 51326 10322 51378 10334
rect 52222 10386 52274 10398
rect 52222 10322 52274 10334
rect 55022 10386 55074 10398
rect 55022 10322 55074 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 12126 10050 12178 10062
rect 8866 9998 8878 10050
rect 8930 9998 8942 10050
rect 10994 9998 11006 10050
rect 11058 9998 11070 10050
rect 12126 9986 12178 9998
rect 14926 10050 14978 10062
rect 14926 9986 14978 9998
rect 15598 10050 15650 10062
rect 15598 9986 15650 9998
rect 15710 10050 15762 10062
rect 15710 9986 15762 9998
rect 20302 10050 20354 10062
rect 23886 10050 23938 10062
rect 22754 9998 22766 10050
rect 22818 9998 22830 10050
rect 20302 9986 20354 9998
rect 23886 9986 23938 9998
rect 29038 10050 29090 10062
rect 29038 9986 29090 9998
rect 31278 10050 31330 10062
rect 31278 9986 31330 9998
rect 36206 10050 36258 10062
rect 42590 10050 42642 10062
rect 37314 9998 37326 10050
rect 37378 9998 37390 10050
rect 41458 9998 41470 10050
rect 41522 9998 41534 10050
rect 36206 9986 36258 9998
rect 42590 9986 42642 9998
rect 43150 10050 43202 10062
rect 43150 9986 43202 9998
rect 47294 10050 47346 10062
rect 47294 9986 47346 9998
rect 47406 10050 47458 10062
rect 47406 9986 47458 9998
rect 51662 10050 51714 10062
rect 56354 9998 56366 10050
rect 56418 9998 56430 10050
rect 51662 9986 51714 9998
rect 4734 9938 4786 9950
rect 3714 9886 3726 9938
rect 3778 9886 3790 9938
rect 4734 9874 4786 9886
rect 6862 9938 6914 9950
rect 8318 9938 8370 9950
rect 7298 9886 7310 9938
rect 7362 9886 7374 9938
rect 6862 9874 6914 9886
rect 8318 9874 8370 9886
rect 9886 9938 9938 9950
rect 9886 9874 9938 9886
rect 12014 9938 12066 9950
rect 12014 9874 12066 9886
rect 12238 9938 12290 9950
rect 12238 9874 12290 9886
rect 12686 9938 12738 9950
rect 12686 9874 12738 9886
rect 12798 9938 12850 9950
rect 16158 9938 16210 9950
rect 13794 9886 13806 9938
rect 13858 9886 13870 9938
rect 12798 9874 12850 9886
rect 16158 9874 16210 9886
rect 17726 9938 17778 9950
rect 36094 9938 36146 9950
rect 19170 9886 19182 9938
rect 19234 9886 19246 9938
rect 27906 9886 27918 9938
rect 27970 9886 27982 9938
rect 30034 9886 30046 9938
rect 30098 9886 30110 9938
rect 33394 9886 33406 9938
rect 33458 9886 33470 9938
rect 44370 9886 44382 9938
rect 44434 9886 44446 9938
rect 48178 9886 48190 9938
rect 48242 9886 48254 9938
rect 48738 9886 48750 9938
rect 48802 9886 48814 9938
rect 51090 9886 51102 9938
rect 51154 9886 51166 9938
rect 52770 9886 52782 9938
rect 52834 9886 52846 9938
rect 54002 9886 54014 9938
rect 54066 9886 54078 9938
rect 17726 9874 17778 9886
rect 36094 9874 36146 9886
rect 3054 9826 3106 9838
rect 9214 9826 9266 9838
rect 1698 9774 1710 9826
rect 1762 9774 1774 9826
rect 2482 9774 2494 9826
rect 2546 9774 2558 9826
rect 3938 9774 3950 9826
rect 4002 9774 4014 9826
rect 4386 9774 4398 9826
rect 4450 9774 4462 9826
rect 5282 9774 5294 9826
rect 5346 9774 5358 9826
rect 6290 9774 6302 9826
rect 6354 9774 6366 9826
rect 7410 9774 7422 9826
rect 7474 9774 7486 9826
rect 7858 9774 7870 9826
rect 7922 9774 7934 9826
rect 3054 9762 3106 9774
rect 9214 9762 9266 9774
rect 15934 9826 15986 9838
rect 15934 9762 15986 9774
rect 16606 9826 16658 9838
rect 16606 9762 16658 9774
rect 16830 9826 16882 9838
rect 16830 9762 16882 9774
rect 16942 9826 16994 9838
rect 16942 9762 16994 9774
rect 17166 9826 17218 9838
rect 17166 9762 17218 9774
rect 17502 9826 17554 9838
rect 17502 9762 17554 9774
rect 17838 9826 17890 9838
rect 17838 9762 17890 9774
rect 18062 9826 18114 9838
rect 34078 9826 34130 9838
rect 48974 9826 49026 9838
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 27458 9774 27470 9826
rect 27522 9774 27534 9826
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 32722 9774 32734 9826
rect 32786 9774 32798 9826
rect 33170 9774 33182 9826
rect 33234 9774 33246 9826
rect 34626 9774 34638 9826
rect 34690 9774 34702 9826
rect 35522 9774 35534 9826
rect 35586 9774 35598 9826
rect 36866 9774 36878 9826
rect 36930 9774 36942 9826
rect 44818 9774 44830 9826
rect 44882 9774 44894 9826
rect 18062 9762 18114 9774
rect 34078 9762 34130 9774
rect 48974 9762 49026 9774
rect 49310 9826 49362 9838
rect 51998 9826 52050 9838
rect 50754 9774 50766 9826
rect 50818 9774 50830 9826
rect 52658 9774 52670 9826
rect 52722 9774 52734 9826
rect 56130 9774 56142 9826
rect 56194 9774 56206 9826
rect 49310 9762 49362 9774
rect 51998 9762 52050 9774
rect 9438 9714 9490 9726
rect 32398 9714 32450 9726
rect 11442 9662 11454 9714
rect 11506 9662 11518 9714
rect 13346 9662 13358 9714
rect 13410 9662 13422 9714
rect 15698 9662 15710 9714
rect 15762 9662 15774 9714
rect 18722 9662 18734 9714
rect 18786 9662 18798 9714
rect 9438 9650 9490 9662
rect 32398 9650 32450 9662
rect 40350 9714 40402 9726
rect 41010 9662 41022 9714
rect 41074 9662 41086 9714
rect 53666 9662 53678 9714
rect 53730 9662 53742 9714
rect 40350 9650 40402 9662
rect 36318 9602 36370 9614
rect 36318 9538 36370 9550
rect 38446 9602 38498 9614
rect 38446 9538 38498 9550
rect 40462 9602 40514 9614
rect 40462 9538 40514 9550
rect 47182 9602 47234 9614
rect 47182 9538 47234 9550
rect 49982 9602 50034 9614
rect 49982 9538 50034 9550
rect 50318 9602 50370 9614
rect 50318 9538 50370 9550
rect 55246 9602 55298 9614
rect 55246 9538 55298 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 4286 9266 4338 9278
rect 4286 9202 4338 9214
rect 6750 9266 6802 9278
rect 6750 9202 6802 9214
rect 11006 9266 11058 9278
rect 11006 9202 11058 9214
rect 11454 9266 11506 9278
rect 11454 9202 11506 9214
rect 20750 9266 20802 9278
rect 20750 9202 20802 9214
rect 40910 9266 40962 9278
rect 40910 9202 40962 9214
rect 44606 9266 44658 9278
rect 44606 9202 44658 9214
rect 50206 9266 50258 9278
rect 50206 9202 50258 9214
rect 50542 9266 50594 9278
rect 50542 9202 50594 9214
rect 15262 9154 15314 9166
rect 5170 9102 5182 9154
rect 5234 9102 5246 9154
rect 9426 9102 9438 9154
rect 9490 9102 9502 9154
rect 13122 9102 13134 9154
rect 13186 9102 13198 9154
rect 15262 9090 15314 9102
rect 37214 9154 37266 9166
rect 37214 9090 37266 9102
rect 43486 9154 43538 9166
rect 43486 9090 43538 9102
rect 44270 9154 44322 9166
rect 44270 9090 44322 9102
rect 46174 9154 46226 9166
rect 46174 9090 46226 9102
rect 7310 9042 7362 9054
rect 11566 9042 11618 9054
rect 14702 9042 14754 9054
rect 16718 9042 16770 9054
rect 33742 9042 33794 9054
rect 38670 9042 38722 9054
rect 43598 9042 43650 9054
rect 52670 9042 52722 9054
rect 1250 8990 1262 9042
rect 1314 8990 1326 9042
rect 1922 8990 1934 9042
rect 1986 8990 1998 9042
rect 2706 8990 2718 9042
rect 2770 8990 2782 9042
rect 7634 8990 7646 9042
rect 7698 8990 7710 9042
rect 7858 8990 7870 9042
rect 7922 8990 7934 9042
rect 11778 8990 11790 9042
rect 11842 8990 11854 9042
rect 15586 8990 15598 9042
rect 15650 8990 15662 9042
rect 16146 8990 16158 9042
rect 16210 8990 16222 9042
rect 17266 8990 17278 9042
rect 17330 8990 17342 9042
rect 17490 8990 17502 9042
rect 17554 8990 17566 9042
rect 18274 8990 18286 9042
rect 18338 8990 18350 9042
rect 22306 8990 22318 9042
rect 22370 8990 22382 9042
rect 23874 8990 23886 9042
rect 23938 8990 23950 9042
rect 32386 8990 32398 9042
rect 32450 8990 32462 9042
rect 32834 8990 32846 9042
rect 32898 8990 32910 9042
rect 34066 8990 34078 9042
rect 34130 8990 34142 9042
rect 35074 8990 35086 9042
rect 35138 8990 35150 9042
rect 36754 8990 36766 9042
rect 36818 8990 36830 9042
rect 37650 8990 37662 9042
rect 37714 8990 37726 9042
rect 37986 8990 37998 9042
rect 38050 8990 38062 9042
rect 39442 8990 39454 9042
rect 39506 8990 39518 9042
rect 40226 8990 40238 9042
rect 40290 8990 40302 9042
rect 42578 8990 42590 9042
rect 42642 8990 42654 9042
rect 46498 8990 46510 9042
rect 46562 8990 46574 9042
rect 46946 8990 46958 9042
rect 47010 8990 47022 9042
rect 47730 8990 47742 9042
rect 47794 8990 47806 9042
rect 48402 8990 48414 9042
rect 48466 8990 48478 9042
rect 49186 8990 49198 9042
rect 49250 8990 49262 9042
rect 53218 8990 53230 9042
rect 53282 8990 53294 9042
rect 55458 8990 55470 9042
rect 55522 8990 55534 9042
rect 7310 8978 7362 8990
rect 11566 8978 11618 8990
rect 14702 8978 14754 8990
rect 16718 8978 16770 8990
rect 33742 8978 33794 8990
rect 38670 8978 38722 8990
rect 43598 8978 43650 8990
rect 52670 8978 52722 8990
rect 7198 8930 7250 8942
rect 8654 8930 8706 8942
rect 12238 8930 12290 8942
rect 32062 8930 32114 8942
rect 56030 8930 56082 8942
rect 1026 8878 1038 8930
rect 1090 8878 1102 8930
rect 1698 8878 1710 8930
rect 1762 8878 1774 8930
rect 3042 8878 3054 8930
rect 3106 8878 3118 8930
rect 5618 8878 5630 8930
rect 5682 8878 5694 8930
rect 8306 8878 8318 8930
rect 8370 8878 8382 8930
rect 9874 8878 9886 8930
rect 9938 8878 9950 8930
rect 16258 8878 16270 8930
rect 16322 8878 16334 8930
rect 38210 8878 38222 8930
rect 38274 8878 38286 8930
rect 42130 8878 42142 8930
rect 42194 8878 42206 8930
rect 44818 8878 44830 8930
rect 44882 8878 44894 8930
rect 45154 8878 45166 8930
rect 45218 8878 45230 8930
rect 47170 8878 47182 8930
rect 47234 8878 47246 8930
rect 50754 8878 50766 8930
rect 50818 8878 50830 8930
rect 51090 8878 51102 8930
rect 51154 8878 51166 8930
rect 52322 8878 52334 8930
rect 52386 8878 52398 8930
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 55234 8878 55246 8930
rect 55298 8878 55310 8930
rect 56354 8878 56366 8930
rect 56418 8878 56430 8930
rect 7198 8866 7250 8878
rect 8654 8866 8706 8878
rect 12238 8866 12290 8878
rect 32062 8866 32114 8878
rect 56030 8866 56082 8878
rect 7422 8818 7474 8830
rect 7422 8754 7474 8766
rect 12126 8818 12178 8830
rect 25454 8818 25506 8830
rect 43150 8818 43202 8830
rect 13570 8766 13582 8818
rect 13634 8766 13646 8818
rect 21858 8766 21870 8818
rect 21922 8766 21934 8818
rect 24322 8766 24334 8818
rect 24386 8766 24398 8818
rect 33058 8766 33070 8818
rect 33122 8766 33134 8818
rect 36530 8766 36542 8818
rect 36594 8766 36606 8818
rect 12126 8754 12178 8766
rect 25454 8754 25506 8766
rect 43150 8754 43202 8766
rect 43374 8818 43426 8830
rect 43374 8754 43426 8766
rect 54798 8818 54850 8830
rect 54798 8754 54850 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 3950 8482 4002 8494
rect 2034 8430 2046 8482
rect 2098 8430 2110 8482
rect 3950 8418 4002 8430
rect 16606 8482 16658 8494
rect 16606 8418 16658 8430
rect 16830 8482 16882 8494
rect 16830 8418 16882 8430
rect 44046 8482 44098 8494
rect 44046 8418 44098 8430
rect 46510 8482 46562 8494
rect 46510 8418 46562 8430
rect 48302 8482 48354 8494
rect 48302 8418 48354 8430
rect 49534 8482 49586 8494
rect 49534 8418 49586 8430
rect 51774 8482 51826 8494
rect 51774 8418 51826 8430
rect 56366 8482 56418 8494
rect 56366 8418 56418 8430
rect 8318 8370 8370 8382
rect 12574 8370 12626 8382
rect 16942 8370 16994 8382
rect 38334 8370 38386 8382
rect 3602 8318 3614 8370
rect 3666 8318 3678 8370
rect 4274 8318 4286 8370
rect 4338 8318 4350 8370
rect 7298 8318 7310 8370
rect 7362 8318 7374 8370
rect 11554 8318 11566 8370
rect 11618 8318 11630 8370
rect 15138 8318 15150 8370
rect 15202 8318 15214 8370
rect 17938 8318 17950 8370
rect 18002 8318 18014 8370
rect 20514 8318 20526 8370
rect 20578 8318 20590 8370
rect 26674 8318 26686 8370
rect 26738 8318 26750 8370
rect 30594 8318 30606 8370
rect 30658 8318 30670 8370
rect 33394 8318 33406 8370
rect 33458 8318 33470 8370
rect 37202 8318 37214 8370
rect 37266 8318 37278 8370
rect 8318 8306 8370 8318
rect 12574 8306 12626 8318
rect 16942 8306 16994 8318
rect 38334 8306 38386 8318
rect 40798 8370 40850 8382
rect 48638 8370 48690 8382
rect 54126 8370 54178 8382
rect 42466 8318 42478 8370
rect 42530 8318 42542 8370
rect 45266 8318 45278 8370
rect 45330 8318 45342 8370
rect 50642 8318 50654 8370
rect 50706 8318 50718 8370
rect 52882 8318 52894 8370
rect 52946 8318 52958 8370
rect 55010 8318 55022 8370
rect 55074 8318 55086 8370
rect 56018 8318 56030 8370
rect 56082 8318 56094 8370
rect 40798 8306 40850 8318
rect 48638 8306 48690 8318
rect 54126 8306 54178 8318
rect 6862 8258 6914 8270
rect 10894 8258 10946 8270
rect 13246 8263 13298 8275
rect 4498 8206 4510 8258
rect 4562 8206 4574 8258
rect 5170 8206 5182 8258
rect 5234 8206 5246 8258
rect 6290 8206 6302 8258
rect 6354 8206 6366 8258
rect 7410 8206 7422 8258
rect 7474 8206 7486 8258
rect 7858 8206 7870 8258
rect 7922 8206 7934 8258
rect 9538 8206 9550 8258
rect 9602 8206 9614 8258
rect 10322 8206 10334 8258
rect 10386 8206 10398 8258
rect 11778 8206 11790 8258
rect 11842 8206 11854 8258
rect 12114 8206 12126 8258
rect 12178 8206 12190 8258
rect 14702 8258 14754 8270
rect 19070 8258 19122 8270
rect 20974 8258 21026 8270
rect 27134 8258 27186 8270
rect 33854 8258 33906 8270
rect 40686 8258 40738 8270
rect 6862 8194 6914 8206
rect 10894 8194 10946 8206
rect 13246 8199 13298 8211
rect 13906 8206 13918 8258
rect 13970 8206 13982 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 15810 8206 15822 8258
rect 15874 8206 15886 8258
rect 17378 8206 17390 8258
rect 17442 8206 17454 8258
rect 19842 8206 19854 8258
rect 19906 8206 19918 8258
rect 20290 8206 20302 8258
rect 20354 8206 20366 8258
rect 21522 8206 21534 8258
rect 21586 8206 21598 8258
rect 22530 8206 22542 8258
rect 22594 8206 22606 8258
rect 26002 8206 26014 8258
rect 26066 8206 26078 8258
rect 26450 8206 26462 8258
rect 26514 8206 26526 8258
rect 27906 8206 27918 8258
rect 27970 8206 27982 8258
rect 28802 8206 28814 8258
rect 28866 8206 28878 8258
rect 32722 8206 32734 8258
rect 32786 8206 32798 8258
rect 33170 8206 33182 8258
rect 33234 8206 33246 8258
rect 34402 8206 34414 8258
rect 34466 8206 34478 8258
rect 35410 8206 35422 8258
rect 35474 8206 35486 8258
rect 36754 8206 36766 8258
rect 36818 8206 36830 8258
rect 14702 8194 14754 8206
rect 19070 8194 19122 8206
rect 20974 8194 21026 8206
rect 27134 8194 27186 8206
rect 33854 8194 33906 8206
rect 40686 8194 40738 8206
rect 41022 8258 41074 8270
rect 44270 8258 44322 8270
rect 47966 8258 48018 8270
rect 43474 8206 43486 8258
rect 43538 8206 43550 8258
rect 43810 8206 43822 8258
rect 43874 8206 43886 8258
rect 44818 8206 44830 8258
rect 44882 8206 44894 8258
rect 41022 8194 41074 8206
rect 44270 8194 44322 8206
rect 47966 8194 48018 8206
rect 48302 8258 48354 8270
rect 48302 8194 48354 8206
rect 54462 8258 54514 8270
rect 54898 8206 54910 8258
rect 54962 8206 54974 8258
rect 54462 8194 54514 8206
rect 8990 8146 9042 8158
rect 1586 8094 1598 8146
rect 1650 8094 1662 8146
rect 8990 8082 9042 8094
rect 16158 8146 16210 8158
rect 19518 8146 19570 8158
rect 17490 8094 17502 8146
rect 17554 8094 17566 8146
rect 16158 8082 16210 8094
rect 19518 8082 19570 8094
rect 25678 8146 25730 8158
rect 32398 8146 32450 8158
rect 30146 8094 30158 8146
rect 30210 8094 30222 8146
rect 42914 8094 42926 8146
rect 42978 8094 42990 8146
rect 43922 8094 43934 8146
rect 43986 8094 43998 8146
rect 51090 8094 51102 8146
rect 51154 8094 51166 8146
rect 53330 8094 53342 8146
rect 53394 8094 53406 8146
rect 25678 8082 25730 8094
rect 32398 8082 32450 8094
rect 3166 8034 3218 8046
rect 3166 7970 3218 7982
rect 8878 8034 8930 8046
rect 8878 7970 8930 7982
rect 31726 8034 31778 8046
rect 31726 7970 31778 7982
rect 41358 8034 41410 8046
rect 41358 7970 41410 7982
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 3166 7698 3218 7710
rect 3166 7634 3218 7646
rect 4958 7698 5010 7710
rect 4958 7634 5010 7646
rect 31838 7698 31890 7710
rect 31838 7634 31890 7646
rect 43374 7698 43426 7710
rect 43374 7634 43426 7646
rect 45950 7698 46002 7710
rect 45950 7634 46002 7646
rect 48190 7698 48242 7710
rect 48190 7634 48242 7646
rect 48750 7698 48802 7710
rect 48750 7634 48802 7646
rect 8654 7586 8706 7598
rect 1586 7534 1598 7586
rect 1650 7534 1662 7586
rect 8654 7522 8706 7534
rect 12238 7586 12290 7598
rect 12238 7522 12290 7534
rect 20638 7586 20690 7598
rect 20638 7522 20690 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 32510 7586 32562 7598
rect 32510 7522 32562 7534
rect 37886 7586 37938 7598
rect 52210 7534 52222 7586
rect 52274 7534 52286 7586
rect 37886 7522 37938 7534
rect 3950 7474 4002 7486
rect 3950 7410 4002 7422
rect 5070 7474 5122 7486
rect 6974 7474 7026 7486
rect 13134 7474 13186 7486
rect 5618 7422 5630 7474
rect 5682 7422 5694 7474
rect 6402 7422 6414 7474
rect 6466 7422 6478 7474
rect 7746 7422 7758 7474
rect 7810 7422 7822 7474
rect 8194 7422 8206 7474
rect 8258 7422 8270 7474
rect 9090 7422 9102 7474
rect 9154 7422 9166 7474
rect 9986 7422 9998 7474
rect 10050 7422 10062 7474
rect 10658 7422 10670 7474
rect 10722 7422 10734 7474
rect 11330 7422 11342 7474
rect 11394 7422 11406 7474
rect 11890 7422 11902 7474
rect 11954 7422 11966 7474
rect 5070 7410 5122 7422
rect 6974 7410 7026 7422
rect 13134 7410 13186 7422
rect 14926 7474 14978 7486
rect 22318 7474 22370 7486
rect 26126 7474 26178 7486
rect 34190 7474 34242 7486
rect 39342 7474 39394 7486
rect 51438 7474 51490 7486
rect 16258 7422 16270 7474
rect 16322 7422 16334 7474
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 17938 7422 17950 7474
rect 18002 7422 18014 7474
rect 18946 7422 18958 7474
rect 19010 7422 19022 7474
rect 20962 7422 20974 7474
rect 21026 7422 21038 7474
rect 21410 7422 21422 7474
rect 21474 7422 21486 7474
rect 22642 7422 22654 7474
rect 22706 7422 22718 7474
rect 23650 7422 23662 7474
rect 23714 7422 23726 7474
rect 24994 7422 25006 7474
rect 25058 7422 25070 7474
rect 25442 7422 25454 7474
rect 25506 7422 25518 7474
rect 26786 7422 26798 7474
rect 26850 7422 26862 7474
rect 27794 7422 27806 7474
rect 27858 7422 27870 7474
rect 30258 7422 30270 7474
rect 30322 7422 30334 7474
rect 32834 7422 32846 7474
rect 32898 7422 32910 7474
rect 33282 7422 33294 7474
rect 33346 7422 33358 7474
rect 34738 7422 34750 7474
rect 34802 7422 34814 7474
rect 35634 7422 35646 7474
rect 35698 7422 35710 7474
rect 38210 7422 38222 7474
rect 38274 7422 38286 7474
rect 38770 7422 38782 7474
rect 38834 7422 38846 7474
rect 39890 7422 39902 7474
rect 39954 7422 39966 7474
rect 40898 7422 40910 7474
rect 40962 7422 40974 7474
rect 41794 7422 41806 7474
rect 41858 7422 41870 7474
rect 44258 7422 44270 7474
rect 44322 7422 44334 7474
rect 46498 7422 46510 7474
rect 46562 7422 46574 7474
rect 50306 7422 50318 7474
rect 50370 7422 50382 7474
rect 54450 7422 54462 7474
rect 54514 7422 54526 7474
rect 14926 7410 14978 7422
rect 22318 7410 22370 7422
rect 26126 7410 26178 7422
rect 34190 7410 34242 7422
rect 39342 7410 39394 7422
rect 51438 7410 51490 7422
rect 4286 7362 4338 7374
rect 2034 7310 2046 7362
rect 2098 7310 2110 7362
rect 3602 7310 3614 7362
rect 3666 7310 3678 7362
rect 4286 7298 4338 7310
rect 4398 7362 4450 7374
rect 14254 7362 14306 7374
rect 12786 7310 12798 7362
rect 12850 7310 12862 7362
rect 13458 7310 13470 7362
rect 13522 7310 13534 7362
rect 4398 7298 4450 7310
rect 14254 7298 14306 7310
rect 14366 7362 14418 7374
rect 14366 7298 14418 7310
rect 14814 7362 14866 7374
rect 14814 7298 14866 7310
rect 15934 7362 15986 7374
rect 15934 7298 15986 7310
rect 17390 7362 17442 7374
rect 30706 7310 30718 7362
rect 30770 7310 30782 7362
rect 38882 7310 38894 7362
rect 38946 7310 38958 7362
rect 42130 7310 42142 7362
rect 42194 7310 42206 7362
rect 44818 7310 44830 7362
rect 44882 7310 44894 7362
rect 46946 7310 46958 7362
rect 47010 7310 47022 7362
rect 49858 7310 49870 7362
rect 49922 7310 49934 7362
rect 52546 7310 52558 7362
rect 52610 7310 52622 7362
rect 54786 7310 54798 7362
rect 54850 7310 54862 7362
rect 17390 7298 17442 7310
rect 13806 7250 13858 7262
rect 7634 7198 7646 7250
rect 7698 7198 7710 7250
rect 11218 7198 11230 7250
rect 11282 7198 11294 7250
rect 13806 7186 13858 7198
rect 14030 7250 14082 7262
rect 14030 7186 14082 7198
rect 14590 7250 14642 7262
rect 53790 7250 53842 7262
rect 16930 7198 16942 7250
rect 16994 7198 17006 7250
rect 21634 7198 21646 7250
rect 21698 7198 21710 7250
rect 25666 7198 25678 7250
rect 25730 7198 25742 7250
rect 33506 7198 33518 7250
rect 33570 7198 33582 7250
rect 51090 7198 51102 7250
rect 51154 7198 51166 7250
rect 14590 7186 14642 7198
rect 53790 7186 53842 7198
rect 56030 7250 56082 7262
rect 56030 7186 56082 7198
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 9326 6914 9378 6926
rect 3826 6862 3838 6914
rect 3890 6862 3902 6914
rect 9326 6850 9378 6862
rect 14478 6914 14530 6926
rect 14478 6850 14530 6862
rect 15822 6914 15874 6926
rect 15822 6850 15874 6862
rect 35422 6914 35474 6926
rect 35422 6850 35474 6862
rect 46174 6914 46226 6926
rect 46174 6850 46226 6862
rect 53118 6914 53170 6926
rect 56254 6914 56306 6926
rect 54114 6862 54126 6914
rect 54178 6862 54190 6914
rect 53118 6850 53170 6862
rect 56254 6850 56306 6862
rect 4398 6802 4450 6814
rect 8318 6802 8370 6814
rect 1922 6750 1934 6802
rect 1986 6750 1998 6802
rect 7298 6750 7310 6802
rect 7362 6750 7374 6802
rect 4398 6738 4450 6750
rect 8318 6738 8370 6750
rect 9102 6802 9154 6814
rect 9102 6738 9154 6750
rect 10110 6802 10162 6814
rect 14590 6802 14642 6814
rect 11778 6750 11790 6802
rect 11842 6750 11854 6802
rect 10110 6738 10162 6750
rect 14590 6738 14642 6750
rect 14926 6802 14978 6814
rect 14926 6738 14978 6750
rect 15038 6802 15090 6814
rect 15038 6738 15090 6750
rect 15262 6802 15314 6814
rect 15262 6738 15314 6750
rect 15934 6802 15986 6814
rect 25566 6802 25618 6814
rect 33070 6802 33122 6814
rect 16706 6750 16718 6802
rect 16770 6750 16782 6802
rect 18050 6750 18062 6802
rect 18114 6750 18126 6802
rect 21858 6750 21870 6802
rect 21922 6750 21934 6802
rect 23650 6750 23662 6802
rect 23714 6750 23726 6802
rect 24546 6750 24558 6802
rect 24610 6750 24622 6802
rect 27234 6750 27246 6802
rect 27298 6750 27310 6802
rect 30482 6750 30494 6802
rect 30546 6750 30558 6802
rect 15934 6738 15986 6750
rect 25566 6738 25618 6750
rect 33070 6738 33122 6750
rect 34414 6802 34466 6814
rect 35646 6802 35698 6814
rect 34738 6750 34750 6802
rect 34802 6750 34814 6802
rect 34414 6738 34466 6750
rect 35646 6738 35698 6750
rect 36430 6802 36482 6814
rect 46286 6802 46338 6814
rect 38434 6750 38446 6802
rect 38498 6750 38510 6802
rect 41234 6750 41246 6802
rect 41298 6750 41310 6802
rect 44370 6750 44382 6802
rect 44434 6750 44446 6802
rect 46610 6750 46622 6802
rect 46674 6750 46686 6802
rect 50530 6750 50542 6802
rect 50594 6750 50606 6802
rect 52770 6750 52782 6802
rect 52834 6750 52846 6802
rect 55906 6750 55918 6802
rect 55970 6750 55982 6802
rect 36430 6738 36482 6750
rect 46286 6738 46338 6750
rect 3054 6690 3106 6702
rect 1474 6638 1486 6690
rect 1538 6638 1550 6690
rect 3054 6626 3106 6638
rect 3502 6690 3554 6702
rect 3502 6626 3554 6638
rect 4286 6690 4338 6702
rect 4286 6626 4338 6638
rect 4622 6690 4674 6702
rect 4622 6626 4674 6638
rect 4846 6690 4898 6702
rect 6638 6690 6690 6702
rect 9214 6690 9266 6702
rect 5282 6638 5294 6690
rect 5346 6638 5358 6690
rect 6178 6638 6190 6690
rect 6242 6638 6254 6690
rect 7522 6638 7534 6690
rect 7586 6638 7598 6690
rect 7970 6638 7982 6690
rect 8034 6638 8046 6690
rect 8866 6638 8878 6690
rect 8930 6638 8942 6690
rect 4846 6626 4898 6638
rect 6638 6626 6690 6638
rect 9214 6626 9266 6638
rect 9438 6690 9490 6702
rect 9438 6626 9490 6638
rect 9998 6690 10050 6702
rect 9998 6626 10050 6638
rect 10558 6690 10610 6702
rect 14254 6690 14306 6702
rect 15710 6690 15762 6702
rect 17054 6690 17106 6702
rect 19182 6690 19234 6702
rect 21198 6690 21250 6702
rect 22878 6690 22930 6702
rect 11106 6638 11118 6690
rect 11170 6638 11182 6690
rect 11554 6638 11566 6690
rect 11618 6638 11630 6690
rect 12338 6638 12350 6690
rect 12402 6638 12414 6690
rect 12786 6638 12798 6690
rect 12850 6638 12862 6690
rect 13794 6638 13806 6690
rect 13858 6638 13870 6690
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 16146 6638 16158 6690
rect 16210 6638 16222 6690
rect 17490 6638 17502 6690
rect 17554 6638 17566 6690
rect 19730 6638 19742 6690
rect 19794 6638 19806 6690
rect 20850 6638 20862 6690
rect 20914 6638 20926 6690
rect 21970 6638 21982 6690
rect 22034 6638 22046 6690
rect 22418 6638 22430 6690
rect 22482 6638 22494 6690
rect 10558 6626 10610 6638
rect 14254 6626 14306 6638
rect 15710 6626 15762 6638
rect 17054 6626 17106 6638
rect 19182 6626 19234 6638
rect 21198 6626 21250 6638
rect 22878 6626 22930 6638
rect 23998 6690 24050 6702
rect 23998 6626 24050 6638
rect 24894 6690 24946 6702
rect 33294 6690 33346 6702
rect 25890 6638 25902 6690
rect 25954 6638 25966 6690
rect 26674 6638 26686 6690
rect 26738 6638 26750 6690
rect 27122 6638 27134 6690
rect 27186 6638 27198 6690
rect 27794 6638 27806 6690
rect 27858 6638 27870 6690
rect 28466 6638 28478 6690
rect 28530 6638 28542 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 24894 6626 24946 6638
rect 33294 6626 33346 6638
rect 34974 6690 35026 6702
rect 34974 6626 35026 6638
rect 35534 6690 35586 6702
rect 39566 6690 39618 6702
rect 41694 6690 41746 6702
rect 46062 6690 46114 6702
rect 35970 6638 35982 6690
rect 36034 6638 36046 6690
rect 40562 6638 40574 6690
rect 40626 6638 40638 6690
rect 41010 6638 41022 6690
rect 41074 6638 41086 6690
rect 42354 6638 42366 6690
rect 42418 6638 42430 6690
rect 43250 6638 43262 6690
rect 43314 6638 43326 6690
rect 46498 6638 46510 6690
rect 46562 6638 46574 6690
rect 50194 6638 50206 6690
rect 50258 6638 50270 6690
rect 35534 6626 35586 6638
rect 39566 6626 39618 6638
rect 41694 6626 41746 6638
rect 46062 6626 46114 6638
rect 10334 6578 10386 6590
rect 10334 6514 10386 6526
rect 10782 6578 10834 6590
rect 23438 6578 23490 6590
rect 15922 6526 15934 6578
rect 15986 6526 15998 6578
rect 10782 6514 10834 6526
rect 23438 6514 23490 6526
rect 26238 6578 26290 6590
rect 32510 6578 32562 6590
rect 30146 6526 30158 6578
rect 30210 6526 30222 6578
rect 26238 6514 26290 6526
rect 32510 6514 32562 6526
rect 33182 6578 33234 6590
rect 33182 6514 33234 6526
rect 33518 6578 33570 6590
rect 33518 6514 33570 6526
rect 34190 6578 34242 6590
rect 40238 6578 40290 6590
rect 35074 6526 35086 6578
rect 35138 6526 35150 6578
rect 37986 6526 37998 6578
rect 38050 6526 38062 6578
rect 44034 6526 44046 6578
rect 44098 6526 44110 6578
rect 53666 6526 53678 6578
rect 53730 6526 53742 6578
rect 34190 6514 34242 6526
rect 40238 6514 40290 6526
rect 25902 6466 25954 6478
rect 25902 6402 25954 6414
rect 31726 6466 31778 6478
rect 31726 6402 31778 6414
rect 32622 6466 32674 6478
rect 32622 6402 32674 6414
rect 33742 6466 33794 6478
rect 33742 6402 33794 6414
rect 34078 6466 34130 6478
rect 34078 6402 34130 6414
rect 36318 6466 36370 6478
rect 36318 6402 36370 6414
rect 45614 6466 45666 6478
rect 45614 6402 45666 6414
rect 51774 6466 51826 6478
rect 51774 6402 51826 6414
rect 55246 6466 55298 6478
rect 55246 6402 55298 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 1262 6130 1314 6142
rect 1262 6066 1314 6078
rect 6750 6130 6802 6142
rect 6750 6066 6802 6078
rect 20078 6130 20130 6142
rect 20078 6066 20130 6078
rect 21870 6130 21922 6142
rect 21870 6066 21922 6078
rect 28478 6130 28530 6142
rect 28478 6066 28530 6078
rect 34190 6130 34242 6142
rect 34190 6066 34242 6078
rect 34638 6130 34690 6142
rect 39006 6130 39058 6142
rect 36866 6078 36878 6130
rect 36930 6078 36942 6130
rect 34638 6066 34690 6078
rect 39006 6066 39058 6078
rect 41246 6130 41298 6142
rect 41246 6066 41298 6078
rect 44270 6130 44322 6142
rect 44270 6066 44322 6078
rect 44606 6130 44658 6142
rect 44606 6066 44658 6078
rect 52110 6130 52162 6142
rect 52110 6066 52162 6078
rect 52446 6130 52498 6142
rect 52446 6066 52498 6078
rect 53790 6130 53842 6142
rect 53790 6066 53842 6078
rect 12910 6018 12962 6030
rect 2818 5966 2830 6018
rect 2882 5966 2894 6018
rect 5170 5966 5182 6018
rect 5234 5966 5246 6018
rect 12002 5966 12014 6018
rect 12066 5966 12078 6018
rect 12910 5954 12962 5966
rect 14478 6018 14530 6030
rect 24670 6018 24722 6030
rect 21522 5966 21534 6018
rect 21586 5966 21598 6018
rect 22642 5966 22654 6018
rect 22706 5966 22718 6018
rect 39666 5966 39678 6018
rect 39730 5966 39742 6018
rect 41906 5966 41918 6018
rect 41970 5966 41982 6018
rect 14478 5954 14530 5966
rect 24670 5954 24722 5966
rect 7086 5906 7138 5918
rect 9214 5906 9266 5918
rect 11678 5906 11730 5918
rect 8082 5854 8094 5906
rect 8146 5854 8158 5906
rect 8530 5854 8542 5906
rect 8594 5854 8606 5906
rect 9874 5854 9886 5906
rect 9938 5854 9950 5906
rect 10882 5854 10894 5906
rect 10946 5854 10958 5906
rect 11442 5854 11454 5906
rect 11506 5854 11518 5906
rect 7086 5842 7138 5854
rect 9214 5842 9266 5854
rect 11678 5842 11730 5854
rect 11902 5906 11954 5918
rect 12686 5906 12738 5918
rect 12114 5854 12126 5906
rect 12178 5854 12190 5906
rect 11902 5842 11954 5854
rect 12686 5842 12738 5854
rect 13246 5906 13298 5918
rect 13246 5842 13298 5854
rect 14142 5906 14194 5918
rect 14142 5842 14194 5854
rect 14366 5906 14418 5918
rect 20750 5906 20802 5918
rect 15250 5854 15262 5906
rect 15314 5854 15326 5906
rect 15810 5854 15822 5906
rect 15874 5854 15886 5906
rect 16482 5854 16494 5906
rect 16546 5854 16558 5906
rect 17154 5854 17166 5906
rect 17218 5854 17230 5906
rect 17938 5854 17950 5906
rect 18002 5854 18014 5906
rect 19730 5854 19742 5906
rect 19794 5854 19806 5906
rect 14366 5842 14418 5854
rect 20750 5842 20802 5854
rect 24222 5906 24274 5918
rect 26126 5906 26178 5918
rect 36318 5906 36370 5918
rect 54126 5906 54178 5918
rect 24994 5854 25006 5906
rect 25058 5854 25070 5906
rect 25442 5854 25454 5906
rect 25506 5854 25518 5906
rect 26674 5854 26686 5906
rect 26738 5854 26750 5906
rect 27682 5854 27694 5906
rect 27746 5854 27758 5906
rect 29474 5854 29486 5906
rect 29538 5854 29550 5906
rect 32610 5854 32622 5906
rect 32674 5854 32686 5906
rect 36530 5854 36542 5906
rect 36594 5854 36606 5906
rect 36978 5854 36990 5906
rect 37042 5854 37054 5906
rect 38994 5854 39006 5906
rect 39058 5854 39070 5906
rect 45042 5854 45054 5906
rect 45106 5854 45118 5906
rect 45378 5854 45390 5906
rect 45442 5854 45454 5906
rect 52882 5854 52894 5906
rect 52946 5854 52958 5906
rect 53106 5854 53118 5906
rect 53170 5854 53182 5906
rect 24222 5842 24274 5854
rect 26126 5842 26178 5854
rect 36318 5842 36370 5854
rect 54126 5842 54178 5854
rect 55806 5906 55858 5918
rect 55806 5842 55858 5854
rect 7310 5794 7362 5806
rect 2370 5742 2382 5794
rect 2434 5742 2446 5794
rect 3490 5742 3502 5794
rect 3554 5742 3566 5794
rect 5506 5742 5518 5794
rect 5570 5742 5582 5794
rect 7310 5730 7362 5742
rect 7422 5794 7474 5806
rect 7422 5730 7474 5742
rect 7758 5794 7810 5806
rect 13134 5794 13186 5806
rect 8754 5742 8766 5794
rect 8818 5742 8830 5794
rect 7758 5730 7810 5742
rect 13134 5730 13186 5742
rect 14590 5794 14642 5806
rect 14590 5730 14642 5742
rect 14926 5794 14978 5806
rect 34862 5794 34914 5806
rect 15922 5742 15934 5794
rect 15986 5742 15998 5794
rect 23090 5742 23102 5794
rect 23154 5742 23166 5794
rect 29922 5742 29934 5794
rect 29986 5742 29998 5794
rect 14926 5730 14978 5742
rect 34862 5730 34914 5742
rect 38670 5794 38722 5806
rect 40114 5742 40126 5794
rect 40178 5742 40190 5794
rect 42242 5742 42254 5794
rect 42306 5742 42318 5794
rect 45154 5742 45166 5794
rect 45218 5742 45230 5794
rect 53218 5742 53230 5794
rect 53282 5742 53294 5794
rect 54338 5742 54350 5794
rect 54402 5742 54414 5794
rect 54898 5742 54910 5794
rect 54962 5742 54974 5794
rect 38670 5730 38722 5742
rect 3838 5682 3890 5694
rect 3838 5618 3890 5630
rect 19854 5682 19906 5694
rect 19854 5618 19906 5630
rect 19966 5682 20018 5694
rect 19966 5618 20018 5630
rect 20638 5682 20690 5694
rect 20638 5618 20690 5630
rect 20862 5682 20914 5694
rect 20862 5618 20914 5630
rect 21086 5682 21138 5694
rect 21086 5618 21138 5630
rect 21646 5682 21698 5694
rect 28590 5682 28642 5694
rect 25666 5630 25678 5682
rect 25730 5630 25742 5682
rect 21646 5618 21698 5630
rect 28590 5618 28642 5630
rect 28702 5682 28754 5694
rect 28702 5618 28754 5630
rect 31166 5682 31218 5694
rect 34750 5682 34802 5694
rect 37886 5682 37938 5694
rect 33058 5630 33070 5682
rect 33122 5630 33134 5682
rect 36754 5630 36766 5682
rect 36818 5630 36830 5682
rect 37538 5630 37550 5682
rect 37602 5630 37614 5682
rect 31166 5618 31218 5630
rect 34750 5618 34802 5630
rect 37886 5618 37938 5630
rect 43486 5682 43538 5694
rect 55458 5630 55470 5682
rect 55522 5630 55534 5682
rect 43486 5618 43538 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 1374 5346 1426 5358
rect 1026 5294 1038 5346
rect 1090 5294 1102 5346
rect 1374 5282 1426 5294
rect 5630 5346 5682 5358
rect 7982 5346 8034 5358
rect 6738 5294 6750 5346
rect 6802 5294 6814 5346
rect 5630 5282 5682 5294
rect 7982 5282 8034 5294
rect 9214 5346 9266 5358
rect 16606 5346 16658 5358
rect 19294 5346 19346 5358
rect 12562 5294 12574 5346
rect 12626 5294 12638 5346
rect 14578 5294 14590 5346
rect 14642 5294 14654 5346
rect 18162 5294 18174 5346
rect 18226 5294 18238 5346
rect 9214 5282 9266 5294
rect 16606 5282 16658 5294
rect 19294 5282 19346 5294
rect 23998 5346 24050 5358
rect 23998 5282 24050 5294
rect 25342 5346 25394 5358
rect 25342 5282 25394 5294
rect 27246 5346 27298 5358
rect 27246 5282 27298 5294
rect 27358 5346 27410 5358
rect 27358 5282 27410 5294
rect 33070 5346 33122 5358
rect 33070 5282 33122 5294
rect 33518 5346 33570 5358
rect 33518 5282 33570 5294
rect 33630 5346 33682 5358
rect 33630 5282 33682 5294
rect 33742 5346 33794 5358
rect 33742 5282 33794 5294
rect 36878 5346 36930 5358
rect 36878 5282 36930 5294
rect 37102 5346 37154 5358
rect 37102 5282 37154 5294
rect 38446 5346 38498 5358
rect 38446 5282 38498 5294
rect 39230 5346 39282 5358
rect 39230 5282 39282 5294
rect 39342 5346 39394 5358
rect 44830 5346 44882 5358
rect 42354 5294 42366 5346
rect 42418 5294 42430 5346
rect 39342 5282 39394 5294
rect 44830 5282 44882 5294
rect 53342 5346 53394 5358
rect 54126 5346 54178 5358
rect 53666 5294 53678 5346
rect 53730 5294 53742 5346
rect 53342 5282 53394 5294
rect 54126 5282 54178 5294
rect 1934 5234 1986 5246
rect 7758 5234 7810 5246
rect 16830 5234 16882 5246
rect 2930 5182 2942 5234
rect 2994 5182 3006 5234
rect 8866 5182 8878 5234
rect 8930 5182 8942 5234
rect 9538 5182 9550 5234
rect 9602 5182 9614 5234
rect 1934 5170 1986 5182
rect 7758 5170 7810 5182
rect 16830 5170 16882 5182
rect 16942 5234 16994 5246
rect 28030 5234 28082 5246
rect 20738 5182 20750 5234
rect 20802 5182 20814 5234
rect 23650 5182 23662 5234
rect 23714 5182 23726 5234
rect 24994 5182 25006 5234
rect 25058 5182 25070 5234
rect 16942 5170 16994 5182
rect 28030 5170 28082 5182
rect 34414 5234 34466 5246
rect 34414 5170 34466 5182
rect 34526 5234 34578 5246
rect 34526 5170 34578 5182
rect 36654 5234 36706 5246
rect 36654 5170 36706 5182
rect 41358 5234 41410 5246
rect 55234 5182 55246 5234
rect 55298 5182 55310 5234
rect 55906 5182 55918 5234
rect 55970 5182 55982 5234
rect 41358 5170 41410 5182
rect 3614 5122 3666 5134
rect 7982 5122 8034 5134
rect 2370 5070 2382 5122
rect 2434 5070 2446 5122
rect 2706 5070 2718 5122
rect 2770 5070 2782 5122
rect 4050 5070 4062 5122
rect 4114 5070 4126 5122
rect 4946 5070 4958 5122
rect 5010 5070 5022 5122
rect 3614 5058 3666 5070
rect 7982 5058 8034 5070
rect 8206 5122 8258 5134
rect 8206 5058 8258 5070
rect 9886 5122 9938 5134
rect 11902 5122 11954 5134
rect 19742 5122 19794 5134
rect 21422 5122 21474 5134
rect 26798 5122 26850 5134
rect 10434 5070 10446 5122
rect 10498 5070 10510 5122
rect 11330 5070 11342 5122
rect 11394 5070 11406 5122
rect 12674 5070 12686 5122
rect 12738 5070 12750 5122
rect 13122 5070 13134 5122
rect 13186 5070 13198 5122
rect 14130 5070 14142 5122
rect 14194 5070 14206 5122
rect 17602 5070 17614 5122
rect 17666 5070 17678 5122
rect 20178 5070 20190 5122
rect 20242 5070 20254 5122
rect 20514 5070 20526 5122
rect 20578 5070 20590 5122
rect 21970 5070 21982 5122
rect 22034 5070 22046 5122
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 25890 5070 25902 5122
rect 25954 5070 25966 5122
rect 9886 5058 9938 5070
rect 11902 5058 11954 5070
rect 19742 5058 19794 5070
rect 21422 5058 21474 5070
rect 26798 5058 26850 5070
rect 27470 5122 27522 5134
rect 27470 5058 27522 5070
rect 27918 5122 27970 5134
rect 34190 5122 34242 5134
rect 32834 5070 32846 5122
rect 32898 5070 32910 5122
rect 27918 5058 27970 5070
rect 34190 5058 34242 5070
rect 38670 5122 38722 5134
rect 43038 5122 43090 5134
rect 56254 5122 56306 5134
rect 41794 5070 41806 5122
rect 41858 5070 41870 5122
rect 42130 5070 42142 5122
rect 42194 5070 42206 5122
rect 43474 5070 43486 5122
rect 43538 5070 43550 5122
rect 44370 5070 44382 5122
rect 44434 5070 44446 5122
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 38670 5058 38722 5070
rect 43038 5058 43090 5070
rect 56254 5058 56306 5070
rect 13582 5010 13634 5022
rect 7186 4958 7198 5010
rect 7250 4958 7262 5010
rect 13582 4946 13634 4958
rect 26126 5010 26178 5022
rect 26126 4946 26178 4958
rect 26238 5010 26290 5022
rect 26238 4946 26290 4958
rect 27022 5010 27074 5022
rect 27022 4946 27074 4958
rect 33182 5010 33234 5022
rect 33182 4946 33234 4958
rect 36990 5010 37042 5022
rect 36990 4946 37042 4958
rect 37998 5010 38050 5022
rect 37998 4946 38050 4958
rect 38222 5010 38274 5022
rect 38222 4946 38274 4958
rect 38558 5010 38610 5022
rect 38558 4946 38610 4958
rect 54462 5010 54514 5022
rect 54462 4946 54514 4958
rect 15710 4898 15762 4910
rect 15710 4834 15762 4846
rect 26574 4898 26626 4910
rect 26574 4834 26626 4846
rect 39118 4898 39170 4910
rect 39118 4834 39170 4846
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 2942 4562 2994 4574
rect 2942 4498 2994 4510
rect 10446 4562 10498 4574
rect 10446 4498 10498 4510
rect 14590 4562 14642 4574
rect 14590 4498 14642 4510
rect 19182 4562 19234 4574
rect 19182 4498 19234 4510
rect 20750 4562 20802 4574
rect 20750 4498 20802 4510
rect 25118 4562 25170 4574
rect 25118 4498 25170 4510
rect 37998 4562 38050 4574
rect 37998 4498 38050 4510
rect 55694 4562 55746 4574
rect 55694 4498 55746 4510
rect 15038 4450 15090 4462
rect 8866 4398 8878 4450
rect 8930 4398 8942 4450
rect 15038 4386 15090 4398
rect 18622 4450 18674 4462
rect 18622 4386 18674 4398
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 26910 4450 26962 4462
rect 26910 4386 26962 4398
rect 30606 4450 30658 4462
rect 40350 4450 40402 4462
rect 38322 4398 38334 4450
rect 38386 4398 38398 4450
rect 30606 4386 30658 4398
rect 40350 4386 40402 4398
rect 44830 4450 44882 4462
rect 44830 4386 44882 4398
rect 3726 4338 3778 4350
rect 1362 4286 1374 4338
rect 1426 4286 1438 4338
rect 3726 4274 3778 4286
rect 4398 4338 4450 4350
rect 5630 4338 5682 4350
rect 19854 4338 19906 4350
rect 5058 4286 5070 4338
rect 5122 4286 5134 4338
rect 6514 4286 6526 4338
rect 6578 4286 6590 4338
rect 7298 4286 7310 4338
rect 7362 4286 7374 4338
rect 8082 4286 8094 4338
rect 8146 4286 8158 4338
rect 12898 4286 12910 4338
rect 12962 4286 12974 4338
rect 15474 4286 15486 4338
rect 15538 4286 15550 4338
rect 15922 4286 15934 4338
rect 15986 4286 15998 4338
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 17266 4286 17278 4338
rect 17330 4286 17342 4338
rect 18050 4286 18062 4338
rect 18114 4286 18126 4338
rect 4398 4274 4450 4286
rect 5630 4274 5682 4286
rect 19854 4274 19906 4286
rect 19966 4338 20018 4350
rect 19966 4274 20018 4286
rect 20078 4338 20130 4350
rect 20078 4274 20130 4286
rect 20638 4338 20690 4350
rect 22990 4338 23042 4350
rect 26798 4338 26850 4350
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 22082 4286 22094 4338
rect 22146 4286 22158 4338
rect 23538 4286 23550 4338
rect 23602 4286 23614 4338
rect 20638 4274 20690 4286
rect 22990 4274 23042 4286
rect 26798 4274 26850 4286
rect 27022 4338 27074 4350
rect 27022 4274 27074 4286
rect 27470 4338 27522 4350
rect 35758 4338 35810 4350
rect 30146 4286 30158 4338
rect 30210 4286 30222 4338
rect 31042 4286 31054 4338
rect 31106 4286 31118 4338
rect 31378 4286 31390 4338
rect 31442 4286 31454 4338
rect 32162 4286 32174 4338
rect 32226 4286 32238 4338
rect 32610 4286 32622 4338
rect 32674 4286 32686 4338
rect 33730 4286 33742 4338
rect 33794 4286 33806 4338
rect 27470 4274 27522 4286
rect 35758 4274 35810 4286
rect 36430 4338 36482 4350
rect 44158 4338 44210 4350
rect 39778 4286 39790 4338
rect 39842 4286 39854 4338
rect 40674 4286 40686 4338
rect 40738 4286 40750 4338
rect 41234 4286 41246 4338
rect 41298 4286 41310 4338
rect 42578 4286 42590 4338
rect 42642 4286 42654 4338
rect 43362 4286 43374 4338
rect 43426 4286 43438 4338
rect 36430 4274 36482 4286
rect 44158 4274 44210 4286
rect 44494 4338 44546 4350
rect 54462 4338 54514 4350
rect 56030 4338 56082 4350
rect 46274 4286 46286 4338
rect 46338 4286 46350 4338
rect 54898 4286 54910 4338
rect 54962 4286 54974 4338
rect 44494 4274 44546 4286
rect 54462 4274 54514 4286
rect 56030 4274 56082 4286
rect 6974 4226 7026 4238
rect 27246 4226 27298 4238
rect 1810 4174 1822 4226
rect 1874 4174 1886 4226
rect 3378 4174 3390 4226
rect 3442 4174 3454 4226
rect 4050 4174 4062 4226
rect 4114 4174 4126 4226
rect 6290 4174 6302 4226
rect 6354 4174 6366 4226
rect 7522 4174 7534 4226
rect 7586 4174 7598 4226
rect 9202 4174 9214 4226
rect 9266 4174 9278 4226
rect 10882 4174 10894 4226
rect 10946 4174 10958 4226
rect 11554 4174 11566 4226
rect 11618 4174 11630 4226
rect 13346 4174 13358 4226
rect 13410 4174 13422 4226
rect 6974 4162 7026 4174
rect 27246 4162 27298 4174
rect 36318 4226 36370 4238
rect 36318 4162 36370 4174
rect 38222 4226 38274 4238
rect 41806 4226 41858 4238
rect 41346 4174 41358 4226
rect 41410 4174 41422 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 38222 4162 38274 4174
rect 41806 4162 41858 4174
rect 11230 4114 11282 4126
rect 5282 4062 5294 4114
rect 5346 4062 5358 4114
rect 5954 4062 5966 4114
rect 6018 4062 6030 4114
rect 7858 4062 7870 4114
rect 7922 4062 7934 4114
rect 11230 4050 11282 4062
rect 11902 4114 11954 4126
rect 18734 4114 18786 4126
rect 16034 4062 16046 4114
rect 16098 4062 16110 4114
rect 11902 4050 11954 4062
rect 18734 4050 18786 4062
rect 19630 4114 19682 4126
rect 19630 4050 19682 4062
rect 21086 4114 21138 4126
rect 21086 4050 21138 4062
rect 21422 4114 21474 4126
rect 26462 4114 26514 4126
rect 28814 4114 28866 4126
rect 34526 4114 34578 4126
rect 44270 4114 44322 4126
rect 22306 4062 22318 4114
rect 22370 4062 22382 4114
rect 22642 4062 22654 4114
rect 22706 4062 22718 4114
rect 23986 4062 23998 4114
rect 24050 4062 24062 4114
rect 26114 4062 26126 4114
rect 26178 4062 26190 4114
rect 28466 4062 28478 4114
rect 28530 4062 28542 4114
rect 29922 4062 29934 4114
rect 29986 4062 29998 4114
rect 31602 4062 31614 4114
rect 31666 4062 31678 4114
rect 34178 4062 34190 4114
rect 34242 4062 34254 4114
rect 35410 4062 35422 4114
rect 35474 4062 35486 4114
rect 40002 4062 40014 4114
rect 40066 4062 40078 4114
rect 46498 4062 46510 4114
rect 46562 4062 46574 4114
rect 54114 4062 54126 4114
rect 54178 4062 54190 4114
rect 21422 4050 21474 4062
rect 26462 4050 26514 4062
rect 28814 4050 28866 4062
rect 34526 4050 34578 4062
rect 44270 4050 44322 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 2830 3778 2882 3790
rect 6750 3778 6802 3790
rect 7982 3778 8034 3790
rect 9102 3778 9154 3790
rect 1362 3726 1374 3778
rect 1426 3726 1438 3778
rect 2034 3726 2046 3778
rect 2098 3726 2110 3778
rect 3938 3726 3950 3778
rect 4002 3726 4014 3778
rect 5618 3726 5630 3778
rect 5682 3726 5694 3778
rect 7298 3726 7310 3778
rect 7362 3726 7374 3778
rect 8306 3726 8318 3778
rect 8370 3726 8382 3778
rect 2830 3714 2882 3726
rect 6750 3714 6802 3726
rect 7982 3714 8034 3726
rect 9102 3714 9154 3726
rect 9774 3778 9826 3790
rect 12238 3778 12290 3790
rect 11106 3726 11118 3778
rect 11170 3726 11182 3778
rect 9774 3714 9826 3726
rect 12238 3714 12290 3726
rect 13022 3778 13074 3790
rect 13022 3714 13074 3726
rect 16942 3778 16994 3790
rect 16942 3714 16994 3726
rect 21646 3778 21698 3790
rect 21646 3714 21698 3726
rect 24894 3778 24946 3790
rect 24894 3714 24946 3726
rect 25566 3778 25618 3790
rect 27694 3778 27746 3790
rect 32398 3778 32450 3790
rect 36766 3778 36818 3790
rect 26562 3726 26574 3778
rect 26626 3726 26638 3778
rect 29138 3726 29150 3778
rect 29202 3726 29214 3778
rect 34290 3726 34302 3778
rect 34354 3726 34366 3778
rect 25566 3714 25618 3726
rect 27694 3714 27746 3726
rect 32398 3714 32450 3726
rect 36766 3714 36818 3726
rect 37550 3778 37602 3790
rect 37550 3714 37602 3726
rect 37998 3778 38050 3790
rect 37998 3714 38050 3726
rect 42142 3778 42194 3790
rect 42142 3714 42194 3726
rect 42814 3778 42866 3790
rect 42814 3714 42866 3726
rect 44830 3778 44882 3790
rect 44830 3714 44882 3726
rect 46174 3778 46226 3790
rect 46174 3714 46226 3726
rect 46846 3778 46898 3790
rect 55358 3778 55410 3790
rect 56366 3778 56418 3790
rect 55010 3726 55022 3778
rect 55074 3726 55086 3778
rect 56018 3726 56030 3778
rect 56082 3726 56094 3778
rect 46846 3714 46898 3726
rect 55358 3714 55410 3726
rect 56366 3714 56418 3726
rect 7646 3666 7698 3678
rect 17054 3666 17106 3678
rect 19854 3666 19906 3678
rect 9426 3614 9438 3666
rect 9490 3614 9502 3666
rect 10098 3614 10110 3666
rect 10162 3614 10174 3666
rect 12674 3614 12686 3666
rect 12738 3614 12750 3666
rect 13682 3614 13694 3666
rect 13746 3614 13758 3666
rect 14914 3614 14926 3666
rect 14978 3614 14990 3666
rect 18722 3614 18734 3666
rect 18786 3614 18798 3666
rect 7646 3602 7698 3614
rect 17054 3602 17106 3614
rect 19854 3602 19906 3614
rect 20974 3666 21026 3678
rect 20974 3602 21026 3614
rect 21758 3666 21810 3678
rect 28142 3666 28194 3678
rect 35870 3666 35922 3678
rect 22642 3614 22654 3666
rect 22706 3614 22718 3666
rect 24546 3614 24558 3666
rect 24610 3614 24622 3666
rect 25218 3614 25230 3666
rect 25282 3614 25294 3666
rect 32722 3614 32734 3666
rect 32786 3614 32798 3666
rect 21758 3602 21810 3614
rect 28142 3602 28194 3614
rect 35870 3602 35922 3614
rect 36094 3666 36146 3678
rect 44158 3666 44210 3678
rect 37202 3614 37214 3666
rect 37266 3614 37278 3666
rect 39666 3614 39678 3666
rect 39730 3614 39742 3666
rect 40898 3614 40910 3666
rect 40962 3614 40974 3666
rect 43026 3614 43038 3666
rect 43090 3614 43102 3666
rect 45154 3614 45166 3666
rect 45218 3614 45230 3666
rect 45490 3614 45502 3666
rect 45554 3614 45566 3666
rect 47058 3614 47070 3666
rect 47122 3614 47134 3666
rect 36094 3602 36146 3614
rect 44158 3602 44210 3614
rect 2382 3554 2434 3566
rect 16606 3554 16658 3566
rect 1586 3502 1598 3554
rect 1650 3502 1662 3554
rect 5170 3502 5182 3554
rect 5234 3502 5246 3554
rect 10658 3502 10670 3554
rect 10722 3502 10734 3554
rect 13458 3502 13470 3554
rect 13522 3502 13534 3554
rect 14466 3502 14478 3554
rect 14530 3502 14542 3554
rect 2382 3490 2434 3502
rect 16606 3490 16658 3502
rect 17166 3554 17218 3566
rect 20526 3554 20578 3566
rect 18162 3502 18174 3554
rect 18226 3502 18238 3554
rect 17166 3490 17218 3502
rect 20526 3490 20578 3502
rect 20750 3554 20802 3566
rect 20750 3490 20802 3502
rect 21198 3554 21250 3566
rect 29822 3554 29874 3566
rect 39342 3554 39394 3566
rect 22306 3502 22318 3554
rect 22370 3502 22382 3554
rect 26114 3502 26126 3554
rect 26178 3502 26190 3554
rect 28466 3502 28478 3554
rect 28530 3502 28542 3554
rect 29026 3502 29038 3554
rect 29090 3502 29102 3554
rect 30146 3502 30158 3554
rect 30210 3502 30222 3554
rect 31154 3502 31166 3554
rect 31218 3502 31230 3554
rect 33842 3502 33854 3554
rect 33906 3502 33918 3554
rect 21198 3490 21250 3502
rect 29822 3490 29874 3502
rect 39342 3490 39394 3502
rect 43374 3554 43426 3566
rect 43374 3490 43426 3502
rect 45838 3554 45890 3566
rect 45838 3490 45890 3502
rect 47406 3554 47458 3566
rect 47406 3490 47458 3502
rect 16046 3442 16098 3454
rect 4386 3390 4398 3442
rect 4450 3390 4462 3442
rect 16046 3378 16098 3390
rect 21086 3442 21138 3454
rect 21086 3378 21138 3390
rect 35422 3442 35474 3454
rect 36542 3442 36594 3454
rect 37886 3442 37938 3454
rect 36194 3390 36206 3442
rect 36258 3390 36270 3442
rect 36866 3390 36878 3442
rect 36930 3390 36942 3442
rect 40562 3390 40574 3442
rect 40626 3390 40638 3442
rect 35422 3378 35474 3390
rect 36542 3378 36594 3390
rect 37886 3378 37938 3390
rect 23886 3330 23938 3342
rect 23886 3266 23938 3278
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 1150 2994 1202 3006
rect 1150 2930 1202 2942
rect 5630 2994 5682 3006
rect 5630 2930 5682 2942
rect 10558 2994 10610 3006
rect 10558 2930 10610 2942
rect 15374 2994 15426 3006
rect 15374 2930 15426 2942
rect 22206 2994 22258 3006
rect 22206 2930 22258 2942
rect 30270 2994 30322 3006
rect 30270 2930 30322 2942
rect 40014 2994 40066 3006
rect 40014 2930 40066 2942
rect 7646 2882 7698 2894
rect 16606 2882 16658 2894
rect 43486 2882 43538 2894
rect 2706 2830 2718 2882
rect 2770 2830 2782 2882
rect 13794 2830 13806 2882
rect 13858 2830 13870 2882
rect 17266 2830 17278 2882
rect 17330 2830 17342 2882
rect 28690 2830 28702 2882
rect 28754 2830 28766 2882
rect 7646 2818 7698 2830
rect 16606 2818 16658 2830
rect 43486 2818 43538 2830
rect 3726 2770 3778 2782
rect 8094 2770 8146 2782
rect 11230 2770 11282 2782
rect 16158 2770 16210 2782
rect 21198 2770 21250 2782
rect 24894 2770 24946 2782
rect 32174 2770 32226 2782
rect 34302 2770 34354 2782
rect 35758 2770 35810 2782
rect 4274 2718 4286 2770
rect 4338 2718 4350 2770
rect 7186 2718 7198 2770
rect 7250 2718 7262 2770
rect 8866 2718 8878 2770
rect 8930 2718 8942 2770
rect 12002 2718 12014 2770
rect 12066 2718 12078 2770
rect 13010 2718 13022 2770
rect 13074 2718 13086 2770
rect 19506 2718 19518 2770
rect 19570 2718 19582 2770
rect 20962 2718 20974 2770
rect 21026 2718 21038 2770
rect 21298 2718 21310 2770
rect 21362 2718 21374 2770
rect 21858 2718 21870 2770
rect 21922 2718 21934 2770
rect 22418 2718 22430 2770
rect 22482 2718 22494 2770
rect 23762 2718 23774 2770
rect 23826 2718 23838 2770
rect 24210 2718 24222 2770
rect 24274 2718 24286 2770
rect 25666 2718 25678 2770
rect 25730 2718 25742 2770
rect 26450 2718 26462 2770
rect 26514 2718 26526 2770
rect 27794 2718 27806 2770
rect 27858 2718 27870 2770
rect 31042 2718 31054 2770
rect 31106 2718 31118 2770
rect 31490 2718 31502 2770
rect 31554 2718 31566 2770
rect 32946 2718 32958 2770
rect 33010 2718 33022 2770
rect 33730 2718 33742 2770
rect 33794 2718 33806 2770
rect 35186 2718 35198 2770
rect 35250 2718 35262 2770
rect 3726 2706 3778 2718
rect 8094 2706 8146 2718
rect 11230 2706 11282 2718
rect 16158 2706 16210 2718
rect 21198 2706 21250 2718
rect 24894 2706 24946 2718
rect 32174 2706 32226 2718
rect 34302 2706 34354 2718
rect 35758 2706 35810 2718
rect 36654 2770 36706 2782
rect 36654 2706 36706 2718
rect 37326 2770 37378 2782
rect 37326 2706 37378 2718
rect 37662 2770 37714 2782
rect 42142 2770 42194 2782
rect 38546 2718 38558 2770
rect 38610 2718 38622 2770
rect 39330 2718 39342 2770
rect 39394 2718 39406 2770
rect 41682 2718 41694 2770
rect 41746 2718 41758 2770
rect 37662 2706 37714 2718
rect 42142 2706 42194 2718
rect 42814 2770 42866 2782
rect 42814 2706 42866 2718
rect 43598 2770 43650 2782
rect 43598 2706 43650 2718
rect 44494 2770 44546 2782
rect 44494 2706 44546 2718
rect 44830 2770 44882 2782
rect 44830 2706 44882 2718
rect 45502 2770 45554 2782
rect 45502 2706 45554 2718
rect 46510 2770 46562 2782
rect 46510 2706 46562 2718
rect 46846 2770 46898 2782
rect 55582 2770 55634 2782
rect 48402 2718 48414 2770
rect 48466 2718 48478 2770
rect 46846 2706 46898 2718
rect 55582 2706 55634 2718
rect 56254 2770 56306 2782
rect 56254 2706 56306 2718
rect 16718 2658 16770 2670
rect 2258 2606 2270 2658
rect 2322 2606 2334 2658
rect 3378 2606 3390 2658
rect 3442 2606 3454 2658
rect 6850 2606 6862 2658
rect 6914 2606 6926 2658
rect 8418 2606 8430 2658
rect 8482 2606 8494 2658
rect 9314 2606 9326 2658
rect 9378 2606 9390 2658
rect 14242 2606 14254 2658
rect 14306 2606 14318 2658
rect 15810 2606 15822 2658
rect 15874 2606 15886 2658
rect 16718 2594 16770 2606
rect 19966 2658 20018 2670
rect 19966 2594 20018 2606
rect 20750 2658 20802 2670
rect 20750 2594 20802 2606
rect 22654 2658 22706 2670
rect 22654 2594 22706 2606
rect 22990 2658 23042 2670
rect 22990 2594 23042 2606
rect 23102 2658 23154 2670
rect 23102 2594 23154 2606
rect 23438 2658 23490 2670
rect 30718 2658 30770 2670
rect 35646 2658 35698 2670
rect 29026 2606 29038 2658
rect 29090 2606 29102 2658
rect 34962 2606 34974 2658
rect 35026 2606 35038 2658
rect 41122 2606 41134 2658
rect 41186 2606 41198 2658
rect 44146 2606 44158 2658
rect 44210 2606 44222 2658
rect 46162 2606 46174 2658
rect 46226 2606 46238 2658
rect 48850 2606 48862 2658
rect 48914 2606 48926 2658
rect 55234 2606 55246 2658
rect 55298 2606 55310 2658
rect 55906 2606 55918 2658
rect 55970 2606 55982 2658
rect 23438 2594 23490 2606
rect 30718 2594 30770 2606
rect 35646 2594 35698 2606
rect 18846 2546 18898 2558
rect 4050 2494 4062 2546
rect 4114 2494 4126 2546
rect 11554 2494 11566 2546
rect 11618 2494 11630 2546
rect 12226 2494 12238 2546
rect 12290 2494 12302 2546
rect 12786 2494 12798 2546
rect 12850 2494 12862 2546
rect 17714 2494 17726 2546
rect 17778 2494 17790 2546
rect 18846 2482 18898 2494
rect 19854 2546 19906 2558
rect 19854 2482 19906 2494
rect 20078 2546 20130 2558
rect 20078 2482 20130 2494
rect 21534 2546 21586 2558
rect 21534 2482 21586 2494
rect 22542 2546 22594 2558
rect 47854 2546 47906 2558
rect 49198 2546 49250 2558
rect 24434 2494 24446 2546
rect 24498 2494 24510 2546
rect 27570 2494 27582 2546
rect 27634 2494 27646 2546
rect 31714 2494 31726 2546
rect 31778 2494 31790 2546
rect 34626 2494 34638 2546
rect 34690 2494 34702 2546
rect 36306 2494 36318 2546
rect 36370 2494 36382 2546
rect 36978 2494 36990 2546
rect 37042 2494 37054 2546
rect 37986 2494 37998 2546
rect 38050 2494 38062 2546
rect 38322 2494 38334 2546
rect 38386 2494 38398 2546
rect 39554 2494 39566 2546
rect 39618 2494 39630 2546
rect 42466 2494 42478 2546
rect 42530 2494 42542 2546
rect 43138 2494 43150 2546
rect 43202 2494 43214 2546
rect 45154 2494 45166 2546
rect 45218 2494 45230 2546
rect 45826 2494 45838 2546
rect 45890 2494 45902 2546
rect 47170 2494 47182 2546
rect 47234 2494 47246 2546
rect 47506 2494 47518 2546
rect 47570 2494 47582 2546
rect 48178 2494 48190 2546
rect 48242 2494 48254 2546
rect 22542 2482 22594 2494
rect 47854 2482 47906 2494
rect 49198 2482 49250 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 2270 2210 2322 2222
rect 1586 2158 1598 2210
rect 1650 2158 1662 2210
rect 2270 2146 2322 2158
rect 5294 2210 5346 2222
rect 10782 2210 10834 2222
rect 6402 2158 6414 2210
rect 6466 2158 6478 2210
rect 7970 2158 7982 2210
rect 8034 2158 8046 2210
rect 9650 2158 9662 2210
rect 9714 2158 9726 2210
rect 5294 2146 5346 2158
rect 10782 2146 10834 2158
rect 11342 2210 11394 2222
rect 13470 2210 13522 2222
rect 14926 2210 14978 2222
rect 15598 2210 15650 2222
rect 12450 2158 12462 2210
rect 12514 2158 12526 2210
rect 13906 2158 13918 2210
rect 13970 2158 13982 2210
rect 15250 2158 15262 2210
rect 15314 2158 15326 2210
rect 11342 2146 11394 2158
rect 13470 2146 13522 2158
rect 14926 2146 14978 2158
rect 15598 2146 15650 2158
rect 17054 2210 17106 2222
rect 23886 2210 23938 2222
rect 19282 2158 19294 2210
rect 19346 2158 19358 2210
rect 17054 2146 17106 2158
rect 23886 2146 23938 2158
rect 24894 2210 24946 2222
rect 24894 2146 24946 2158
rect 25230 2210 25282 2222
rect 27694 2210 27746 2222
rect 26562 2158 26574 2210
rect 26626 2158 26638 2210
rect 25230 2146 25282 2158
rect 27694 2146 27746 2158
rect 28590 2210 28642 2222
rect 29262 2210 29314 2222
rect 31726 2210 31778 2222
rect 28914 2158 28926 2210
rect 28978 2158 28990 2210
rect 30594 2158 30606 2210
rect 30658 2158 30670 2210
rect 28590 2146 28642 2158
rect 29262 2146 29314 2158
rect 31726 2146 31778 2158
rect 33630 2210 33682 2222
rect 33630 2146 33682 2158
rect 34414 2210 34466 2222
rect 34414 2146 34466 2158
rect 35086 2210 35138 2222
rect 37550 2210 37602 2222
rect 36194 2158 36206 2210
rect 36258 2158 36270 2210
rect 35086 2146 35138 2158
rect 37550 2146 37602 2158
rect 38222 2210 38274 2222
rect 38222 2146 38274 2158
rect 38558 2210 38610 2222
rect 39230 2210 39282 2222
rect 38882 2158 38894 2210
rect 38946 2158 38958 2210
rect 38558 2146 38610 2158
rect 39230 2146 39282 2158
rect 40798 2210 40850 2222
rect 40798 2146 40850 2158
rect 41470 2210 41522 2222
rect 41470 2146 41522 2158
rect 42142 2210 42194 2222
rect 42142 2146 42194 2158
rect 42926 2210 42978 2222
rect 42926 2146 42978 2158
rect 43934 2210 43986 2222
rect 43934 2146 43986 2158
rect 44270 2210 44322 2222
rect 44270 2146 44322 2158
rect 44942 2210 44994 2222
rect 46286 2210 46338 2222
rect 45602 2158 45614 2210
rect 45666 2158 45678 2210
rect 44942 2146 44994 2158
rect 46286 2146 46338 2158
rect 47294 2210 47346 2222
rect 47294 2146 47346 2158
rect 48078 2210 48130 2222
rect 49086 2210 49138 2222
rect 48402 2158 48414 2210
rect 48466 2158 48478 2210
rect 48738 2158 48750 2210
rect 48802 2158 48814 2210
rect 48078 2146 48130 2158
rect 49086 2146 49138 2158
rect 49758 2210 49810 2222
rect 55906 2158 55918 2210
rect 55970 2158 55982 2210
rect 49758 2146 49810 2158
rect 4734 2098 4786 2110
rect 2594 2046 2606 2098
rect 2658 2046 2670 2098
rect 3490 2046 3502 2098
rect 3554 2046 3566 2098
rect 4734 2034 4786 2046
rect 13582 2098 13634 2110
rect 16158 2098 16210 2110
rect 17726 2098 17778 2110
rect 14578 2046 14590 2098
rect 14642 2046 14654 2098
rect 16706 2046 16718 2098
rect 16770 2046 16782 2098
rect 13582 2034 13634 2046
rect 16158 2034 16210 2046
rect 17726 2034 17778 2046
rect 18286 2098 18338 2110
rect 22642 2046 22654 2098
rect 22706 2046 22718 2098
rect 24546 2046 24558 2098
rect 24610 2046 24622 2098
rect 25554 2046 25566 2098
rect 25618 2046 25630 2098
rect 29586 2046 29598 2098
rect 29650 2046 29662 2098
rect 32498 2046 32510 2098
rect 32562 2046 32574 2098
rect 33058 2046 33070 2098
rect 33122 2046 33134 2098
rect 34066 2046 34078 2098
rect 34130 2046 34142 2098
rect 37202 2046 37214 2098
rect 37266 2046 37278 2098
rect 37874 2046 37886 2098
rect 37938 2046 37950 2098
rect 39554 2046 39566 2098
rect 39618 2046 39630 2098
rect 40450 2046 40462 2098
rect 40514 2046 40526 2098
rect 41122 2046 41134 2098
rect 41186 2046 41198 2098
rect 43250 2046 43262 2098
rect 43314 2046 43326 2098
rect 43586 2046 43598 2098
rect 43650 2046 43662 2098
rect 44594 2046 44606 2098
rect 44658 2046 44670 2098
rect 45266 2046 45278 2098
rect 45330 2046 45342 2098
rect 46610 2046 46622 2098
rect 46674 2046 46686 2098
rect 46946 2046 46958 2098
rect 47010 2046 47022 2098
rect 49410 2046 49422 2098
rect 49474 2046 49486 2098
rect 18286 2034 18338 2046
rect 1934 1986 1986 1998
rect 17950 1986 18002 1998
rect 33294 1986 33346 1998
rect 3154 1934 3166 1986
rect 3218 1934 3230 1986
rect 6962 1934 6974 1986
rect 7026 1934 7038 1986
rect 8194 1934 8206 1986
rect 8258 1934 8270 1986
rect 9090 1934 9102 1986
rect 9154 1934 9166 1986
rect 12898 1934 12910 1986
rect 12962 1934 12974 1986
rect 14130 1934 14142 1986
rect 14194 1934 14206 1986
rect 18722 1934 18734 1986
rect 18786 1934 18798 1986
rect 19058 1934 19070 1986
rect 19122 1934 19134 1986
rect 19842 1934 19854 1986
rect 19906 1934 19918 1986
rect 20290 1934 20302 1986
rect 20354 1934 20366 1986
rect 21410 1934 21422 1986
rect 21474 1934 21486 1986
rect 22306 1934 22318 1986
rect 22370 1934 22382 1986
rect 26002 1934 26014 1986
rect 26066 1934 26078 1986
rect 30034 1934 30046 1986
rect 30098 1934 30110 1986
rect 36754 1934 36766 1986
rect 36818 1934 36830 1986
rect 45826 1934 45838 1986
rect 45890 1934 45902 1986
rect 56130 1934 56142 1986
rect 56194 1934 56206 1986
rect 1934 1922 1986 1934
rect 17950 1922 18002 1934
rect 33294 1922 33346 1934
rect 1374 1874 1426 1886
rect 17602 1822 17614 1874
rect 17666 1822 17678 1874
rect 1374 1810 1426 1822
rect 16046 1762 16098 1774
rect 16046 1698 16098 1710
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 2494 1426 2546 1438
rect 2494 1362 2546 1374
rect 5630 1426 5682 1438
rect 5630 1362 5682 1374
rect 8766 1426 8818 1438
rect 8766 1362 8818 1374
rect 19182 1426 19234 1438
rect 19182 1362 19234 1374
rect 33294 1426 33346 1438
rect 33294 1362 33346 1374
rect 42254 1426 42306 1438
rect 42254 1362 42306 1374
rect 42926 1314 42978 1326
rect 31714 1262 31726 1314
rect 31778 1262 31790 1314
rect 40674 1262 40686 1314
rect 40738 1262 40750 1314
rect 42926 1250 42978 1262
rect 44270 1314 44322 1326
rect 44270 1250 44322 1262
rect 44830 1314 44882 1326
rect 44830 1250 44882 1262
rect 46286 1314 46338 1326
rect 46286 1250 46338 1262
rect 48078 1314 48130 1326
rect 48078 1250 48130 1262
rect 1038 1202 1090 1214
rect 4846 1202 4898 1214
rect 12574 1202 12626 1214
rect 15486 1202 15538 1214
rect 20302 1202 20354 1214
rect 21646 1202 21698 1214
rect 25454 1202 25506 1214
rect 1810 1150 1822 1202
rect 1874 1150 1886 1202
rect 4162 1150 4174 1202
rect 4226 1150 4238 1202
rect 7186 1150 7198 1202
rect 7250 1150 7262 1202
rect 10322 1150 10334 1202
rect 10386 1150 10398 1202
rect 11778 1150 11790 1202
rect 11842 1150 11854 1202
rect 14242 1150 14254 1202
rect 14306 1150 14318 1202
rect 16482 1150 16494 1202
rect 16546 1150 16558 1202
rect 17490 1150 17502 1202
rect 17554 1150 17566 1202
rect 21074 1150 21086 1202
rect 21138 1150 21150 1202
rect 23090 1150 23102 1202
rect 23154 1150 23166 1202
rect 24210 1150 24222 1202
rect 24274 1150 24286 1202
rect 24882 1150 24894 1202
rect 24946 1150 24958 1202
rect 1038 1138 1090 1150
rect 4846 1138 4898 1150
rect 12574 1138 12626 1150
rect 15486 1138 15538 1150
rect 20302 1138 20354 1150
rect 21646 1138 21698 1150
rect 25454 1138 25506 1150
rect 26126 1202 26178 1214
rect 28030 1202 28082 1214
rect 26898 1150 26910 1202
rect 26962 1150 26974 1202
rect 26126 1138 26178 1150
rect 28030 1138 28082 1150
rect 28702 1202 28754 1214
rect 28702 1138 28754 1150
rect 29374 1202 29426 1214
rect 36318 1202 36370 1214
rect 37662 1202 37714 1214
rect 39454 1202 39506 1214
rect 43486 1202 43538 1214
rect 48638 1202 48690 1214
rect 30146 1150 30158 1202
rect 30210 1150 30222 1202
rect 35522 1150 35534 1202
rect 35586 1150 35598 1202
rect 36866 1150 36878 1202
rect 36930 1150 36942 1202
rect 38210 1150 38222 1202
rect 38274 1150 38286 1202
rect 40002 1150 40014 1202
rect 40066 1150 40078 1202
rect 45266 1150 45278 1202
rect 45330 1150 45342 1202
rect 46946 1150 46958 1202
rect 47010 1150 47022 1202
rect 47618 1150 47630 1202
rect 47682 1150 47694 1202
rect 49186 1150 49198 1202
rect 49250 1150 49262 1202
rect 49858 1150 49870 1202
rect 49922 1150 49934 1202
rect 50754 1150 50766 1202
rect 50818 1150 50830 1202
rect 29374 1138 29426 1150
rect 36318 1138 36370 1150
rect 37662 1138 37714 1150
rect 39454 1138 39506 1150
rect 43486 1138 43538 1150
rect 48638 1138 48690 1150
rect 11230 1090 11282 1102
rect 22318 1090 22370 1102
rect 34750 1090 34802 1102
rect 1362 1038 1374 1090
rect 1426 1038 1438 1090
rect 2034 1038 2046 1090
rect 2098 1038 2110 1090
rect 3602 1038 3614 1090
rect 3666 1038 3678 1090
rect 6850 1038 6862 1090
rect 6914 1038 6926 1090
rect 9874 1038 9886 1090
rect 9938 1038 9950 1090
rect 13682 1038 13694 1090
rect 13746 1038 13758 1090
rect 18050 1038 18062 1090
rect 18114 1038 18126 1090
rect 21970 1038 21982 1090
rect 22034 1038 22046 1090
rect 24434 1038 24446 1090
rect 24498 1038 24510 1090
rect 25778 1038 25790 1090
rect 25842 1038 25854 1090
rect 29026 1038 29038 1090
rect 29090 1038 29102 1090
rect 29698 1038 29710 1090
rect 29762 1038 29774 1090
rect 32050 1038 32062 1090
rect 32114 1038 32126 1090
rect 35298 1038 35310 1090
rect 35362 1038 35374 1090
rect 41010 1038 41022 1090
rect 41074 1038 41086 1090
rect 47394 1038 47406 1090
rect 47458 1038 47470 1090
rect 11230 1026 11282 1038
rect 22318 1026 22370 1038
rect 34750 1026 34802 1038
rect 8094 978 8146 990
rect 34078 978 34130 990
rect 5170 926 5182 978
rect 5234 926 5246 978
rect 7746 926 7758 978
rect 7810 926 7822 978
rect 10882 926 10894 978
rect 10946 926 10958 978
rect 11554 926 11566 978
rect 11618 926 11630 978
rect 15138 926 15150 978
rect 15202 926 15214 978
rect 16258 926 16270 978
rect 16322 926 16334 978
rect 20626 926 20638 978
rect 20690 926 20702 978
rect 21298 926 21310 978
rect 21362 926 21374 978
rect 22642 926 22654 978
rect 22706 926 22718 978
rect 23314 926 23326 978
rect 23378 926 23390 978
rect 25106 926 25118 978
rect 25170 926 25182 978
rect 26450 926 26462 978
rect 26514 926 26526 978
rect 27122 926 27134 978
rect 27186 926 27198 978
rect 28354 926 28366 978
rect 28418 926 28430 978
rect 30370 926 30382 978
rect 30434 926 30446 978
rect 33730 926 33742 978
rect 33794 926 33806 978
rect 34402 926 34414 978
rect 34466 926 34478 978
rect 35970 926 35982 978
rect 36034 926 36046 978
rect 36642 926 36654 978
rect 36706 926 36718 978
rect 37314 926 37326 978
rect 37378 926 37390 978
rect 37986 926 37998 978
rect 38050 926 38062 978
rect 39106 926 39118 978
rect 39170 926 39182 978
rect 39778 926 39790 978
rect 39842 926 39854 978
rect 43138 926 43150 978
rect 43202 926 43214 978
rect 45042 926 45054 978
rect 45106 926 45118 978
rect 46722 926 46734 978
rect 46786 926 46798 978
rect 48290 926 48302 978
rect 48354 926 48366 978
rect 48962 926 48974 978
rect 49026 926 49038 978
rect 49634 926 49646 978
rect 49698 926 49710 978
rect 50530 926 50542 978
rect 50594 926 50606 978
rect 8094 914 8146 926
rect 34078 914 34130 926
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 43806 56422 43858 56474
rect 43910 56422 43962 56474
rect 44014 56422 44066 56474
rect 8094 56142 8146 56194
rect 3390 56030 3442 56082
rect 6750 56030 6802 56082
rect 7422 56030 7474 56082
rect 7982 56030 8034 56082
rect 9886 56030 9938 56082
rect 13246 56030 13298 56082
rect 14030 56030 14082 56082
rect 17390 56030 17442 56082
rect 17950 56030 18002 56082
rect 19294 56030 19346 56082
rect 20638 56030 20690 56082
rect 21646 56030 21698 56082
rect 24558 56030 24610 56082
rect 25118 56030 25170 56082
rect 26910 56030 26962 56082
rect 28702 56030 28754 56082
rect 30606 56030 30658 56082
rect 33182 56030 33234 56082
rect 34526 56030 34578 56082
rect 35534 56030 35586 56082
rect 36430 56030 36482 56082
rect 36878 56030 36930 56082
rect 37550 56030 37602 56082
rect 38446 56030 38498 56082
rect 39454 56030 39506 56082
rect 42142 56030 42194 56082
rect 43262 56030 43314 56082
rect 43822 56030 43874 56082
rect 45166 56030 45218 56082
rect 45838 56030 45890 56082
rect 54574 56030 54626 56082
rect 55022 56030 55074 56082
rect 2270 55918 2322 55970
rect 3614 55918 3666 55970
rect 3950 55918 4002 55970
rect 4846 55918 4898 55970
rect 6302 55918 6354 55970
rect 10110 55918 10162 55970
rect 10782 55918 10834 55970
rect 11902 55918 11954 55970
rect 13470 55918 13522 55970
rect 14366 55918 14418 55970
rect 16830 55918 16882 55970
rect 18174 55918 18226 55970
rect 18846 55918 18898 55970
rect 20414 55918 20466 55970
rect 21982 55918 22034 55970
rect 22654 55918 22706 55970
rect 23326 55918 23378 55970
rect 24222 55918 24274 55970
rect 24894 55918 24946 55970
rect 25790 55918 25842 55970
rect 28254 55918 28306 55970
rect 29934 55918 29986 55970
rect 32734 55918 32786 55970
rect 41022 55918 41074 55970
rect 43486 55918 43538 55970
rect 44158 55918 44210 55970
rect 46174 55918 46226 55970
rect 47070 55918 47122 55970
rect 47742 55918 47794 55970
rect 49086 55918 49138 55970
rect 49758 55918 49810 55970
rect 50542 55918 50594 55970
rect 51886 55918 51938 55970
rect 52558 55918 52610 55970
rect 53230 55918 53282 55970
rect 53566 55918 53618 55970
rect 1262 55806 1314 55858
rect 1598 55806 1650 55858
rect 1934 55806 1986 55858
rect 2606 55806 2658 55858
rect 2942 55806 2994 55858
rect 4286 55806 4338 55858
rect 4958 55806 5010 55858
rect 5294 55806 5346 55858
rect 5630 55806 5682 55858
rect 5966 55806 6018 55858
rect 6974 55806 7026 55858
rect 7646 55806 7698 55858
rect 9102 55806 9154 55858
rect 10446 55806 10498 55858
rect 11118 55806 11170 55858
rect 11566 55806 11618 55858
rect 12462 55806 12514 55858
rect 15598 55806 15650 55858
rect 16494 55806 16546 55858
rect 17166 55806 17218 55858
rect 18510 55806 18562 55858
rect 19518 55806 19570 55858
rect 20190 55806 20242 55858
rect 21534 55806 21586 55858
rect 21870 55806 21922 55858
rect 22318 55806 22370 55858
rect 22990 55806 23042 55858
rect 25454 55806 25506 55858
rect 25678 55806 25730 55858
rect 26126 55806 26178 55858
rect 26462 55806 26514 55858
rect 27134 55806 27186 55858
rect 27918 55806 27970 55858
rect 28926 55806 28978 55858
rect 29262 55806 29314 55858
rect 29598 55806 29650 55858
rect 30270 55806 30322 55858
rect 30942 55806 30994 55858
rect 31726 55806 31778 55858
rect 32062 55806 32114 55858
rect 32398 55806 32450 55858
rect 33406 55806 33458 55858
rect 33742 55806 33794 55858
rect 34078 55806 34130 55858
rect 34750 55806 34802 55858
rect 35758 55806 35810 55858
rect 36094 55806 36146 55858
rect 37102 55806 37154 55858
rect 37774 55806 37826 55858
rect 38110 55806 38162 55858
rect 39118 55806 39170 55858
rect 40014 55806 40066 55858
rect 40350 55806 40402 55858
rect 40686 55806 40738 55858
rect 41358 55806 41410 55858
rect 41694 55806 41746 55858
rect 42366 55806 42418 55858
rect 44494 55806 44546 55858
rect 44830 55806 44882 55858
rect 45502 55806 45554 55858
rect 46734 55806 46786 55858
rect 47406 55806 47458 55858
rect 48078 55806 48130 55858
rect 48414 55806 48466 55858
rect 48750 55806 48802 55858
rect 49422 55806 49474 55858
rect 50878 55806 50930 55858
rect 51214 55806 51266 55858
rect 51550 55806 51602 55858
rect 52222 55806 52274 55858
rect 52894 55806 52946 55858
rect 54350 55806 54402 55858
rect 55358 55806 55410 55858
rect 55694 55806 55746 55858
rect 56030 55806 56082 55858
rect 56254 55806 56306 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 44466 55638 44518 55690
rect 44570 55638 44622 55690
rect 44674 55638 44726 55690
rect 7310 55470 7362 55522
rect 20190 55470 20242 55522
rect 20526 55470 20578 55522
rect 22206 55470 22258 55522
rect 38558 55470 38610 55522
rect 39230 55470 39282 55522
rect 40238 55470 40290 55522
rect 43486 55470 43538 55522
rect 1710 55358 1762 55410
rect 3390 55358 3442 55410
rect 3502 55358 3554 55410
rect 4510 55358 4562 55410
rect 6190 55358 6242 55410
rect 6974 55358 7026 55410
rect 8318 55358 8370 55410
rect 9438 55358 9490 55410
rect 9774 55358 9826 55410
rect 10782 55358 10834 55410
rect 11118 55358 11170 55410
rect 12126 55358 12178 55410
rect 12462 55358 12514 55410
rect 13470 55358 13522 55410
rect 14478 55358 14530 55410
rect 15486 55358 15538 55410
rect 15822 55358 15874 55410
rect 17502 55358 17554 55410
rect 17838 55358 17890 55410
rect 18510 55358 18562 55410
rect 19182 55358 19234 55410
rect 19518 55358 19570 55410
rect 20862 55358 20914 55410
rect 21534 55358 21586 55410
rect 22878 55358 22930 55410
rect 23550 55358 23602 55410
rect 24558 55358 24610 55410
rect 25342 55358 25394 55410
rect 26574 55358 26626 55410
rect 27246 55358 27298 55410
rect 27918 55358 27970 55410
rect 28254 55358 28306 55410
rect 29038 55358 29090 55410
rect 29822 55358 29874 55410
rect 30494 55358 30546 55410
rect 30830 55358 30882 55410
rect 31502 55358 31554 55410
rect 31838 55358 31890 55410
rect 33182 55358 33234 55410
rect 33854 55358 33906 55410
rect 35646 55358 35698 55410
rect 35982 55358 36034 55410
rect 36318 55358 36370 55410
rect 37214 55358 37266 55410
rect 37550 55358 37602 55410
rect 38894 55358 38946 55410
rect 39566 55358 39618 55410
rect 40574 55358 40626 55410
rect 41134 55358 41186 55410
rect 41470 55358 41522 55410
rect 42142 55358 42194 55410
rect 42814 55358 42866 55410
rect 43822 55358 43874 55410
rect 44494 55358 44546 55410
rect 45166 55358 45218 55410
rect 46062 55358 46114 55410
rect 46734 55358 46786 55410
rect 53678 55358 53730 55410
rect 54686 55358 54738 55410
rect 55918 55358 55970 55410
rect 3166 55246 3218 55298
rect 6078 55246 6130 55298
rect 6414 55246 6466 55298
rect 6638 55246 6690 55298
rect 7646 55246 7698 55298
rect 8094 55246 8146 55298
rect 9102 55246 9154 55298
rect 9998 55246 10050 55298
rect 10446 55246 10498 55298
rect 11454 55246 11506 55298
rect 11902 55246 11954 55298
rect 12798 55246 12850 55298
rect 13022 55246 13074 55298
rect 13582 55246 13634 55298
rect 14702 55246 14754 55298
rect 15150 55246 15202 55298
rect 16158 55246 16210 55298
rect 18286 55246 18338 55298
rect 18958 55246 19010 55298
rect 19742 55246 19794 55298
rect 20302 55246 20354 55298
rect 21086 55246 21138 55298
rect 21758 55246 21810 55298
rect 22542 55246 22594 55298
rect 23102 55246 23154 55298
rect 23774 55246 23826 55298
rect 24782 55246 24834 55298
rect 25678 55246 25730 55298
rect 26350 55246 26402 55298
rect 26910 55246 26962 55298
rect 27582 55246 27634 55298
rect 28590 55246 28642 55298
rect 28926 55246 28978 55298
rect 29598 55246 29650 55298
rect 30270 55246 30322 55298
rect 31166 55246 31218 55298
rect 32510 55246 32562 55298
rect 32958 55246 33010 55298
rect 33630 55246 33682 55298
rect 34526 55246 34578 55298
rect 34638 55246 34690 55298
rect 34750 55246 34802 55298
rect 34862 55246 34914 55298
rect 35422 55246 35474 55298
rect 41918 55246 41970 55298
rect 42590 55246 42642 55298
rect 43150 55246 43202 55298
rect 44158 55246 44210 55298
rect 44830 55246 44882 55298
rect 45390 55246 45442 55298
rect 46398 55246 46450 55298
rect 46958 55246 47010 55298
rect 48862 55246 48914 55298
rect 54014 55246 54066 55298
rect 54910 55246 54962 55298
rect 56254 55246 56306 55298
rect 1262 55134 1314 55186
rect 4062 55134 4114 55186
rect 13246 55134 13298 55186
rect 16718 55134 16770 55186
rect 17166 55134 17218 55186
rect 50430 55134 50482 55186
rect 2830 55022 2882 55074
rect 5630 55022 5682 55074
rect 16830 55022 16882 55074
rect 29038 55022 29090 55074
rect 32398 55022 32450 55074
rect 34190 55022 34242 55074
rect 37774 55022 37826 55074
rect 38110 55022 38162 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 43806 54854 43858 54906
rect 43910 54854 43962 54906
rect 44014 54854 44066 54906
rect 29150 54686 29202 54738
rect 33966 54686 34018 54738
rect 38670 54686 38722 54738
rect 12126 54574 12178 54626
rect 48862 54574 48914 54626
rect 2718 54462 2770 54514
rect 4286 54462 4338 54514
rect 5854 54462 5906 54514
rect 6414 54462 6466 54514
rect 7086 54462 7138 54514
rect 7870 54462 7922 54514
rect 8430 54462 8482 54514
rect 9214 54462 9266 54514
rect 11902 54462 11954 54514
rect 12798 54462 12850 54514
rect 13022 54462 13074 54514
rect 13358 54462 13410 54514
rect 16046 54462 16098 54514
rect 18846 54462 18898 54514
rect 19966 54462 20018 54514
rect 21758 54462 21810 54514
rect 23774 54462 23826 54514
rect 26126 54462 26178 54514
rect 27022 54462 27074 54514
rect 29486 54462 29538 54514
rect 30158 54462 30210 54514
rect 30942 54462 30994 54514
rect 32398 54462 32450 54514
rect 34750 54462 34802 54514
rect 34974 54462 35026 54514
rect 36542 54462 36594 54514
rect 39006 54462 39058 54514
rect 41134 54462 41186 54514
rect 42478 54462 42530 54514
rect 42702 54462 42754 54514
rect 44158 54462 44210 54514
rect 44494 54462 44546 54514
rect 45614 54462 45666 54514
rect 46174 54462 46226 54514
rect 53006 54462 53058 54514
rect 1486 54350 1538 54402
rect 2158 54350 2210 54402
rect 3166 54350 3218 54402
rect 5966 54350 6018 54402
rect 8990 54350 9042 54402
rect 10334 54350 10386 54402
rect 11006 54350 11058 54402
rect 11678 54350 11730 54402
rect 12238 54350 12290 54402
rect 13806 54350 13858 54402
rect 16382 54350 16434 54402
rect 18510 54350 18562 54402
rect 19742 54350 19794 54402
rect 21198 54350 21250 54402
rect 22094 54350 22146 54402
rect 22430 54350 22482 54402
rect 28478 54350 28530 54402
rect 30046 54350 30098 54402
rect 31166 54350 31218 54402
rect 31838 54350 31890 54402
rect 35198 54350 35250 54402
rect 35422 54350 35474 54402
rect 36878 54350 36930 54402
rect 39230 54350 39282 54402
rect 39566 54350 39618 54402
rect 40798 54350 40850 54402
rect 42142 54350 42194 54402
rect 43374 54350 43426 54402
rect 44270 54350 44322 54402
rect 45390 54350 45442 54402
rect 51998 54350 52050 54402
rect 52670 54350 52722 54402
rect 54014 54350 54066 54402
rect 1150 54238 1202 54290
rect 1822 54238 1874 54290
rect 5070 54238 5122 54290
rect 5406 54238 5458 54290
rect 6190 54238 6242 54290
rect 6638 54238 6690 54290
rect 7310 54238 7362 54290
rect 7646 54238 7698 54290
rect 8654 54238 8706 54290
rect 9774 54238 9826 54290
rect 10670 54238 10722 54290
rect 11342 54238 11394 54290
rect 13134 54238 13186 54290
rect 13246 54238 13298 54290
rect 14142 54238 14194 54290
rect 14478 54238 14530 54290
rect 15150 54238 15202 54290
rect 15822 54238 15874 54290
rect 17278 54238 17330 54290
rect 19518 54238 19570 54290
rect 20862 54238 20914 54290
rect 21534 54238 21586 54290
rect 21982 54238 22034 54290
rect 22766 54238 22818 54290
rect 23102 54238 23154 54290
rect 23438 54238 23490 54290
rect 23886 54238 23938 54290
rect 24110 54238 24162 54290
rect 24446 54238 24498 54290
rect 25566 54238 25618 54290
rect 27246 54238 27298 54290
rect 27582 54238 27634 54290
rect 27918 54238 27970 54290
rect 28590 54238 28642 54290
rect 28814 54238 28866 54290
rect 31502 54238 31554 54290
rect 32846 54238 32898 54290
rect 35086 54238 35138 54290
rect 38110 54238 38162 54290
rect 40462 54238 40514 54290
rect 41470 54238 41522 54290
rect 41806 54238 41858 54290
rect 43038 54238 43090 54290
rect 43486 54238 43538 54290
rect 43710 54238 43762 54290
rect 44718 54238 44770 54290
rect 45054 54238 45106 54290
rect 52334 54238 52386 54290
rect 53342 54238 53394 54290
rect 53678 54238 53730 54290
rect 54350 54238 54402 54290
rect 55022 54238 55074 54290
rect 55358 54238 55410 54290
rect 56030 54238 56082 54290
rect 56366 54238 56418 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 44466 54070 44518 54122
rect 44570 54070 44622 54122
rect 44674 54070 44726 54122
rect 2158 53902 2210 53954
rect 6078 53902 6130 53954
rect 16158 53902 16210 53954
rect 19294 53902 19346 53954
rect 20862 53902 20914 53954
rect 25678 53902 25730 53954
rect 30158 53902 30210 53954
rect 32510 53902 32562 53954
rect 34190 53902 34242 53954
rect 49422 53902 49474 53954
rect 53230 53902 53282 53954
rect 1486 53790 1538 53842
rect 2494 53790 2546 53842
rect 3726 53790 3778 53842
rect 9662 53790 9714 53842
rect 13694 53790 13746 53842
rect 15150 53790 15202 53842
rect 17390 53790 17442 53842
rect 20078 53790 20130 53842
rect 21758 53790 21810 53842
rect 22654 53790 22706 53842
rect 23326 53790 23378 53842
rect 28030 53790 28082 53842
rect 29038 53790 29090 53842
rect 30830 53790 30882 53842
rect 31838 53790 31890 53842
rect 32398 53790 32450 53842
rect 35758 53790 35810 53842
rect 38222 53790 38274 53842
rect 41582 53790 41634 53842
rect 43150 53790 43202 53842
rect 45502 53790 45554 53842
rect 46174 53790 46226 53842
rect 46510 53790 46562 53842
rect 47182 53790 47234 53842
rect 48414 53790 48466 53842
rect 49086 53790 49138 53842
rect 50206 53790 50258 53842
rect 50542 53790 50594 53842
rect 51214 53790 51266 53842
rect 51886 53790 51938 53842
rect 52894 53790 52946 53842
rect 54238 53790 54290 53842
rect 55358 53790 55410 53842
rect 56366 53790 56418 53842
rect 1150 53678 1202 53730
rect 1934 53678 1986 53730
rect 2718 53678 2770 53730
rect 9998 53678 10050 53730
rect 11678 53678 11730 53730
rect 12462 53678 12514 53730
rect 13022 53678 13074 53730
rect 13918 53678 13970 53730
rect 14254 53678 14306 53730
rect 15486 53678 15538 53730
rect 15822 53678 15874 53730
rect 19518 53678 19570 53730
rect 19966 53678 20018 53730
rect 20638 53678 20690 53730
rect 22094 53678 22146 53730
rect 22990 53678 23042 53730
rect 23550 53678 23602 53730
rect 24446 53678 24498 53730
rect 24670 53678 24722 53730
rect 24782 53678 24834 53730
rect 25006 53678 25058 53730
rect 25454 53678 25506 53730
rect 25902 53678 25954 53730
rect 26126 53678 26178 53730
rect 26350 53678 26402 53730
rect 26798 53678 26850 53730
rect 27022 53678 27074 53730
rect 27806 53678 27858 53730
rect 31166 53678 31218 53730
rect 31502 53678 31554 53730
rect 32734 53678 32786 53730
rect 41806 53678 41858 53730
rect 44718 53678 44770 53730
rect 45278 53678 45330 53730
rect 45950 53678 46002 53730
rect 46734 53678 46786 53730
rect 47518 53678 47570 53730
rect 48190 53678 48242 53730
rect 49870 53678 49922 53730
rect 50766 53678 50818 53730
rect 51550 53678 51602 53730
rect 52110 53678 52162 53730
rect 52558 53678 52610 53730
rect 53566 53678 53618 53730
rect 53902 53678 53954 53730
rect 55022 53678 55074 53730
rect 56030 53678 56082 53730
rect 3390 53566 3442 53618
rect 5630 53566 5682 53618
rect 7646 53566 7698 53618
rect 7982 53566 8034 53618
rect 8318 53566 8370 53618
rect 8990 53566 9042 53618
rect 10334 53566 10386 53618
rect 11006 53566 11058 53618
rect 14702 53566 14754 53618
rect 16942 53566 16994 53618
rect 21198 53566 21250 53618
rect 22430 53566 22482 53618
rect 25790 53566 25842 53618
rect 26574 53566 26626 53618
rect 28590 53566 28642 53618
rect 34638 53566 34690 53618
rect 35422 53566 35474 53618
rect 37774 53566 37826 53618
rect 42702 53566 42754 53618
rect 44830 53566 44882 53618
rect 4958 53454 5010 53506
rect 7198 53454 7250 53506
rect 7870 53454 7922 53506
rect 18510 53454 18562 53506
rect 20078 53454 20130 53506
rect 33070 53454 33122 53506
rect 36990 53454 37042 53506
rect 39342 53454 39394 53506
rect 40686 53454 40738 53506
rect 41022 53454 41074 53506
rect 44270 53454 44322 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 43806 53286 43858 53338
rect 43910 53286 43962 53338
rect 44014 53286 44066 53338
rect 9886 53118 9938 53170
rect 20078 53118 20130 53170
rect 23102 53118 23154 53170
rect 31726 53118 31778 53170
rect 32062 53118 32114 53170
rect 32174 53118 32226 53170
rect 34302 53118 34354 53170
rect 52670 53118 52722 53170
rect 1262 53006 1314 53058
rect 6190 53006 6242 53058
rect 10558 53006 10610 53058
rect 15710 53006 15762 53058
rect 19966 53006 20018 53058
rect 25230 53006 25282 53058
rect 27358 53006 27410 53058
rect 32734 53006 32786 53058
rect 37102 53006 37154 53058
rect 6526 52894 6578 52946
rect 7086 52894 7138 52946
rect 7646 52894 7698 52946
rect 8318 52894 8370 52946
rect 9326 52894 9378 52946
rect 12126 52894 12178 52946
rect 13134 52894 13186 52946
rect 16046 52894 16098 52946
rect 16494 52894 16546 52946
rect 17390 52894 17442 52946
rect 17726 52894 17778 52946
rect 18734 52894 18786 52946
rect 20862 52894 20914 52946
rect 21646 52894 21698 52946
rect 24670 52894 24722 52946
rect 30270 52894 30322 52946
rect 31614 52894 31666 52946
rect 31838 52894 31890 52946
rect 34750 52894 34802 52946
rect 35086 52894 35138 52946
rect 35198 52894 35250 52946
rect 37438 52894 37490 52946
rect 37998 52894 38050 52946
rect 38670 52894 38722 52946
rect 39342 52894 39394 52946
rect 40126 52894 40178 52946
rect 43374 52894 43426 52946
rect 44158 52894 44210 52946
rect 44382 52894 44434 52946
rect 44718 52894 44770 52946
rect 46062 52894 46114 52946
rect 54686 52894 54738 52946
rect 1598 52782 1650 52834
rect 3726 52782 3778 52834
rect 4062 52782 4114 52834
rect 5294 52782 5346 52834
rect 5518 52782 5570 52834
rect 5854 52782 5906 52834
rect 9998 52782 10050 52834
rect 10894 52782 10946 52834
rect 21982 52782 22034 52834
rect 30942 52782 30994 52834
rect 41022 52782 41074 52834
rect 42926 52782 42978 52834
rect 45054 52782 45106 52834
rect 45278 52782 45330 52834
rect 48414 52782 48466 52834
rect 52334 52782 52386 52834
rect 2830 52670 2882 52722
rect 3390 52670 3442 52722
rect 4398 52670 4450 52722
rect 5630 52670 5682 52722
rect 7198 52670 7250 52722
rect 9886 52670 9938 52722
rect 13582 52670 13634 52722
rect 14702 52670 14754 52722
rect 15150 52670 15202 52722
rect 16718 52670 16770 52722
rect 19294 52670 19346 52722
rect 19742 52670 19794 52722
rect 20638 52670 20690 52722
rect 21310 52670 21362 52722
rect 22318 52670 22370 52722
rect 24222 52670 24274 52722
rect 25342 52670 25394 52722
rect 25790 52670 25842 52722
rect 26910 52670 26962 52722
rect 28590 52670 28642 52722
rect 29710 52670 29762 52722
rect 31278 52670 31330 52722
rect 33182 52670 33234 52722
rect 35310 52670 35362 52722
rect 35422 52670 35474 52722
rect 36430 52670 36482 52722
rect 36766 52670 36818 52722
rect 38110 52670 38162 52722
rect 41358 52670 41410 52722
rect 41806 52670 41858 52722
rect 44606 52670 44658 52722
rect 45166 52670 45218 52722
rect 46622 52670 46674 52722
rect 47742 52670 47794 52722
rect 48750 52670 48802 52722
rect 49198 52670 49250 52722
rect 49534 52670 49586 52722
rect 50206 52670 50258 52722
rect 50542 52670 50594 52722
rect 50878 52670 50930 52722
rect 51214 52670 51266 52722
rect 51998 52670 52050 52722
rect 52782 52670 52834 52722
rect 52894 52670 52946 52722
rect 53342 52670 53394 52722
rect 53678 52670 53730 52722
rect 54350 52670 54402 52722
rect 55022 52670 55074 52722
rect 55358 52670 55410 52722
rect 56030 52670 56082 52722
rect 56366 52670 56418 52722
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 44466 52502 44518 52554
rect 44570 52502 44622 52554
rect 44674 52502 44726 52554
rect 3502 52334 3554 52386
rect 3838 52334 3890 52386
rect 5966 52334 6018 52386
rect 7086 52334 7138 52386
rect 8990 52334 9042 52386
rect 11118 52334 11170 52386
rect 12574 52334 12626 52386
rect 15262 52334 15314 52386
rect 22766 52334 22818 52386
rect 25902 52334 25954 52386
rect 31166 52334 31218 52386
rect 39566 52334 39618 52386
rect 42030 52334 42082 52386
rect 46510 52334 46562 52386
rect 50654 52334 50706 52386
rect 56030 52334 56082 52386
rect 1598 52222 1650 52274
rect 4734 52222 4786 52274
rect 8878 52222 8930 52274
rect 9998 52222 10050 52274
rect 15598 52222 15650 52274
rect 18958 52222 19010 52274
rect 20862 52222 20914 52274
rect 21198 52222 21250 52274
rect 23886 52222 23938 52274
rect 24894 52222 24946 52274
rect 29486 52222 29538 52274
rect 31502 52222 31554 52274
rect 31838 52222 31890 52274
rect 33742 52222 33794 52274
rect 34638 52222 34690 52274
rect 34750 52222 34802 52274
rect 35870 52222 35922 52274
rect 38334 52222 38386 52274
rect 40910 52222 40962 52274
rect 42926 52222 42978 52274
rect 46846 52222 46898 52274
rect 47518 52222 47570 52274
rect 49534 52222 49586 52274
rect 50094 52222 50146 52274
rect 50206 52222 50258 52274
rect 51886 52222 51938 52274
rect 53118 52222 53170 52274
rect 53678 52222 53730 52274
rect 54350 52222 54402 52274
rect 55358 52222 55410 52274
rect 56366 52222 56418 52274
rect 1262 52110 1314 52162
rect 4286 52110 4338 52162
rect 6638 52110 6690 52162
rect 8206 52110 8258 52162
rect 12014 52110 12066 52162
rect 12462 52110 12514 52162
rect 13246 52110 13298 52162
rect 13694 52110 13746 52162
rect 14702 52110 14754 52162
rect 15150 52110 15202 52162
rect 15934 52110 15986 52162
rect 16270 52110 16322 52162
rect 16830 52110 16882 52162
rect 17950 52110 18002 52162
rect 18286 52110 18338 52162
rect 19182 52110 19234 52162
rect 19518 52110 19570 52162
rect 19966 52110 20018 52162
rect 20414 52110 20466 52162
rect 20526 52110 20578 52162
rect 21534 52110 21586 52162
rect 22318 52110 22370 52162
rect 25230 52110 25282 52162
rect 25678 52110 25730 52162
rect 26350 52110 26402 52162
rect 26910 52110 26962 52162
rect 27918 52110 27970 52162
rect 28926 52110 28978 52162
rect 31054 52110 31106 52162
rect 32510 52110 32562 52162
rect 34078 52110 34130 52162
rect 40462 52110 40514 52162
rect 42590 52110 42642 52162
rect 45390 52110 45442 52162
rect 46174 52110 46226 52162
rect 47294 52110 47346 52162
rect 48190 52110 48242 52162
rect 49870 52110 49922 52162
rect 52894 52110 52946 52162
rect 54014 52110 54066 52162
rect 54686 52110 54738 52162
rect 55134 52110 55186 52162
rect 9550 51998 9602 52050
rect 11566 51998 11618 52050
rect 16046 51998 16098 52050
rect 20750 51998 20802 52050
rect 35422 51998 35474 52050
rect 37998 51998 38050 52050
rect 43262 51998 43314 52050
rect 49422 51998 49474 52050
rect 52222 51998 52274 52050
rect 2830 51886 2882 51938
rect 30606 51886 30658 51938
rect 34750 51886 34802 51938
rect 36990 51886 37042 51938
rect 48414 51886 48466 51938
rect 48750 51886 48802 51938
rect 49310 51886 49362 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 43806 51718 43858 51770
rect 43910 51718 43962 51770
rect 44014 51718 44066 51770
rect 3838 51550 3890 51602
rect 11678 51550 11730 51602
rect 28702 51550 28754 51602
rect 34638 51550 34690 51602
rect 42254 51550 42306 51602
rect 42702 51550 42754 51602
rect 43262 51550 43314 51602
rect 43486 51550 43538 51602
rect 49646 51550 49698 51602
rect 50430 51550 50482 51602
rect 4398 51438 4450 51490
rect 10110 51438 10162 51490
rect 12126 51438 12178 51490
rect 20974 51438 21026 51490
rect 21870 51438 21922 51490
rect 33070 51438 33122 51490
rect 36430 51438 36482 51490
rect 36654 51438 36706 51490
rect 37662 51438 37714 51490
rect 46398 51438 46450 51490
rect 48526 51438 48578 51490
rect 49870 51438 49922 51490
rect 1262 51326 1314 51378
rect 1374 51326 1426 51378
rect 4174 51326 4226 51378
rect 5406 51326 5458 51378
rect 5518 51326 5570 51378
rect 5966 51326 6018 51378
rect 6750 51326 6802 51378
rect 7086 51326 7138 51378
rect 7758 51326 7810 51378
rect 8430 51326 8482 51378
rect 9326 51326 9378 51378
rect 13134 51326 13186 51378
rect 13582 51326 13634 51378
rect 14254 51326 14306 51378
rect 15038 51326 15090 51378
rect 15822 51326 15874 51378
rect 17166 51326 17218 51378
rect 17614 51326 17666 51378
rect 18398 51326 18450 51378
rect 18846 51326 18898 51378
rect 19854 51326 19906 51378
rect 20638 51326 20690 51378
rect 23998 51326 24050 51378
rect 24670 51326 24722 51378
rect 25118 51326 25170 51378
rect 25454 51326 25506 51378
rect 26350 51326 26402 51378
rect 26798 51326 26850 51378
rect 27694 51326 27746 51378
rect 28590 51326 28642 51378
rect 29486 51326 29538 51378
rect 30046 51326 30098 51378
rect 30606 51326 30658 51378
rect 31166 51326 31218 51378
rect 32174 51326 32226 51378
rect 35086 51326 35138 51378
rect 35422 51326 35474 51378
rect 40686 51326 40738 51378
rect 42814 51326 42866 51378
rect 44494 51326 44546 51378
rect 44718 51326 44770 51378
rect 44942 51326 44994 51378
rect 45278 51326 45330 51378
rect 45726 51326 45778 51378
rect 49198 51326 49250 51378
rect 50206 51326 50258 51378
rect 50990 51326 51042 51378
rect 51102 51326 51154 51378
rect 51326 51326 51378 51378
rect 51438 51326 51490 51378
rect 52110 51326 52162 51378
rect 52670 51326 52722 51378
rect 53342 51326 53394 51378
rect 1822 51214 1874 51266
rect 3390 51214 3442 51266
rect 6302 51214 6354 51266
rect 7310 51214 7362 51266
rect 10558 51214 10610 51266
rect 12798 51214 12850 51266
rect 13806 51214 13858 51266
rect 16494 51214 16546 51266
rect 16830 51214 16882 51266
rect 17838 51214 17890 51266
rect 24222 51214 24274 51266
rect 24334 51214 24386 51266
rect 25678 51214 25730 51266
rect 29150 51214 29202 51266
rect 30158 51214 30210 51266
rect 36318 51214 36370 51266
rect 36542 51214 36594 51266
rect 38110 51214 38162 51266
rect 39790 51214 39842 51266
rect 41134 51214 41186 51266
rect 49870 51214 49922 51266
rect 52334 51214 52386 51266
rect 53006 51214 53058 51266
rect 54574 51214 54626 51266
rect 54910 51214 54962 51266
rect 2942 51102 2994 51154
rect 3502 51102 3554 51154
rect 5630 51102 5682 51154
rect 5742 51102 5794 51154
rect 12238 51102 12290 51154
rect 16382 51102 16434 51154
rect 20862 51102 20914 51154
rect 21086 51102 21138 51154
rect 21198 51102 21250 51154
rect 22318 51102 22370 51154
rect 23438 51102 23490 51154
rect 28702 51102 28754 51154
rect 33518 51102 33570 51154
rect 35198 51102 35250 51154
rect 35534 51102 35586 51154
rect 35646 51102 35698 51154
rect 39230 51102 39282 51154
rect 40126 51102 40178 51154
rect 43598 51102 43650 51154
rect 44270 51102 44322 51154
rect 44382 51102 44434 51154
rect 45614 51102 45666 51154
rect 45838 51102 45890 51154
rect 52894 51102 52946 51154
rect 53678 51102 53730 51154
rect 54238 51102 54290 51154
rect 55246 51102 55298 51154
rect 55582 51102 55634 51154
rect 56030 51102 56082 51154
rect 56366 51102 56418 51154
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 44466 50934 44518 50986
rect 44570 50934 44622 50986
rect 44674 50934 44726 50986
rect 9550 50766 9602 50818
rect 12350 50766 12402 50818
rect 25566 50766 25618 50818
rect 29598 50766 29650 50818
rect 35982 50766 36034 50818
rect 42814 50766 42866 50818
rect 46286 50766 46338 50818
rect 51998 50766 52050 50818
rect 53454 50766 53506 50818
rect 54462 50766 54514 50818
rect 55358 50766 55410 50818
rect 1598 50654 1650 50706
rect 4734 50654 4786 50706
rect 6862 50654 6914 50706
rect 7310 50654 7362 50706
rect 14926 50654 14978 50706
rect 18062 50654 18114 50706
rect 18510 50654 18562 50706
rect 20750 50654 20802 50706
rect 21758 50654 21810 50706
rect 28590 50654 28642 50706
rect 33742 50654 33794 50706
rect 35086 50654 35138 50706
rect 35422 50654 35474 50706
rect 36430 50654 36482 50706
rect 37438 50654 37490 50706
rect 37886 50654 37938 50706
rect 41582 50654 41634 50706
rect 43934 50654 43986 50706
rect 45054 50654 45106 50706
rect 47406 50654 47458 50706
rect 49086 50654 49138 50706
rect 49646 50654 49698 50706
rect 50766 50654 50818 50706
rect 52894 50654 52946 50706
rect 56366 50654 56418 50706
rect 3502 50542 3554 50594
rect 3838 50542 3890 50594
rect 3950 50542 4002 50594
rect 4510 50542 4562 50594
rect 5294 50542 5346 50594
rect 6078 50542 6130 50594
rect 7534 50542 7586 50594
rect 7982 50542 8034 50594
rect 8318 50542 8370 50594
rect 9102 50542 9154 50594
rect 11342 50542 11394 50594
rect 11790 50542 11842 50594
rect 12238 50542 12290 50594
rect 13022 50542 13074 50594
rect 13470 50542 13522 50594
rect 14478 50542 14530 50594
rect 15262 50542 15314 50594
rect 15598 50542 15650 50594
rect 15822 50542 15874 50594
rect 16158 50542 16210 50594
rect 17390 50542 17442 50594
rect 17838 50542 17890 50594
rect 19070 50542 19122 50594
rect 20078 50542 20130 50594
rect 21198 50542 21250 50594
rect 21534 50542 21586 50594
rect 22430 50542 22482 50594
rect 22766 50542 22818 50594
rect 23774 50542 23826 50594
rect 25006 50542 25058 50594
rect 25342 50542 25394 50594
rect 26238 50542 26290 50594
rect 26574 50542 26626 50594
rect 27582 50542 27634 50594
rect 28926 50542 28978 50594
rect 29374 50542 29426 50594
rect 30270 50542 30322 50594
rect 30830 50542 30882 50594
rect 31726 50542 31778 50594
rect 34078 50542 34130 50594
rect 35646 50542 35698 50594
rect 36766 50542 36818 50594
rect 37214 50542 37266 50594
rect 38670 50542 38722 50594
rect 39566 50542 39618 50594
rect 40350 50542 40402 50594
rect 41918 50542 41970 50594
rect 45278 50542 45330 50594
rect 48526 50542 48578 50594
rect 48862 50542 48914 50594
rect 53678 50542 53730 50594
rect 55022 50542 55074 50594
rect 56142 50542 56194 50594
rect 1262 50430 1314 50482
rect 2830 50430 2882 50482
rect 3614 50430 3666 50482
rect 16046 50430 16098 50482
rect 17054 50430 17106 50482
rect 24558 50430 24610 50482
rect 44382 50430 44434 50482
rect 44942 50430 44994 50482
rect 45838 50430 45890 50482
rect 50430 50430 50482 50482
rect 52782 50430 52834 50482
rect 54238 50430 54290 50482
rect 54574 50430 54626 50482
rect 10670 50318 10722 50370
rect 32510 50318 32562 50370
rect 53118 50318 53170 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 43806 50150 43858 50202
rect 43910 50150 43962 50202
rect 44014 50150 44066 50202
rect 22654 49982 22706 50034
rect 35086 49982 35138 50034
rect 35422 49982 35474 50034
rect 36430 49982 36482 50034
rect 43374 49982 43426 50034
rect 47518 49982 47570 50034
rect 48750 49982 48802 50034
rect 13134 49870 13186 49922
rect 21086 49870 21138 49922
rect 32286 49870 32338 49922
rect 39230 49870 39282 49922
rect 44606 49870 44658 49922
rect 1262 49758 1314 49810
rect 3166 49758 3218 49810
rect 4398 49758 4450 49810
rect 5630 49758 5682 49810
rect 5966 49758 6018 49810
rect 6750 49758 6802 49810
rect 7198 49758 7250 49810
rect 8318 49758 8370 49810
rect 9214 49758 9266 49810
rect 10110 49758 10162 49810
rect 10558 49758 10610 49810
rect 11342 49758 11394 49810
rect 11790 49758 11842 49810
rect 14702 49758 14754 49810
rect 15486 49758 15538 49810
rect 15934 49758 15986 49810
rect 16718 49758 16770 49810
rect 17390 49758 17442 49810
rect 18174 49758 18226 49810
rect 19182 49758 19234 49810
rect 23774 49758 23826 49810
rect 24222 49758 24274 49810
rect 25118 49758 25170 49810
rect 25566 49758 25618 49810
rect 26462 49758 26514 49810
rect 29822 49758 29874 49810
rect 30046 49758 30098 49810
rect 30270 49758 30322 49810
rect 32958 49758 33010 49810
rect 34526 49758 34578 49810
rect 35646 49758 35698 49810
rect 38110 49758 38162 49810
rect 41694 49758 41746 49810
rect 44494 49758 44546 49810
rect 44718 49758 44770 49810
rect 45278 49758 45330 49810
rect 46846 49758 46898 49810
rect 47294 49758 47346 49810
rect 47854 49758 47906 49810
rect 48078 49758 48130 49810
rect 48974 49758 49026 49810
rect 50206 49758 50258 49810
rect 50990 49758 51042 49810
rect 51214 49758 51266 49810
rect 51326 49758 51378 49810
rect 53006 49758 53058 49810
rect 1598 49646 1650 49698
rect 3502 49646 3554 49698
rect 3838 49646 3890 49698
rect 4174 49646 4226 49698
rect 5182 49646 5234 49698
rect 6190 49646 6242 49698
rect 12238 49646 12290 49698
rect 15150 49646 15202 49698
rect 16158 49646 16210 49698
rect 19406 49646 19458 49698
rect 19966 49646 20018 49698
rect 21534 49646 21586 49698
rect 23438 49646 23490 49698
rect 24446 49646 24498 49698
rect 29598 49646 29650 49698
rect 30718 49646 30770 49698
rect 31838 49646 31890 49698
rect 37662 49646 37714 49698
rect 38558 49646 38610 49698
rect 42142 49646 42194 49698
rect 44158 49646 44210 49698
rect 47966 49646 48018 49698
rect 49646 49646 49698 49698
rect 50430 49646 50482 49698
rect 50878 49646 50930 49698
rect 2830 49534 2882 49586
rect 3390 49534 3442 49586
rect 4062 49534 4114 49586
rect 11230 49534 11282 49586
rect 13582 49534 13634 49586
rect 18846 49534 18898 49586
rect 29710 49534 29762 49586
rect 34078 49534 34130 49586
rect 38670 49534 38722 49586
rect 39678 49534 39730 49586
rect 40798 49534 40850 49586
rect 45726 49534 45778 49586
rect 48414 49534 48466 49586
rect 49422 49534 49474 49586
rect 49534 49534 49586 49586
rect 51998 49534 52050 49586
rect 52334 49534 52386 49586
rect 53566 49534 53618 49586
rect 54686 49534 54738 49586
rect 55246 49534 55298 49586
rect 55582 49534 55634 49586
rect 55918 49534 55970 49586
rect 56254 49534 56306 49586
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 44466 49366 44518 49418
rect 44570 49366 44622 49418
rect 44674 49366 44726 49418
rect 1150 49198 1202 49250
rect 1486 49198 1538 49250
rect 1822 49198 1874 49250
rect 2158 49198 2210 49250
rect 3502 49198 3554 49250
rect 7086 49198 7138 49250
rect 16046 49198 16098 49250
rect 25118 49198 25170 49250
rect 30606 49198 30658 49250
rect 30830 49198 30882 49250
rect 31390 49198 31442 49250
rect 34750 49198 34802 49250
rect 35870 49198 35922 49250
rect 39678 49198 39730 49250
rect 40910 49198 40962 49250
rect 47182 49198 47234 49250
rect 48974 49198 49026 49250
rect 55358 49198 55410 49250
rect 56366 49198 56418 49250
rect 3950 49086 4002 49138
rect 9326 49086 9378 49138
rect 10334 49086 10386 49138
rect 13806 49086 13858 49138
rect 18062 49086 18114 49138
rect 19182 49086 19234 49138
rect 21758 49086 21810 49138
rect 25790 49086 25842 49138
rect 26238 49086 26290 49138
rect 27694 49086 27746 49138
rect 33630 49086 33682 49138
rect 37438 49086 37490 49138
rect 45278 49086 45330 49138
rect 46510 49086 46562 49138
rect 50094 49086 50146 49138
rect 53006 49086 53058 49138
rect 54350 49086 54402 49138
rect 2942 48974 2994 49026
rect 3390 48974 3442 49026
rect 4510 48974 4562 49026
rect 5518 48974 5570 49026
rect 8206 48974 8258 49026
rect 9774 48974 9826 49026
rect 10110 48974 10162 49026
rect 10782 48974 10834 49026
rect 11342 48974 11394 49026
rect 12462 48974 12514 49026
rect 13246 48974 13298 49026
rect 15486 48974 15538 49026
rect 15710 48974 15762 49026
rect 15934 48974 15986 49026
rect 17278 48974 17330 49026
rect 17950 48974 18002 49026
rect 18734 48974 18786 49026
rect 21086 48974 21138 49026
rect 21534 48974 21586 49026
rect 22430 48974 22482 49026
rect 22766 48974 22818 49026
rect 23774 48974 23826 49026
rect 27022 48974 27074 49026
rect 27582 48974 27634 49026
rect 28366 48974 28418 49026
rect 28702 48974 28754 49026
rect 29710 48974 29762 49026
rect 30494 48974 30546 49026
rect 31166 48974 31218 49026
rect 34190 48974 34242 49026
rect 37102 48974 37154 49026
rect 39454 48974 39506 49026
rect 40350 48974 40402 49026
rect 42478 48974 42530 49026
rect 46062 48974 46114 49026
rect 46622 48974 46674 49026
rect 46734 48974 46786 49026
rect 48302 48974 48354 49026
rect 48638 48974 48690 49026
rect 48862 48974 48914 49026
rect 53454 48974 53506 49026
rect 54014 48974 54066 49026
rect 55022 48974 55074 49026
rect 56030 48974 56082 49026
rect 2494 48862 2546 48914
rect 6638 48862 6690 48914
rect 8990 48862 9042 48914
rect 14926 48862 14978 48914
rect 16046 48862 16098 48914
rect 20750 48862 20802 48914
rect 26686 48862 26738 48914
rect 31278 48862 31330 48914
rect 31614 48862 31666 48914
rect 36318 48862 36370 48914
rect 43150 48862 43202 48914
rect 49758 48862 49810 48914
rect 8878 48750 8930 48802
rect 16942 48750 16994 48802
rect 20302 48750 20354 48802
rect 25454 48750 25506 48802
rect 31838 48750 31890 48802
rect 32510 48750 32562 48802
rect 38670 48750 38722 48802
rect 42030 48750 42082 48802
rect 42478 48750 42530 48802
rect 42814 48750 42866 48802
rect 48078 48750 48130 48802
rect 51326 48750 51378 48802
rect 51886 48750 51938 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 43806 48582 43858 48634
rect 43910 48582 43962 48634
rect 44014 48582 44066 48634
rect 20750 48414 20802 48466
rect 36654 48414 36706 48466
rect 43038 48414 43090 48466
rect 1150 48302 1202 48354
rect 4958 48302 5010 48354
rect 13246 48302 13298 48354
rect 15262 48302 15314 48354
rect 33966 48302 34018 48354
rect 35086 48302 35138 48354
rect 46958 48302 47010 48354
rect 49086 48302 49138 48354
rect 1598 48190 1650 48242
rect 1934 48190 1986 48242
rect 2718 48190 2770 48242
rect 3166 48190 3218 48242
rect 4174 48185 4226 48237
rect 5294 48190 5346 48242
rect 5742 48190 5794 48242
rect 6414 48190 6466 48242
rect 6974 48190 7026 48242
rect 7198 48190 7250 48242
rect 7982 48190 8034 48242
rect 9438 48190 9490 48242
rect 9774 48190 9826 48242
rect 10558 48190 10610 48242
rect 11230 48190 11282 48242
rect 12126 48190 12178 48242
rect 15598 48190 15650 48242
rect 16046 48190 16098 48242
rect 16830 48190 16882 48242
rect 17278 48190 17330 48242
rect 18286 48190 18338 48242
rect 20638 48190 20690 48242
rect 21646 48190 21698 48242
rect 23998 48190 24050 48242
rect 26238 48190 26290 48242
rect 30270 48190 30322 48242
rect 34862 48190 34914 48242
rect 35534 48190 35586 48242
rect 36430 48190 36482 48242
rect 37102 48190 37154 48242
rect 38110 48190 38162 48242
rect 38558 48190 38610 48242
rect 39790 48190 39842 48242
rect 40798 48190 40850 48242
rect 41358 48190 41410 48242
rect 43598 48190 43650 48242
rect 44382 48190 44434 48242
rect 44942 48190 44994 48242
rect 49870 48190 49922 48242
rect 50654 48190 50706 48242
rect 50878 48190 50930 48242
rect 51102 48190 51154 48242
rect 52110 48190 52162 48242
rect 54798 48190 54850 48242
rect 55582 48190 55634 48242
rect 56142 48190 56194 48242
rect 2158 48078 2210 48130
rect 5966 48078 6018 48130
rect 8654 48078 8706 48130
rect 8990 48078 9042 48130
rect 9998 48078 10050 48130
rect 22094 48078 22146 48130
rect 24334 48078 24386 48130
rect 26574 48078 26626 48130
rect 30718 48078 30770 48130
rect 36878 48078 36930 48130
rect 37214 48078 37266 48130
rect 37662 48078 37714 48130
rect 39118 48078 39170 48130
rect 41806 48078 41858 48130
rect 45278 48078 45330 48130
rect 50206 48078 50258 48130
rect 50318 48078 50370 48130
rect 54238 48078 54290 48130
rect 55022 48078 55074 48130
rect 8542 47966 8594 48018
rect 13694 47966 13746 48018
rect 14814 47966 14866 48018
rect 16270 47966 16322 48018
rect 18846 47966 18898 48018
rect 19182 47966 19234 48018
rect 19518 47966 19570 48018
rect 19854 47966 19906 48018
rect 20078 47966 20130 48018
rect 20750 47966 20802 48018
rect 23326 47966 23378 48018
rect 25566 47966 25618 48018
rect 27806 47966 27858 48018
rect 31838 47966 31890 48018
rect 32398 47966 32450 48018
rect 33518 47966 33570 48018
rect 35310 47966 35362 48018
rect 35422 47966 35474 48018
rect 38670 47966 38722 48018
rect 43486 47966 43538 48018
rect 44046 47966 44098 48018
rect 44270 47966 44322 48018
rect 46510 47966 46562 48018
rect 51550 47966 51602 48018
rect 52670 47966 52722 48018
rect 53790 47966 53842 48018
rect 54350 47966 54402 48018
rect 55358 47966 55410 48018
rect 56366 47966 56418 48018
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 44466 47798 44518 47850
rect 44570 47798 44622 47850
rect 44674 47798 44726 47850
rect 2830 47630 2882 47682
rect 3390 47630 3442 47682
rect 18062 47630 18114 47682
rect 27694 47630 27746 47682
rect 31390 47630 31442 47682
rect 37886 47630 37938 47682
rect 41022 47630 41074 47682
rect 41358 47630 41410 47682
rect 44270 47630 44322 47682
rect 45726 47630 45778 47682
rect 48078 47630 48130 47682
rect 50766 47630 50818 47682
rect 55134 47630 55186 47682
rect 1598 47518 1650 47570
rect 3726 47518 3778 47570
rect 5070 47518 5122 47570
rect 7758 47518 7810 47570
rect 8318 47518 8370 47570
rect 9102 47518 9154 47570
rect 10110 47518 10162 47570
rect 10558 47518 10610 47570
rect 15150 47518 15202 47570
rect 17166 47518 17218 47570
rect 19070 47518 19122 47570
rect 20302 47518 20354 47570
rect 21758 47518 21810 47570
rect 25342 47518 25394 47570
rect 25678 47518 25730 47570
rect 28142 47518 28194 47570
rect 30382 47518 30434 47570
rect 33070 47518 33122 47570
rect 33406 47518 33458 47570
rect 33966 47518 34018 47570
rect 34526 47518 34578 47570
rect 35646 47518 35698 47570
rect 36654 47518 36706 47570
rect 38334 47518 38386 47570
rect 38446 47518 38498 47570
rect 38558 47518 38610 47570
rect 41694 47518 41746 47570
rect 42030 47518 42082 47570
rect 46846 47518 46898 47570
rect 49534 47518 49586 47570
rect 51214 47518 51266 47570
rect 52222 47518 52274 47570
rect 56366 47518 56418 47570
rect 4398 47406 4450 47458
rect 4958 47406 5010 47458
rect 5630 47406 5682 47458
rect 6190 47406 6242 47458
rect 7086 47406 7138 47458
rect 7982 47406 8034 47458
rect 9438 47406 9490 47458
rect 9886 47406 9938 47458
rect 11342 47406 11394 47458
rect 12126 47406 12178 47458
rect 13022 47406 13074 47458
rect 13918 47406 13970 47458
rect 14702 47406 14754 47458
rect 15262 47406 15314 47458
rect 15710 47406 15762 47458
rect 17278 47406 17330 47458
rect 17726 47406 17778 47458
rect 18734 47406 18786 47458
rect 21086 47406 21138 47458
rect 21646 47406 21698 47458
rect 22430 47406 22482 47458
rect 22766 47406 22818 47458
rect 23774 47406 23826 47458
rect 25006 47406 25058 47458
rect 27022 47406 27074 47458
rect 27582 47406 27634 47458
rect 28366 47406 28418 47458
rect 28702 47406 28754 47458
rect 29710 47406 29762 47458
rect 30718 47406 30770 47458
rect 31166 47406 31218 47458
rect 31278 47406 31330 47458
rect 31614 47406 31666 47458
rect 31838 47406 31890 47458
rect 33630 47406 33682 47458
rect 35310 47406 35362 47458
rect 39118 47406 39170 47458
rect 39454 47406 39506 47458
rect 39566 47406 39618 47458
rect 40238 47406 40290 47458
rect 40798 47406 40850 47458
rect 42366 47406 42418 47458
rect 42478 47406 42530 47458
rect 44830 47406 44882 47458
rect 47406 47406 47458 47458
rect 48302 47406 48354 47458
rect 48638 47406 48690 47458
rect 51550 47406 51602 47458
rect 51998 47406 52050 47458
rect 52894 47406 52946 47458
rect 53454 47406 53506 47458
rect 54350 47406 54402 47458
rect 54798 47406 54850 47458
rect 56030 47406 56082 47458
rect 1262 47294 1314 47346
rect 4062 47294 4114 47346
rect 8206 47294 8258 47346
rect 16158 47294 16210 47346
rect 20750 47294 20802 47346
rect 26686 47294 26738 47346
rect 36318 47294 36370 47346
rect 39230 47294 39282 47346
rect 40350 47294 40402 47346
rect 42142 47294 42194 47346
rect 48190 47294 48242 47346
rect 49198 47294 49250 47346
rect 24670 47182 24722 47234
rect 30718 47182 30770 47234
rect 34862 47182 34914 47234
rect 43150 47182 43202 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 43806 47014 43858 47066
rect 43910 47014 43962 47066
rect 44014 47014 44066 47066
rect 19182 46846 19234 46898
rect 20750 46846 20802 46898
rect 23326 46846 23378 46898
rect 29262 46846 29314 46898
rect 35086 46846 35138 46898
rect 36430 46846 36482 46898
rect 39790 46846 39842 46898
rect 48750 46846 48802 46898
rect 51326 46846 51378 46898
rect 1262 46734 1314 46786
rect 15150 46734 15202 46786
rect 26238 46734 26290 46786
rect 29150 46734 29202 46786
rect 32958 46734 33010 46786
rect 36766 46734 36818 46786
rect 42702 46734 42754 46786
rect 42926 46734 42978 46786
rect 49758 46734 49810 46786
rect 3838 46622 3890 46674
rect 4286 46622 4338 46674
rect 5294 46622 5346 46674
rect 7534 46622 7586 46674
rect 9886 46622 9938 46674
rect 10110 46622 10162 46674
rect 11118 46622 11170 46674
rect 11790 46622 11842 46674
rect 13134 46622 13186 46674
rect 15486 46622 15538 46674
rect 15934 46622 15986 46674
rect 16606 46622 16658 46674
rect 17278 46622 17330 46674
rect 18174 46622 18226 46674
rect 19854 46622 19906 46674
rect 20862 46622 20914 46674
rect 21646 46622 21698 46674
rect 23886 46622 23938 46674
rect 29598 46622 29650 46674
rect 30270 46622 30322 46674
rect 33406 46622 33458 46674
rect 38222 46622 38274 46674
rect 40686 46622 40738 46674
rect 43150 46622 43202 46674
rect 45950 46622 46002 46674
rect 46398 46622 46450 46674
rect 46734 46622 46786 46674
rect 47070 46622 47122 46674
rect 49646 46622 49698 46674
rect 52334 46622 52386 46674
rect 52446 46622 52498 46674
rect 53342 46622 53394 46674
rect 53790 46622 53842 46674
rect 55358 46622 55410 46674
rect 1598 46510 1650 46562
rect 3278 46510 3330 46562
rect 3390 46510 3442 46562
rect 3950 46510 4002 46562
rect 6862 46510 6914 46562
rect 7982 46510 8034 46562
rect 10558 46510 10610 46562
rect 11006 46510 11058 46562
rect 13582 46510 13634 46562
rect 19966 46510 20018 46562
rect 20750 46510 20802 46562
rect 22094 46510 22146 46562
rect 24446 46510 24498 46562
rect 30718 46510 30770 46562
rect 32622 46510 32674 46562
rect 33854 46510 33906 46562
rect 35758 46510 35810 46562
rect 36990 46510 37042 46562
rect 37326 46510 37378 46562
rect 38558 46510 38610 46562
rect 45502 46510 45554 46562
rect 52670 46510 52722 46562
rect 53006 46510 53058 46562
rect 2830 46398 2882 46450
rect 4062 46398 4114 46450
rect 4174 46398 4226 46450
rect 5742 46398 5794 46450
rect 9102 46398 9154 46450
rect 10222 46398 10274 46450
rect 10334 46398 10386 46450
rect 12126 46398 12178 46450
rect 14702 46398 14754 46450
rect 16158 46398 16210 46450
rect 18846 46398 18898 46450
rect 25566 46398 25618 46450
rect 26686 46398 26738 46450
rect 27806 46398 27858 46450
rect 29710 46398 29762 46450
rect 29934 46398 29986 46450
rect 31950 46398 32002 46450
rect 32846 46398 32898 46450
rect 35422 46398 35474 46450
rect 35646 46398 35698 46450
rect 41134 46398 41186 46450
rect 42254 46398 42306 46450
rect 43262 46398 43314 46450
rect 43374 46398 43426 46450
rect 44270 46398 44322 46450
rect 46510 46398 46562 46450
rect 47630 46398 47682 46450
rect 50206 46398 50258 46450
rect 53118 46398 53170 46450
rect 54910 46398 54962 46450
rect 56030 46398 56082 46450
rect 56366 46398 56418 46450
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 44466 46230 44518 46282
rect 44570 46230 44622 46282
rect 44674 46230 44726 46282
rect 1374 46062 1426 46114
rect 18510 46062 18562 46114
rect 20302 46062 20354 46114
rect 21758 46062 21810 46114
rect 25342 46062 25394 46114
rect 27918 46062 27970 46114
rect 31166 46062 31218 46114
rect 31278 46062 31330 46114
rect 34750 46062 34802 46114
rect 39118 46062 39170 46114
rect 42590 46062 42642 46114
rect 43822 46062 43874 46114
rect 46062 46062 46114 46114
rect 51438 46062 51490 46114
rect 52446 46062 52498 46114
rect 53566 46062 53618 46114
rect 2046 45950 2098 46002
rect 2718 45950 2770 46002
rect 3054 45950 3106 46002
rect 4062 45950 4114 46002
rect 4510 45950 4562 46002
rect 7982 45950 8034 46002
rect 9886 45950 9938 46002
rect 11566 45950 11618 46002
rect 12462 45950 12514 46002
rect 14590 45950 14642 46002
rect 17390 45950 17442 46002
rect 19294 45950 19346 46002
rect 20750 45950 20802 46002
rect 30606 45950 30658 46002
rect 33630 45950 33682 46002
rect 35870 45950 35922 46002
rect 37438 45950 37490 46002
rect 40798 45950 40850 46002
rect 47406 45950 47458 46002
rect 49086 45950 49138 46002
rect 55918 45950 55970 46002
rect 1038 45838 1090 45890
rect 1710 45838 1762 45890
rect 2382 45838 2434 45890
rect 3390 45838 3442 45890
rect 3838 45838 3890 45890
rect 4734 45838 4786 45890
rect 5070 45838 5122 45890
rect 6190 45838 6242 45890
rect 8206 45838 8258 45890
rect 9998 45838 10050 45890
rect 11006 45838 11058 45890
rect 11454 45838 11506 45890
rect 12350 45838 12402 45890
rect 14030 45838 14082 45890
rect 19406 45838 19458 45890
rect 19966 45838 20018 45890
rect 21086 45838 21138 45890
rect 21646 45838 21698 45890
rect 22430 45838 22482 45890
rect 22766 45838 22818 45890
rect 23886 45838 23938 45890
rect 27246 45838 27298 45890
rect 27694 45838 27746 45890
rect 28366 45838 28418 45890
rect 28926 45838 28978 45890
rect 29934 45838 29986 45890
rect 30494 45838 30546 45890
rect 31390 45838 31442 45890
rect 31614 45838 31666 45890
rect 36990 45838 37042 45890
rect 39230 45838 39282 45890
rect 39342 45838 39394 45890
rect 39790 45838 39842 45890
rect 45614 45838 45666 45890
rect 45950 45838 46002 45890
rect 46286 45838 46338 45890
rect 47182 45838 47234 45890
rect 50318 45838 50370 45890
rect 50766 45838 50818 45890
rect 50990 45838 51042 45890
rect 51214 45838 51266 45890
rect 54574 45838 54626 45890
rect 54798 45838 54850 45890
rect 55134 45838 55186 45890
rect 56254 45838 56306 45890
rect 16942 45726 16994 45778
rect 24894 45726 24946 45778
rect 26910 45726 26962 45778
rect 34078 45726 34130 45778
rect 36318 45726 36370 45778
rect 40462 45726 40514 45778
rect 42702 45726 42754 45778
rect 43374 45726 43426 45778
rect 46174 45726 46226 45778
rect 46958 45726 47010 45778
rect 47294 45726 47346 45778
rect 48750 45726 48802 45778
rect 51326 45726 51378 45778
rect 51998 45726 52050 45778
rect 54014 45726 54066 45778
rect 54686 45726 54738 45778
rect 7086 45614 7138 45666
rect 7422 45614 7474 45666
rect 8990 45614 9042 45666
rect 9326 45614 9378 45666
rect 10670 45614 10722 45666
rect 13134 45614 13186 45666
rect 13470 45614 13522 45666
rect 15710 45614 15762 45666
rect 26462 45614 26514 45666
rect 30606 45614 30658 45666
rect 31838 45614 31890 45666
rect 32510 45614 32562 45666
rect 38670 45614 38722 45666
rect 42030 45614 42082 45666
rect 42814 45614 42866 45666
rect 44942 45614 44994 45666
rect 46734 45614 46786 45666
rect 51886 45614 51938 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 43806 45446 43858 45498
rect 43910 45446 43962 45498
rect 44014 45446 44066 45498
rect 11006 45278 11058 45330
rect 17726 45278 17778 45330
rect 35310 45278 35362 45330
rect 35646 45278 35698 45330
rect 39118 45278 39170 45330
rect 42590 45278 42642 45330
rect 45950 45278 46002 45330
rect 50878 45278 50930 45330
rect 52446 45278 52498 45330
rect 53790 45278 53842 45330
rect 4398 45166 4450 45218
rect 6526 45166 6578 45218
rect 8878 45166 8930 45218
rect 12910 45166 12962 45218
rect 14030 45166 14082 45218
rect 24222 45166 24274 45218
rect 40014 45166 40066 45218
rect 43150 45166 43202 45218
rect 44382 45166 44434 45218
rect 46510 45166 46562 45218
rect 47070 45166 47122 45218
rect 49310 45166 49362 45218
rect 55358 45166 55410 45218
rect 55806 45166 55858 45218
rect 1262 45054 1314 45106
rect 2158 45054 2210 45106
rect 2830 45054 2882 45106
rect 3502 45054 3554 45106
rect 3950 45054 4002 45106
rect 5294 45054 5346 45106
rect 5518 45054 5570 45106
rect 10110 45054 10162 45106
rect 11342 45054 11394 45106
rect 12686 45054 12738 45106
rect 13022 45054 13074 45106
rect 13246 45054 13298 45106
rect 14478 45054 14530 45106
rect 14814 45057 14866 45109
rect 15710 45054 15762 45106
rect 16046 45054 16098 45106
rect 17054 45054 17106 45106
rect 19294 45054 19346 45106
rect 22206 45054 22258 45106
rect 24670 45054 24722 45106
rect 25006 45054 25058 45106
rect 25678 45054 25730 45106
rect 26350 45054 26402 45106
rect 27358 45054 27410 45106
rect 30158 45054 30210 45106
rect 30942 45054 30994 45106
rect 33182 45054 33234 45106
rect 37438 45054 37490 45106
rect 40574 45054 40626 45106
rect 42142 45054 42194 45106
rect 42926 45054 42978 45106
rect 43038 45054 43090 45106
rect 46398 45054 46450 45106
rect 49198 45054 49250 45106
rect 52894 45054 52946 45106
rect 56030 45054 56082 45106
rect 3390 44942 3442 44994
rect 4958 44942 5010 44994
rect 5966 44942 6018 44994
rect 6862 44942 6914 44994
rect 8542 44942 8594 44994
rect 8766 44942 8818 44994
rect 9326 44942 9378 44994
rect 9886 44942 9938 44994
rect 11566 44942 11618 44994
rect 12126 44942 12178 44994
rect 22542 44942 22594 44994
rect 29822 44942 29874 44994
rect 33518 44942 33570 44994
rect 37886 44942 37938 44994
rect 39678 44942 39730 44994
rect 39902 44942 39954 44994
rect 51326 44942 51378 44994
rect 53230 44942 53282 44994
rect 56366 44942 56418 44994
rect 5070 44830 5122 44882
rect 5854 44830 5906 44882
rect 8094 44830 8146 44882
rect 10446 44830 10498 44882
rect 15038 44830 15090 44882
rect 18846 44830 18898 44882
rect 23774 44830 23826 44882
rect 25230 44830 25282 44882
rect 28590 44830 28642 44882
rect 31390 44830 31442 44882
rect 32510 44830 32562 44882
rect 34750 44830 34802 44882
rect 35534 44830 35586 44882
rect 36654 44830 36706 44882
rect 36990 44830 37042 44882
rect 41022 44830 41074 44882
rect 43262 44830 43314 44882
rect 44830 44830 44882 44882
rect 47518 44830 47570 44882
rect 48638 44830 48690 44882
rect 49758 44830 49810 44882
rect 51438 44830 51490 44882
rect 52110 44830 52162 44882
rect 54910 44830 54962 44882
rect 56254 44830 56306 44882
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 44466 44662 44518 44714
rect 44570 44662 44622 44714
rect 44674 44662 44726 44714
rect 5518 44494 5570 44546
rect 16606 44494 16658 44546
rect 16830 44494 16882 44546
rect 18286 44494 18338 44546
rect 19406 44494 19458 44546
rect 21646 44494 21698 44546
rect 27918 44494 27970 44546
rect 31278 44494 31330 44546
rect 31390 44494 31442 44546
rect 37326 44494 37378 44546
rect 37438 44494 37490 44546
rect 38782 44494 38834 44546
rect 42366 44494 42418 44546
rect 50094 44494 50146 44546
rect 50654 44494 50706 44546
rect 1822 44382 1874 44434
rect 4510 44382 4562 44434
rect 8206 44382 8258 44434
rect 9550 44382 9602 44434
rect 12686 44382 12738 44434
rect 14814 44382 14866 44434
rect 16942 44382 16994 44434
rect 20526 44382 20578 44434
rect 22766 44382 22818 44434
rect 23886 44382 23938 44434
rect 25230 44382 25282 44434
rect 30606 44382 30658 44434
rect 31166 44382 31218 44434
rect 33630 44382 33682 44434
rect 35198 44382 35250 44434
rect 37550 44382 37602 44434
rect 38446 44382 38498 44434
rect 38670 44382 38722 44434
rect 41134 44382 41186 44434
rect 42926 44382 42978 44434
rect 43822 44382 43874 44434
rect 46286 44382 46338 44434
rect 48974 44382 49026 44434
rect 51774 44382 51826 44434
rect 52894 44382 52946 44434
rect 53454 44382 53506 44434
rect 55358 44382 55410 44434
rect 56366 44382 56418 44434
rect 3726 44270 3778 44322
rect 3950 44270 4002 44322
rect 4286 44270 4338 44322
rect 4846 44270 4898 44322
rect 5294 44270 5346 44322
rect 6190 44270 6242 44322
rect 6638 44270 6690 44322
rect 7534 44270 7586 44322
rect 8094 44270 8146 44322
rect 11342 44270 11394 44322
rect 14366 44270 14418 44322
rect 17838 44270 17890 44322
rect 22206 44270 22258 44322
rect 27246 44270 27298 44322
rect 27694 44270 27746 44322
rect 28478 44270 28530 44322
rect 28926 44270 28978 44322
rect 29934 44270 29986 44322
rect 30494 44270 30546 44322
rect 31614 44270 31666 44322
rect 31838 44270 31890 44322
rect 34078 44270 34130 44322
rect 34862 44270 34914 44322
rect 37102 44270 37154 44322
rect 38894 44270 38946 44322
rect 39342 44270 39394 44322
rect 40686 44270 40738 44322
rect 45838 44270 45890 44322
rect 50990 44270 51042 44322
rect 51438 44270 51490 44322
rect 54350 44270 54402 44322
rect 54574 44270 54626 44322
rect 55022 44270 55074 44322
rect 56142 44270 56194 44322
rect 1486 44158 1538 44210
rect 4062 44158 4114 44210
rect 9102 44158 9154 44210
rect 12238 44158 12290 44210
rect 20078 44158 20130 44210
rect 24894 44158 24946 44210
rect 26910 44158 26962 44210
rect 3054 44046 3106 44098
rect 8206 44046 8258 44098
rect 11118 44102 11170 44154
rect 38110 44158 38162 44210
rect 39118 44158 39170 44210
rect 43486 44158 43538 44210
rect 48526 44158 48578 44210
rect 54126 44158 54178 44210
rect 54462 44158 54514 44210
rect 10670 44046 10722 44098
rect 11678 44046 11730 44098
rect 13806 44046 13858 44098
rect 16046 44046 16098 44098
rect 26462 44046 26514 44098
rect 30606 44046 30658 44098
rect 32510 44046 32562 44098
rect 36430 44046 36482 44098
rect 36878 44046 36930 44098
rect 37998 44046 38050 44098
rect 42814 44046 42866 44098
rect 45054 44046 45106 44098
rect 47406 44046 47458 44098
rect 52334 44046 52386 44098
rect 52670 44046 52722 44098
rect 53902 44046 53954 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 43806 43878 43858 43930
rect 43910 43878 43962 43930
rect 44014 43878 44066 43930
rect 45054 43710 45106 43762
rect 3166 43598 3218 43650
rect 5182 43598 5234 43650
rect 10782 43598 10834 43650
rect 11342 43598 11394 43650
rect 12238 43598 12290 43650
rect 15598 43598 15650 43650
rect 16382 43598 16434 43650
rect 16830 43598 16882 43650
rect 28702 43598 28754 43650
rect 33182 43598 33234 43650
rect 34750 43598 34802 43650
rect 39678 43598 39730 43650
rect 41246 43598 41298 43650
rect 41694 43598 41746 43650
rect 43374 43598 43426 43650
rect 43598 43598 43650 43650
rect 48190 43598 48242 43650
rect 1486 43486 1538 43538
rect 3614 43486 3666 43538
rect 4062 43486 4114 43538
rect 4286 43486 4338 43538
rect 5518 43486 5570 43538
rect 6190 43486 6242 43538
rect 6974 43486 7026 43538
rect 9102 43486 9154 43538
rect 11790 43486 11842 43538
rect 13246 43486 13298 43538
rect 15374 43486 15426 43538
rect 15822 43486 15874 43538
rect 17166 43486 17218 43538
rect 17726 43486 17778 43538
rect 19070 43486 19122 43538
rect 19854 43486 19906 43538
rect 22206 43486 22258 43538
rect 24558 43486 24610 43538
rect 25006 43486 25058 43538
rect 26350 43486 26402 43538
rect 27246 43486 27298 43538
rect 32510 43486 32562 43538
rect 35198 43486 35250 43538
rect 35534 43486 35586 43538
rect 37326 43486 37378 43538
rect 42254 43486 42306 43538
rect 44494 43486 44546 43538
rect 44830 43486 44882 43538
rect 45166 43486 45218 43538
rect 49198 43486 49250 43538
rect 50542 43486 50594 43538
rect 50766 43486 50818 43538
rect 52110 43486 52162 43538
rect 52558 43486 52610 43538
rect 52782 43486 52834 43538
rect 54126 43486 54178 43538
rect 6302 43374 6354 43426
rect 7422 43374 7474 43426
rect 11230 43374 11282 43426
rect 11566 43374 11618 43426
rect 13694 43374 13746 43426
rect 16046 43374 16098 43426
rect 16494 43374 16546 43426
rect 18286 43374 18338 43426
rect 24222 43374 24274 43426
rect 25678 43374 25730 43426
rect 32062 43374 32114 43426
rect 33518 43374 33570 43426
rect 35646 43374 35698 43426
rect 36766 43374 36818 43426
rect 39342 43374 39394 43426
rect 39678 43374 39730 43426
rect 39790 43374 39842 43426
rect 40462 43374 40514 43426
rect 40798 43374 40850 43426
rect 40910 43374 40962 43426
rect 41918 43374 41970 43426
rect 43150 43374 43202 43426
rect 44158 43374 44210 43426
rect 45502 43374 45554 43426
rect 47854 43374 47906 43426
rect 49422 43374 49474 43426
rect 49758 43374 49810 43426
rect 51102 43374 51154 43426
rect 51326 43374 51378 43426
rect 51998 43374 52050 43426
rect 52334 43374 52386 43426
rect 54574 43374 54626 43426
rect 55806 43374 55858 43426
rect 56366 43374 56418 43426
rect 2046 43262 2098 43314
rect 3838 43262 3890 43314
rect 3950 43262 4002 43314
rect 8542 43262 8594 43314
rect 9662 43262 9714 43314
rect 12126 43262 12178 43314
rect 14926 43262 14978 43314
rect 17838 43262 17890 43314
rect 22654 43262 22706 43314
rect 23774 43262 23826 43314
rect 25230 43262 25282 43314
rect 29150 43262 29202 43314
rect 30270 43262 30322 43314
rect 30830 43262 30882 43314
rect 35758 43262 35810 43314
rect 36430 43262 36482 43314
rect 37774 43262 37826 43314
rect 38894 43262 38946 43314
rect 39566 43262 39618 43314
rect 40686 43262 40738 43314
rect 41582 43262 41634 43314
rect 41806 43262 41858 43314
rect 42926 43262 42978 43314
rect 43038 43262 43090 43314
rect 44270 43262 44322 43314
rect 45390 43262 45442 43314
rect 45838 43262 45890 43314
rect 46174 43262 46226 43314
rect 46622 43262 46674 43314
rect 48862 43262 48914 43314
rect 50430 43262 50482 43314
rect 53230 43262 53282 43314
rect 53566 43262 53618 43314
rect 56254 43262 56306 43314
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 44466 43094 44518 43146
rect 44570 43094 44622 43146
rect 44674 43094 44726 43146
rect 1822 42926 1874 42978
rect 4398 42926 4450 42978
rect 8206 42926 8258 42978
rect 10446 42926 10498 42978
rect 12686 42926 12738 42978
rect 27470 42926 27522 42978
rect 35310 42926 35362 42978
rect 36430 42926 36482 42978
rect 37550 42926 37602 42978
rect 39118 42926 39170 42978
rect 43934 42926 43986 42978
rect 45054 42926 45106 42978
rect 46286 42926 46338 42978
rect 55246 42926 55298 42978
rect 4846 42814 4898 42866
rect 7198 42814 7250 42866
rect 7534 42814 7586 42866
rect 9550 42814 9602 42866
rect 9774 42814 9826 42866
rect 11006 42814 11058 42866
rect 11454 42814 11506 42866
rect 14926 42814 14978 42866
rect 18062 42814 18114 42866
rect 19742 42814 19794 42866
rect 20750 42814 20802 42866
rect 27918 42814 27970 42866
rect 30718 42814 30770 42866
rect 33630 42814 33682 42866
rect 41246 42814 41298 42866
rect 45726 42814 45778 42866
rect 47406 42814 47458 42866
rect 49982 42814 50034 42866
rect 53678 42814 53730 42866
rect 53902 42814 53954 42866
rect 56366 42814 56418 42866
rect 3726 42702 3778 42754
rect 4286 42702 4338 42754
rect 5406 42702 5458 42754
rect 6414 42702 6466 42754
rect 7870 42702 7922 42754
rect 8990 42702 9042 42754
rect 11566 42702 11618 42754
rect 14366 42702 14418 42754
rect 17614 42702 17666 42754
rect 20078 42702 20130 42754
rect 20526 42702 20578 42754
rect 21422 42702 21474 42754
rect 21758 42702 21810 42754
rect 22766 42702 22818 42754
rect 26798 42702 26850 42754
rect 27246 42702 27298 42754
rect 28702 42702 28754 42754
rect 29486 42702 29538 42754
rect 30830 42702 30882 42754
rect 34862 42702 34914 42754
rect 37102 42702 37154 42754
rect 38670 42702 38722 42754
rect 39454 42702 39506 42754
rect 43374 42702 43426 42754
rect 45502 42702 45554 42754
rect 45950 42702 46002 42754
rect 46062 42702 46114 42754
rect 46622 42702 46674 42754
rect 46846 42702 46898 42754
rect 47070 42702 47122 42754
rect 47294 42702 47346 42754
rect 52110 42702 52162 42754
rect 54126 42702 54178 42754
rect 54350 42702 54402 42754
rect 1374 42590 1426 42642
rect 3390 42590 3442 42642
rect 12238 42590 12290 42642
rect 16046 42590 16098 42642
rect 17726 42590 17778 42642
rect 26462 42590 26514 42642
rect 34078 42590 34130 42642
rect 39678 42590 39730 42642
rect 40798 42590 40850 42642
rect 42814 42590 42866 42642
rect 54462 42590 54514 42642
rect 54574 42646 54626 42698
rect 54910 42702 54962 42754
rect 56030 42702 56082 42754
rect 2942 42478 2994 42530
rect 9214 42478 9266 42530
rect 9662 42478 9714 42530
rect 10782 42478 10834 42530
rect 13806 42478 13858 42530
rect 19294 42478 19346 42530
rect 31390 42478 31442 42530
rect 31726 42478 31778 42530
rect 32510 42478 32562 42530
rect 42366 42478 42418 42530
rect 42926 42478 42978 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 43806 42310 43858 42362
rect 43910 42310 43962 42362
rect 44014 42310 44066 42362
rect 5854 42142 5906 42194
rect 6190 42142 6242 42194
rect 8990 42142 9042 42194
rect 36766 42142 36818 42194
rect 43262 42142 43314 42194
rect 43598 42142 43650 42194
rect 50430 42142 50482 42194
rect 54014 42142 54066 42194
rect 54574 42142 54626 42194
rect 6862 42030 6914 42082
rect 9214 42030 9266 42082
rect 30606 42030 30658 42082
rect 35758 42030 35810 42082
rect 38110 42030 38162 42082
rect 39230 42030 39282 42082
rect 42254 42030 42306 42082
rect 51214 42030 51266 42082
rect 56142 42030 56194 42082
rect 1262 41918 1314 41970
rect 3278 41918 3330 41970
rect 3614 41918 3666 41970
rect 3726 41918 3778 41970
rect 4062 41918 4114 41970
rect 4286 41918 4338 41970
rect 9326 41918 9378 41970
rect 10446 41918 10498 41970
rect 12126 41918 12178 41970
rect 12798 41918 12850 41970
rect 12910 41918 12962 41970
rect 13358 41918 13410 41970
rect 14254 41918 14306 41970
rect 14814 41918 14866 41970
rect 15710 41918 15762 41970
rect 16158 41918 16210 41970
rect 16830 41918 16882 41970
rect 17166 41918 17218 41970
rect 17614 41918 17666 41970
rect 18286 41918 18338 41970
rect 19070 41918 19122 41970
rect 19966 41918 20018 41970
rect 21646 41918 21698 41970
rect 21982 41918 22034 41970
rect 22542 41918 22594 41970
rect 23662 41918 23714 41970
rect 24782 41918 24834 41970
rect 25454 41918 25506 41970
rect 31054 41918 31106 41970
rect 31502 41918 31554 41970
rect 32286 41918 32338 41970
rect 32622 41918 32674 41970
rect 33630 41918 33682 41970
rect 34974 41918 35026 41970
rect 35422 41918 35474 41970
rect 35646 41918 35698 41970
rect 38222 41918 38274 41970
rect 38558 41918 38610 41970
rect 45950 41918 46002 41970
rect 48078 41918 48130 41970
rect 48750 41918 48802 41970
rect 52446 41918 52498 41970
rect 1598 41806 1650 41858
rect 3390 41806 3442 41858
rect 5294 41806 5346 41858
rect 5630 41806 5682 41858
rect 9998 41806 10050 41858
rect 10894 41806 10946 41858
rect 15486 41806 15538 41858
rect 16494 41806 16546 41858
rect 23102 41806 23154 41858
rect 31614 41806 31666 41858
rect 34414 41806 34466 41858
rect 34526 41806 34578 41858
rect 35198 41806 35250 41858
rect 36990 41806 37042 41858
rect 37438 41806 37490 41858
rect 41582 41806 41634 41858
rect 41918 41806 41970 41858
rect 42590 41806 42642 41858
rect 43038 41806 43090 41858
rect 51438 41806 51490 41858
rect 2830 41694 2882 41746
rect 4062 41694 4114 41746
rect 7310 41694 7362 41746
rect 8430 41694 8482 41746
rect 9662 41694 9714 41746
rect 11006 41694 11058 41746
rect 17838 41694 17890 41746
rect 22654 41694 22706 41746
rect 25902 41694 25954 41746
rect 27022 41694 27074 41746
rect 34750 41694 34802 41746
rect 36430 41694 36482 41746
rect 37998 41694 38050 41746
rect 39678 41694 39730 41746
rect 40798 41694 40850 41746
rect 44270 41694 44322 41746
rect 45390 41694 45442 41746
rect 46510 41694 46562 41746
rect 47630 41694 47682 41746
rect 49310 41694 49362 41746
rect 51214 41694 51266 41746
rect 52894 41694 52946 41746
rect 55694 41694 55746 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 44466 41526 44518 41578
rect 44570 41526 44622 41578
rect 44674 41526 44726 41578
rect 2270 41358 2322 41410
rect 7086 41358 7138 41410
rect 8094 41358 8146 41410
rect 12462 41358 12514 41410
rect 12798 41358 12850 41410
rect 13134 41358 13186 41410
rect 20190 41358 20242 41410
rect 26350 41358 26402 41410
rect 28926 41358 28978 41410
rect 33406 41358 33458 41410
rect 37102 41358 37154 41410
rect 37326 41358 37378 41410
rect 38446 41358 38498 41410
rect 40910 41358 40962 41410
rect 42590 41358 42642 41410
rect 43262 41358 43314 41410
rect 43822 41358 43874 41410
rect 46286 41358 46338 41410
rect 48190 41358 48242 41410
rect 48302 41358 48354 41410
rect 48526 41358 48578 41410
rect 49982 41358 50034 41410
rect 56254 41358 56306 41410
rect 4510 41246 4562 41298
rect 9886 41246 9938 41298
rect 10334 41246 10386 41298
rect 14814 41246 14866 41298
rect 16046 41246 16098 41298
rect 17390 41246 17442 41298
rect 17950 41246 18002 41298
rect 18958 41246 19010 41298
rect 20638 41246 20690 41298
rect 21646 41246 21698 41298
rect 22094 41246 22146 41298
rect 26238 41246 26290 41298
rect 35646 41246 35698 41298
rect 44942 41246 44994 41298
rect 47182 41246 47234 41298
rect 48078 41246 48130 41298
rect 50206 41246 50258 41298
rect 51326 41246 51378 41298
rect 53566 41246 53618 41298
rect 2718 41134 2770 41186
rect 3838 41134 3890 41186
rect 4286 41134 4338 41186
rect 5070 41134 5122 41186
rect 5518 41134 5570 41186
rect 6526 41134 6578 41186
rect 7310 41134 7362 41186
rect 7758 41134 7810 41186
rect 9326 41134 9378 41186
rect 9774 41134 9826 41186
rect 10446 41134 10498 41186
rect 11118 41134 11170 41186
rect 12014 41134 12066 41186
rect 13358 41134 13410 41186
rect 14366 41134 14418 41186
rect 18510 41134 18562 41186
rect 20974 41134 21026 41186
rect 21534 41134 21586 41186
rect 22654 41134 22706 41186
rect 23662 41134 23714 41186
rect 25790 41134 25842 41186
rect 28366 41134 28418 41186
rect 28702 41134 28754 41186
rect 29598 41134 29650 41186
rect 30046 41134 30098 41186
rect 30942 41134 30994 41186
rect 32958 41134 33010 41186
rect 35086 41134 35138 41186
rect 37438 41134 37490 41186
rect 37886 41134 37938 41186
rect 40350 41134 40402 41186
rect 42478 41134 42530 41186
rect 42814 41134 42866 41186
rect 43038 41134 43090 41186
rect 45390 41134 45442 41186
rect 46622 41134 46674 41186
rect 47406 41134 47458 41186
rect 49310 41134 49362 41186
rect 49646 41134 49698 41186
rect 50430 41134 50482 41186
rect 50878 41134 50930 41186
rect 55358 41134 55410 41186
rect 55918 41134 55970 41186
rect 3502 41022 3554 41074
rect 8878 41022 8930 41074
rect 27918 41022 27970 41074
rect 49198 41022 49250 41074
rect 49982 41022 50034 41074
rect 52558 41022 52610 41074
rect 53230 41022 53282 41074
rect 1150 40910 1202 40962
rect 16830 40910 16882 40962
rect 17166 40910 17218 40962
rect 27470 40910 27522 40962
rect 34526 40910 34578 40962
rect 36766 40910 36818 40962
rect 39566 40910 39618 40962
rect 42030 40910 42082 40962
rect 43374 40910 43426 40962
rect 48974 40910 49026 40962
rect 54798 40910 54850 40962
rect 55246 40910 55298 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 43806 40742 43858 40794
rect 43910 40742 43962 40794
rect 44014 40742 44066 40794
rect 30494 40574 30546 40626
rect 42926 40574 42978 40626
rect 5406 40462 5458 40514
rect 6302 40462 6354 40514
rect 8318 40462 8370 40514
rect 18398 40462 18450 40514
rect 21982 40462 22034 40514
rect 28926 40462 28978 40514
rect 30942 40462 30994 40514
rect 42814 40462 42866 40514
rect 46622 40462 46674 40514
rect 51214 40462 51266 40514
rect 52222 40462 52274 40514
rect 55918 40462 55970 40514
rect 1598 40350 1650 40402
rect 1934 40350 1986 40402
rect 2606 40350 2658 40402
rect 3166 40350 3218 40402
rect 4174 40350 4226 40402
rect 4958 40350 5010 40402
rect 5518 40350 5570 40402
rect 8766 40350 8818 40402
rect 9102 40350 9154 40402
rect 9774 40350 9826 40402
rect 10334 40350 10386 40402
rect 11342 40350 11394 40402
rect 12238 40350 12290 40402
rect 13918 40350 13970 40402
rect 14478 40350 14530 40402
rect 15150 40350 15202 40402
rect 15598 40350 15650 40402
rect 16718 40350 16770 40402
rect 19966 40350 20018 40402
rect 22318 40350 22370 40402
rect 22766 40350 22818 40402
rect 23438 40350 23490 40402
rect 24110 40350 24162 40402
rect 25006 40350 25058 40402
rect 26238 40350 26290 40402
rect 31278 40350 31330 40402
rect 31726 40350 31778 40402
rect 32398 40350 32450 40402
rect 32958 40350 33010 40402
rect 33966 40350 34018 40402
rect 35086 40350 35138 40402
rect 36318 40350 36370 40402
rect 36654 40350 36706 40402
rect 37214 40350 37266 40402
rect 38782 40350 38834 40402
rect 39566 40350 39618 40402
rect 40126 40344 40178 40396
rect 40798 40350 40850 40402
rect 41246 40350 41298 40402
rect 42366 40350 42418 40402
rect 43374 40350 43426 40402
rect 44382 40350 44434 40402
rect 48862 40350 48914 40402
rect 1150 40238 1202 40290
rect 5182 40238 5234 40290
rect 9326 40238 9378 40290
rect 11902 40238 11954 40290
rect 12798 40238 12850 40290
rect 13582 40238 13634 40290
rect 14590 40238 14642 40290
rect 18846 40238 18898 40290
rect 22990 40238 23042 40290
rect 29374 40238 29426 40290
rect 31950 40238 32002 40290
rect 35422 40238 35474 40290
rect 35758 40238 35810 40290
rect 36430 40238 36482 40290
rect 37550 40238 37602 40290
rect 39230 40238 39282 40290
rect 40238 40238 40290 40290
rect 49310 40238 49362 40290
rect 51326 40238 51378 40290
rect 2158 40126 2210 40178
rect 5406 40126 5458 40178
rect 6750 40126 6802 40178
rect 7870 40126 7922 40178
rect 13134 40126 13186 40178
rect 26686 40126 26738 40178
rect 27806 40126 27858 40178
rect 35534 40126 35586 40178
rect 35646 40126 35698 40178
rect 43598 40126 43650 40178
rect 44830 40126 44882 40178
rect 45950 40126 46002 40178
rect 47070 40126 47122 40178
rect 48190 40126 48242 40178
rect 50430 40126 50482 40178
rect 50878 40126 50930 40178
rect 51102 40126 51154 40178
rect 52670 40126 52722 40178
rect 53790 40126 53842 40178
rect 54350 40126 54402 40178
rect 55470 40126 55522 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 44466 39958 44518 40010
rect 44570 39958 44622 40010
rect 44674 39958 44726 40010
rect 1038 39790 1090 39842
rect 1374 39790 1426 39842
rect 1710 39790 1762 39842
rect 2046 39790 2098 39842
rect 2718 39790 2770 39842
rect 3950 39790 4002 39842
rect 6526 39790 6578 39842
rect 6862 39790 6914 39842
rect 7310 39790 7362 39842
rect 13470 39790 13522 39842
rect 16158 39790 16210 39842
rect 20078 39790 20130 39842
rect 21534 39790 21586 39842
rect 27470 39790 27522 39842
rect 33630 39790 33682 39842
rect 36430 39790 36482 39842
rect 39566 39790 39618 39842
rect 39790 39790 39842 39842
rect 41246 39790 41298 39842
rect 45054 39790 45106 39842
rect 47518 39790 47570 39842
rect 48414 39790 48466 39842
rect 49310 39790 49362 39842
rect 53566 39790 53618 39842
rect 54574 39790 54626 39842
rect 56254 39790 56306 39842
rect 2382 39678 2434 39730
rect 2494 39678 2546 39730
rect 7198 39678 7250 39730
rect 8878 39678 8930 39730
rect 9886 39678 9938 39730
rect 18846 39678 18898 39730
rect 30158 39678 30210 39730
rect 35198 39678 35250 39730
rect 37774 39678 37826 39730
rect 39454 39678 39506 39730
rect 40238 39678 40290 39730
rect 48190 39678 48242 39730
rect 51550 39678 51602 39730
rect 3278 39566 3330 39618
rect 3726 39566 3778 39618
rect 4622 39566 4674 39618
rect 4958 39566 5010 39618
rect 6078 39566 6130 39618
rect 7870 39566 7922 39618
rect 7982 39566 8034 39618
rect 8430 39566 8482 39618
rect 9214 39566 9266 39618
rect 9774 39566 9826 39618
rect 10446 39566 10498 39618
rect 10894 39566 10946 39618
rect 11902 39566 11954 39618
rect 12910 39566 12962 39618
rect 18510 39566 18562 39618
rect 20862 39566 20914 39618
rect 21422 39566 21474 39618
rect 22094 39566 22146 39618
rect 22542 39566 22594 39618
rect 23550 39566 23602 39618
rect 26910 39566 26962 39618
rect 27246 39566 27298 39618
rect 28030 39566 28082 39618
rect 28702 39566 28754 39618
rect 29486 39566 29538 39618
rect 30382 39566 30434 39618
rect 34078 39566 34130 39618
rect 34862 39566 34914 39618
rect 37326 39566 37378 39618
rect 40574 39566 40626 39618
rect 41022 39566 41074 39618
rect 41918 39566 41970 39618
rect 42254 39566 42306 39618
rect 43262 39566 43314 39618
rect 45502 39566 45554 39618
rect 46174 39566 46226 39618
rect 46398 39566 46450 39618
rect 47182 39566 47234 39618
rect 48078 39566 48130 39618
rect 48862 39566 48914 39618
rect 50990 39566 51042 39618
rect 53678 39566 53730 39618
rect 53790 39566 53842 39618
rect 54350 39566 54402 39618
rect 54798 39566 54850 39618
rect 55022 39566 55074 39618
rect 56030 39566 56082 39618
rect 2942 39454 2994 39506
rect 8206 39454 8258 39506
rect 16046 39454 16098 39506
rect 20526 39454 20578 39506
rect 26462 39454 26514 39506
rect 53342 39454 53394 39506
rect 54462 39454 54514 39506
rect 7310 39342 7362 39394
rect 14590 39342 14642 39394
rect 30942 39342 30994 39394
rect 31278 39342 31330 39394
rect 32510 39342 32562 39394
rect 39006 39342 39058 39394
rect 43934 39342 43986 39394
rect 46734 39342 46786 39394
rect 50430 39342 50482 39394
rect 52670 39342 52722 39394
rect 53118 39342 53170 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 43806 39174 43858 39226
rect 43910 39174 43962 39226
rect 44014 39174 44066 39226
rect 11790 39006 11842 39058
rect 30382 39006 30434 39058
rect 35646 39006 35698 39058
rect 43486 39006 43538 39058
rect 48190 39006 48242 39058
rect 51998 39006 52050 39058
rect 53342 39006 53394 39058
rect 1262 38894 1314 38946
rect 11902 38894 11954 38946
rect 14366 38894 14418 38946
rect 21310 38894 21362 38946
rect 23550 38894 23602 38946
rect 31390 38894 31442 38946
rect 35086 38894 35138 38946
rect 35758 38894 35810 38946
rect 36766 38894 36818 38946
rect 39678 38894 39730 38946
rect 44382 38894 44434 38946
rect 46622 38894 46674 38946
rect 50766 38894 50818 38946
rect 52222 38894 52274 38946
rect 53118 38894 53170 38946
rect 53678 38894 53730 38946
rect 55694 38894 55746 38946
rect 3278 38782 3330 38834
rect 3838 38782 3890 38834
rect 4174 38782 4226 38834
rect 4398 38782 4450 38834
rect 5294 38782 5346 38834
rect 6078 38782 6130 38834
rect 8206 38782 8258 38834
rect 8654 38782 8706 38834
rect 9102 38782 9154 38834
rect 9662 38782 9714 38834
rect 10334 38782 10386 38834
rect 11342 38782 11394 38834
rect 12686 38782 12738 38834
rect 13022 38782 13074 38834
rect 14814 38782 14866 38834
rect 15262 38782 15314 38834
rect 15822 38782 15874 38834
rect 16606 38782 16658 38834
rect 17502 38782 17554 38834
rect 18286 38782 18338 38834
rect 26238 38782 26290 38834
rect 28702 38782 28754 38834
rect 36206 38782 36258 38834
rect 36654 38782 36706 38834
rect 36878 38782 36930 38834
rect 37326 38782 37378 38834
rect 41918 38782 41970 38834
rect 49086 38782 49138 38834
rect 50542 38782 50594 38834
rect 51214 38782 51266 38834
rect 52446 38782 52498 38834
rect 52670 38782 52722 38834
rect 54014 38782 54066 38834
rect 55582 38782 55634 38834
rect 55806 38782 55858 38834
rect 1710 38670 1762 38722
rect 3390 38670 3442 38722
rect 4958 38670 5010 38722
rect 6638 38670 6690 38722
rect 9214 38670 9266 38722
rect 18846 38670 18898 38722
rect 21646 38670 21698 38722
rect 23998 38670 24050 38722
rect 26686 38670 26738 38722
rect 29262 38670 29314 38722
rect 34638 38670 34690 38722
rect 37886 38670 37938 38722
rect 40014 38670 40066 38722
rect 42366 38670 42418 38722
rect 44718 38670 44770 38722
rect 46958 38670 47010 38722
rect 49422 38670 49474 38722
rect 49870 38670 49922 38722
rect 54350 38670 54402 38722
rect 54910 38670 54962 38722
rect 55246 38670 55298 38722
rect 2830 38558 2882 38610
rect 3614 38558 3666 38610
rect 4062 38558 4114 38610
rect 7758 38558 7810 38610
rect 12910 38558 12962 38610
rect 15374 38558 15426 38610
rect 19966 38558 20018 38610
rect 22878 38558 22930 38610
rect 25118 38558 25170 38610
rect 27806 38558 27858 38610
rect 31838 38558 31890 38610
rect 32958 38558 33010 38610
rect 33518 38558 33570 38610
rect 39006 38558 39058 38610
rect 41246 38558 41298 38610
rect 45950 38558 46002 38610
rect 48750 38558 48802 38610
rect 50990 38558 51042 38610
rect 51102 38558 51154 38610
rect 52558 38558 52610 38610
rect 54686 38558 54738 38610
rect 56030 38558 56082 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 44466 38390 44518 38442
rect 44570 38390 44622 38442
rect 44674 38390 44726 38442
rect 7086 38222 7138 38274
rect 7310 38222 7362 38274
rect 9550 38222 9602 38274
rect 12126 38222 12178 38274
rect 13246 38222 13298 38274
rect 22766 38222 22818 38274
rect 26462 38222 26514 38274
rect 29262 38222 29314 38274
rect 33630 38222 33682 38274
rect 41470 38222 41522 38274
rect 44942 38222 44994 38274
rect 48190 38222 48242 38274
rect 50430 38222 50482 38274
rect 1598 38110 1650 38162
rect 4622 38110 4674 38162
rect 7422 38110 7474 38162
rect 7758 38110 7810 38162
rect 8318 38110 8370 38162
rect 8878 38110 8930 38162
rect 8990 38110 9042 38162
rect 11006 38110 11058 38162
rect 15150 38110 15202 38162
rect 18846 38110 18898 38162
rect 19854 38110 19906 38162
rect 20302 38110 20354 38162
rect 23886 38110 23938 38162
rect 29710 38110 29762 38162
rect 34078 38110 34130 38162
rect 37550 38110 37602 38162
rect 47294 38110 47346 38162
rect 48078 38110 48130 38162
rect 49310 38110 49362 38162
rect 51774 38110 51826 38162
rect 54126 38110 54178 38162
rect 56366 38110 56418 38162
rect 1262 37998 1314 38050
rect 3614 37998 3666 38050
rect 3950 37998 4002 38050
rect 4510 37998 4562 38050
rect 5182 37998 5234 38050
rect 5630 37998 5682 38050
rect 6638 37998 6690 38050
rect 8094 37998 8146 38050
rect 8206 37998 8258 38050
rect 9326 37998 9378 38050
rect 9774 37998 9826 38050
rect 9886 37998 9938 38050
rect 10558 37998 10610 38050
rect 15038 37998 15090 38050
rect 15710 37998 15762 38050
rect 19294 37998 19346 38050
rect 19630 37998 19682 38050
rect 21086 37998 21138 38050
rect 21870 37998 21922 38050
rect 23550 37998 23602 38050
rect 26014 37998 26066 38050
rect 28702 37998 28754 38050
rect 29038 37998 29090 38050
rect 29934 37998 29986 38050
rect 30494 37998 30546 38050
rect 31278 37998 31330 38050
rect 32958 37998 33010 38050
rect 33406 37998 33458 38050
rect 34638 37998 34690 38050
rect 35646 37998 35698 38050
rect 37886 37998 37938 38050
rect 42814 37998 42866 38050
rect 43710 37998 43762 38050
rect 44270 37998 44322 38050
rect 45054 37998 45106 38050
rect 45614 37998 45666 38050
rect 53566 37998 53618 38050
rect 56030 37998 56082 38050
rect 9662 37886 9714 37938
rect 12798 37886 12850 37938
rect 28254 37886 28306 37938
rect 32622 37886 32674 37938
rect 41918 37886 41970 37938
rect 42478 37886 42530 37938
rect 45950 37886 46002 37938
rect 46734 37886 46786 37938
rect 47294 37886 47346 37938
rect 48862 37886 48914 37938
rect 51438 37886 51490 37938
rect 2830 37774 2882 37826
rect 14366 37774 14418 37826
rect 16046 37774 16098 37826
rect 23102 37774 23154 37826
rect 27582 37774 27634 37826
rect 36318 37774 36370 37826
rect 40350 37774 40402 37826
rect 46958 37774 47010 37826
rect 47518 37774 47570 37826
rect 48190 37774 48242 37826
rect 53006 37774 53058 37826
rect 55246 37774 55298 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 43806 37606 43858 37658
rect 43910 37606 43962 37658
rect 44014 37606 44066 37658
rect 19966 37438 20018 37490
rect 50654 37438 50706 37490
rect 8094 37326 8146 37378
rect 28478 37326 28530 37378
rect 46286 37326 46338 37378
rect 48414 37326 48466 37378
rect 49086 37326 49138 37378
rect 52446 37326 52498 37378
rect 1374 37214 1426 37266
rect 2158 37214 2210 37266
rect 2942 37214 2994 37266
rect 3502 37214 3554 37266
rect 3950 37214 4002 37266
rect 5070 37214 5122 37266
rect 5854 37214 5906 37266
rect 10334 37214 10386 37266
rect 14926 37214 14978 37266
rect 15374 37214 15426 37266
rect 15934 37214 15986 37266
rect 16494 37214 16546 37266
rect 17614 37214 17666 37266
rect 18286 37214 18338 37266
rect 22206 37214 22258 37266
rect 24558 37214 24610 37266
rect 25006 37214 25058 37266
rect 25678 37214 25730 37266
rect 26462 37214 26514 37266
rect 27246 37214 27298 37266
rect 28814 37214 28866 37266
rect 29374 37214 29426 37266
rect 29934 37214 29986 37266
rect 30494 37214 30546 37266
rect 31390 37209 31442 37261
rect 32846 37214 32898 37266
rect 33406 37214 33458 37266
rect 34190 37214 34242 37266
rect 34638 37214 34690 37266
rect 35646 37214 35698 37266
rect 36766 37214 36818 37266
rect 39118 37214 39170 37266
rect 39678 37214 39730 37266
rect 40350 37214 40402 37266
rect 40910 37214 40962 37266
rect 41918 37214 41970 37266
rect 43262 37214 43314 37266
rect 45614 37214 45666 37266
rect 51102 37214 51154 37266
rect 54574 37214 54626 37266
rect 3390 37102 3442 37154
rect 4398 37102 4450 37154
rect 5294 37102 5346 37154
rect 6190 37102 6242 37154
rect 8430 37102 8482 37154
rect 10782 37102 10834 37154
rect 14478 37102 14530 37154
rect 18846 37102 18898 37154
rect 22542 37102 22594 37154
rect 24222 37102 24274 37154
rect 25230 37102 25282 37154
rect 29486 37102 29538 37154
rect 32510 37102 32562 37154
rect 33518 37102 33570 37154
rect 37214 37102 37266 37154
rect 38782 37102 38834 37154
rect 39790 37102 39842 37154
rect 42702 37102 42754 37154
rect 43598 37102 43650 37154
rect 44158 37102 44210 37154
rect 44494 37102 44546 37154
rect 44718 37102 44770 37154
rect 7422 36990 7474 37042
rect 9662 36990 9714 37042
rect 11902 36990 11954 37042
rect 15486 36990 15538 37042
rect 23774 36990 23826 37042
rect 38334 36990 38386 37042
rect 42814 36990 42866 37042
rect 43038 36990 43090 37042
rect 49534 36990 49586 37042
rect 51438 36990 51490 37042
rect 52894 36990 52946 37042
rect 54014 36990 54066 37042
rect 55134 36990 55186 37042
rect 56254 36990 56306 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 44466 36822 44518 36874
rect 44570 36822 44622 36874
rect 44674 36822 44726 36874
rect 6862 36654 6914 36706
rect 7198 36654 7250 36706
rect 7534 36654 7586 36706
rect 9214 36654 9266 36706
rect 9438 36654 9490 36706
rect 9662 36654 9714 36706
rect 16046 36654 16098 36706
rect 17390 36654 17442 36706
rect 25566 36654 25618 36706
rect 36206 36654 36258 36706
rect 42142 36654 42194 36706
rect 47070 36654 47122 36706
rect 54126 36654 54178 36706
rect 54238 36654 54290 36706
rect 54798 36654 54850 36706
rect 1598 36542 1650 36594
rect 3782 36542 3834 36594
rect 4286 36542 4338 36594
rect 7870 36542 7922 36594
rect 8318 36542 8370 36594
rect 8878 36542 8930 36594
rect 9774 36542 9826 36594
rect 11118 36542 11170 36594
rect 14926 36542 14978 36594
rect 18958 36542 19010 36594
rect 19966 36542 20018 36594
rect 20414 36542 20466 36594
rect 24558 36542 24610 36594
rect 26014 36542 26066 36594
rect 30158 36542 30210 36594
rect 33518 36542 33570 36594
rect 35198 36542 35250 36594
rect 36654 36542 36706 36594
rect 42590 36542 42642 36594
rect 45278 36542 45330 36594
rect 47294 36542 47346 36594
rect 55918 36542 55970 36594
rect 56142 36542 56194 36594
rect 1262 36430 1314 36482
rect 2830 36430 2882 36482
rect 4062 36430 4114 36482
rect 4734 36430 4786 36482
rect 5518 36430 5570 36482
rect 6302 36430 6354 36482
rect 10446 36430 10498 36482
rect 11006 36430 11058 36482
rect 11678 36430 11730 36482
rect 12126 36430 12178 36482
rect 12350 36430 12402 36482
rect 13134 36430 13186 36482
rect 14478 36430 14530 36482
rect 19406 36430 19458 36482
rect 19742 36430 19794 36482
rect 20974 36430 21026 36482
rect 22094 36430 22146 36482
rect 25006 36430 25058 36482
rect 25454 36430 25506 36482
rect 26798 36430 26850 36482
rect 27582 36430 27634 36482
rect 33182 36430 33234 36482
rect 34750 36430 34802 36482
rect 35534 36430 35586 36482
rect 35982 36430 36034 36482
rect 37438 36430 37490 36482
rect 38222 36430 38274 36482
rect 41582 36430 41634 36482
rect 41918 36430 41970 36482
rect 43150 36430 43202 36482
rect 44158 36430 44210 36482
rect 46958 36430 47010 36482
rect 47518 36430 47570 36482
rect 49534 36430 49586 36482
rect 53678 36430 53730 36482
rect 53902 36430 53954 36482
rect 54350 36430 54402 36482
rect 3278 36318 3330 36370
rect 8206 36318 8258 36370
rect 10110 36318 10162 36370
rect 16942 36318 16994 36370
rect 29822 36318 29874 36370
rect 41134 36318 41186 36370
rect 44942 36318 44994 36370
rect 52222 36318 52274 36370
rect 55358 36318 55410 36370
rect 18510 36206 18562 36258
rect 31390 36206 31442 36258
rect 46510 36206 46562 36258
rect 55134 36206 55186 36258
rect 56254 36206 56306 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 43806 36038 43858 36090
rect 43910 36038 43962 36090
rect 44014 36038 44066 36090
rect 23326 35870 23378 35922
rect 44270 35870 44322 35922
rect 48190 35870 48242 35922
rect 55358 35870 55410 35922
rect 4398 35758 4450 35810
rect 4958 35758 5010 35810
rect 21758 35758 21810 35810
rect 30606 35758 30658 35810
rect 38894 35758 38946 35810
rect 48862 35758 48914 35810
rect 52558 35758 52610 35810
rect 53230 35758 53282 35810
rect 54238 35758 54290 35810
rect 54798 35758 54850 35810
rect 55806 35758 55858 35810
rect 1486 35641 1538 35693
rect 2382 35646 2434 35698
rect 2830 35646 2882 35698
rect 3614 35646 3666 35698
rect 3950 35646 4002 35698
rect 5294 35646 5346 35698
rect 5742 35646 5794 35698
rect 6974 35646 7026 35698
rect 7982 35646 8034 35698
rect 9326 35646 9378 35698
rect 9774 35646 9826 35698
rect 10446 35646 10498 35698
rect 11230 35646 11282 35698
rect 12126 35646 12178 35698
rect 13918 35646 13970 35698
rect 20078 35646 20130 35698
rect 23998 35646 24050 35698
rect 26126 35646 26178 35698
rect 28702 35646 28754 35698
rect 31054 35646 31106 35698
rect 32174 35646 32226 35698
rect 32510 35646 32562 35698
rect 33294 35646 33346 35698
rect 33742 35646 33794 35698
rect 37998 35646 38050 35698
rect 39230 35646 39282 35698
rect 39790 35646 39842 35698
rect 40574 35646 40626 35698
rect 40910 35646 40962 35698
rect 42030 35646 42082 35698
rect 43374 35646 43426 35698
rect 45838 35646 45890 35698
rect 46622 35646 46674 35698
rect 52110 35646 52162 35698
rect 52334 35646 52386 35698
rect 52670 35646 52722 35698
rect 53454 35646 53506 35698
rect 54126 35646 54178 35698
rect 54910 35646 54962 35698
rect 55134 35646 55186 35698
rect 55694 35646 55746 35698
rect 6414 35534 6466 35586
rect 8990 35534 9042 35586
rect 9998 35534 10050 35586
rect 14366 35534 14418 35586
rect 19518 35534 19570 35586
rect 19742 35534 19794 35586
rect 22094 35534 22146 35586
rect 26686 35534 26738 35586
rect 33182 35534 33234 35586
rect 34190 35534 34242 35586
rect 37550 35534 37602 35586
rect 42926 35534 42978 35586
rect 43486 35534 43538 35586
rect 43710 35534 43762 35586
rect 45390 35534 45442 35586
rect 46958 35534 47010 35586
rect 49198 35534 49250 35586
rect 50878 35534 50930 35586
rect 51214 35534 51266 35586
rect 51438 35534 51490 35586
rect 52894 35534 52946 35586
rect 3390 35422 3442 35474
rect 5966 35422 6018 35474
rect 15486 35422 15538 35474
rect 19854 35422 19906 35474
rect 24446 35422 24498 35474
rect 25566 35422 25618 35474
rect 27806 35422 27858 35474
rect 29150 35422 29202 35474
rect 30270 35422 30322 35474
rect 36430 35422 36482 35474
rect 39902 35422 39954 35474
rect 43038 35422 43090 35474
rect 50430 35422 50482 35474
rect 50990 35422 51042 35474
rect 53790 35422 53842 35474
rect 54686 35422 54738 35474
rect 55918 35422 55970 35474
rect 56142 35422 56194 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 44466 35254 44518 35306
rect 44570 35254 44622 35306
rect 44674 35254 44726 35306
rect 19630 35086 19682 35138
rect 32510 35086 32562 35138
rect 33630 35086 33682 35138
rect 35646 35086 35698 35138
rect 44830 35086 44882 35138
rect 47182 35086 47234 35138
rect 54798 35086 54850 35138
rect 55246 35086 55298 35138
rect 1598 34974 1650 35026
rect 2830 34974 2882 35026
rect 3390 34974 3442 35026
rect 5294 34974 5346 35026
rect 7982 34974 8034 35026
rect 8094 34974 8146 35026
rect 11006 34974 11058 35026
rect 14814 34974 14866 35026
rect 17278 34974 17330 35026
rect 19070 34974 19122 35026
rect 19182 34974 19234 35026
rect 21758 34974 21810 35026
rect 22206 34974 22258 35026
rect 25678 34974 25730 35026
rect 28254 34974 28306 35026
rect 28702 34974 28754 35026
rect 41582 34974 41634 35026
rect 43150 34974 43202 35026
rect 45950 34974 46002 35026
rect 47406 34974 47458 35026
rect 49982 34974 50034 35026
rect 51326 34974 51378 35026
rect 54686 34974 54738 35026
rect 56142 34974 56194 35026
rect 3502 34862 3554 34914
rect 3614 34862 3666 34914
rect 3726 34862 3778 34914
rect 3950 34862 4002 34914
rect 4622 34862 4674 34914
rect 5070 34862 5122 34914
rect 5854 34862 5906 34914
rect 6302 34862 6354 34914
rect 7310 34862 7362 34914
rect 7758 34862 7810 34914
rect 10334 34862 10386 34914
rect 10894 34862 10946 34914
rect 11678 34862 11730 34914
rect 12014 34862 12066 34914
rect 13022 34862 13074 34914
rect 15374 34862 15426 34914
rect 19742 34862 19794 34914
rect 19966 34862 20018 34914
rect 20190 34862 20242 34914
rect 21086 34862 21138 34914
rect 21646 34862 21698 34914
rect 22766 34862 22818 34914
rect 23886 34862 23938 34914
rect 25230 34862 25282 34914
rect 27694 34862 27746 34914
rect 28030 34862 28082 34914
rect 29486 34862 29538 34914
rect 30382 34862 30434 34914
rect 35086 34862 35138 34914
rect 35422 34862 35474 34914
rect 36318 34862 36370 34914
rect 36878 34862 36930 34914
rect 37774 34862 37826 34914
rect 42030 34862 42082 34914
rect 46398 34862 46450 34914
rect 46958 34862 47010 34914
rect 52222 34862 52274 34914
rect 54574 34862 54626 34914
rect 1262 34750 1314 34802
rect 4286 34750 4338 34802
rect 9998 34750 10050 34802
rect 16942 34750 16994 34802
rect 19854 34750 19906 34802
rect 20750 34750 20802 34802
rect 27246 34750 27298 34802
rect 34078 34750 34130 34802
rect 34638 34750 34690 34802
rect 42702 34750 42754 34802
rect 47070 34750 47122 34802
rect 54350 34750 54402 34802
rect 55358 34750 55410 34802
rect 56142 34750 56194 34802
rect 13694 34638 13746 34690
rect 18510 34638 18562 34690
rect 19070 34638 19122 34690
rect 26798 34638 26850 34690
rect 40350 34638 40402 34690
rect 44270 34638 44322 34690
rect 54126 34638 54178 34690
rect 55918 34638 55970 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 43806 34470 43858 34522
rect 43910 34470 43962 34522
rect 44014 34470 44066 34522
rect 19070 34302 19122 34354
rect 35198 34302 35250 34354
rect 45614 34302 45666 34354
rect 50318 34302 50370 34354
rect 54686 34302 54738 34354
rect 5070 34190 5122 34242
rect 10558 34190 10610 34242
rect 14030 34190 14082 34242
rect 29822 34190 29874 34242
rect 33630 34190 33682 34242
rect 37326 34190 37378 34242
rect 46286 34190 46338 34242
rect 48302 34190 48354 34242
rect 50878 34190 50930 34242
rect 52558 34190 52610 34242
rect 55694 34190 55746 34242
rect 1262 34078 1314 34130
rect 3838 34078 3890 34130
rect 3950 34078 4002 34130
rect 4174 34078 4226 34130
rect 4846 34078 4898 34130
rect 6078 34078 6130 34130
rect 9886 34078 9938 34130
rect 14478 34078 14530 34130
rect 14814 34078 14866 34130
rect 15486 34078 15538 34130
rect 16158 34078 16210 34130
rect 17054 34078 17106 34130
rect 18622 34078 18674 34130
rect 19630 34078 19682 34130
rect 20078 34078 20130 34130
rect 20526 34078 20578 34130
rect 20862 34078 20914 34130
rect 22430 34078 22482 34130
rect 24894 34078 24946 34130
rect 25342 34078 25394 34130
rect 26014 34078 26066 34130
rect 26686 34078 26738 34130
rect 27582 34078 27634 34130
rect 30270 34078 30322 34130
rect 30606 34078 30658 34130
rect 31278 34078 31330 34130
rect 32062 34078 32114 34130
rect 32846 34078 32898 34130
rect 36766 34078 36818 34130
rect 38110 34078 38162 34130
rect 39006 34078 39058 34130
rect 39566 34078 39618 34130
rect 40350 34078 40402 34130
rect 40798 34078 40850 34130
rect 43374 34078 43426 34130
rect 44830 34078 44882 34130
rect 45278 34078 45330 34130
rect 46062 34078 46114 34130
rect 47854 34078 47906 34130
rect 50542 34078 50594 34130
rect 52222 34078 52274 34130
rect 53118 34078 53170 34130
rect 55358 34078 55410 34130
rect 55918 34078 55970 34130
rect 3278 33966 3330 34018
rect 4398 33966 4450 34018
rect 5294 33966 5346 34018
rect 5518 33966 5570 34018
rect 6526 33966 6578 34018
rect 15038 33966 15090 34018
rect 18510 33966 18562 34018
rect 18958 33966 19010 34018
rect 19406 33966 19458 34018
rect 20750 33966 20802 34018
rect 24558 33966 24610 34018
rect 25566 33966 25618 34018
rect 30830 33966 30882 34018
rect 34078 33966 34130 34018
rect 37438 33966 37490 34018
rect 40238 33966 40290 34018
rect 41246 33966 41298 34018
rect 42814 33966 42866 34018
rect 44718 33966 44770 34018
rect 46286 33966 46338 34018
rect 46398 33966 46450 34018
rect 46622 33966 46674 34018
rect 47182 33966 47234 34018
rect 47294 33966 47346 34018
rect 48638 33966 48690 34018
rect 50766 33966 50818 34018
rect 50990 33966 51042 34018
rect 51998 33966 52050 34018
rect 53566 33966 53618 34018
rect 1710 33854 1762 33906
rect 2830 33854 2882 33906
rect 3390 33854 3442 33906
rect 3614 33854 3666 33906
rect 7646 33854 7698 33906
rect 8206 33854 8258 33906
rect 9326 33854 9378 33906
rect 11006 33854 11058 33906
rect 12126 33854 12178 33906
rect 19854 33854 19906 33906
rect 22990 33854 23042 33906
rect 24110 33854 24162 33906
rect 37214 33854 37266 33906
rect 41694 33854 41746 33906
rect 47406 33854 47458 33906
rect 49870 33854 49922 33906
rect 55246 33854 55298 33906
rect 55470 33854 55522 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 44466 33686 44518 33738
rect 44570 33686 44622 33738
rect 44674 33686 44726 33738
rect 1374 33518 1426 33570
rect 2494 33518 2546 33570
rect 2718 33518 2770 33570
rect 3950 33518 4002 33570
rect 6526 33518 6578 33570
rect 13918 33518 13970 33570
rect 18510 33518 18562 33570
rect 20526 33518 20578 33570
rect 33070 33518 33122 33570
rect 38446 33518 38498 33570
rect 39566 33518 39618 33570
rect 40910 33518 40962 33570
rect 53902 33518 53954 33570
rect 55022 33518 55074 33570
rect 2046 33406 2098 33458
rect 2382 33406 2434 33458
rect 6638 33406 6690 33458
rect 8094 33406 8146 33458
rect 9886 33406 9938 33458
rect 14366 33406 14418 33458
rect 17390 33406 17442 33458
rect 19518 33406 19570 33458
rect 20974 33406 21026 33458
rect 27582 33406 27634 33458
rect 28030 33406 28082 33458
rect 32958 33406 33010 33458
rect 35870 33406 35922 33458
rect 40798 33406 40850 33458
rect 44606 33406 44658 33458
rect 47518 33406 47570 33458
rect 48750 33406 48802 33458
rect 52670 33406 52722 33458
rect 56030 33406 56082 33458
rect 56366 33406 56418 33458
rect 1150 33294 1202 33346
rect 1822 33294 1874 33346
rect 3390 33294 3442 33346
rect 3726 33294 3778 33346
rect 4398 33294 4450 33346
rect 5070 33294 5122 33346
rect 5966 33294 6018 33346
rect 7086 33294 7138 33346
rect 7422 33294 7474 33346
rect 8206 33294 8258 33346
rect 9214 33294 9266 33346
rect 9774 33294 9826 33346
rect 10334 33294 10386 33346
rect 10894 33294 10946 33346
rect 12014 33294 12066 33346
rect 13246 33294 13298 33346
rect 13806 33294 13858 33346
rect 14926 33294 14978 33346
rect 16046 33294 16098 33346
rect 19966 33294 20018 33346
rect 20414 33282 20466 33334
rect 21758 33294 21810 33346
rect 22654 33294 22706 33346
rect 27022 33294 27074 33346
rect 27358 33294 27410 33346
rect 28590 33294 28642 33346
rect 29710 33294 29762 33346
rect 32510 33294 32562 33346
rect 35422 33294 35474 33346
rect 36990 33294 37042 33346
rect 37998 33294 38050 33346
rect 44046 33294 44098 33346
rect 44382 33294 44434 33346
rect 45278 33294 45330 33346
rect 45614 33294 45666 33346
rect 46622 33294 46674 33346
rect 47182 33294 47234 33346
rect 50654 33294 50706 33346
rect 51326 33294 51378 33346
rect 51550 33294 51602 33346
rect 51886 33294 51938 33346
rect 52222 33294 52274 33346
rect 52446 33294 52498 33346
rect 2942 33182 2994 33234
rect 8878 33182 8930 33234
rect 12910 33182 12962 33234
rect 16942 33182 16994 33234
rect 26574 33182 26626 33234
rect 40462 33182 40514 33234
rect 43598 33182 43650 33234
rect 48414 33182 48466 33234
rect 50430 33182 50482 33234
rect 51438 33182 51490 33234
rect 52334 33182 52386 33234
rect 53454 33182 53506 33234
rect 34190 33070 34242 33122
rect 42030 33070 42082 33122
rect 49982 33070 50034 33122
rect 50990 33070 51042 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 43806 32902 43858 32954
rect 43910 32902 43962 32954
rect 44014 32902 44066 32954
rect 7982 32734 8034 32786
rect 45950 32734 46002 32786
rect 50094 32734 50146 32786
rect 1262 32622 1314 32674
rect 4174 32622 4226 32674
rect 8430 32622 8482 32674
rect 15486 32622 15538 32674
rect 20862 32622 20914 32674
rect 26126 32622 26178 32674
rect 28814 32622 28866 32674
rect 37998 32622 38050 32674
rect 40350 32622 40402 32674
rect 44382 32622 44434 32674
rect 3838 32510 3890 32562
rect 6414 32510 6466 32562
rect 8766 32510 8818 32562
rect 9214 32510 9266 32562
rect 9886 32510 9938 32562
rect 10670 32510 10722 32562
rect 11454 32510 11506 32562
rect 13470 32510 13522 32562
rect 15038 32510 15090 32562
rect 15822 32510 15874 32562
rect 16270 32510 16322 32562
rect 17502 32510 17554 32562
rect 18510 32510 18562 32562
rect 23102 32510 23154 32562
rect 23886 32510 23938 32562
rect 24110 32510 24162 32562
rect 24446 32510 24498 32562
rect 25342 32510 25394 32562
rect 25678 32510 25730 32562
rect 29934 32510 29986 32562
rect 32286 32510 32338 32562
rect 33070 32510 33122 32562
rect 34414 32510 34466 32562
rect 34862 32510 34914 32562
rect 38558 32510 38610 32562
rect 39230 32510 39282 32562
rect 40686 32510 40738 32562
rect 41134 32510 41186 32562
rect 41806 32510 41858 32562
rect 42478 32510 42530 32562
rect 43486 32510 43538 32562
rect 46622 32510 46674 32562
rect 48638 32510 48690 32562
rect 48974 32510 49026 32562
rect 50878 32510 50930 32562
rect 51102 32510 51154 32562
rect 51998 32510 52050 32562
rect 52670 32510 52722 32562
rect 52894 32510 52946 32562
rect 54574 32510 54626 32562
rect 54798 32510 54850 32562
rect 1710 32398 1762 32450
rect 3278 32398 3330 32450
rect 3390 32398 3442 32450
rect 4958 32398 5010 32450
rect 5854 32398 5906 32450
rect 6750 32398 6802 32450
rect 9438 32398 9490 32450
rect 16942 32398 16994 32450
rect 21310 32398 21362 32450
rect 29262 32398 29314 32450
rect 30494 32398 30546 32450
rect 33854 32398 33906 32450
rect 34302 32398 34354 32450
rect 35310 32398 35362 32450
rect 38782 32398 38834 32450
rect 38894 32398 38946 32450
rect 46958 32398 47010 32450
rect 48750 32398 48802 32450
rect 49310 32398 49362 32450
rect 49870 32398 49922 32450
rect 53342 32398 53394 32450
rect 53790 32398 53842 32450
rect 55694 32398 55746 32450
rect 56030 32398 56082 32450
rect 2830 32286 2882 32338
rect 3950 32286 4002 32338
rect 4174 32286 4226 32338
rect 4286 32286 4338 32338
rect 5294 32286 5346 32338
rect 5518 32286 5570 32338
rect 5742 32286 5794 32338
rect 13918 32286 13970 32338
rect 16494 32286 16546 32338
rect 22430 32286 22482 32338
rect 25118 32286 25170 32338
rect 28926 32286 28978 32338
rect 29374 32286 29426 32338
rect 29598 32286 29650 32338
rect 31614 32286 31666 32338
rect 36430 32286 36482 32338
rect 37550 32286 37602 32338
rect 38670 32286 38722 32338
rect 41358 32286 41410 32338
rect 44830 32286 44882 32338
rect 48190 32286 48242 32338
rect 50430 32286 50482 32338
rect 51438 32286 51490 32338
rect 52334 32286 52386 32338
rect 53118 32286 53170 32338
rect 53230 32286 53282 32338
rect 54126 32286 54178 32338
rect 55022 32286 55074 32338
rect 55134 32286 55186 32338
rect 55246 32286 55298 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 44466 32118 44518 32170
rect 44570 32118 44622 32170
rect 44674 32118 44726 32170
rect 2830 31950 2882 32002
rect 34190 31950 34242 32002
rect 50206 31950 50258 32002
rect 52894 31950 52946 32002
rect 1598 31838 1650 31890
rect 3614 31838 3666 31890
rect 4958 31838 5010 31890
rect 7534 31838 7586 31890
rect 7646 31838 7698 31890
rect 8206 31838 8258 31890
rect 9886 31838 9938 31890
rect 10334 31838 10386 31890
rect 14926 31838 14978 31890
rect 16046 31838 16098 31890
rect 20414 31838 20466 31890
rect 22654 31838 22706 31890
rect 25230 31838 25282 31890
rect 25566 31838 25618 31890
rect 27470 31838 27522 31890
rect 33070 31838 33122 31890
rect 34750 31838 34802 31890
rect 34974 31838 35026 31890
rect 35422 31838 35474 31890
rect 35534 31838 35586 31890
rect 37326 31838 37378 31890
rect 41246 31838 41298 31890
rect 42254 31838 42306 31890
rect 45390 31838 45442 31890
rect 47182 31838 47234 31890
rect 47406 31838 47458 31890
rect 48190 31838 48242 31890
rect 49422 31838 49474 31890
rect 50654 31838 50706 31890
rect 51774 31838 51826 31890
rect 54126 31838 54178 31890
rect 55246 31838 55298 31890
rect 56366 31838 56418 31890
rect 1262 31726 1314 31778
rect 3390 31726 3442 31778
rect 4286 31726 4338 31778
rect 4846 31726 4898 31778
rect 5406 31726 5458 31778
rect 6190 31726 6242 31778
rect 7086 31726 7138 31778
rect 7870 31726 7922 31778
rect 8318 31726 8370 31778
rect 9214 31726 9266 31778
rect 9774 31726 9826 31778
rect 10894 31726 10946 31778
rect 11902 31726 11954 31778
rect 18286 31726 18338 31778
rect 19406 31726 19458 31778
rect 19966 31726 20018 31778
rect 20638 31726 20690 31778
rect 20974 31726 21026 31778
rect 23886 31726 23938 31778
rect 25006 31726 25058 31778
rect 26910 31726 26962 31778
rect 27358 31726 27410 31778
rect 27918 31726 27970 31778
rect 28590 31726 28642 31778
rect 29598 31726 29650 31778
rect 32510 31726 32562 31778
rect 34638 31726 34690 31778
rect 35198 31726 35250 31778
rect 35310 31726 35362 31778
rect 35870 31726 35922 31778
rect 36766 31726 36818 31778
rect 37102 31726 37154 31778
rect 37886 31726 37938 31778
rect 38446 31726 38498 31778
rect 39342 31726 39394 31778
rect 41694 31726 41746 31778
rect 42030 31726 42082 31778
rect 42814 31726 42866 31778
rect 43262 31726 43314 31778
rect 44270 31726 44322 31778
rect 45054 31726 45106 31778
rect 48078 31726 48130 31778
rect 48414 31726 48466 31778
rect 48526 31726 48578 31778
rect 49086 31726 49138 31778
rect 49758 31726 49810 31778
rect 50094 31726 50146 31778
rect 50430 31726 50482 31778
rect 56030 31726 56082 31778
rect 3950 31614 4002 31666
rect 8878 31614 8930 31666
rect 14478 31614 14530 31666
rect 21422 31614 21474 31666
rect 22318 31614 22370 31666
rect 24670 31614 24722 31666
rect 26462 31614 26514 31666
rect 36318 31614 36370 31666
rect 51326 31614 51378 31666
rect 53678 31614 53730 31666
rect 8206 31502 8258 31554
rect 46622 31502 46674 31554
rect 47070 31502 47122 31554
rect 50206 31502 50258 31554
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 43806 31334 43858 31386
rect 43910 31334 43962 31386
rect 44014 31334 44066 31386
rect 22430 31166 22482 31218
rect 42814 31166 42866 31218
rect 48526 31166 48578 31218
rect 51326 31166 51378 31218
rect 53790 31166 53842 31218
rect 56030 31166 56082 31218
rect 5070 31054 5122 31106
rect 6190 31054 6242 31106
rect 8206 31054 8258 31106
rect 16830 31054 16882 31106
rect 20862 31054 20914 31106
rect 26126 31054 26178 31106
rect 28926 31054 28978 31106
rect 29934 31054 29986 31106
rect 36542 31054 36594 31106
rect 38782 31054 38834 31106
rect 43486 31054 43538 31106
rect 47518 31054 47570 31106
rect 1374 30942 1426 30994
rect 2382 30942 2434 30994
rect 3614 30942 3666 30994
rect 3950 30942 4002 30994
rect 4958 30942 5010 30994
rect 5182 30942 5234 30994
rect 8542 30942 8594 30994
rect 8990 30942 9042 30994
rect 9886 30942 9938 30994
rect 10334 30942 10386 30994
rect 11342 30942 11394 30994
rect 13470 30942 13522 30994
rect 13918 30942 13970 30994
rect 15150 30942 15202 30994
rect 16270 30942 16322 30994
rect 17166 30942 17218 30994
rect 17614 30942 17666 30994
rect 18510 30942 18562 30994
rect 18846 30942 18898 30994
rect 19854 30942 19906 30994
rect 23102 30942 23154 30994
rect 23886 30942 23938 30994
rect 24110 30942 24162 30994
rect 24558 30942 24610 30994
rect 25230 30942 25282 30994
rect 25678 30942 25730 30994
rect 26798 30942 26850 30994
rect 27470 30942 27522 30994
rect 32398 30942 32450 30994
rect 32734 30942 32786 30994
rect 34078 30942 34130 30994
rect 34974 30942 35026 30994
rect 35870 30942 35922 30994
rect 41134 30942 41186 30994
rect 45166 30942 45218 30994
rect 47854 30942 47906 30994
rect 48414 30942 48466 30994
rect 49198 30942 49250 30994
rect 51214 30942 51266 30994
rect 52222 30942 52274 30994
rect 54350 30942 54402 30994
rect 2942 30830 2994 30882
rect 4398 30830 4450 30882
rect 5518 30830 5570 30882
rect 13134 30830 13186 30882
rect 14142 30830 14194 30882
rect 14590 30830 14642 30882
rect 17838 30830 17890 30882
rect 21198 30830 21250 30882
rect 25118 30830 25170 30882
rect 26686 30830 26738 30882
rect 30382 30830 30434 30882
rect 31950 30830 32002 30882
rect 33406 30830 33458 30882
rect 35534 30830 35586 30882
rect 35646 30830 35698 30882
rect 39118 30830 39170 30882
rect 41582 30830 41634 30882
rect 44382 30830 44434 30882
rect 44494 30830 44546 30882
rect 44718 30830 44770 30882
rect 47406 30830 47458 30882
rect 47518 30830 47570 30882
rect 48526 30830 48578 30882
rect 52670 30830 52722 30882
rect 3390 30718 3442 30770
rect 6638 30718 6690 30770
rect 7758 30718 7810 30770
rect 9214 30718 9266 30770
rect 21310 30718 21362 30770
rect 27806 30718 27858 30770
rect 28814 30718 28866 30770
rect 29038 30718 29090 30770
rect 29262 30718 29314 30770
rect 31502 30718 31554 30770
rect 32958 30718 33010 30770
rect 36990 30718 37042 30770
rect 38110 30718 38162 30770
rect 40350 30718 40402 30770
rect 43598 30718 43650 30770
rect 45614 30718 45666 30770
rect 46734 30718 46786 30770
rect 47182 30718 47234 30770
rect 49646 30718 49698 30770
rect 50766 30718 50818 30770
rect 51326 30718 51378 30770
rect 54910 30718 54962 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 44466 30550 44518 30602
rect 44570 30550 44622 30602
rect 44674 30550 44726 30602
rect 2830 30382 2882 30434
rect 9326 30382 9378 30434
rect 9550 30382 9602 30434
rect 13806 30382 13858 30434
rect 14926 30382 14978 30434
rect 17950 30382 18002 30434
rect 19070 30382 19122 30434
rect 27246 30382 27298 30434
rect 29934 30382 29986 30434
rect 30046 30382 30098 30434
rect 30158 30382 30210 30434
rect 36654 30382 36706 30434
rect 38446 30382 38498 30434
rect 38670 30382 38722 30434
rect 50094 30382 50146 30434
rect 52222 30382 52274 30434
rect 1598 30270 1650 30322
rect 4622 30270 4674 30322
rect 12686 30270 12738 30322
rect 16830 30270 16882 30322
rect 16942 30270 16994 30322
rect 20526 30270 20578 30322
rect 26014 30270 26066 30322
rect 28366 30270 28418 30322
rect 30494 30270 30546 30322
rect 33406 30270 33458 30322
rect 38222 30270 38274 30322
rect 39230 30270 39282 30322
rect 39342 30326 39394 30378
rect 52334 30382 52386 30434
rect 56142 30382 56194 30434
rect 41246 30270 41298 30322
rect 45054 30270 45106 30322
rect 47182 30270 47234 30322
rect 47406 30270 47458 30322
rect 48974 30270 49026 30322
rect 51214 30270 51266 30322
rect 52110 30270 52162 30322
rect 53678 30270 53730 30322
rect 55918 30270 55970 30322
rect 1262 30158 1314 30210
rect 4062 30158 4114 30210
rect 4510 30158 4562 30210
rect 5294 30158 5346 30210
rect 5630 30158 5682 30210
rect 6638 30158 6690 30210
rect 7758 30158 7810 30210
rect 9102 30158 9154 30210
rect 9438 30158 9490 30210
rect 9774 30158 9826 30210
rect 10110 30158 10162 30210
rect 10222 30158 10274 30210
rect 10334 30158 10386 30210
rect 10558 30158 10610 30210
rect 12238 30158 12290 30210
rect 14478 30158 14530 30210
rect 16046 30158 16098 30210
rect 17390 30158 17442 30210
rect 19966 30158 20018 30210
rect 20414 30158 20466 30210
rect 20974 30158 21026 30210
rect 21534 30158 21586 30210
rect 22654 30158 22706 30210
rect 29486 30158 29538 30210
rect 30382 30158 30434 30210
rect 31502 30158 31554 30210
rect 32734 30158 32786 30210
rect 33182 30158 33234 30210
rect 33966 30158 34018 30210
rect 34526 30158 34578 30210
rect 35534 30158 35586 30210
rect 40238 30158 40290 30210
rect 40574 30158 40626 30210
rect 41022 30158 41074 30210
rect 41918 30158 41970 30210
rect 42366 30158 42418 30210
rect 43262 30158 43314 30210
rect 44494 30158 44546 30210
rect 46174 30158 46226 30210
rect 46734 30158 46786 30210
rect 46958 30158 47010 30210
rect 47294 30158 47346 30210
rect 48302 30158 48354 30210
rect 49534 30158 49586 30210
rect 51662 30158 51714 30210
rect 51886 30158 51938 30210
rect 54910 30158 54962 30210
rect 3614 30046 3666 30098
rect 8206 30046 8258 30098
rect 19518 30046 19570 30098
rect 25678 30046 25730 30098
rect 27918 30046 27970 30098
rect 31278 30046 31330 30098
rect 32398 30046 32450 30098
rect 36206 30046 36258 30098
rect 38334 30046 38386 30098
rect 53342 30046 53394 30098
rect 56030 30046 56082 30098
rect 7870 29934 7922 29986
rect 8318 29934 8370 29986
rect 16830 29934 16882 29986
rect 31838 29934 31890 29986
rect 37774 29934 37826 29986
rect 39230 29934 39282 29986
rect 48190 29934 48242 29986
rect 48526 29934 48578 29986
rect 48638 29934 48690 29986
rect 49086 29934 49138 29986
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 43806 29766 43858 29818
rect 43910 29766 43962 29818
rect 44014 29766 44066 29818
rect 5854 29598 5906 29650
rect 6302 29598 6354 29650
rect 8990 29598 9042 29650
rect 12910 29598 12962 29650
rect 23326 29598 23378 29650
rect 27806 29598 27858 29650
rect 34750 29598 34802 29650
rect 36430 29598 36482 29650
rect 42142 29598 42194 29650
rect 53230 29598 53282 29650
rect 55470 29598 55522 29650
rect 1262 29486 1314 29538
rect 4174 29486 4226 29538
rect 6414 29486 6466 29538
rect 20078 29486 20130 29538
rect 21758 29486 21810 29538
rect 23998 29486 24050 29538
rect 26238 29486 26290 29538
rect 33966 29486 34018 29538
rect 46846 29486 46898 29538
rect 52558 29486 52610 29538
rect 2830 29374 2882 29426
rect 3838 29374 3890 29426
rect 4062 29374 4114 29426
rect 4398 29374 4450 29426
rect 5182 29374 5234 29426
rect 5406 29374 5458 29426
rect 5966 29374 6018 29426
rect 7422 29374 7474 29426
rect 9326 29374 9378 29426
rect 9662 29374 9714 29426
rect 9886 29374 9938 29426
rect 11678 29374 11730 29426
rect 14478 29374 14530 29426
rect 17166 29369 17218 29421
rect 17838 29374 17890 29426
rect 18510 29374 18562 29426
rect 19182 29374 19234 29426
rect 19630 29374 19682 29426
rect 20862 29374 20914 29426
rect 21086 29374 21138 29426
rect 28702 29374 28754 29426
rect 30830 29374 30882 29426
rect 31838 29374 31890 29426
rect 32510 29374 32562 29426
rect 33070 29374 33122 29426
rect 33630 29374 33682 29426
rect 34862 29374 34914 29426
rect 35646 29374 35698 29426
rect 37214 29374 37266 29426
rect 37662 29374 37714 29426
rect 38334 29374 38386 29426
rect 38782 29374 38834 29426
rect 39790 29374 39842 29426
rect 40462 29374 40514 29426
rect 45838 29374 45890 29426
rect 46622 29374 46674 29426
rect 47518 29374 47570 29426
rect 49534 29374 49586 29426
rect 50318 29374 50370 29426
rect 50766 29374 50818 29426
rect 50990 29374 51042 29426
rect 52110 29374 52162 29426
rect 52782 29374 52834 29426
rect 53342 29374 53394 29426
rect 53902 29374 53954 29426
rect 1598 29262 1650 29314
rect 3278 29262 3330 29314
rect 4958 29262 5010 29314
rect 7758 29262 7810 29314
rect 11230 29262 11282 29314
rect 11902 29262 11954 29314
rect 12238 29262 12290 29314
rect 14142 29262 14194 29314
rect 16382 29262 16434 29314
rect 19070 29262 19122 29314
rect 20638 29262 20690 29314
rect 22094 29262 22146 29314
rect 24446 29262 24498 29314
rect 26574 29262 26626 29314
rect 32958 29262 33010 29314
rect 34302 29262 34354 29314
rect 34526 29262 34578 29314
rect 35534 29262 35586 29314
rect 36318 29262 36370 29314
rect 36766 29262 36818 29314
rect 37774 29262 37826 29314
rect 45502 29262 45554 29314
rect 46398 29262 46450 29314
rect 46958 29262 47010 29314
rect 49870 29262 49922 29314
rect 50206 29262 50258 29314
rect 52446 29262 52498 29314
rect 54238 29262 54290 29314
rect 3390 29150 3442 29202
rect 5070 29150 5122 29202
rect 9550 29150 9602 29202
rect 11342 29150 11394 29202
rect 12126 29150 12178 29202
rect 16494 29150 16546 29202
rect 20750 29150 20802 29202
rect 25566 29150 25618 29202
rect 29150 29150 29202 29202
rect 30270 29150 30322 29202
rect 35086 29150 35138 29202
rect 35310 29150 35362 29202
rect 41022 29150 41074 29202
rect 44270 29150 44322 29202
rect 47966 29150 48018 29202
rect 49086 29150 49138 29202
rect 49758 29150 49810 29202
rect 51102 29150 51154 29202
rect 52558 29150 52610 29202
rect 53230 29150 53282 29202
rect 55918 29150 55970 29202
rect 56254 29150 56306 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 44466 28982 44518 29034
rect 44570 28982 44622 29034
rect 44674 28982 44726 29034
rect 2830 28814 2882 28866
rect 11902 28814 11954 28866
rect 18510 28814 18562 28866
rect 19070 28814 19122 28866
rect 19182 28814 19234 28866
rect 19406 28814 19458 28866
rect 19854 28814 19906 28866
rect 20078 28814 20130 28866
rect 26462 28814 26514 28866
rect 29038 28814 29090 28866
rect 31726 28814 31778 28866
rect 38334 28814 38386 28866
rect 38782 28814 38834 28866
rect 40910 28814 40962 28866
rect 46286 28814 46338 28866
rect 46398 28814 46450 28866
rect 46510 28814 46562 28866
rect 46734 28814 46786 28866
rect 51102 28814 51154 28866
rect 53342 28814 53394 28866
rect 55022 28814 55074 28866
rect 55918 28814 55970 28866
rect 56254 28814 56306 28866
rect 1598 28702 1650 28754
rect 3502 28702 3554 28754
rect 4958 28702 5010 28754
rect 7534 28702 7586 28754
rect 9326 28702 9378 28754
rect 10782 28702 10834 28754
rect 13582 28702 13634 28754
rect 17390 28702 17442 28754
rect 20190 28702 20242 28754
rect 20638 28702 20690 28754
rect 21646 28702 21698 28754
rect 27582 28702 27634 28754
rect 28030 28702 28082 28754
rect 31614 28702 31666 28754
rect 32398 28702 32450 28754
rect 33406 28702 33458 28754
rect 36094 28702 36146 28754
rect 37214 28702 37266 28754
rect 43710 28702 43762 28754
rect 47406 28702 47458 28754
rect 47630 28702 47682 28754
rect 49310 28702 49362 28754
rect 50094 28702 50146 28754
rect 3278 28590 3330 28642
rect 3614 28590 3666 28642
rect 3950 28590 4002 28642
rect 4398 28590 4450 28642
rect 4846 28590 4898 28642
rect 5406 28590 5458 28642
rect 6078 28590 6130 28642
rect 7086 28590 7138 28642
rect 7758 28590 7810 28642
rect 8206 28590 8258 28642
rect 8878 28590 8930 28642
rect 9102 28590 9154 28642
rect 12574 28590 12626 28642
rect 13022 28590 13074 28642
rect 13358 28590 13410 28642
rect 14254 28590 14306 28642
rect 14590 28590 14642 28642
rect 15598 28590 15650 28642
rect 16942 28590 16994 28642
rect 19630 28590 19682 28642
rect 20974 28590 21026 28642
rect 21422 28590 21474 28642
rect 22094 28590 22146 28642
rect 22654 28590 22706 28642
rect 23662 28590 23714 28642
rect 28366 28590 28418 28642
rect 28926 28590 28978 28642
rect 29710 28590 29762 28642
rect 30046 28590 30098 28642
rect 31054 28590 31106 28642
rect 32734 28590 32786 28642
rect 33182 28590 33234 28642
rect 34078 28590 34130 28642
rect 34414 28590 34466 28642
rect 35534 28590 35586 28642
rect 35982 28590 36034 28642
rect 36318 28590 36370 28642
rect 36654 28590 36706 28642
rect 39006 28590 39058 28642
rect 39454 28590 39506 28642
rect 40462 28590 40514 28642
rect 43150 28590 43202 28642
rect 43486 28590 43538 28642
rect 44270 28590 44322 28642
rect 44718 28590 44770 28642
rect 45726 28590 45778 28642
rect 47294 28590 47346 28642
rect 48190 28590 48242 28642
rect 48974 28590 49026 28642
rect 49758 28590 49810 28642
rect 52894 28590 52946 28642
rect 53118 28590 53170 28642
rect 53902 28590 53954 28642
rect 54126 28590 54178 28642
rect 54350 28590 54402 28642
rect 1262 28478 1314 28530
rect 8990 28478 9042 28530
rect 10334 28478 10386 28530
rect 19294 28478 19346 28530
rect 26014 28478 26066 28530
rect 38894 28478 38946 28530
rect 42702 28478 42754 28530
rect 50654 28478 50706 28530
rect 53230 28478 53282 28530
rect 54014 28478 54066 28530
rect 8318 28366 8370 28418
rect 31726 28366 31778 28418
rect 42030 28366 42082 28418
rect 48526 28366 48578 28418
rect 52222 28366 52274 28418
rect 52670 28366 52722 28418
rect 54574 28366 54626 28418
rect 54910 28366 54962 28418
rect 55246 28366 55298 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 43806 28198 43858 28250
rect 43910 28198 43962 28250
rect 44014 28198 44066 28250
rect 11454 28030 11506 28082
rect 20750 28030 20802 28082
rect 32510 28030 32562 28082
rect 33070 28030 33122 28082
rect 38110 28030 38162 28082
rect 43374 28030 43426 28082
rect 44606 28030 44658 28082
rect 51998 28030 52050 28082
rect 53342 28030 53394 28082
rect 53902 28030 53954 28082
rect 4398 27918 4450 27970
rect 9326 27918 9378 27970
rect 9886 27918 9938 27970
rect 13694 27918 13746 27970
rect 17502 27918 17554 27970
rect 21870 27918 21922 27970
rect 38894 27918 38946 27970
rect 39790 27918 39842 27970
rect 44494 27918 44546 27970
rect 46398 27918 46450 27970
rect 52222 27918 52274 27970
rect 1374 27806 1426 27858
rect 2382 27806 2434 27858
rect 3502 27806 3554 27858
rect 3950 27806 4002 27858
rect 5294 27806 5346 27858
rect 5854 27806 5906 27858
rect 7198 27806 7250 27858
rect 7982 27806 8034 27858
rect 9214 27806 9266 27858
rect 12798 27806 12850 27858
rect 13358 27806 13410 27858
rect 14030 27806 14082 27858
rect 14590 27806 14642 27858
rect 15710 27806 15762 27858
rect 16718 27806 16770 27858
rect 19070 27806 19122 27858
rect 19630 27806 19682 27858
rect 19742 27806 19794 27858
rect 20078 27806 20130 27858
rect 20638 27806 20690 27858
rect 23438 27806 23490 27858
rect 24222 27806 24274 27858
rect 24782 27806 24834 27858
rect 25566 27806 25618 27858
rect 25902 27806 25954 27858
rect 27022 27806 27074 27858
rect 27694 27806 27746 27858
rect 30158 27806 30210 27858
rect 30830 27806 30882 27858
rect 34638 27806 34690 27858
rect 35198 27806 35250 27858
rect 35758 27806 35810 27858
rect 36542 27806 36594 27858
rect 38558 27806 38610 27858
rect 39230 27806 39282 27858
rect 39678 27806 39730 27858
rect 40014 27806 40066 27858
rect 40126 27806 40178 27858
rect 40910 27806 40962 27858
rect 41806 27806 41858 27858
rect 44942 27806 44994 27858
rect 45054 27806 45106 27858
rect 45502 27806 45554 27858
rect 50318 27806 50370 27858
rect 52110 27806 52162 27858
rect 52558 27806 52610 27858
rect 52782 27806 52834 27858
rect 55582 27806 55634 27858
rect 2942 27694 2994 27746
rect 3390 27694 3442 27746
rect 4958 27694 5010 27746
rect 6414 27694 6466 27746
rect 8542 27694 8594 27746
rect 8878 27694 8930 27746
rect 10222 27694 10274 27746
rect 12126 27694 12178 27746
rect 12238 27694 12290 27746
rect 13022 27694 13074 27746
rect 14702 27694 14754 27746
rect 15150 27694 15202 27746
rect 21310 27694 21362 27746
rect 23886 27694 23938 27746
rect 24894 27694 24946 27746
rect 27918 27694 27970 27746
rect 31390 27694 31442 27746
rect 34190 27694 34242 27746
rect 35422 27694 35474 27746
rect 36990 27694 37042 27746
rect 38894 27694 38946 27746
rect 42142 27694 42194 27746
rect 45278 27694 45330 27746
rect 48078 27694 48130 27746
rect 53342 27694 53394 27746
rect 53454 27694 53506 27746
rect 55022 27694 55074 27746
rect 56366 27694 56418 27746
rect 5966 27582 6018 27634
rect 8766 27582 8818 27634
rect 11902 27582 11954 27634
rect 13246 27582 13298 27634
rect 17950 27582 18002 27634
rect 19854 27582 19906 27634
rect 20974 27582 21026 27634
rect 21198 27582 21250 27634
rect 22318 27582 22370 27634
rect 30382 27582 30434 27634
rect 35646 27582 35698 27634
rect 38782 27582 38834 27634
rect 40686 27582 40738 27634
rect 40798 27582 40850 27634
rect 41134 27582 41186 27634
rect 56030 27582 56082 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 44466 27414 44518 27466
rect 44570 27414 44622 27466
rect 44674 27414 44726 27466
rect 1710 27246 1762 27298
rect 2830 27246 2882 27298
rect 3502 27246 3554 27298
rect 7758 27246 7810 27298
rect 7870 27246 7922 27298
rect 10110 27246 10162 27298
rect 12014 27246 12066 27298
rect 13918 27246 13970 27298
rect 19182 27246 19234 27298
rect 20302 27246 20354 27298
rect 27582 27246 27634 27298
rect 31838 27246 31890 27298
rect 37550 27246 37602 27298
rect 38670 27246 38722 27298
rect 41694 27246 41746 27298
rect 45502 27246 45554 27298
rect 47294 27246 47346 27298
rect 53790 27246 53842 27298
rect 54910 27246 54962 27298
rect 55022 27246 55074 27298
rect 56142 27246 56194 27298
rect 3614 27134 3666 27186
rect 3950 27134 4002 27186
rect 4958 27134 5010 27186
rect 5406 27134 5458 27186
rect 7982 27134 8034 27186
rect 11902 27134 11954 27186
rect 12462 27134 12514 27186
rect 12910 27134 12962 27186
rect 14366 27134 14418 27186
rect 21758 27134 21810 27186
rect 22206 27134 22258 27186
rect 26574 27134 26626 27186
rect 31726 27134 31778 27186
rect 33742 27134 33794 27186
rect 35198 27134 35250 27186
rect 40910 27134 40962 27186
rect 41806 27134 41858 27186
rect 42254 27134 42306 27186
rect 43262 27134 43314 27186
rect 47406 27134 47458 27186
rect 49422 27134 49474 27186
rect 50878 27134 50930 27186
rect 52670 27134 52722 27186
rect 1150 27022 1202 27074
rect 4398 27022 4450 27074
rect 4734 27022 4786 27074
rect 6078 27022 6130 27074
rect 6974 27022 7026 27074
rect 8430 27022 8482 27074
rect 10670 27022 10722 27074
rect 12350 27022 12402 27074
rect 12686 27022 12738 27074
rect 13246 27022 13298 27074
rect 13694 27022 13746 27074
rect 15038 27022 15090 27074
rect 16046 27022 16098 27074
rect 18734 27022 18786 27074
rect 20750 27022 20802 27074
rect 21086 27022 21138 27074
rect 21534 27022 21586 27074
rect 22430 27022 22482 27074
rect 22766 27022 22818 27074
rect 23774 27022 23826 27074
rect 26910 27022 26962 27074
rect 27358 27010 27410 27062
rect 28030 27022 28082 27074
rect 28590 27022 28642 27074
rect 29598 27022 29650 27074
rect 34750 27022 34802 27074
rect 37102 27022 37154 27074
rect 39118 27022 39170 27074
rect 40238 27022 40290 27074
rect 40574 27022 40626 27074
rect 41134 27022 41186 27074
rect 41582 27022 41634 27074
rect 42814 27022 42866 27074
rect 45054 27022 45106 27074
rect 49870 27022 49922 27074
rect 50430 27022 50482 27074
rect 31278 26910 31330 26962
rect 31390 26910 31442 26962
rect 34078 26910 34130 26962
rect 39342 26910 39394 26962
rect 40462 26910 40514 26962
rect 48190 26910 48242 26962
rect 54238 26910 54290 26962
rect 55918 26910 55970 26962
rect 56142 26910 56194 26962
rect 3502 26798 3554 26850
rect 8990 26798 9042 26850
rect 32510 26798 32562 26850
rect 36430 26798 36482 26850
rect 39678 26798 39730 26850
rect 42142 26798 42194 26850
rect 44382 26798 44434 26850
rect 46622 26798 46674 26850
rect 47182 26798 47234 26850
rect 52110 26798 52162 26850
rect 54798 26798 54850 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 43806 26630 43858 26682
rect 43910 26630 43962 26682
rect 44014 26630 44066 26682
rect 2830 26462 2882 26514
rect 9214 26462 9266 26514
rect 9774 26462 9826 26514
rect 10334 26462 10386 26514
rect 35758 26462 35810 26514
rect 43150 26462 43202 26514
rect 49758 26462 49810 26514
rect 51998 26462 52050 26514
rect 55246 26462 55298 26514
rect 3278 26350 3330 26402
rect 6638 26350 6690 26402
rect 7646 26350 7698 26402
rect 17278 26350 17330 26402
rect 18398 26350 18450 26402
rect 21310 26350 21362 26402
rect 26238 26350 26290 26402
rect 28702 26350 28754 26402
rect 35646 26350 35698 26402
rect 37886 26350 37938 26402
rect 46622 26350 46674 26402
rect 48750 26350 48802 26402
rect 49198 26350 49250 26402
rect 49422 26350 49474 26402
rect 52558 26350 52610 26402
rect 1262 26238 1314 26290
rect 3950 26238 4002 26290
rect 4174 26238 4226 26290
rect 4398 26238 4450 26290
rect 9662 26238 9714 26290
rect 12798 26238 12850 26290
rect 13022 26238 13074 26290
rect 13246 26238 13298 26290
rect 13470 26238 13522 26290
rect 16830 26238 16882 26290
rect 17054 26238 17106 26290
rect 20974 26238 21026 26290
rect 21646 26238 21698 26290
rect 22206 26238 22258 26290
rect 23326 26238 23378 26290
rect 24334 26238 24386 26290
rect 26126 26238 26178 26290
rect 27806 26238 27858 26290
rect 29038 26238 29090 26290
rect 29598 26238 29650 26290
rect 30382 26238 30434 26290
rect 30942 26238 30994 26290
rect 31838 26238 31890 26290
rect 32398 26238 32450 26290
rect 34526 26238 34578 26290
rect 40126 26238 40178 26290
rect 40798 26238 40850 26290
rect 41470 26238 41522 26290
rect 42926 26238 42978 26290
rect 43262 26238 43314 26290
rect 45614 26238 45666 26290
rect 45950 26238 46002 26290
rect 50542 26238 50594 26290
rect 51214 26238 51266 26290
rect 52222 26238 52274 26290
rect 52446 26238 52498 26290
rect 52670 26238 52722 26290
rect 53566 26238 53618 26290
rect 56142 26238 56194 26290
rect 6302 26126 6354 26178
rect 8094 26126 8146 26178
rect 9774 26126 9826 26178
rect 10222 26126 10274 26178
rect 10334 26126 10386 26178
rect 17614 26126 17666 26178
rect 18846 26126 18898 26178
rect 20862 26126 20914 26178
rect 22766 26126 22818 26178
rect 25006 26126 25058 26178
rect 26574 26126 26626 26178
rect 29710 26126 29762 26178
rect 34974 26126 35026 26178
rect 36542 26126 36594 26178
rect 36654 26126 36706 26178
rect 36766 26126 36818 26178
rect 38334 26126 38386 26178
rect 40574 26126 40626 26178
rect 41246 26126 41298 26178
rect 41358 26126 41410 26178
rect 41918 26126 41970 26178
rect 42254 26126 42306 26178
rect 42478 26126 42530 26178
rect 43374 26126 43426 26178
rect 45278 26126 45330 26178
rect 45390 26126 45442 26178
rect 51326 26126 51378 26178
rect 54014 26126 54066 26178
rect 55918 26126 55970 26178
rect 1710 26014 1762 26066
rect 3390 26014 3442 26066
rect 3838 26014 3890 26066
rect 4062 26014 4114 26066
rect 5070 26014 5122 26066
rect 6190 26014 6242 26066
rect 13134 26014 13186 26066
rect 17502 26014 17554 26066
rect 17726 26014 17778 26066
rect 19966 26014 20018 26066
rect 20638 26014 20690 26066
rect 22318 26014 22370 26066
rect 24894 26014 24946 26066
rect 32958 26014 33010 26066
rect 34078 26014 34130 26066
rect 35086 26014 35138 26066
rect 35198 26014 35250 26066
rect 35310 26014 35362 26066
rect 36318 26014 36370 26066
rect 36430 26014 36482 26066
rect 39454 26014 39506 26066
rect 40462 26014 40514 26066
rect 42702 26014 42754 26066
rect 50206 26014 50258 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 44466 25846 44518 25898
rect 44570 25846 44622 25898
rect 44674 25846 44726 25898
rect 1822 25678 1874 25730
rect 2942 25678 2994 25730
rect 4398 25678 4450 25730
rect 10782 25678 10834 25730
rect 12238 25678 12290 25730
rect 24782 25678 24834 25730
rect 26574 25678 26626 25730
rect 27694 25678 27746 25730
rect 29262 25678 29314 25730
rect 30382 25678 30434 25730
rect 4062 25566 4114 25618
rect 5854 25566 5906 25618
rect 6974 25566 7026 25618
rect 7646 25566 7698 25618
rect 21646 25622 21698 25674
rect 36542 25678 36594 25730
rect 39678 25678 39730 25730
rect 40686 25678 40738 25730
rect 41918 25678 41970 25730
rect 42030 25678 42082 25730
rect 47294 25678 47346 25730
rect 48190 25678 48242 25730
rect 49310 25678 49362 25730
rect 52110 25678 52162 25730
rect 52670 25678 52722 25730
rect 7758 25566 7810 25618
rect 7870 25566 7922 25618
rect 9662 25566 9714 25618
rect 11230 25566 11282 25618
rect 17726 25566 17778 25618
rect 31614 25566 31666 25618
rect 31726 25566 31778 25618
rect 33630 25566 33682 25618
rect 34862 25566 34914 25618
rect 37550 25566 37602 25618
rect 40798 25566 40850 25618
rect 41022 25566 41074 25618
rect 42702 25566 42754 25618
rect 43150 25566 43202 25618
rect 44158 25566 44210 25618
rect 50990 25566 51042 25618
rect 53006 25566 53058 25618
rect 53902 25566 53954 25618
rect 56254 25566 56306 25618
rect 1262 25454 1314 25506
rect 4398 25454 4450 25506
rect 4734 25454 4786 25506
rect 7422 25454 7474 25506
rect 11678 25454 11730 25506
rect 12014 25454 12066 25506
rect 12910 25454 12962 25506
rect 13246 25454 13298 25506
rect 14366 25454 14418 25506
rect 17054 25454 17106 25506
rect 17614 25454 17666 25506
rect 18174 25454 18226 25506
rect 18734 25454 18786 25506
rect 19742 25454 19794 25506
rect 20638 25454 20690 25506
rect 20974 25454 21026 25506
rect 21422 25442 21474 25494
rect 22318 25454 22370 25506
rect 22654 25454 22706 25506
rect 23662 25454 23714 25506
rect 24558 25454 24610 25506
rect 25006 25454 25058 25506
rect 25230 25454 25282 25506
rect 26126 25454 26178 25506
rect 28814 25454 28866 25506
rect 33742 25454 33794 25506
rect 34414 25454 34466 25506
rect 36990 25454 37042 25506
rect 39118 25454 39170 25506
rect 40462 25454 40514 25506
rect 41134 25454 41186 25506
rect 41470 25454 41522 25506
rect 42142 25454 42194 25506
rect 43598 25454 43650 25506
rect 44046 25454 44098 25506
rect 44606 25454 44658 25506
rect 45390 25454 45442 25506
rect 46174 25454 46226 25506
rect 46734 25454 46786 25506
rect 50542 25454 50594 25506
rect 55918 25454 55970 25506
rect 5406 25342 5458 25394
rect 7534 25342 7586 25394
rect 9214 25342 9266 25394
rect 16718 25342 16770 25394
rect 24894 25342 24946 25394
rect 36430 25342 36482 25394
rect 41246 25342 41298 25394
rect 42702 25342 42754 25394
rect 49758 25342 49810 25394
rect 53566 25342 53618 25394
rect 31726 25230 31778 25282
rect 32622 25230 32674 25282
rect 32958 25230 33010 25282
rect 35982 25230 36034 25282
rect 38670 25230 38722 25282
rect 39342 25230 39394 25282
rect 42478 25230 42530 25282
rect 46958 25230 47010 25282
rect 55134 25230 55186 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 43806 25062 43858 25114
rect 43910 25062 43962 25114
rect 44014 25062 44066 25114
rect 5070 24894 5122 24946
rect 5518 24894 5570 24946
rect 25566 24894 25618 24946
rect 41246 24894 41298 24946
rect 44270 24894 44322 24946
rect 48974 24894 49026 24946
rect 52446 24894 52498 24946
rect 6414 24782 6466 24834
rect 6862 24782 6914 24834
rect 21086 24782 21138 24834
rect 23998 24782 24050 24834
rect 26238 24782 26290 24834
rect 34078 24782 34130 24834
rect 36542 24782 36594 24834
rect 39678 24782 39730 24834
rect 41918 24782 41970 24834
rect 47406 24782 47458 24834
rect 51102 24782 51154 24834
rect 1486 24670 1538 24722
rect 1934 24670 1986 24722
rect 2830 24670 2882 24722
rect 3278 24670 3330 24722
rect 4174 24670 4226 24722
rect 6302 24670 6354 24722
rect 7310 24670 7362 24722
rect 7646 24670 7698 24722
rect 8430 24670 8482 24722
rect 9102 24670 9154 24722
rect 9998 24670 10050 24722
rect 14030 24670 14082 24722
rect 17054 24670 17106 24722
rect 17390 24670 17442 24722
rect 18174 24670 18226 24722
rect 18846 24670 18898 24722
rect 19630 24670 19682 24722
rect 21310 24670 21362 24722
rect 21646 24670 21698 24722
rect 28814 24670 28866 24722
rect 29262 24670 29314 24722
rect 30718 24670 30770 24722
rect 31502 24670 31554 24722
rect 32734 24670 32786 24722
rect 32958 24670 33010 24722
rect 33294 24670 33346 24722
rect 39230 24670 39282 24722
rect 42030 24670 42082 24722
rect 45838 24670 45890 24722
rect 53902 24670 53954 24722
rect 56142 24670 56194 24722
rect 1150 24558 1202 24610
rect 2158 24558 2210 24610
rect 4958 24558 5010 24610
rect 5406 24558 5458 24610
rect 5518 24558 5570 24610
rect 6078 24558 6130 24610
rect 16606 24558 16658 24610
rect 20638 24558 20690 24610
rect 20862 24558 20914 24610
rect 24446 24558 24498 24610
rect 27806 24558 27858 24610
rect 28478 24558 28530 24610
rect 29934 24558 29986 24610
rect 34414 24558 34466 24610
rect 38894 24558 38946 24610
rect 39006 24558 39058 24610
rect 41694 24558 41746 24610
rect 47854 24558 47906 24610
rect 50654 24558 50706 24610
rect 52782 24558 52834 24610
rect 53230 24558 53282 24610
rect 54238 24558 54290 24610
rect 56366 24558 56418 24610
rect 6526 24446 6578 24498
rect 7870 24446 7922 24498
rect 14590 24446 14642 24498
rect 15710 24446 15762 24498
rect 17614 24446 17666 24498
rect 22206 24446 22258 24498
rect 23326 24446 23378 24498
rect 26686 24446 26738 24498
rect 29486 24446 29538 24498
rect 32846 24446 32898 24498
rect 35646 24446 35698 24498
rect 36990 24446 37042 24498
rect 38110 24446 38162 24498
rect 40126 24446 40178 24498
rect 45390 24446 45442 24498
rect 46510 24446 46562 24498
rect 46846 24446 46898 24498
rect 49534 24446 49586 24498
rect 52110 24446 52162 24498
rect 55470 24446 55522 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 44466 24278 44518 24330
rect 44570 24278 44622 24330
rect 44674 24278 44726 24330
rect 3726 24110 3778 24162
rect 6078 24110 6130 24162
rect 8990 24110 9042 24162
rect 12910 24110 12962 24162
rect 20862 24110 20914 24162
rect 21646 24110 21698 24162
rect 22766 24110 22818 24162
rect 30270 24110 30322 24162
rect 32510 24110 32562 24162
rect 33630 24110 33682 24162
rect 41470 24110 41522 24162
rect 52558 24110 52610 24162
rect 53678 24110 53730 24162
rect 55918 24110 55970 24162
rect 5070 23998 5122 24050
rect 9550 23998 9602 24050
rect 9886 23998 9938 24050
rect 11678 23998 11730 24050
rect 14702 23998 14754 24050
rect 16718 23998 16770 24050
rect 17726 23998 17778 24050
rect 20750 23998 20802 24050
rect 21422 23998 21474 24050
rect 21758 23998 21810 24050
rect 26574 23998 26626 24050
rect 34862 23998 34914 24050
rect 37438 23998 37490 24050
rect 43150 23998 43202 24050
rect 45278 23998 45330 24050
rect 48862 23998 48914 24050
rect 54238 23998 54290 24050
rect 54574 23998 54626 24050
rect 56254 23998 56306 24050
rect 1710 23886 1762 23938
rect 2606 23886 2658 23938
rect 3054 23886 3106 23938
rect 3838 23886 3890 23938
rect 4286 23886 4338 23938
rect 5406 23886 5458 23938
rect 5966 23886 6018 23938
rect 6750 23886 6802 23938
rect 7086 23886 7138 23938
rect 8094 23886 8146 23938
rect 9326 23886 9378 23938
rect 11342 23886 11394 23938
rect 14254 23886 14306 23938
rect 17054 23886 17106 23938
rect 17502 23886 17554 23938
rect 18174 23886 18226 23938
rect 18846 23886 18898 23938
rect 19742 23886 19794 23938
rect 21310 23886 21362 23938
rect 22206 23886 22258 23938
rect 23886 23886 23938 23938
rect 25902 23892 25954 23944
rect 26350 23886 26402 23938
rect 27022 23886 27074 23938
rect 27694 23886 27746 23938
rect 28702 23886 28754 23938
rect 29710 23886 29762 23938
rect 35086 23886 35138 23938
rect 35646 23886 35698 23938
rect 36766 23886 36818 23938
rect 37214 23886 37266 23938
rect 38110 23886 38162 23938
rect 38446 23886 38498 23938
rect 39566 23886 39618 23938
rect 44942 23886 44994 23938
rect 48078 23886 48130 23938
rect 53006 23886 53058 23938
rect 54014 23886 54066 23938
rect 4734 23774 4786 23826
rect 22318 23774 22370 23826
rect 25566 23774 25618 23826
rect 34078 23774 34130 23826
rect 36430 23774 36482 23826
rect 41918 23774 41970 23826
rect 42702 23774 42754 23826
rect 50990 23774 51042 23826
rect 15934 23662 15986 23714
rect 31390 23662 31442 23714
rect 35982 23662 36034 23714
rect 40350 23662 40402 23714
rect 44270 23662 44322 23714
rect 46510 23662 46562 23714
rect 51438 23662 51490 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 43806 23494 43858 23546
rect 43910 23494 43962 23546
rect 44014 23494 44066 23546
rect 2942 23326 2994 23378
rect 6750 23326 6802 23378
rect 19406 23326 19458 23378
rect 51214 23326 51266 23378
rect 54574 23326 54626 23378
rect 4062 23214 4114 23266
rect 14478 23214 14530 23266
rect 15374 23214 15426 23266
rect 21534 23214 21586 23266
rect 35646 23214 35698 23266
rect 36318 23214 36370 23266
rect 49646 23214 49698 23266
rect 52222 23214 52274 23266
rect 53790 23214 53842 23266
rect 55134 23214 55186 23266
rect 1262 23102 1314 23154
rect 5182 23102 5234 23154
rect 7870 23102 7922 23154
rect 8318 23102 8370 23154
rect 8990 23102 9042 23154
rect 9774 23102 9826 23154
rect 10670 23102 10722 23154
rect 16270 23102 16322 23154
rect 16606 23102 16658 23154
rect 17278 23102 17330 23154
rect 18062 23102 18114 23154
rect 18958 23102 19010 23154
rect 23102 23102 23154 23154
rect 23886 23102 23938 23154
rect 24446 23102 24498 23154
rect 25006 23102 25058 23154
rect 25678 23102 25730 23154
rect 26686 23102 26738 23154
rect 29038 23102 29090 23154
rect 30606 23102 30658 23154
rect 31166 23102 31218 23154
rect 32062 23102 32114 23154
rect 32622 23102 32674 23154
rect 33406 23102 33458 23154
rect 33854 23102 33906 23154
rect 35198 23102 35250 23154
rect 35758 23102 35810 23154
rect 36654 23102 36706 23154
rect 36990 23102 37042 23154
rect 37214 23102 37266 23154
rect 37662 23102 37714 23154
rect 38670 23102 38722 23154
rect 39006 23102 39058 23154
rect 39902 23102 39954 23154
rect 40238 23102 40290 23154
rect 41358 23102 41410 23154
rect 45726 23102 45778 23154
rect 46510 23102 46562 23154
rect 47070 23102 47122 23154
rect 47854 23102 47906 23154
rect 48302 23102 48354 23154
rect 54798 23102 54850 23154
rect 55022 23102 55074 23154
rect 55246 23102 55298 23154
rect 55918 23102 55970 23154
rect 5518 22990 5570 23042
rect 7534 22990 7586 23042
rect 8542 22990 8594 23042
rect 14142 22990 14194 23042
rect 15486 22990 15538 23042
rect 15822 22990 15874 23042
rect 21870 22990 21922 23042
rect 23550 22990 23602 23042
rect 29486 22990 29538 23042
rect 34302 22990 34354 23042
rect 35534 22990 35586 23042
rect 38222 22990 38274 23042
rect 48750 22990 48802 23042
rect 52670 22990 52722 23042
rect 56254 22990 56306 23042
rect 1822 22878 1874 22930
rect 3390 22878 3442 22930
rect 3726 22878 3778 22930
rect 4174 22878 4226 22930
rect 12910 22878 12962 22930
rect 15262 22878 15314 22930
rect 16830 22878 16882 22930
rect 19518 22878 19570 22930
rect 19630 22878 19682 22930
rect 24558 22878 24610 22930
rect 33294 22878 33346 22930
rect 36430 22878 36482 22930
rect 37102 22878 37154 22930
rect 39230 22878 39282 22930
rect 47742 22878 47794 22930
rect 50094 22878 50146 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 44466 22710 44518 22762
rect 44570 22710 44622 22762
rect 44674 22710 44726 22762
rect 10222 22542 10274 22594
rect 16046 22542 16098 22594
rect 17278 22542 17330 22594
rect 17390 22542 17442 22594
rect 18398 22542 18450 22594
rect 20974 22542 21026 22594
rect 27694 22542 27746 22594
rect 1374 22430 1426 22482
rect 3726 22430 3778 22482
rect 6974 22430 7026 22482
rect 11790 22430 11842 22482
rect 12798 22430 12850 22482
rect 13246 22430 13298 22482
rect 16158 22430 16210 22482
rect 16942 22430 16994 22482
rect 19966 22430 20018 22482
rect 26574 22430 26626 22482
rect 28142 22430 28194 22482
rect 29150 22430 29202 22482
rect 32846 22430 32898 22482
rect 33854 22430 33906 22482
rect 37102 22430 37154 22482
rect 40462 22430 40514 22482
rect 40798 22430 40850 22482
rect 41022 22430 41074 22482
rect 41470 22486 41522 22538
rect 47182 22542 47234 22594
rect 49310 22542 49362 22594
rect 51326 22542 51378 22594
rect 54126 22542 54178 22594
rect 56254 22542 56306 22594
rect 41582 22430 41634 22482
rect 43150 22430 43202 22482
rect 46062 22430 46114 22482
rect 46846 22430 46898 22482
rect 47518 22430 47570 22482
rect 48190 22430 48242 22482
rect 53006 22430 53058 22482
rect 1150 22318 1202 22370
rect 1934 22318 1986 22370
rect 3054 22318 3106 22370
rect 3614 22318 3666 22370
rect 4174 22318 4226 22370
rect 4958 22318 5010 22370
rect 5854 22318 5906 22370
rect 9774 22318 9826 22370
rect 11342 22318 11394 22370
rect 12126 22318 12178 22370
rect 12574 22318 12626 22370
rect 13806 22318 13858 22370
rect 14814 22318 14866 22370
rect 15822 22318 15874 22370
rect 17166 22318 17218 22370
rect 19518 22318 19570 22370
rect 20302 22318 20354 22370
rect 20750 22318 20802 22370
rect 21422 22318 21474 22370
rect 21982 22318 22034 22370
rect 22990 22318 23042 22370
rect 26126 22318 26178 22370
rect 28590 22318 28642 22370
rect 28926 22318 28978 22370
rect 29822 22318 29874 22370
rect 30382 22318 30434 22370
rect 31166 22318 31218 22370
rect 33182 22318 33234 22370
rect 33630 22318 33682 22370
rect 34526 22318 34578 22370
rect 34862 22318 34914 22370
rect 35982 22318 36034 22370
rect 36542 22318 36594 22370
rect 42590 22318 42642 22370
rect 42926 22318 42978 22370
rect 43822 22318 43874 22370
rect 44158 22318 44210 22370
rect 45166 22318 45218 22370
rect 45950 22318 46002 22370
rect 46622 22318 46674 22370
rect 50766 22318 50818 22370
rect 53118 22318 53170 22370
rect 53566 22318 53618 22370
rect 56030 22318 56082 22370
rect 2718 22206 2770 22258
rect 6526 22206 6578 22258
rect 17950 22206 18002 22258
rect 40910 22206 40962 22258
rect 42142 22206 42194 22258
rect 49758 22206 49810 22258
rect 53678 22206 53730 22258
rect 2270 22094 2322 22146
rect 8094 22094 8146 22146
rect 38222 22094 38274 22146
rect 40350 22094 40402 22146
rect 41582 22094 41634 22146
rect 46062 22094 46114 22146
rect 52446 22094 52498 22146
rect 53006 22094 53058 22146
rect 55246 22094 55298 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 43806 21926 43858 21978
rect 43910 21926 43962 21978
rect 44014 21926 44066 21978
rect 12126 21758 12178 21810
rect 19966 21758 20018 21810
rect 22430 21758 22482 21810
rect 27022 21758 27074 21810
rect 32510 21758 32562 21810
rect 34638 21758 34690 21810
rect 40574 21758 40626 21810
rect 42926 21758 42978 21810
rect 47070 21758 47122 21810
rect 2718 21646 2770 21698
rect 4286 21646 4338 21698
rect 10558 21646 10610 21698
rect 28478 21646 28530 21698
rect 32398 21646 32450 21698
rect 41358 21646 41410 21698
rect 55694 21646 55746 21698
rect 7198 21534 7250 21586
rect 7534 21534 7586 21586
rect 8206 21534 8258 21586
rect 8430 21534 8482 21586
rect 8766 21534 8818 21586
rect 9774 21534 9826 21586
rect 13134 21534 13186 21586
rect 13694 21534 13746 21586
rect 14814 21534 14866 21586
rect 15822 21534 15874 21586
rect 16830 21534 16882 21586
rect 17278 21534 17330 21586
rect 18398 21534 18450 21586
rect 20750 21534 20802 21586
rect 23102 21534 23154 21586
rect 24782 21534 24834 21586
rect 25454 21534 25506 21586
rect 28814 21534 28866 21586
rect 29262 21534 29314 21586
rect 29934 21534 29986 21586
rect 30718 21534 30770 21586
rect 31614 21534 31666 21586
rect 32958 21534 33010 21586
rect 36430 21534 36482 21586
rect 37326 21534 37378 21586
rect 38110 21534 38162 21586
rect 38670 21534 38722 21586
rect 39230 21534 39282 21586
rect 39566 21534 39618 21586
rect 40014 21534 40066 21586
rect 40574 21534 40626 21586
rect 45390 21534 45442 21586
rect 49198 21534 49250 21586
rect 49982 21534 50034 21586
rect 51214 21534 51266 21586
rect 51550 21534 51602 21586
rect 53006 21534 53058 21586
rect 53454 21534 53506 21586
rect 55470 21534 55522 21586
rect 55918 21534 55970 21586
rect 1374 21422 1426 21474
rect 1710 21422 1762 21474
rect 6750 21422 6802 21474
rect 7758 21422 7810 21474
rect 10894 21422 10946 21474
rect 12798 21422 12850 21474
rect 13806 21422 13858 21474
rect 14254 21422 14306 21474
rect 16494 21422 16546 21474
rect 21198 21422 21250 21474
rect 23550 21422 23602 21474
rect 33518 21422 33570 21474
rect 40238 21422 40290 21474
rect 48750 21422 48802 21474
rect 50766 21422 50818 21474
rect 51326 21422 51378 21474
rect 53790 21422 53842 21474
rect 1038 21310 1090 21362
rect 2046 21310 2098 21362
rect 3166 21310 3218 21362
rect 4958 21310 5010 21362
rect 5294 21310 5346 21362
rect 17614 21310 17666 21362
rect 18846 21310 18898 21362
rect 25902 21310 25954 21362
rect 29486 21310 29538 21362
rect 38558 21310 38610 21362
rect 40798 21310 40850 21362
rect 41806 21310 41858 21362
rect 45950 21310 46002 21362
rect 47630 21310 47682 21362
rect 49758 21310 49810 21362
rect 50430 21310 50482 21362
rect 52334 21310 52386 21362
rect 52446 21310 52498 21362
rect 52558 21310 52610 21362
rect 55022 21310 55074 21362
rect 56030 21310 56082 21362
rect 56142 21310 56194 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 44466 21142 44518 21194
rect 44570 21142 44622 21194
rect 44674 21142 44726 21194
rect 1710 20974 1762 21026
rect 2830 20974 2882 21026
rect 4286 20974 4338 21026
rect 13806 20974 13858 21026
rect 20526 20974 20578 21026
rect 21646 20974 21698 21026
rect 22766 20974 22818 21026
rect 29934 20974 29986 21026
rect 33406 20974 33458 21026
rect 36654 20974 36706 21026
rect 37774 20974 37826 21026
rect 41246 20974 41298 21026
rect 41358 20974 41410 21026
rect 41470 20974 41522 21026
rect 44158 20974 44210 21026
rect 47182 20974 47234 21026
rect 47518 20974 47570 21026
rect 49198 20974 49250 21026
rect 50206 20974 50258 21026
rect 54126 20974 54178 21026
rect 55246 20974 55298 21026
rect 56030 20974 56082 21026
rect 56366 20974 56418 21026
rect 3278 20862 3330 20914
rect 4734 20862 4786 20914
rect 9438 20862 9490 20914
rect 10670 20862 10722 20914
rect 11342 20862 11394 20914
rect 11566 20862 11618 20914
rect 12686 20862 12738 20914
rect 14814 20862 14866 20914
rect 16046 20862 16098 20914
rect 17166 20862 17218 20914
rect 18174 20862 18226 20914
rect 25566 20862 25618 20914
rect 28702 20862 28754 20914
rect 30606 20862 30658 20914
rect 39118 20862 39170 20914
rect 39230 20862 39282 20914
rect 40350 20862 40402 20914
rect 40686 20862 40738 20914
rect 43038 20862 43090 20914
rect 46510 20862 46562 20914
rect 46846 20862 46898 20914
rect 52334 20862 52386 20914
rect 52782 20862 52834 20914
rect 1262 20750 1314 20802
rect 3614 20750 3666 20802
rect 4174 20750 4226 20802
rect 5518 20750 5570 20802
rect 6302 20750 6354 20802
rect 11118 20750 11170 20802
rect 12126 20750 12178 20802
rect 17838 20750 17890 20802
rect 19966 20750 20018 20802
rect 23886 20750 23938 20802
rect 24894 20750 24946 20802
rect 25342 20750 25394 20802
rect 26126 20750 26178 20802
rect 26574 20750 26626 20802
rect 27582 20750 27634 20802
rect 30494 20750 30546 20802
rect 31278 20750 31330 20802
rect 32398 20750 32450 20802
rect 32734 20750 32786 20802
rect 33294 20750 33346 20802
rect 33854 20750 33906 20802
rect 34414 20750 34466 20802
rect 35422 20750 35474 20802
rect 38894 20750 38946 20802
rect 39678 20750 39730 20802
rect 40574 20750 40626 20802
rect 40798 20750 40850 20802
rect 41582 20750 41634 20802
rect 42366 20750 42418 20802
rect 42814 20750 42866 20802
rect 43598 20750 43650 20802
rect 48862 20750 48914 20802
rect 52558 20750 52610 20802
rect 53678 20750 53730 20802
rect 9102 20638 9154 20690
rect 11230 20638 11282 20690
rect 14478 20638 14530 20690
rect 17278 20638 17330 20690
rect 22318 20638 22370 20690
rect 24558 20638 24610 20690
rect 28366 20638 28418 20690
rect 36206 20638 36258 20690
rect 39230 20638 39282 20690
rect 42590 20638 42642 20690
rect 48638 20638 48690 20690
rect 49758 20638 49810 20690
rect 52894 20638 52946 20690
rect 19406 20526 19458 20578
rect 31614 20526 31666 20578
rect 41918 20526 41970 20578
rect 42142 20526 42194 20578
rect 45278 20526 45330 20578
rect 51326 20526 51378 20578
rect 51886 20526 51938 20578
rect 51998 20526 52050 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 43806 20358 43858 20410
rect 43910 20358 43962 20410
rect 44014 20358 44066 20410
rect 32622 20190 32674 20242
rect 33182 20190 33234 20242
rect 38670 20190 38722 20242
rect 51326 20190 51378 20242
rect 52894 20190 52946 20242
rect 2718 20078 2770 20130
rect 4958 20078 5010 20130
rect 11566 20078 11618 20130
rect 18510 20078 18562 20130
rect 21086 20078 21138 20130
rect 22654 20078 22706 20130
rect 34750 20078 34802 20130
rect 41470 20078 41522 20130
rect 53230 20078 53282 20130
rect 3614 19966 3666 20018
rect 5406 19966 5458 20018
rect 5742 19966 5794 20018
rect 6526 19966 6578 20018
rect 7198 19966 7250 20018
rect 7982 19966 8034 20018
rect 8766 19966 8818 20018
rect 13134 19966 13186 20018
rect 14814 19966 14866 20018
rect 15374 19966 15426 20018
rect 16494 19966 16546 20018
rect 16830 19966 16882 20018
rect 17614 19966 17666 20018
rect 18062 19966 18114 20018
rect 23438 19966 23490 20018
rect 23998 19966 24050 20018
rect 24782 19966 24834 20018
rect 25342 19966 25394 20018
rect 26238 19966 26290 20018
rect 28702 19966 28754 20018
rect 31054 19966 31106 20018
rect 37102 19966 37154 20018
rect 39342 19966 39394 20018
rect 41358 19966 41410 20018
rect 42702 19966 42754 20018
rect 45390 19966 45442 20018
rect 45838 19966 45890 20018
rect 46734 19966 46786 20018
rect 47070 19966 47122 20018
rect 48078 19966 48130 20018
rect 48750 19966 48802 20018
rect 49758 19966 49810 20018
rect 53902 19966 53954 20018
rect 2382 19854 2434 19906
rect 3278 19854 3330 19906
rect 3950 19854 4002 19906
rect 9214 19854 9266 19906
rect 10782 19854 10834 19906
rect 11118 19854 11170 19906
rect 11342 19854 11394 19906
rect 11790 19854 11842 19906
rect 12126 19854 12178 19906
rect 13582 19854 13634 19906
rect 17502 19854 17554 19906
rect 21422 19854 21474 19906
rect 23102 19854 23154 19906
rect 29150 19854 29202 19906
rect 30270 19854 30322 19906
rect 37550 19854 37602 19906
rect 42142 19854 42194 19906
rect 42366 19854 42418 19906
rect 45054 19854 45106 19906
rect 48974 19854 49026 19906
rect 50094 19854 50146 19906
rect 52110 19854 52162 19906
rect 52670 19854 52722 19906
rect 56254 19854 56306 19906
rect 1150 19742 1202 19794
rect 4286 19742 4338 19794
rect 5966 19742 6018 19794
rect 10334 19742 10386 19794
rect 11006 19742 11058 19794
rect 12014 19742 12066 19794
rect 24110 19742 24162 19794
rect 31502 19742 31554 19794
rect 34302 19742 34354 19794
rect 39790 19742 39842 19794
rect 40910 19742 40962 19794
rect 43038 19742 43090 19794
rect 46062 19742 46114 19794
rect 54350 19742 54402 19794
rect 55470 19742 55522 19794
rect 55918 19742 55970 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 44466 19574 44518 19626
rect 44570 19574 44622 19626
rect 44674 19574 44726 19626
rect 9214 19406 9266 19458
rect 9326 19406 9378 19458
rect 13358 19406 13410 19458
rect 14926 19406 14978 19458
rect 16046 19406 16098 19458
rect 20302 19406 20354 19458
rect 25342 19406 25394 19458
rect 27918 19406 27970 19458
rect 33070 19406 33122 19458
rect 37550 19406 37602 19458
rect 39566 19406 39618 19458
rect 42142 19406 42194 19458
rect 42814 19406 42866 19458
rect 48414 19406 48466 19458
rect 49198 19406 49250 19458
rect 52446 19406 52498 19458
rect 54126 19406 54178 19458
rect 55022 19406 55074 19458
rect 56030 19406 56082 19458
rect 56366 19406 56418 19458
rect 1486 19294 1538 19346
rect 2494 19294 2546 19346
rect 5070 19294 5122 19346
rect 6078 19294 6130 19346
rect 9774 19294 9826 19346
rect 10782 19294 10834 19346
rect 13470 19294 13522 19346
rect 18062 19294 18114 19346
rect 20750 19294 20802 19346
rect 26910 19294 26962 19346
rect 30718 19294 30770 19346
rect 30830 19294 30882 19346
rect 31054 19294 31106 19346
rect 35198 19294 35250 19346
rect 41022 19294 41074 19346
rect 44270 19294 44322 19346
rect 45278 19294 45330 19346
rect 48078 19294 48130 19346
rect 50206 19294 50258 19346
rect 53566 19294 53618 19346
rect 54238 19294 54290 19346
rect 55246 19294 55298 19346
rect 1934 19182 1986 19234
rect 2382 19182 2434 19234
rect 3166 19182 3218 19234
rect 3614 19182 3666 19234
rect 4622 19182 4674 19234
rect 5406 19182 5458 19234
rect 5854 19182 5906 19234
rect 6526 19182 6578 19234
rect 7086 19182 7138 19234
rect 8206 19182 8258 19234
rect 8878 19182 8930 19234
rect 9438 19182 9490 19234
rect 10222 19182 10274 19234
rect 10558 19170 10610 19222
rect 11230 19182 11282 19234
rect 11790 19182 11842 19234
rect 12014 19182 12066 19234
rect 12798 19182 12850 19234
rect 14478 19182 14530 19234
rect 16830 19182 16882 19234
rect 18398 19182 18450 19234
rect 19742 19182 19794 19234
rect 20078 19182 20130 19234
rect 21310 19182 21362 19234
rect 21534 19182 21586 19234
rect 22318 19182 22370 19234
rect 26462 19182 26514 19234
rect 27246 19182 27298 19234
rect 27694 19182 27746 19234
rect 28366 19182 28418 19234
rect 28926 19182 28978 19234
rect 29934 19182 29986 19234
rect 31166 19182 31218 19234
rect 31614 19182 31666 19234
rect 31838 19182 31890 19234
rect 36990 19182 37042 19234
rect 42590 19182 42642 19234
rect 43038 19182 43090 19234
rect 43262 19182 43314 19234
rect 44606 19182 44658 19234
rect 45166 19182 45218 19234
rect 45838 19182 45890 19234
rect 46398 19182 46450 19234
rect 47406 19182 47458 19234
rect 48974 19182 49026 19234
rect 51886 19182 51938 19234
rect 54014 19182 54066 19234
rect 54462 19182 54514 19234
rect 54686 19182 54738 19234
rect 55358 19182 55410 19234
rect 19294 19070 19346 19122
rect 24894 19070 24946 19122
rect 31726 19070 31778 19122
rect 32622 19070 32674 19122
rect 34862 19070 34914 19122
rect 40574 19070 40626 19122
rect 42926 19070 42978 19122
rect 49758 19070 49810 19122
rect 34190 18958 34242 19010
rect 36430 18958 36482 19010
rect 38670 18958 38722 19010
rect 39342 18958 39394 19010
rect 39678 18958 39730 19010
rect 51326 18958 51378 19010
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 43806 18790 43858 18842
rect 43910 18790 43962 18842
rect 44014 18790 44066 18842
rect 24670 18622 24722 18674
rect 27806 18622 27858 18674
rect 40574 18622 40626 18674
rect 43262 18622 43314 18674
rect 44270 18622 44322 18674
rect 53006 18622 53058 18674
rect 20862 18510 20914 18562
rect 23102 18510 23154 18562
rect 28702 18510 28754 18562
rect 34302 18510 34354 18562
rect 41022 18510 41074 18562
rect 45838 18510 45890 18562
rect 49086 18510 49138 18562
rect 51214 18510 51266 18562
rect 52110 18510 52162 18562
rect 2046 18398 2098 18450
rect 2718 18398 2770 18450
rect 4286 18398 4338 18450
rect 5406 18398 5458 18450
rect 5854 18398 5906 18450
rect 6526 18398 6578 18450
rect 7310 18398 7362 18450
rect 8206 18398 8258 18450
rect 9326 18398 9378 18450
rect 9886 18398 9938 18450
rect 10670 18398 10722 18450
rect 11006 18398 11058 18450
rect 12126 18398 12178 18450
rect 13022 18398 13074 18450
rect 14590 18398 14642 18450
rect 15038 18398 15090 18450
rect 15486 18398 15538 18450
rect 15822 18398 15874 18450
rect 16718 18398 16770 18450
rect 17166 18398 17218 18450
rect 18062 18398 18114 18450
rect 22430 18398 22482 18450
rect 26238 18398 26290 18450
rect 30270 18398 30322 18450
rect 30830 18398 30882 18450
rect 31726 18398 31778 18450
rect 32510 18398 32562 18450
rect 33070 18398 33122 18450
rect 33518 18398 33570 18450
rect 33966 18398 34018 18450
rect 34414 18398 34466 18450
rect 34638 18398 34690 18450
rect 35086 18398 35138 18450
rect 36654 18398 36706 18450
rect 37102 18398 37154 18450
rect 37998 18398 38050 18450
rect 38558 18398 38610 18450
rect 39342 18398 39394 18450
rect 40574 18398 40626 18450
rect 40910 18398 40962 18450
rect 41582 18398 41634 18450
rect 45950 18398 46002 18450
rect 46958 18398 47010 18450
rect 49646 18398 49698 18450
rect 50318 18398 50370 18450
rect 51326 18398 51378 18450
rect 51998 18398 52050 18450
rect 52894 18398 52946 18450
rect 54126 18398 54178 18450
rect 56254 18398 56306 18450
rect 1038 18286 1090 18338
rect 3166 18286 3218 18338
rect 5070 18286 5122 18338
rect 6078 18286 6130 18338
rect 8990 18286 9042 18338
rect 9998 18286 10050 18338
rect 13358 18286 13410 18338
rect 16046 18286 16098 18338
rect 26686 18286 26738 18338
rect 29038 18286 29090 18338
rect 34862 18286 34914 18338
rect 35422 18286 35474 18338
rect 35534 18286 35586 18338
rect 36318 18286 36370 18338
rect 37326 18286 37378 18338
rect 41134 18286 41186 18338
rect 46734 18286 46786 18338
rect 48750 18286 48802 18338
rect 49982 18286 50034 18338
rect 50878 18286 50930 18338
rect 52334 18286 52386 18338
rect 52558 18286 52610 18338
rect 56366 18286 56418 18338
rect 1374 18174 1426 18226
rect 1710 18174 1762 18226
rect 21310 18174 21362 18226
rect 23550 18174 23602 18226
rect 32958 18174 33010 18226
rect 42142 18174 42194 18226
rect 45390 18174 45442 18226
rect 47518 18174 47570 18226
rect 49758 18174 49810 18226
rect 49870 18174 49922 18226
rect 51102 18174 51154 18226
rect 53342 18174 53394 18226
rect 53678 18174 53730 18226
rect 54686 18174 54738 18226
rect 55806 18174 55858 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 44466 18006 44518 18058
rect 44570 18006 44622 18058
rect 44674 18006 44726 18058
rect 3390 17838 3442 17890
rect 5742 17838 5794 17890
rect 11230 17838 11282 17890
rect 11454 17838 11506 17890
rect 12686 17838 12738 17890
rect 14926 17838 14978 17890
rect 20190 17838 20242 17890
rect 31726 17838 31778 17890
rect 33070 17838 33122 17890
rect 34974 17838 35026 17890
rect 35086 17838 35138 17890
rect 37326 17838 37378 17890
rect 43710 17838 43762 17890
rect 43934 17838 43986 17890
rect 46622 17838 46674 17890
rect 47182 17838 47234 17890
rect 51998 17838 52050 17890
rect 53678 17838 53730 17890
rect 56366 17838 56418 17890
rect 6190 17726 6242 17778
rect 9550 17726 9602 17778
rect 16942 17726 16994 17778
rect 17054 17726 17106 17778
rect 17166 17726 17218 17778
rect 25902 17726 25954 17778
rect 29038 17726 29090 17778
rect 36318 17726 36370 17778
rect 41246 17726 41298 17778
rect 45502 17726 45554 17778
rect 47070 17726 47122 17778
rect 54910 17726 54962 17778
rect 1374 17614 1426 17666
rect 2158 17614 2210 17666
rect 2942 17614 2994 17666
rect 3614 17614 3666 17666
rect 3950 17614 4002 17666
rect 5070 17614 5122 17666
rect 5518 17614 5570 17666
rect 6974 17614 7026 17666
rect 7870 17614 7922 17666
rect 9102 17614 9154 17666
rect 11118 17614 11170 17666
rect 12238 17614 12290 17666
rect 14478 17614 14530 17666
rect 16046 17614 16098 17666
rect 16718 17614 16770 17666
rect 18062 17614 18114 17666
rect 18958 17614 19010 17666
rect 19518 17614 19570 17666
rect 20414 17614 20466 17666
rect 20750 17614 20802 17666
rect 26238 17614 26290 17666
rect 28366 17614 28418 17666
rect 28926 17614 28978 17666
rect 29710 17614 29762 17666
rect 30158 17614 30210 17666
rect 31054 17614 31106 17666
rect 31614 17614 31666 17666
rect 34526 17614 34578 17666
rect 35198 17614 35250 17666
rect 36654 17614 36706 17666
rect 37102 17614 37154 17666
rect 37998 17614 38050 17666
rect 38558 17614 38610 17666
rect 39342 17614 39394 17666
rect 40574 17614 40626 17666
rect 41022 17614 41074 17666
rect 41918 17614 41970 17666
rect 42254 17614 42306 17666
rect 43262 17614 43314 17666
rect 44046 17614 44098 17666
rect 45054 17614 45106 17666
rect 47406 17614 47458 17666
rect 48190 17614 48242 17666
rect 54238 17614 54290 17666
rect 55022 17614 55074 17666
rect 55358 17614 55410 17666
rect 56142 17614 56194 17666
rect 4398 17502 4450 17554
rect 4734 17502 4786 17554
rect 16942 17502 16994 17554
rect 21198 17502 21250 17554
rect 28030 17502 28082 17554
rect 32622 17502 32674 17554
rect 40238 17502 40290 17554
rect 48862 17502 48914 17554
rect 50990 17502 51042 17554
rect 51550 17502 51602 17554
rect 53566 17502 53618 17554
rect 54014 17502 54066 17554
rect 10670 17390 10722 17442
rect 13806 17390 13858 17442
rect 24670 17390 24722 17442
rect 31726 17390 31778 17442
rect 34190 17390 34242 17442
rect 53118 17390 53170 17442
rect 54350 17390 54402 17442
rect 54798 17390 54850 17442
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 43806 17222 43858 17274
rect 43910 17222 43962 17274
rect 44014 17222 44066 17274
rect 3390 17054 3442 17106
rect 8542 17054 8594 17106
rect 14926 17054 14978 17106
rect 15486 17054 15538 17106
rect 17726 17054 17778 17106
rect 19966 17054 20018 17106
rect 30270 17054 30322 17106
rect 38110 17054 38162 17106
rect 40350 17054 40402 17106
rect 42590 17054 42642 17106
rect 50318 17054 50370 17106
rect 51326 17054 51378 17106
rect 53566 17054 53618 17106
rect 1822 16942 1874 16994
rect 5406 16942 5458 16994
rect 6974 16942 7026 16994
rect 8990 16942 9042 16994
rect 13358 16942 13410 16994
rect 16158 16942 16210 16994
rect 18398 16942 18450 16994
rect 21758 16942 21810 16994
rect 23774 16942 23826 16994
rect 28702 16942 28754 16994
rect 32846 16942 32898 16994
rect 43486 16942 43538 16994
rect 48190 16942 48242 16994
rect 52334 16942 52386 16994
rect 55134 16942 55186 16994
rect 3726 16830 3778 16882
rect 4286 16830 4338 16882
rect 5966 16830 6018 16882
rect 9326 16830 9378 16882
rect 9774 16830 9826 16882
rect 10558 16830 10610 16882
rect 11230 16830 11282 16882
rect 12014 16830 12066 16882
rect 15374 16830 15426 16882
rect 23326 16830 23378 16882
rect 24110 16830 24162 16882
rect 24558 16830 24610 16882
rect 25230 16830 25282 16882
rect 25790 16830 25842 16882
rect 26798 16830 26850 16882
rect 32958 16830 33010 16882
rect 33294 16830 33346 16882
rect 33854 16830 33906 16882
rect 36542 16830 36594 16882
rect 38782 16830 38834 16882
rect 40910 16830 40962 16882
rect 42926 16830 42978 16882
rect 43374 16830 43426 16882
rect 45950 16830 46002 16882
rect 46286 16830 46338 16882
rect 46958 16830 47010 16882
rect 47630 16830 47682 16882
rect 50206 16830 50258 16882
rect 50766 16830 50818 16882
rect 50990 16830 51042 16882
rect 52446 16830 52498 16882
rect 55694 16830 55746 16882
rect 2270 16718 2322 16770
rect 5630 16718 5682 16770
rect 9998 16718 10050 16770
rect 13806 16718 13858 16770
rect 16494 16718 16546 16770
rect 18846 16718 18898 16770
rect 22206 16718 22258 16770
rect 24782 16718 24834 16770
rect 32510 16718 32562 16770
rect 32734 16718 32786 16770
rect 36990 16718 37042 16770
rect 43598 16718 43650 16770
rect 45390 16718 45442 16770
rect 47294 16718 47346 16770
rect 48638 16718 48690 16770
rect 49758 16718 49810 16770
rect 52782 16718 52834 16770
rect 52894 16718 52946 16770
rect 53118 16718 53170 16770
rect 54686 16718 54738 16770
rect 4174 16606 4226 16658
rect 4398 16606 4450 16658
rect 7422 16606 7474 16658
rect 15486 16606 15538 16658
rect 29150 16606 29202 16658
rect 34302 16606 34354 16658
rect 35422 16606 35474 16658
rect 39230 16606 39282 16658
rect 41470 16606 41522 16658
rect 44270 16606 44322 16658
rect 46622 16606 46674 16658
rect 46846 16606 46898 16658
rect 47406 16606 47458 16658
rect 50318 16606 50370 16658
rect 56030 16606 56082 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 44466 16438 44518 16490
rect 44570 16438 44622 16490
rect 44674 16438 44726 16490
rect 2830 16270 2882 16322
rect 4286 16270 4338 16322
rect 6862 16270 6914 16322
rect 7086 16270 7138 16322
rect 7422 16270 7474 16322
rect 7758 16270 7810 16322
rect 8990 16270 9042 16322
rect 10334 16270 10386 16322
rect 13022 16270 13074 16322
rect 13582 16270 13634 16322
rect 21198 16270 21250 16322
rect 28366 16270 28418 16322
rect 30606 16270 30658 16322
rect 35534 16270 35586 16322
rect 36654 16270 36706 16322
rect 38334 16270 38386 16322
rect 40574 16270 40626 16322
rect 42702 16270 42754 16322
rect 46398 16270 46450 16322
rect 48862 16270 48914 16322
rect 49198 16270 49250 16322
rect 49310 16270 49362 16322
rect 49646 16270 49698 16322
rect 53454 16270 53506 16322
rect 54798 16270 54850 16322
rect 56030 16270 56082 16322
rect 56366 16270 56418 16322
rect 1598 16158 1650 16210
rect 8094 16158 8146 16210
rect 8878 16158 8930 16210
rect 10782 16158 10834 16210
rect 14814 16158 14866 16210
rect 16046 16158 16098 16210
rect 18510 16158 18562 16210
rect 20190 16158 20242 16210
rect 27246 16158 27298 16210
rect 32958 16158 33010 16210
rect 41470 16158 41522 16210
rect 44382 16158 44434 16210
rect 45390 16158 45442 16210
rect 45502 16158 45554 16210
rect 47182 16158 47234 16210
rect 47406 16158 47458 16210
rect 49422 16158 49474 16210
rect 51550 16158 51602 16210
rect 1262 16046 1314 16098
rect 3614 16046 3666 16098
rect 4062 16046 4114 16098
rect 4958 16046 5010 16098
rect 5518 16046 5570 16098
rect 6302 16046 6354 16098
rect 9662 16046 9714 16098
rect 10110 16046 10162 16098
rect 11342 16046 11394 16098
rect 12462 16046 12514 16098
rect 13358 16046 13410 16098
rect 14030 16046 14082 16098
rect 14366 16046 14418 16098
rect 19742 16046 19794 16098
rect 20526 16046 20578 16098
rect 20974 16046 21026 16098
rect 21870 16046 21922 16098
rect 22430 16046 22482 16098
rect 23214 16046 23266 16098
rect 26686 16046 26738 16098
rect 30046 16046 30098 16098
rect 32622 16046 32674 16098
rect 34974 16046 35026 16098
rect 38894 16046 38946 16098
rect 41022 16046 41074 16098
rect 44830 16046 44882 16098
rect 45614 16046 45666 16098
rect 46062 16046 46114 16098
rect 46174 16046 46226 16098
rect 46622 16046 46674 16098
rect 46734 16046 46786 16098
rect 48190 16046 48242 16098
rect 48638 16046 48690 16098
rect 51438 16046 51490 16098
rect 51998 16046 52050 16098
rect 52334 16046 52386 16098
rect 54574 16046 54626 16098
rect 54686 16046 54738 16098
rect 54910 16046 54962 16098
rect 55246 16046 55298 16098
rect 3278 15934 3330 15986
rect 9326 15934 9378 15986
rect 12910 15934 12962 15986
rect 13470 15934 13522 15986
rect 18174 15934 18226 15986
rect 37214 15934 37266 15986
rect 40462 15934 40514 15986
rect 48750 15934 48802 15986
rect 50094 15934 50146 15986
rect 50206 15934 50258 15986
rect 50542 15934 50594 15986
rect 53902 15934 53954 15986
rect 31726 15822 31778 15874
rect 34190 15822 34242 15874
rect 43262 15822 43314 15874
rect 47518 15822 47570 15874
rect 50766 15822 50818 15874
rect 50878 15822 50930 15874
rect 51886 15822 51938 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 43806 15654 43858 15706
rect 43910 15654 43962 15706
rect 44014 15654 44066 15706
rect 1150 15486 1202 15538
rect 22430 15486 22482 15538
rect 43486 15486 43538 15538
rect 46286 15486 46338 15538
rect 48302 15486 48354 15538
rect 52110 15486 52162 15538
rect 56142 15486 56194 15538
rect 2718 15374 2770 15426
rect 3726 15374 3778 15426
rect 5742 15374 5794 15426
rect 10558 15374 10610 15426
rect 31950 15374 32002 15426
rect 37550 15374 37602 15426
rect 42814 15374 42866 15426
rect 53678 15374 53730 15426
rect 54574 15374 54626 15426
rect 3278 15262 3330 15314
rect 3502 15262 3554 15314
rect 4174 15262 4226 15314
rect 4958 15262 5010 15314
rect 6078 15262 6130 15314
rect 6638 15262 6690 15314
rect 7982 15262 8034 15314
rect 8878 15262 8930 15314
rect 13134 15262 13186 15314
rect 13582 15262 13634 15314
rect 14366 15262 14418 15314
rect 14814 15262 14866 15314
rect 15822 15262 15874 15314
rect 17166 15262 17218 15314
rect 17726 15262 17778 15314
rect 18510 15262 18562 15314
rect 18846 15262 18898 15314
rect 19854 15262 19906 15314
rect 20750 15262 20802 15314
rect 24446 15262 24498 15314
rect 32286 15262 32338 15314
rect 32734 15262 32786 15314
rect 33630 15262 33682 15314
rect 34190 15262 34242 15314
rect 34974 15262 35026 15314
rect 37886 15262 37938 15314
rect 38446 15262 38498 15314
rect 39118 15262 39170 15314
rect 39566 15262 39618 15314
rect 40686 15262 40738 15314
rect 44718 15262 44770 15314
rect 46846 15262 46898 15314
rect 47182 15262 47234 15314
rect 47406 15262 47458 15314
rect 47742 15262 47794 15314
rect 49982 15262 50034 15314
rect 50654 15262 50706 15314
rect 51438 15262 51490 15314
rect 2382 15150 2434 15202
rect 3950 15150 4002 15202
rect 5294 15150 5346 15202
rect 7198 15150 7250 15202
rect 9326 15150 9378 15202
rect 9662 15150 9714 15202
rect 10894 15150 10946 15202
rect 12126 15150 12178 15202
rect 12798 15150 12850 15202
rect 13806 15150 13858 15202
rect 16830 15150 16882 15202
rect 17838 15150 17890 15202
rect 21310 15150 21362 15202
rect 24894 15150 24946 15202
rect 38558 15150 38610 15202
rect 42366 15150 42418 15202
rect 43374 15150 43426 15202
rect 43486 15150 43538 15202
rect 45166 15150 45218 15202
rect 46958 15150 47010 15202
rect 47518 15150 47570 15202
rect 49422 15150 49474 15202
rect 50430 15150 50482 15202
rect 51102 15150 51154 15202
rect 53342 15150 53394 15202
rect 54910 15150 54962 15202
rect 4062 15038 4114 15090
rect 6750 15038 6802 15090
rect 26126 15038 26178 15090
rect 32958 15038 33010 15090
rect 41246 15038 41298 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 44466 14870 44518 14922
rect 44570 14870 44622 14922
rect 44674 14870 44726 14922
rect 2382 14702 2434 14754
rect 4622 14702 4674 14754
rect 8878 14702 8930 14754
rect 17502 14702 17554 14754
rect 18622 14702 18674 14754
rect 29598 14702 29650 14754
rect 35982 14702 36034 14754
rect 42030 14702 42082 14754
rect 44942 14702 44994 14754
rect 45166 14702 45218 14754
rect 49870 14702 49922 14754
rect 50878 14702 50930 14754
rect 52558 14702 52610 14754
rect 53342 14702 53394 14754
rect 56030 14702 56082 14754
rect 56366 14702 56418 14754
rect 1598 14590 1650 14642
rect 1822 14590 1874 14642
rect 2494 14590 2546 14642
rect 3502 14590 3554 14642
rect 6078 14590 6130 14642
rect 9886 14590 9938 14642
rect 10894 14590 10946 14642
rect 14814 14590 14866 14642
rect 19070 14590 19122 14642
rect 20078 14590 20130 14642
rect 24670 14590 24722 14642
rect 25678 14590 25730 14642
rect 26126 14590 26178 14642
rect 41022 14590 41074 14642
rect 46174 14590 46226 14642
rect 48638 14590 48690 14642
rect 48750 14590 48802 14642
rect 48974 14590 49026 14642
rect 49534 14590 49586 14642
rect 54462 14590 54514 14642
rect 1150 14478 1202 14530
rect 2158 14478 2210 14530
rect 3054 14478 3106 14530
rect 5406 14478 5458 14530
rect 5854 14478 5906 14530
rect 6638 14478 6690 14530
rect 7310 14478 7362 14530
rect 8094 14478 8146 14530
rect 9102 14478 9154 14530
rect 10334 14478 10386 14530
rect 10670 14478 10722 14530
rect 11342 14478 11394 14530
rect 11902 14478 11954 14530
rect 12126 14478 12178 14530
rect 12910 14478 12962 14530
rect 14478 14478 14530 14530
rect 17054 14478 17106 14530
rect 19518 14478 19570 14530
rect 19966 14478 20018 14530
rect 20750 14478 20802 14530
rect 21086 14478 21138 14530
rect 21310 14478 21362 14530
rect 22094 14478 22146 14530
rect 25006 14478 25058 14530
rect 25566 14478 25618 14530
rect 26798 14478 26850 14530
rect 27806 14478 27858 14530
rect 28926 14478 28978 14530
rect 29486 14478 29538 14530
rect 30270 14478 30322 14530
rect 30606 14478 30658 14530
rect 31614 14478 31666 14530
rect 35422 14478 35474 14530
rect 35870 14478 35922 14530
rect 36654 14478 36706 14530
rect 36990 14478 37042 14530
rect 37998 14478 38050 14530
rect 41358 14478 41410 14530
rect 41806 14478 41858 14530
rect 42702 14478 42754 14530
rect 43038 14478 43090 14530
rect 44046 14478 44098 14530
rect 44830 14478 44882 14530
rect 45726 14478 45778 14530
rect 52894 14478 52946 14530
rect 54910 14478 54962 14530
rect 1038 14366 1090 14418
rect 1486 14366 1538 14418
rect 5070 14366 5122 14418
rect 28590 14366 28642 14418
rect 34974 14366 35026 14418
rect 48414 14366 48466 14418
rect 50430 14366 50482 14418
rect 16046 14254 16098 14306
rect 47294 14254 47346 14306
rect 48190 14254 48242 14306
rect 51998 14254 52050 14306
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 43806 14086 43858 14138
rect 43910 14086 43962 14138
rect 44014 14086 44066 14138
rect 4958 13918 5010 13970
rect 12126 13918 12178 13970
rect 13246 13918 13298 13970
rect 13582 13918 13634 13970
rect 19070 13918 19122 13970
rect 24334 13918 24386 13970
rect 30494 13918 30546 13970
rect 39118 13918 39170 13970
rect 43486 13918 43538 13970
rect 48526 13918 48578 13970
rect 55582 13918 55634 13970
rect 1710 13806 1762 13858
rect 2158 13806 2210 13858
rect 5966 13806 6018 13858
rect 10558 13806 10610 13858
rect 14814 13806 14866 13858
rect 18622 13806 18674 13858
rect 19854 13806 19906 13858
rect 20638 13806 20690 13858
rect 28926 13806 28978 13858
rect 32286 13806 32338 13858
rect 37550 13806 37602 13858
rect 44158 13806 44210 13858
rect 52894 13806 52946 13858
rect 55694 13806 55746 13858
rect 6302 13694 6354 13746
rect 6862 13694 6914 13746
rect 7422 13694 7474 13746
rect 7982 13694 8034 13746
rect 8206 13694 8258 13746
rect 8990 13694 9042 13746
rect 9774 13694 9826 13746
rect 15262 13694 15314 13746
rect 15598 13694 15650 13746
rect 16270 13694 16322 13746
rect 16830 13694 16882 13746
rect 17838 13694 17890 13746
rect 19294 13694 19346 13746
rect 19630 13694 19682 13746
rect 20974 13694 21026 13746
rect 21422 13694 21474 13746
rect 22766 13694 22818 13746
rect 23662 13694 23714 13746
rect 25902 13694 25954 13746
rect 32734 13694 32786 13746
rect 33070 13694 33122 13746
rect 33966 13694 34018 13746
rect 34414 13694 34466 13746
rect 35310 13694 35362 13746
rect 39790 13694 39842 13746
rect 44494 13694 44546 13746
rect 44942 13694 44994 13746
rect 46174 13694 46226 13746
rect 47182 13694 47234 13746
rect 47966 13694 48018 13746
rect 50094 13694 50146 13746
rect 51102 13694 51154 13746
rect 52334 13694 52386 13746
rect 55022 13694 55074 13746
rect 56142 13694 56194 13746
rect 1038 13582 1090 13634
rect 5070 13582 5122 13634
rect 5294 13582 5346 13634
rect 9550 13582 9602 13634
rect 11006 13582 11058 13634
rect 13918 13582 13970 13634
rect 14366 13582 14418 13634
rect 15822 13582 15874 13634
rect 18734 13582 18786 13634
rect 22094 13582 22146 13634
rect 29262 13582 29314 13634
rect 33294 13582 33346 13634
rect 37998 13582 38050 13634
rect 40238 13582 40290 13634
rect 43598 13582 43650 13634
rect 45614 13582 45666 13634
rect 50878 13582 50930 13634
rect 51998 13582 52050 13634
rect 52558 13582 52610 13634
rect 53006 13582 53058 13634
rect 54574 13582 54626 13634
rect 56366 13582 56418 13634
rect 1374 13470 1426 13522
rect 2606 13470 2658 13522
rect 3726 13470 3778 13522
rect 6974 13470 7026 13522
rect 18510 13470 18562 13522
rect 19742 13470 19794 13522
rect 19966 13470 20018 13522
rect 21646 13470 21698 13522
rect 25454 13470 25506 13522
rect 41358 13470 41410 13522
rect 45166 13470 45218 13522
rect 48078 13470 48130 13522
rect 49646 13470 49698 13522
rect 51438 13470 51490 13522
rect 52110 13470 52162 13522
rect 53454 13470 53506 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 1150 13134 1202 13186
rect 2270 13134 2322 13186
rect 4510 13134 4562 13186
rect 7982 13134 8034 13186
rect 15486 13134 15538 13186
rect 17838 13134 17890 13186
rect 23102 13134 23154 13186
rect 25790 13134 25842 13186
rect 28814 13134 28866 13186
rect 34190 13134 34242 13186
rect 35534 13134 35586 13186
rect 36654 13134 36706 13186
rect 37774 13134 37826 13186
rect 41246 13134 41298 13186
rect 45614 13134 45666 13186
rect 46622 13134 46674 13186
rect 46958 13134 47010 13186
rect 47182 13134 47234 13186
rect 47406 13134 47458 13186
rect 48862 13134 48914 13186
rect 52110 13134 52162 13186
rect 52446 13134 52498 13186
rect 53006 13134 53058 13186
rect 53230 13134 53282 13186
rect 54686 13134 54738 13186
rect 56254 13134 56306 13186
rect 3502 13022 3554 13074
rect 8990 13022 9042 13074
rect 9550 13022 9602 13074
rect 11118 13022 11170 13074
rect 14254 13022 14306 13074
rect 16046 13022 16098 13074
rect 20414 13022 20466 13074
rect 22990 13022 23042 13074
rect 23214 13022 23266 13074
rect 27694 13022 27746 13074
rect 33070 13022 33122 13074
rect 44494 13022 44546 13074
rect 46062 13022 46114 13074
rect 46174 13022 46226 13074
rect 50206 13022 50258 13074
rect 51886 13022 51938 13074
rect 52894 13022 52946 13074
rect 2718 12910 2770 12962
rect 3838 12910 3890 12962
rect 4398 12910 4450 12962
rect 5070 12910 5122 12962
rect 5742 12910 5794 12962
rect 6638 12910 6690 12962
rect 6974 12910 7026 12962
rect 7422 12910 7474 12962
rect 7534 12910 7586 12962
rect 7646 12910 7698 12962
rect 8206 12910 8258 12962
rect 9102 12910 9154 12962
rect 10558 12910 10610 12962
rect 10894 12910 10946 12962
rect 11678 12910 11730 12962
rect 12350 12910 12402 12962
rect 13134 12910 13186 12962
rect 13918 12910 13970 12962
rect 15822 12910 15874 12962
rect 16158 12910 16210 12962
rect 17278 12910 17330 12962
rect 19742 12910 19794 12962
rect 20190 12910 20242 12962
rect 20862 12910 20914 12962
rect 21086 12910 21138 12962
rect 21534 12910 21586 12962
rect 22542 12910 22594 12962
rect 32622 12910 32674 12962
rect 34974 12910 35026 12962
rect 37326 12910 37378 12962
rect 40686 12910 40738 12962
rect 41022 12910 41074 12962
rect 41694 12910 41746 12962
rect 42254 12910 42306 12962
rect 43374 12910 43426 12962
rect 44046 12910 44098 12962
rect 46510 12910 46562 12962
rect 48638 12910 48690 12962
rect 48750 12910 48802 12962
rect 48974 12910 49026 12962
rect 52334 12910 52386 12962
rect 55918 12910 55970 12962
rect 10110 12798 10162 12850
rect 16718 12798 16770 12850
rect 18958 12798 19010 12850
rect 19406 12798 19458 12850
rect 26238 12798 26290 12850
rect 27246 12798 27298 12850
rect 40238 12798 40290 12850
rect 47070 12798 47122 12850
rect 49870 12798 49922 12850
rect 52446 12798 52498 12850
rect 55134 12798 55186 12850
rect 8990 12686 9042 12738
rect 9438 12686 9490 12738
rect 9774 12686 9826 12738
rect 16830 12686 16882 12738
rect 24670 12686 24722 12738
rect 38894 12686 38946 12738
rect 48078 12686 48130 12738
rect 48302 12686 48354 12738
rect 51438 12686 51490 12738
rect 53566 12686 53618 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 19070 12350 19122 12402
rect 20638 12350 20690 12402
rect 32734 12350 32786 12402
rect 41694 12350 41746 12402
rect 50990 12350 51042 12402
rect 52110 12350 52162 12402
rect 1150 12238 1202 12290
rect 4958 12238 5010 12290
rect 5406 12238 5458 12290
rect 8990 12238 9042 12290
rect 13358 12238 13410 12290
rect 19966 12238 20018 12290
rect 20750 12238 20802 12290
rect 30158 12238 30210 12290
rect 31166 12238 31218 12290
rect 48302 12238 48354 12290
rect 1486 12126 1538 12178
rect 1934 12126 1986 12178
rect 3278 12126 3330 12178
rect 4174 12126 4226 12178
rect 5742 12126 5794 12178
rect 6302 12126 6354 12178
rect 7086 12126 7138 12178
rect 7422 12126 7474 12178
rect 8542 12126 8594 12178
rect 9326 12126 9378 12178
rect 9886 12126 9938 12178
rect 10558 12126 10610 12178
rect 11230 12126 11282 12178
rect 12014 12126 12066 12178
rect 15710 12126 15762 12178
rect 16158 12126 16210 12178
rect 17502 12126 17554 12178
rect 18398 12126 18450 12178
rect 19854 12126 19906 12178
rect 20078 12126 20130 12178
rect 20974 12126 21026 12178
rect 21422 12126 21474 12178
rect 23102 12126 23154 12178
rect 23886 12126 23938 12178
rect 24446 12126 24498 12178
rect 25006 12126 25058 12178
rect 25566 12126 25618 12178
rect 26574 12126 26626 12178
rect 33966 12126 34018 12178
rect 38222 12126 38274 12178
rect 39230 12126 39282 12178
rect 40350 12126 40402 12178
rect 40798 12126 40850 12178
rect 43262 12126 43314 12178
rect 47294 12126 47346 12178
rect 47966 12126 48018 12178
rect 49758 12126 49810 12178
rect 52446 12126 52498 12178
rect 54014 12126 54066 12178
rect 56030 12126 56082 12178
rect 2158 12014 2210 12066
rect 2606 12014 2658 12066
rect 6862 12014 6914 12066
rect 15374 12014 15426 12066
rect 16382 12014 16434 12066
rect 16830 12014 16882 12066
rect 19182 12014 19234 12066
rect 21982 12014 22034 12066
rect 23550 12014 23602 12066
rect 29822 12014 29874 12066
rect 31614 12014 31666 12066
rect 34526 12014 34578 12066
rect 36766 12014 36818 12066
rect 39790 12014 39842 12066
rect 41246 12014 41298 12066
rect 47518 12014 47570 12066
rect 47742 12014 47794 12066
rect 48638 12014 48690 12066
rect 49422 12014 49474 12066
rect 50318 12014 50370 12066
rect 50654 12014 50706 12066
rect 52670 12014 52722 12066
rect 53006 12014 53058 12066
rect 54462 12014 54514 12066
rect 56366 12014 56418 12066
rect 5070 11902 5122 11954
rect 6414 11902 6466 11954
rect 9998 11902 10050 11954
rect 13806 11902 13858 11954
rect 14926 11902 14978 11954
rect 19630 11902 19682 11954
rect 24558 11902 24610 11954
rect 28590 11902 28642 11954
rect 35646 11902 35698 11954
rect 36318 11902 36370 11954
rect 36430 11902 36482 11954
rect 36542 11902 36594 11954
rect 40238 11902 40290 11954
rect 42814 11902 42866 11954
rect 48190 11902 48242 11954
rect 48414 11902 48466 11954
rect 51326 11902 51378 11954
rect 55582 11902 55634 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 2830 11566 2882 11618
rect 3390 11566 3442 11618
rect 4510 11566 4562 11618
rect 8206 11566 8258 11618
rect 20190 11566 20242 11618
rect 36542 11566 36594 11618
rect 43038 11566 43090 11618
rect 48190 11566 48242 11618
rect 50766 11566 50818 11618
rect 51886 11566 51938 11618
rect 52446 11566 52498 11618
rect 55022 11566 55074 11618
rect 56366 11566 56418 11618
rect 1598 11454 1650 11506
rect 5854 11454 5906 11506
rect 6974 11454 7026 11506
rect 10222 11454 10274 11506
rect 11230 11454 11282 11506
rect 14814 11454 14866 11506
rect 17614 11454 17666 11506
rect 25566 11454 25618 11506
rect 28254 11454 28306 11506
rect 28702 11454 28754 11506
rect 36094 11454 36146 11506
rect 37550 11454 37602 11506
rect 38446 11454 38498 11506
rect 39006 11454 39058 11506
rect 42030 11454 42082 11506
rect 46286 11454 46338 11506
rect 47406 11454 47458 11506
rect 48750 11454 48802 11506
rect 49086 11454 49138 11506
rect 53678 11454 53730 11506
rect 55358 11454 55410 11506
rect 1262 11342 1314 11394
rect 4958 11342 5010 11394
rect 5406 11342 5458 11394
rect 5630 11342 5682 11394
rect 5966 11342 6018 11394
rect 6638 11342 6690 11394
rect 8878 11342 8930 11394
rect 9550 11342 9602 11394
rect 9774 11342 9826 11394
rect 10558 11342 10610 11394
rect 11118 11342 11170 11394
rect 11902 11342 11954 11394
rect 12238 11342 12290 11394
rect 13246 11342 13298 11394
rect 14366 11342 14418 11394
rect 18734 11342 18786 11394
rect 19518 11342 19570 11394
rect 19966 11342 20018 11394
rect 20862 11342 20914 11394
rect 21198 11342 21250 11394
rect 22206 11342 22258 11394
rect 25230 11342 25282 11394
rect 26798 11342 26850 11394
rect 27582 11342 27634 11394
rect 28030 11342 28082 11394
rect 29486 11342 29538 11394
rect 30270 11342 30322 11394
rect 34414 11342 34466 11394
rect 35310 11342 35362 11394
rect 35534 11342 35586 11394
rect 35870 11342 35922 11394
rect 36654 11342 36706 11394
rect 37102 11342 37154 11394
rect 42478 11342 42530 11394
rect 42814 11342 42866 11394
rect 43486 11342 43538 11394
rect 44158 11342 44210 11394
rect 45054 11342 45106 11394
rect 45726 11342 45778 11394
rect 48526 11342 48578 11394
rect 54014 11342 54066 11394
rect 56030 11342 56082 11394
rect 9326 11230 9378 11282
rect 9662 11230 9714 11282
rect 13806 11230 13858 11282
rect 17166 11230 17218 11282
rect 19182 11230 19234 11282
rect 27246 11230 27298 11282
rect 50318 11230 50370 11282
rect 9102 11118 9154 11170
rect 13918 11118 13970 11170
rect 16046 11118 16098 11170
rect 39230 11118 39282 11170
rect 39566 11118 39618 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 10894 10782 10946 10834
rect 22542 10782 22594 10834
rect 36654 10782 36706 10834
rect 39790 10782 39842 10834
rect 43150 10782 43202 10834
rect 52334 10782 52386 10834
rect 52670 10782 52722 10834
rect 4398 10670 4450 10722
rect 11454 10670 11506 10722
rect 16382 10670 16434 10722
rect 20974 10670 21026 10722
rect 29262 10670 29314 10722
rect 35646 10670 35698 10722
rect 38222 10670 38274 10722
rect 44270 10670 44322 10722
rect 49534 10670 49586 10722
rect 52782 10670 52834 10722
rect 1374 10558 1426 10610
rect 2158 10558 2210 10610
rect 2942 10558 2994 10610
rect 3614 10558 3666 10610
rect 4062 10558 4114 10610
rect 5518 10558 5570 10610
rect 5966 10558 6018 10610
rect 6302 10558 6354 10610
rect 7198 10558 7250 10610
rect 7646 10558 7698 10610
rect 8542 10558 8594 10610
rect 9214 10558 9266 10610
rect 11342 10558 11394 10610
rect 11566 10558 11618 10610
rect 12910 10558 12962 10610
rect 14030 10558 14082 10610
rect 14590 10558 14642 10610
rect 15262 10558 15314 10610
rect 15710 10558 15762 10610
rect 16718 10558 16770 10610
rect 17278 10570 17330 10622
rect 17838 10558 17890 10610
rect 18510 10558 18562 10610
rect 19406 10558 19458 10610
rect 23326 10558 23378 10610
rect 23774 10558 23826 10610
rect 24446 10558 24498 10610
rect 25006 10558 25058 10610
rect 26014 10558 26066 10610
rect 29598 10558 29650 10610
rect 30158 10558 30210 10610
rect 30942 10558 30994 10610
rect 31278 10558 31330 10610
rect 32286 10558 32338 10610
rect 32958 10558 33010 10610
rect 35758 10558 35810 10610
rect 36318 10558 36370 10610
rect 36766 10558 36818 10610
rect 41582 10558 41634 10610
rect 44158 10558 44210 10610
rect 47742 10558 47794 10610
rect 48414 10558 48466 10610
rect 48750 10558 48802 10610
rect 48974 10558 49026 10610
rect 49310 10558 49362 10610
rect 50430 10558 50482 10610
rect 50990 10558 51042 10610
rect 51998 10558 52050 10610
rect 53454 10558 53506 10610
rect 56030 10558 56082 10610
rect 4958 10446 5010 10498
rect 6974 10446 7026 10498
rect 16046 10446 16098 10498
rect 22990 10446 23042 10498
rect 37102 10446 37154 10498
rect 38670 10446 38722 10498
rect 42030 10446 42082 10498
rect 44382 10446 44434 10498
rect 47966 10446 48018 10498
rect 48078 10446 48130 10498
rect 48526 10446 48578 10498
rect 50206 10446 50258 10498
rect 50654 10446 50706 10498
rect 53790 10446 53842 10498
rect 56366 10446 56418 10498
rect 3390 10334 3442 10386
rect 5070 10334 5122 10386
rect 5294 10334 5346 10386
rect 6526 10334 6578 10386
rect 9774 10334 9826 10386
rect 11790 10334 11842 10386
rect 15038 10334 15090 10386
rect 17390 10334 17442 10386
rect 21422 10334 21474 10386
rect 23998 10334 24050 10386
rect 30270 10334 30322 10386
rect 33518 10334 33570 10386
rect 34638 10334 34690 10386
rect 36654 10334 36706 10386
rect 44606 10334 44658 10386
rect 49422 10334 49474 10386
rect 49646 10334 49698 10386
rect 51326 10334 51378 10386
rect 52222 10334 52274 10386
rect 55022 10334 55074 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 8878 9998 8930 10050
rect 11006 9998 11058 10050
rect 12126 9998 12178 10050
rect 14926 9998 14978 10050
rect 15598 9998 15650 10050
rect 15710 9998 15762 10050
rect 20302 9998 20354 10050
rect 22766 9998 22818 10050
rect 23886 9998 23938 10050
rect 29038 9998 29090 10050
rect 31278 9998 31330 10050
rect 36206 9998 36258 10050
rect 37326 9998 37378 10050
rect 41470 9998 41522 10050
rect 42590 9998 42642 10050
rect 43150 9998 43202 10050
rect 47294 9998 47346 10050
rect 47406 9998 47458 10050
rect 51662 9998 51714 10050
rect 56366 9998 56418 10050
rect 3726 9886 3778 9938
rect 4734 9886 4786 9938
rect 6862 9886 6914 9938
rect 7310 9886 7362 9938
rect 8318 9886 8370 9938
rect 9886 9886 9938 9938
rect 12014 9886 12066 9938
rect 12238 9886 12290 9938
rect 12686 9886 12738 9938
rect 12798 9886 12850 9938
rect 13806 9886 13858 9938
rect 16158 9886 16210 9938
rect 17726 9886 17778 9938
rect 19182 9886 19234 9938
rect 27918 9886 27970 9938
rect 30046 9886 30098 9938
rect 33406 9886 33458 9938
rect 36094 9886 36146 9938
rect 44382 9886 44434 9938
rect 48190 9886 48242 9938
rect 48750 9886 48802 9938
rect 51102 9886 51154 9938
rect 52782 9886 52834 9938
rect 54014 9886 54066 9938
rect 1710 9774 1762 9826
rect 2494 9774 2546 9826
rect 3054 9774 3106 9826
rect 3950 9774 4002 9826
rect 4398 9774 4450 9826
rect 5294 9774 5346 9826
rect 6302 9774 6354 9826
rect 7422 9774 7474 9826
rect 7870 9774 7922 9826
rect 9214 9774 9266 9826
rect 15934 9774 15986 9826
rect 16606 9774 16658 9826
rect 16830 9774 16882 9826
rect 16942 9774 16994 9826
rect 17166 9774 17218 9826
rect 17502 9774 17554 9826
rect 17838 9774 17890 9826
rect 18062 9774 18114 9826
rect 22206 9774 22258 9826
rect 27470 9774 27522 9826
rect 29598 9774 29650 9826
rect 32734 9774 32786 9826
rect 33182 9774 33234 9826
rect 34078 9774 34130 9826
rect 34638 9774 34690 9826
rect 35534 9774 35586 9826
rect 36878 9774 36930 9826
rect 44830 9774 44882 9826
rect 48974 9774 49026 9826
rect 49310 9774 49362 9826
rect 50766 9774 50818 9826
rect 51998 9774 52050 9826
rect 52670 9774 52722 9826
rect 56142 9774 56194 9826
rect 9438 9662 9490 9714
rect 11454 9662 11506 9714
rect 13358 9662 13410 9714
rect 15710 9662 15762 9714
rect 18734 9662 18786 9714
rect 32398 9662 32450 9714
rect 40350 9662 40402 9714
rect 41022 9662 41074 9714
rect 53678 9662 53730 9714
rect 36318 9550 36370 9602
rect 38446 9550 38498 9602
rect 40462 9550 40514 9602
rect 47182 9550 47234 9602
rect 49982 9550 50034 9602
rect 50318 9550 50370 9602
rect 55246 9550 55298 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 4286 9214 4338 9266
rect 6750 9214 6802 9266
rect 11006 9214 11058 9266
rect 11454 9214 11506 9266
rect 20750 9214 20802 9266
rect 40910 9214 40962 9266
rect 44606 9214 44658 9266
rect 50206 9214 50258 9266
rect 50542 9214 50594 9266
rect 5182 9102 5234 9154
rect 9438 9102 9490 9154
rect 13134 9102 13186 9154
rect 15262 9102 15314 9154
rect 37214 9102 37266 9154
rect 43486 9102 43538 9154
rect 44270 9102 44322 9154
rect 46174 9102 46226 9154
rect 1262 8990 1314 9042
rect 1934 8990 1986 9042
rect 2718 8990 2770 9042
rect 7310 8990 7362 9042
rect 7646 8990 7698 9042
rect 7870 8990 7922 9042
rect 11566 8990 11618 9042
rect 11790 8990 11842 9042
rect 14702 8990 14754 9042
rect 15598 8990 15650 9042
rect 16158 8990 16210 9042
rect 16718 8990 16770 9042
rect 17278 8990 17330 9042
rect 17502 8990 17554 9042
rect 18286 8990 18338 9042
rect 22318 8990 22370 9042
rect 23886 8990 23938 9042
rect 32398 8990 32450 9042
rect 32846 8990 32898 9042
rect 33742 8990 33794 9042
rect 34078 8990 34130 9042
rect 35086 8990 35138 9042
rect 36766 8990 36818 9042
rect 37662 8990 37714 9042
rect 37998 8990 38050 9042
rect 38670 8990 38722 9042
rect 39454 8990 39506 9042
rect 40238 8990 40290 9042
rect 42590 8990 42642 9042
rect 43598 8990 43650 9042
rect 46510 8990 46562 9042
rect 46958 8990 47010 9042
rect 47742 8990 47794 9042
rect 48414 8990 48466 9042
rect 49198 8990 49250 9042
rect 52670 8990 52722 9042
rect 53230 8990 53282 9042
rect 55470 8990 55522 9042
rect 1038 8878 1090 8930
rect 1710 8878 1762 8930
rect 3054 8878 3106 8930
rect 5630 8878 5682 8930
rect 7198 8878 7250 8930
rect 8318 8878 8370 8930
rect 8654 8878 8706 8930
rect 9886 8878 9938 8930
rect 12238 8878 12290 8930
rect 16270 8878 16322 8930
rect 32062 8878 32114 8930
rect 38222 8878 38274 8930
rect 42142 8878 42194 8930
rect 44830 8878 44882 8930
rect 45166 8878 45218 8930
rect 47182 8878 47234 8930
rect 50766 8878 50818 8930
rect 51102 8878 51154 8930
rect 52334 8878 52386 8930
rect 53566 8878 53618 8930
rect 55246 8878 55298 8930
rect 56030 8878 56082 8930
rect 56366 8878 56418 8930
rect 7422 8766 7474 8818
rect 12126 8766 12178 8818
rect 13582 8766 13634 8818
rect 21870 8766 21922 8818
rect 24334 8766 24386 8818
rect 25454 8766 25506 8818
rect 33070 8766 33122 8818
rect 36542 8766 36594 8818
rect 43150 8766 43202 8818
rect 43374 8766 43426 8818
rect 54798 8766 54850 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 2046 8430 2098 8482
rect 3950 8430 4002 8482
rect 16606 8430 16658 8482
rect 16830 8430 16882 8482
rect 44046 8430 44098 8482
rect 46510 8430 46562 8482
rect 48302 8430 48354 8482
rect 49534 8430 49586 8482
rect 51774 8430 51826 8482
rect 56366 8430 56418 8482
rect 3614 8318 3666 8370
rect 4286 8318 4338 8370
rect 7310 8318 7362 8370
rect 8318 8318 8370 8370
rect 11566 8318 11618 8370
rect 12574 8318 12626 8370
rect 15150 8318 15202 8370
rect 16942 8318 16994 8370
rect 17950 8318 18002 8370
rect 20526 8318 20578 8370
rect 26686 8318 26738 8370
rect 30606 8318 30658 8370
rect 33406 8318 33458 8370
rect 37214 8318 37266 8370
rect 38334 8318 38386 8370
rect 40798 8318 40850 8370
rect 42478 8318 42530 8370
rect 45278 8318 45330 8370
rect 48638 8318 48690 8370
rect 50654 8318 50706 8370
rect 52894 8318 52946 8370
rect 54126 8318 54178 8370
rect 55022 8318 55074 8370
rect 56030 8318 56082 8370
rect 4510 8206 4562 8258
rect 5182 8206 5234 8258
rect 6302 8206 6354 8258
rect 6862 8206 6914 8258
rect 7422 8206 7474 8258
rect 7870 8206 7922 8258
rect 9550 8206 9602 8258
rect 10334 8206 10386 8258
rect 10894 8206 10946 8258
rect 11790 8206 11842 8258
rect 12126 8206 12178 8258
rect 13246 8211 13298 8263
rect 13918 8206 13970 8258
rect 14702 8206 14754 8258
rect 15374 8206 15426 8258
rect 15822 8206 15874 8258
rect 17390 8206 17442 8258
rect 19070 8206 19122 8258
rect 19854 8206 19906 8258
rect 20302 8206 20354 8258
rect 20974 8206 21026 8258
rect 21534 8206 21586 8258
rect 22542 8206 22594 8258
rect 26014 8206 26066 8258
rect 26462 8206 26514 8258
rect 27134 8206 27186 8258
rect 27918 8206 27970 8258
rect 28814 8206 28866 8258
rect 32734 8206 32786 8258
rect 33182 8206 33234 8258
rect 33854 8206 33906 8258
rect 34414 8206 34466 8258
rect 35422 8206 35474 8258
rect 36766 8206 36818 8258
rect 40686 8206 40738 8258
rect 41022 8206 41074 8258
rect 43486 8206 43538 8258
rect 43822 8206 43874 8258
rect 44270 8206 44322 8258
rect 44830 8206 44882 8258
rect 47966 8206 48018 8258
rect 48302 8206 48354 8258
rect 54462 8206 54514 8258
rect 54910 8206 54962 8258
rect 1598 8094 1650 8146
rect 8990 8094 9042 8146
rect 16158 8094 16210 8146
rect 17502 8094 17554 8146
rect 19518 8094 19570 8146
rect 25678 8094 25730 8146
rect 30158 8094 30210 8146
rect 32398 8094 32450 8146
rect 42926 8094 42978 8146
rect 43934 8094 43986 8146
rect 51102 8094 51154 8146
rect 53342 8094 53394 8146
rect 3166 7982 3218 8034
rect 8878 7982 8930 8034
rect 31726 7982 31778 8034
rect 41358 7982 41410 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 3166 7646 3218 7698
rect 4958 7646 5010 7698
rect 31838 7646 31890 7698
rect 43374 7646 43426 7698
rect 45950 7646 46002 7698
rect 48190 7646 48242 7698
rect 48750 7646 48802 7698
rect 1598 7534 1650 7586
rect 8654 7534 8706 7586
rect 12238 7534 12290 7586
rect 20638 7534 20690 7586
rect 24670 7534 24722 7586
rect 32510 7534 32562 7586
rect 37886 7534 37938 7586
rect 52222 7534 52274 7586
rect 3950 7422 4002 7474
rect 5070 7422 5122 7474
rect 5630 7422 5682 7474
rect 6414 7422 6466 7474
rect 6974 7422 7026 7474
rect 7758 7422 7810 7474
rect 8206 7422 8258 7474
rect 9102 7422 9154 7474
rect 9998 7422 10050 7474
rect 10670 7422 10722 7474
rect 11342 7422 11394 7474
rect 11902 7422 11954 7474
rect 13134 7422 13186 7474
rect 14926 7422 14978 7474
rect 16270 7422 16322 7474
rect 16718 7422 16770 7474
rect 17950 7422 18002 7474
rect 18958 7422 19010 7474
rect 20974 7422 21026 7474
rect 21422 7422 21474 7474
rect 22318 7422 22370 7474
rect 22654 7422 22706 7474
rect 23662 7422 23714 7474
rect 25006 7422 25058 7474
rect 25454 7422 25506 7474
rect 26126 7422 26178 7474
rect 26798 7422 26850 7474
rect 27806 7422 27858 7474
rect 30270 7422 30322 7474
rect 32846 7422 32898 7474
rect 33294 7422 33346 7474
rect 34190 7422 34242 7474
rect 34750 7422 34802 7474
rect 35646 7422 35698 7474
rect 38222 7422 38274 7474
rect 38782 7422 38834 7474
rect 39342 7422 39394 7474
rect 39902 7422 39954 7474
rect 40910 7422 40962 7474
rect 41806 7422 41858 7474
rect 44270 7422 44322 7474
rect 46510 7422 46562 7474
rect 50318 7422 50370 7474
rect 51438 7422 51490 7474
rect 54462 7422 54514 7474
rect 2046 7310 2098 7362
rect 3614 7310 3666 7362
rect 4286 7310 4338 7362
rect 4398 7310 4450 7362
rect 12798 7310 12850 7362
rect 13470 7310 13522 7362
rect 14254 7310 14306 7362
rect 14366 7310 14418 7362
rect 14814 7310 14866 7362
rect 15934 7310 15986 7362
rect 17390 7310 17442 7362
rect 30718 7310 30770 7362
rect 38894 7310 38946 7362
rect 42142 7310 42194 7362
rect 44830 7310 44882 7362
rect 46958 7310 47010 7362
rect 49870 7310 49922 7362
rect 52558 7310 52610 7362
rect 54798 7310 54850 7362
rect 7646 7198 7698 7250
rect 11230 7198 11282 7250
rect 13806 7198 13858 7250
rect 14030 7198 14082 7250
rect 14590 7198 14642 7250
rect 16942 7198 16994 7250
rect 21646 7198 21698 7250
rect 25678 7198 25730 7250
rect 33518 7198 33570 7250
rect 51102 7198 51154 7250
rect 53790 7198 53842 7250
rect 56030 7198 56082 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 3838 6862 3890 6914
rect 9326 6862 9378 6914
rect 14478 6862 14530 6914
rect 15822 6862 15874 6914
rect 35422 6862 35474 6914
rect 46174 6862 46226 6914
rect 53118 6862 53170 6914
rect 54126 6862 54178 6914
rect 56254 6862 56306 6914
rect 1934 6750 1986 6802
rect 4398 6750 4450 6802
rect 7310 6750 7362 6802
rect 8318 6750 8370 6802
rect 9102 6750 9154 6802
rect 10110 6750 10162 6802
rect 11790 6750 11842 6802
rect 14590 6750 14642 6802
rect 14926 6750 14978 6802
rect 15038 6750 15090 6802
rect 15262 6750 15314 6802
rect 15934 6750 15986 6802
rect 16718 6750 16770 6802
rect 18062 6750 18114 6802
rect 21870 6750 21922 6802
rect 23662 6750 23714 6802
rect 24558 6750 24610 6802
rect 25566 6750 25618 6802
rect 27246 6750 27298 6802
rect 30494 6750 30546 6802
rect 33070 6750 33122 6802
rect 34414 6750 34466 6802
rect 34750 6750 34802 6802
rect 35646 6750 35698 6802
rect 36430 6750 36482 6802
rect 38446 6750 38498 6802
rect 41246 6750 41298 6802
rect 44382 6750 44434 6802
rect 46286 6750 46338 6802
rect 46622 6750 46674 6802
rect 50542 6750 50594 6802
rect 52782 6750 52834 6802
rect 55918 6750 55970 6802
rect 1486 6638 1538 6690
rect 3054 6638 3106 6690
rect 3502 6638 3554 6690
rect 4286 6638 4338 6690
rect 4622 6638 4674 6690
rect 4846 6638 4898 6690
rect 5294 6638 5346 6690
rect 6190 6638 6242 6690
rect 6638 6638 6690 6690
rect 7534 6638 7586 6690
rect 7982 6638 8034 6690
rect 8878 6638 8930 6690
rect 9214 6638 9266 6690
rect 9438 6638 9490 6690
rect 9998 6638 10050 6690
rect 10558 6638 10610 6690
rect 11118 6638 11170 6690
rect 11566 6638 11618 6690
rect 12350 6638 12402 6690
rect 12798 6638 12850 6690
rect 13806 6638 13858 6690
rect 14254 6638 14306 6690
rect 15486 6638 15538 6690
rect 15710 6638 15762 6690
rect 16158 6638 16210 6690
rect 17054 6638 17106 6690
rect 17502 6638 17554 6690
rect 19182 6638 19234 6690
rect 19742 6638 19794 6690
rect 20862 6638 20914 6690
rect 21198 6638 21250 6690
rect 21982 6638 22034 6690
rect 22430 6638 22482 6690
rect 22878 6638 22930 6690
rect 23998 6638 24050 6690
rect 24894 6638 24946 6690
rect 25902 6638 25954 6690
rect 26686 6638 26738 6690
rect 27134 6638 27186 6690
rect 27806 6638 27858 6690
rect 28478 6638 28530 6690
rect 29374 6638 29426 6690
rect 33294 6638 33346 6690
rect 34974 6638 35026 6690
rect 35534 6638 35586 6690
rect 35982 6638 36034 6690
rect 39566 6638 39618 6690
rect 40574 6638 40626 6690
rect 41022 6638 41074 6690
rect 41694 6638 41746 6690
rect 42366 6638 42418 6690
rect 43262 6638 43314 6690
rect 46062 6638 46114 6690
rect 46510 6638 46562 6690
rect 50206 6638 50258 6690
rect 10334 6526 10386 6578
rect 10782 6526 10834 6578
rect 15934 6526 15986 6578
rect 23438 6526 23490 6578
rect 26238 6526 26290 6578
rect 30158 6526 30210 6578
rect 32510 6526 32562 6578
rect 33182 6526 33234 6578
rect 33518 6526 33570 6578
rect 34190 6526 34242 6578
rect 35086 6526 35138 6578
rect 37998 6526 38050 6578
rect 40238 6526 40290 6578
rect 44046 6526 44098 6578
rect 53678 6526 53730 6578
rect 25902 6414 25954 6466
rect 31726 6414 31778 6466
rect 32622 6414 32674 6466
rect 33742 6414 33794 6466
rect 34078 6414 34130 6466
rect 36318 6414 36370 6466
rect 45614 6414 45666 6466
rect 51774 6414 51826 6466
rect 55246 6414 55298 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 1262 6078 1314 6130
rect 6750 6078 6802 6130
rect 20078 6078 20130 6130
rect 21870 6078 21922 6130
rect 28478 6078 28530 6130
rect 34190 6078 34242 6130
rect 34638 6078 34690 6130
rect 36878 6078 36930 6130
rect 39006 6078 39058 6130
rect 41246 6078 41298 6130
rect 44270 6078 44322 6130
rect 44606 6078 44658 6130
rect 52110 6078 52162 6130
rect 52446 6078 52498 6130
rect 53790 6078 53842 6130
rect 2830 5966 2882 6018
rect 5182 5966 5234 6018
rect 12014 5966 12066 6018
rect 12910 5966 12962 6018
rect 14478 5966 14530 6018
rect 21534 5966 21586 6018
rect 22654 5966 22706 6018
rect 24670 5966 24722 6018
rect 39678 5966 39730 6018
rect 41918 5966 41970 6018
rect 7086 5854 7138 5906
rect 8094 5854 8146 5906
rect 8542 5854 8594 5906
rect 9214 5854 9266 5906
rect 9886 5854 9938 5906
rect 10894 5854 10946 5906
rect 11454 5854 11506 5906
rect 11678 5854 11730 5906
rect 11902 5854 11954 5906
rect 12126 5854 12178 5906
rect 12686 5854 12738 5906
rect 13246 5854 13298 5906
rect 14142 5854 14194 5906
rect 14366 5854 14418 5906
rect 15262 5854 15314 5906
rect 15822 5854 15874 5906
rect 16494 5854 16546 5906
rect 17166 5854 17218 5906
rect 17950 5854 18002 5906
rect 19742 5854 19794 5906
rect 20750 5854 20802 5906
rect 24222 5854 24274 5906
rect 25006 5854 25058 5906
rect 25454 5854 25506 5906
rect 26126 5854 26178 5906
rect 26686 5854 26738 5906
rect 27694 5854 27746 5906
rect 29486 5854 29538 5906
rect 32622 5854 32674 5906
rect 36318 5854 36370 5906
rect 36542 5854 36594 5906
rect 36990 5854 37042 5906
rect 39006 5854 39058 5906
rect 45054 5854 45106 5906
rect 45390 5854 45442 5906
rect 52894 5854 52946 5906
rect 53118 5854 53170 5906
rect 54126 5854 54178 5906
rect 55806 5854 55858 5906
rect 2382 5742 2434 5794
rect 3502 5742 3554 5794
rect 5518 5742 5570 5794
rect 7310 5742 7362 5794
rect 7422 5742 7474 5794
rect 7758 5742 7810 5794
rect 8766 5742 8818 5794
rect 13134 5742 13186 5794
rect 14590 5742 14642 5794
rect 14926 5742 14978 5794
rect 15934 5742 15986 5794
rect 23102 5742 23154 5794
rect 29934 5742 29986 5794
rect 34862 5742 34914 5794
rect 38670 5742 38722 5794
rect 40126 5742 40178 5794
rect 42254 5742 42306 5794
rect 45166 5742 45218 5794
rect 53230 5742 53282 5794
rect 54350 5742 54402 5794
rect 54910 5742 54962 5794
rect 3838 5630 3890 5682
rect 19854 5630 19906 5682
rect 19966 5630 20018 5682
rect 20638 5630 20690 5682
rect 20862 5630 20914 5682
rect 21086 5630 21138 5682
rect 21646 5630 21698 5682
rect 25678 5630 25730 5682
rect 28590 5630 28642 5682
rect 28702 5630 28754 5682
rect 31166 5630 31218 5682
rect 33070 5630 33122 5682
rect 34750 5630 34802 5682
rect 36766 5630 36818 5682
rect 37550 5630 37602 5682
rect 37886 5630 37938 5682
rect 43486 5630 43538 5682
rect 55470 5630 55522 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 1038 5294 1090 5346
rect 1374 5294 1426 5346
rect 5630 5294 5682 5346
rect 6750 5294 6802 5346
rect 7982 5294 8034 5346
rect 9214 5294 9266 5346
rect 12574 5294 12626 5346
rect 14590 5294 14642 5346
rect 16606 5294 16658 5346
rect 18174 5294 18226 5346
rect 19294 5294 19346 5346
rect 23998 5294 24050 5346
rect 25342 5294 25394 5346
rect 27246 5294 27298 5346
rect 27358 5294 27410 5346
rect 33070 5294 33122 5346
rect 33518 5294 33570 5346
rect 33630 5294 33682 5346
rect 33742 5294 33794 5346
rect 36878 5294 36930 5346
rect 37102 5294 37154 5346
rect 38446 5294 38498 5346
rect 39230 5294 39282 5346
rect 39342 5294 39394 5346
rect 42366 5294 42418 5346
rect 44830 5294 44882 5346
rect 53342 5294 53394 5346
rect 53678 5294 53730 5346
rect 54126 5294 54178 5346
rect 1934 5182 1986 5234
rect 2942 5182 2994 5234
rect 7758 5182 7810 5234
rect 8878 5182 8930 5234
rect 9550 5182 9602 5234
rect 16830 5182 16882 5234
rect 16942 5182 16994 5234
rect 20750 5182 20802 5234
rect 23662 5182 23714 5234
rect 25006 5182 25058 5234
rect 28030 5182 28082 5234
rect 34414 5182 34466 5234
rect 34526 5182 34578 5234
rect 36654 5182 36706 5234
rect 41358 5182 41410 5234
rect 55246 5182 55298 5234
rect 55918 5182 55970 5234
rect 2382 5070 2434 5122
rect 2718 5070 2770 5122
rect 3614 5070 3666 5122
rect 4062 5070 4114 5122
rect 4958 5070 5010 5122
rect 7982 5070 8034 5122
rect 8206 5070 8258 5122
rect 9886 5070 9938 5122
rect 10446 5070 10498 5122
rect 11342 5070 11394 5122
rect 11902 5070 11954 5122
rect 12686 5070 12738 5122
rect 13134 5070 13186 5122
rect 14142 5070 14194 5122
rect 17614 5070 17666 5122
rect 19742 5070 19794 5122
rect 20190 5070 20242 5122
rect 20526 5070 20578 5122
rect 21422 5070 21474 5122
rect 21982 5070 22034 5122
rect 22766 5070 22818 5122
rect 25902 5070 25954 5122
rect 26798 5070 26850 5122
rect 27470 5070 27522 5122
rect 27918 5070 27970 5122
rect 32846 5070 32898 5122
rect 34190 5070 34242 5122
rect 38670 5070 38722 5122
rect 41806 5070 41858 5122
rect 42142 5070 42194 5122
rect 43038 5070 43090 5122
rect 43486 5070 43538 5122
rect 44382 5070 44434 5122
rect 54910 5070 54962 5122
rect 56254 5070 56306 5122
rect 7198 4958 7250 5010
rect 13582 4958 13634 5010
rect 26126 4958 26178 5010
rect 26238 4958 26290 5010
rect 27022 4958 27074 5010
rect 33182 4958 33234 5010
rect 36990 4958 37042 5010
rect 37998 4958 38050 5010
rect 38222 4958 38274 5010
rect 38558 4958 38610 5010
rect 54462 4958 54514 5010
rect 15710 4846 15762 4898
rect 26574 4846 26626 4898
rect 39118 4846 39170 4898
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 2942 4510 2994 4562
rect 10446 4510 10498 4562
rect 14590 4510 14642 4562
rect 19182 4510 19234 4562
rect 20750 4510 20802 4562
rect 25118 4510 25170 4562
rect 37998 4510 38050 4562
rect 55694 4510 55746 4562
rect 8878 4398 8930 4450
rect 15038 4398 15090 4450
rect 18622 4398 18674 4450
rect 19070 4398 19122 4450
rect 26910 4398 26962 4450
rect 30606 4398 30658 4450
rect 38334 4398 38386 4450
rect 40350 4398 40402 4450
rect 44830 4398 44882 4450
rect 1374 4286 1426 4338
rect 3726 4286 3778 4338
rect 4398 4286 4450 4338
rect 5070 4286 5122 4338
rect 5630 4286 5682 4338
rect 6526 4286 6578 4338
rect 7310 4286 7362 4338
rect 8094 4286 8146 4338
rect 12910 4286 12962 4338
rect 15486 4286 15538 4338
rect 15934 4286 15986 4338
rect 16606 4286 16658 4338
rect 17278 4286 17330 4338
rect 18062 4286 18114 4338
rect 19854 4286 19906 4338
rect 19966 4286 20018 4338
rect 20078 4286 20130 4338
rect 20638 4286 20690 4338
rect 21310 4286 21362 4338
rect 21646 4286 21698 4338
rect 22094 4286 22146 4338
rect 22990 4286 23042 4338
rect 23550 4286 23602 4338
rect 26798 4286 26850 4338
rect 27022 4286 27074 4338
rect 27470 4286 27522 4338
rect 30158 4286 30210 4338
rect 31054 4286 31106 4338
rect 31390 4286 31442 4338
rect 32174 4286 32226 4338
rect 32622 4286 32674 4338
rect 33742 4286 33794 4338
rect 35758 4286 35810 4338
rect 36430 4286 36482 4338
rect 39790 4286 39842 4338
rect 40686 4286 40738 4338
rect 41246 4286 41298 4338
rect 42590 4286 42642 4338
rect 43374 4286 43426 4338
rect 44158 4286 44210 4338
rect 44494 4286 44546 4338
rect 46286 4286 46338 4338
rect 54462 4286 54514 4338
rect 54910 4286 54962 4338
rect 56030 4286 56082 4338
rect 1822 4174 1874 4226
rect 3390 4174 3442 4226
rect 4062 4174 4114 4226
rect 6302 4174 6354 4226
rect 6974 4174 7026 4226
rect 7534 4174 7586 4226
rect 9214 4174 9266 4226
rect 10894 4174 10946 4226
rect 11566 4174 11618 4226
rect 13358 4174 13410 4226
rect 27246 4174 27298 4226
rect 36318 4174 36370 4226
rect 38222 4174 38274 4226
rect 41358 4174 41410 4226
rect 41806 4174 41858 4226
rect 55134 4174 55186 4226
rect 5294 4062 5346 4114
rect 5966 4062 6018 4114
rect 7870 4062 7922 4114
rect 11230 4062 11282 4114
rect 11902 4062 11954 4114
rect 16046 4062 16098 4114
rect 18734 4062 18786 4114
rect 19630 4062 19682 4114
rect 21086 4062 21138 4114
rect 21422 4062 21474 4114
rect 22318 4062 22370 4114
rect 22654 4062 22706 4114
rect 23998 4062 24050 4114
rect 26126 4062 26178 4114
rect 26462 4062 26514 4114
rect 28478 4062 28530 4114
rect 28814 4062 28866 4114
rect 29934 4062 29986 4114
rect 31614 4062 31666 4114
rect 34190 4062 34242 4114
rect 34526 4062 34578 4114
rect 35422 4062 35474 4114
rect 40014 4062 40066 4114
rect 44270 4062 44322 4114
rect 46510 4062 46562 4114
rect 54126 4062 54178 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 1374 3726 1426 3778
rect 2046 3726 2098 3778
rect 2830 3726 2882 3778
rect 3950 3726 4002 3778
rect 5630 3726 5682 3778
rect 6750 3726 6802 3778
rect 7310 3726 7362 3778
rect 7982 3726 8034 3778
rect 8318 3726 8370 3778
rect 9102 3726 9154 3778
rect 9774 3726 9826 3778
rect 11118 3726 11170 3778
rect 12238 3726 12290 3778
rect 13022 3726 13074 3778
rect 16942 3726 16994 3778
rect 21646 3726 21698 3778
rect 24894 3726 24946 3778
rect 25566 3726 25618 3778
rect 26574 3726 26626 3778
rect 27694 3726 27746 3778
rect 29150 3726 29202 3778
rect 32398 3726 32450 3778
rect 34302 3726 34354 3778
rect 36766 3726 36818 3778
rect 37550 3726 37602 3778
rect 37998 3726 38050 3778
rect 42142 3726 42194 3778
rect 42814 3726 42866 3778
rect 44830 3726 44882 3778
rect 46174 3726 46226 3778
rect 46846 3726 46898 3778
rect 55022 3726 55074 3778
rect 55358 3726 55410 3778
rect 56030 3726 56082 3778
rect 56366 3726 56418 3778
rect 7646 3614 7698 3666
rect 9438 3614 9490 3666
rect 10110 3614 10162 3666
rect 12686 3614 12738 3666
rect 13694 3614 13746 3666
rect 14926 3614 14978 3666
rect 17054 3614 17106 3666
rect 18734 3614 18786 3666
rect 19854 3614 19906 3666
rect 20974 3614 21026 3666
rect 21758 3614 21810 3666
rect 22654 3614 22706 3666
rect 24558 3614 24610 3666
rect 25230 3614 25282 3666
rect 28142 3614 28194 3666
rect 32734 3614 32786 3666
rect 35870 3614 35922 3666
rect 36094 3614 36146 3666
rect 37214 3614 37266 3666
rect 39678 3614 39730 3666
rect 40910 3614 40962 3666
rect 43038 3614 43090 3666
rect 44158 3614 44210 3666
rect 45166 3614 45218 3666
rect 45502 3614 45554 3666
rect 47070 3614 47122 3666
rect 1598 3502 1650 3554
rect 2382 3502 2434 3554
rect 5182 3502 5234 3554
rect 10670 3502 10722 3554
rect 13470 3502 13522 3554
rect 14478 3502 14530 3554
rect 16606 3502 16658 3554
rect 17166 3502 17218 3554
rect 18174 3502 18226 3554
rect 20526 3502 20578 3554
rect 20750 3502 20802 3554
rect 21198 3502 21250 3554
rect 22318 3502 22370 3554
rect 26126 3502 26178 3554
rect 28478 3502 28530 3554
rect 29038 3502 29090 3554
rect 29822 3502 29874 3554
rect 30158 3502 30210 3554
rect 31166 3502 31218 3554
rect 33854 3502 33906 3554
rect 39342 3502 39394 3554
rect 43374 3502 43426 3554
rect 45838 3502 45890 3554
rect 47406 3502 47458 3554
rect 4398 3390 4450 3442
rect 16046 3390 16098 3442
rect 21086 3390 21138 3442
rect 35422 3390 35474 3442
rect 36206 3390 36258 3442
rect 36542 3390 36594 3442
rect 36878 3390 36930 3442
rect 37886 3390 37938 3442
rect 40574 3390 40626 3442
rect 23886 3278 23938 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 1150 2942 1202 2994
rect 5630 2942 5682 2994
rect 10558 2942 10610 2994
rect 15374 2942 15426 2994
rect 22206 2942 22258 2994
rect 30270 2942 30322 2994
rect 40014 2942 40066 2994
rect 2718 2830 2770 2882
rect 7646 2830 7698 2882
rect 13806 2830 13858 2882
rect 16606 2830 16658 2882
rect 17278 2830 17330 2882
rect 28702 2830 28754 2882
rect 43486 2830 43538 2882
rect 3726 2718 3778 2770
rect 4286 2718 4338 2770
rect 7198 2718 7250 2770
rect 8094 2718 8146 2770
rect 8878 2718 8930 2770
rect 11230 2718 11282 2770
rect 12014 2718 12066 2770
rect 13022 2718 13074 2770
rect 16158 2718 16210 2770
rect 19518 2718 19570 2770
rect 20974 2718 21026 2770
rect 21198 2718 21250 2770
rect 21310 2718 21362 2770
rect 21870 2718 21922 2770
rect 22430 2718 22482 2770
rect 23774 2718 23826 2770
rect 24222 2718 24274 2770
rect 24894 2718 24946 2770
rect 25678 2718 25730 2770
rect 26462 2718 26514 2770
rect 27806 2718 27858 2770
rect 31054 2718 31106 2770
rect 31502 2718 31554 2770
rect 32174 2718 32226 2770
rect 32958 2718 33010 2770
rect 33742 2718 33794 2770
rect 34302 2718 34354 2770
rect 35198 2718 35250 2770
rect 35758 2718 35810 2770
rect 36654 2718 36706 2770
rect 37326 2718 37378 2770
rect 37662 2718 37714 2770
rect 38558 2718 38610 2770
rect 39342 2718 39394 2770
rect 41694 2718 41746 2770
rect 42142 2718 42194 2770
rect 42814 2718 42866 2770
rect 43598 2718 43650 2770
rect 44494 2718 44546 2770
rect 44830 2718 44882 2770
rect 45502 2718 45554 2770
rect 46510 2718 46562 2770
rect 46846 2718 46898 2770
rect 48414 2718 48466 2770
rect 55582 2718 55634 2770
rect 56254 2718 56306 2770
rect 2270 2606 2322 2658
rect 3390 2606 3442 2658
rect 6862 2606 6914 2658
rect 8430 2606 8482 2658
rect 9326 2606 9378 2658
rect 14254 2606 14306 2658
rect 15822 2606 15874 2658
rect 16718 2606 16770 2658
rect 19966 2606 20018 2658
rect 20750 2606 20802 2658
rect 22654 2606 22706 2658
rect 22990 2606 23042 2658
rect 23102 2606 23154 2658
rect 23438 2606 23490 2658
rect 29038 2606 29090 2658
rect 30718 2606 30770 2658
rect 34974 2606 35026 2658
rect 35646 2606 35698 2658
rect 41134 2606 41186 2658
rect 44158 2606 44210 2658
rect 46174 2606 46226 2658
rect 48862 2606 48914 2658
rect 55246 2606 55298 2658
rect 55918 2606 55970 2658
rect 4062 2494 4114 2546
rect 11566 2494 11618 2546
rect 12238 2494 12290 2546
rect 12798 2494 12850 2546
rect 17726 2494 17778 2546
rect 18846 2494 18898 2546
rect 19854 2494 19906 2546
rect 20078 2494 20130 2546
rect 21534 2494 21586 2546
rect 22542 2494 22594 2546
rect 24446 2494 24498 2546
rect 27582 2494 27634 2546
rect 31726 2494 31778 2546
rect 34638 2494 34690 2546
rect 36318 2494 36370 2546
rect 36990 2494 37042 2546
rect 37998 2494 38050 2546
rect 38334 2494 38386 2546
rect 39566 2494 39618 2546
rect 42478 2494 42530 2546
rect 43150 2494 43202 2546
rect 45166 2494 45218 2546
rect 45838 2494 45890 2546
rect 47182 2494 47234 2546
rect 47518 2494 47570 2546
rect 47854 2494 47906 2546
rect 48190 2494 48242 2546
rect 49198 2494 49250 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 1598 2158 1650 2210
rect 2270 2158 2322 2210
rect 5294 2158 5346 2210
rect 6414 2158 6466 2210
rect 7982 2158 8034 2210
rect 9662 2158 9714 2210
rect 10782 2158 10834 2210
rect 11342 2158 11394 2210
rect 12462 2158 12514 2210
rect 13470 2158 13522 2210
rect 13918 2158 13970 2210
rect 14926 2158 14978 2210
rect 15262 2158 15314 2210
rect 15598 2158 15650 2210
rect 17054 2158 17106 2210
rect 19294 2158 19346 2210
rect 23886 2158 23938 2210
rect 24894 2158 24946 2210
rect 25230 2158 25282 2210
rect 26574 2158 26626 2210
rect 27694 2158 27746 2210
rect 28590 2158 28642 2210
rect 28926 2158 28978 2210
rect 29262 2158 29314 2210
rect 30606 2158 30658 2210
rect 31726 2158 31778 2210
rect 33630 2158 33682 2210
rect 34414 2158 34466 2210
rect 35086 2158 35138 2210
rect 36206 2158 36258 2210
rect 37550 2158 37602 2210
rect 38222 2158 38274 2210
rect 38558 2158 38610 2210
rect 38894 2158 38946 2210
rect 39230 2158 39282 2210
rect 40798 2158 40850 2210
rect 41470 2158 41522 2210
rect 42142 2158 42194 2210
rect 42926 2158 42978 2210
rect 43934 2158 43986 2210
rect 44270 2158 44322 2210
rect 44942 2158 44994 2210
rect 45614 2158 45666 2210
rect 46286 2158 46338 2210
rect 47294 2158 47346 2210
rect 48078 2158 48130 2210
rect 48414 2158 48466 2210
rect 48750 2158 48802 2210
rect 49086 2158 49138 2210
rect 49758 2158 49810 2210
rect 55918 2158 55970 2210
rect 2606 2046 2658 2098
rect 3502 2046 3554 2098
rect 4734 2046 4786 2098
rect 13582 2046 13634 2098
rect 14590 2046 14642 2098
rect 16158 2046 16210 2098
rect 16718 2046 16770 2098
rect 17726 2046 17778 2098
rect 18286 2046 18338 2098
rect 22654 2046 22706 2098
rect 24558 2046 24610 2098
rect 25566 2046 25618 2098
rect 29598 2046 29650 2098
rect 32510 2046 32562 2098
rect 33070 2046 33122 2098
rect 34078 2046 34130 2098
rect 37214 2046 37266 2098
rect 37886 2046 37938 2098
rect 39566 2046 39618 2098
rect 40462 2046 40514 2098
rect 41134 2046 41186 2098
rect 43262 2046 43314 2098
rect 43598 2046 43650 2098
rect 44606 2046 44658 2098
rect 45278 2046 45330 2098
rect 46622 2046 46674 2098
rect 46958 2046 47010 2098
rect 49422 2046 49474 2098
rect 1934 1934 1986 1986
rect 3166 1934 3218 1986
rect 6974 1934 7026 1986
rect 8206 1934 8258 1986
rect 9102 1934 9154 1986
rect 12910 1934 12962 1986
rect 14142 1934 14194 1986
rect 17950 1934 18002 1986
rect 18734 1934 18786 1986
rect 19070 1934 19122 1986
rect 19854 1934 19906 1986
rect 20302 1934 20354 1986
rect 21422 1934 21474 1986
rect 22318 1934 22370 1986
rect 26014 1934 26066 1986
rect 30046 1934 30098 1986
rect 33294 1934 33346 1986
rect 36766 1934 36818 1986
rect 45838 1934 45890 1986
rect 56142 1934 56194 1986
rect 1374 1822 1426 1874
rect 17614 1822 17666 1874
rect 16046 1710 16098 1762
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 2494 1374 2546 1426
rect 5630 1374 5682 1426
rect 8766 1374 8818 1426
rect 19182 1374 19234 1426
rect 33294 1374 33346 1426
rect 42254 1374 42306 1426
rect 31726 1262 31778 1314
rect 40686 1262 40738 1314
rect 42926 1262 42978 1314
rect 44270 1262 44322 1314
rect 44830 1262 44882 1314
rect 46286 1262 46338 1314
rect 48078 1262 48130 1314
rect 1038 1150 1090 1202
rect 1822 1150 1874 1202
rect 4174 1150 4226 1202
rect 4846 1150 4898 1202
rect 7198 1150 7250 1202
rect 10334 1150 10386 1202
rect 11790 1150 11842 1202
rect 12574 1150 12626 1202
rect 14254 1150 14306 1202
rect 15486 1150 15538 1202
rect 16494 1150 16546 1202
rect 17502 1150 17554 1202
rect 20302 1150 20354 1202
rect 21086 1150 21138 1202
rect 21646 1150 21698 1202
rect 23102 1150 23154 1202
rect 24222 1150 24274 1202
rect 24894 1150 24946 1202
rect 25454 1150 25506 1202
rect 26126 1150 26178 1202
rect 26910 1150 26962 1202
rect 28030 1150 28082 1202
rect 28702 1150 28754 1202
rect 29374 1150 29426 1202
rect 30158 1150 30210 1202
rect 35534 1150 35586 1202
rect 36318 1150 36370 1202
rect 36878 1150 36930 1202
rect 37662 1150 37714 1202
rect 38222 1150 38274 1202
rect 39454 1150 39506 1202
rect 40014 1150 40066 1202
rect 43486 1150 43538 1202
rect 45278 1150 45330 1202
rect 46958 1150 47010 1202
rect 47630 1150 47682 1202
rect 48638 1150 48690 1202
rect 49198 1150 49250 1202
rect 49870 1150 49922 1202
rect 50766 1150 50818 1202
rect 1374 1038 1426 1090
rect 2046 1038 2098 1090
rect 3614 1038 3666 1090
rect 6862 1038 6914 1090
rect 9886 1038 9938 1090
rect 11230 1038 11282 1090
rect 13694 1038 13746 1090
rect 18062 1038 18114 1090
rect 21982 1038 22034 1090
rect 22318 1038 22370 1090
rect 24446 1038 24498 1090
rect 25790 1038 25842 1090
rect 29038 1038 29090 1090
rect 29710 1038 29762 1090
rect 32062 1038 32114 1090
rect 34750 1038 34802 1090
rect 35310 1038 35362 1090
rect 41022 1038 41074 1090
rect 47406 1038 47458 1090
rect 5182 926 5234 978
rect 7758 926 7810 978
rect 8094 926 8146 978
rect 10894 926 10946 978
rect 11566 926 11618 978
rect 15150 926 15202 978
rect 16270 926 16322 978
rect 20638 926 20690 978
rect 21310 926 21362 978
rect 22654 926 22706 978
rect 23326 926 23378 978
rect 25118 926 25170 978
rect 26462 926 26514 978
rect 27134 926 27186 978
rect 28366 926 28418 978
rect 30382 926 30434 978
rect 33742 926 33794 978
rect 34078 926 34130 978
rect 34414 926 34466 978
rect 35982 926 36034 978
rect 36654 926 36706 978
rect 37326 926 37378 978
rect 37998 926 38050 978
rect 39118 926 39170 978
rect 39790 926 39842 978
rect 43150 926 43202 978
rect 45054 926 45106 978
rect 46734 926 46786 978
rect 48302 926 48354 978
rect 48974 926 49026 978
rect 49646 926 49698 978
rect 50542 926 50594 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 672 57344 784 57456
rect 1120 57344 1232 57456
rect 1568 57344 1680 57456
rect 2016 57344 2128 57456
rect 2464 57344 2576 57456
rect 2912 57344 3024 57456
rect 3360 57344 3472 57456
rect 3808 57344 3920 57456
rect 4256 57344 4368 57456
rect 4704 57344 4816 57456
rect 5152 57344 5264 57456
rect 5600 57344 5712 57456
rect 6048 57344 6160 57456
rect 6496 57344 6608 57456
rect 6944 57344 7056 57456
rect 7392 57344 7504 57456
rect 7840 57344 7952 57456
rect 8288 57344 8400 57456
rect 8736 57344 8848 57456
rect 9184 57344 9296 57456
rect 9632 57344 9744 57456
rect 10080 57344 10192 57456
rect 10528 57344 10640 57456
rect 10976 57344 11088 57456
rect 11424 57344 11536 57456
rect 11872 57344 11984 57456
rect 12320 57344 12432 57456
rect 12768 57344 12880 57456
rect 13216 57344 13328 57456
rect 13664 57344 13776 57456
rect 14112 57344 14224 57456
rect 14560 57344 14672 57456
rect 15008 57344 15120 57456
rect 15456 57344 15568 57456
rect 15904 57344 16016 57456
rect 16352 57344 16464 57456
rect 16800 57344 16912 57456
rect 17248 57344 17360 57456
rect 17696 57344 17808 57456
rect 18144 57344 18256 57456
rect 18592 57344 18704 57456
rect 19040 57344 19152 57456
rect 19488 57344 19600 57456
rect 19936 57344 20048 57456
rect 20384 57344 20496 57456
rect 20832 57344 20944 57456
rect 21280 57344 21392 57456
rect 21728 57344 21840 57456
rect 22176 57344 22288 57456
rect 22624 57344 22736 57456
rect 23072 57344 23184 57456
rect 23520 57344 23632 57456
rect 23968 57344 24080 57456
rect 24416 57344 24528 57456
rect 24864 57344 24976 57456
rect 25312 57344 25424 57456
rect 25760 57344 25872 57456
rect 26208 57344 26320 57456
rect 26656 57344 26768 57456
rect 27104 57344 27216 57456
rect 27552 57344 27664 57456
rect 28000 57344 28112 57456
rect 28448 57344 28560 57456
rect 28896 57344 29008 57456
rect 29344 57344 29456 57456
rect 29792 57344 29904 57456
rect 30240 57344 30352 57456
rect 30688 57344 30800 57456
rect 31136 57344 31248 57456
rect 31584 57344 31696 57456
rect 32032 57344 32144 57456
rect 32480 57344 32592 57456
rect 32928 57344 33040 57456
rect 33376 57344 33488 57456
rect 33824 57344 33936 57456
rect 34272 57344 34384 57456
rect 34720 57344 34832 57456
rect 35168 57344 35280 57456
rect 35616 57344 35728 57456
rect 36064 57344 36176 57456
rect 36512 57344 36624 57456
rect 36960 57344 37072 57456
rect 37408 57344 37520 57456
rect 37856 57344 37968 57456
rect 38304 57344 38416 57456
rect 38752 57344 38864 57456
rect 39200 57344 39312 57456
rect 39648 57344 39760 57456
rect 40096 57344 40208 57456
rect 40544 57344 40656 57456
rect 40992 57344 41104 57456
rect 41440 57344 41552 57456
rect 41888 57344 42000 57456
rect 42336 57344 42448 57456
rect 42784 57344 42896 57456
rect 43232 57344 43344 57456
rect 43680 57344 43792 57456
rect 44128 57344 44240 57456
rect 44576 57344 44688 57456
rect 45024 57344 45136 57456
rect 45472 57344 45584 57456
rect 45920 57344 46032 57456
rect 46368 57344 46480 57456
rect 46816 57344 46928 57456
rect 47264 57344 47376 57456
rect 47712 57344 47824 57456
rect 48160 57344 48272 57456
rect 48608 57344 48720 57456
rect 49056 57344 49168 57456
rect 49504 57344 49616 57456
rect 49952 57344 50064 57456
rect 50400 57344 50512 57456
rect 50848 57344 50960 57456
rect 51296 57344 51408 57456
rect 51744 57344 51856 57456
rect 52192 57344 52304 57456
rect 52640 57344 52752 57456
rect 53088 57344 53200 57456
rect 53536 57344 53648 57456
rect 53984 57344 54096 57456
rect 54432 57344 54544 57456
rect 54880 57344 54992 57456
rect 55328 57344 55440 57456
rect 55776 57344 55888 57456
rect 56224 57344 56336 57456
rect 56672 57344 56784 57456
rect 588 56868 644 56878
rect 476 52724 532 52734
rect 140 51380 196 51390
rect 140 43988 196 51324
rect 140 43922 196 43932
rect 252 49588 308 49598
rect 140 43764 196 43774
rect 140 43316 196 43708
rect 252 43428 308 49532
rect 364 48244 420 48254
rect 364 46564 420 48188
rect 364 46498 420 46508
rect 364 43428 420 43438
rect 252 43372 364 43428
rect 364 43362 420 43372
rect 140 43260 308 43316
rect 140 43092 196 43102
rect 140 29428 196 43036
rect 252 39172 308 43260
rect 476 39172 532 52668
rect 588 50596 644 56812
rect 700 56756 756 57344
rect 700 56690 756 56700
rect 924 57204 980 57214
rect 700 55748 756 55758
rect 700 54180 756 55692
rect 924 54404 980 57148
rect 1148 55748 1204 57344
rect 1596 57092 1652 57344
rect 1596 57026 1652 57036
rect 1708 56980 1764 56990
rect 1148 55682 1204 55692
rect 1260 55858 1316 55870
rect 1260 55806 1262 55858
rect 1314 55806 1316 55858
rect 1260 55412 1316 55806
rect 1596 55858 1652 55870
rect 1596 55806 1598 55858
rect 1650 55806 1652 55858
rect 1596 55748 1652 55806
rect 1260 55346 1316 55356
rect 1372 55692 1652 55748
rect 924 54338 980 54348
rect 1260 55186 1316 55198
rect 1260 55134 1262 55186
rect 1314 55134 1316 55186
rect 700 54114 756 54124
rect 1148 54290 1204 54302
rect 1148 54238 1150 54290
rect 1202 54238 1204 54290
rect 1148 53956 1204 54238
rect 1148 53890 1204 53900
rect 1148 53730 1204 53742
rect 1148 53678 1150 53730
rect 1202 53678 1204 53730
rect 924 53620 980 53630
rect 812 53172 868 53182
rect 588 50530 644 50540
rect 700 50932 756 50942
rect 588 48804 644 48814
rect 588 43540 644 48748
rect 700 43652 756 50876
rect 700 43586 756 43596
rect 588 43474 644 43484
rect 476 39116 756 39172
rect 252 39106 308 39116
rect 476 38948 532 38958
rect 140 29362 196 29372
rect 252 38388 308 38398
rect 252 19012 308 38332
rect 252 18946 308 18956
rect 364 31892 420 31902
rect 252 18676 308 18686
rect 140 12852 196 12862
rect 28 12180 84 12190
rect 28 6244 84 12124
rect 140 7364 196 12796
rect 252 10276 308 18620
rect 364 18564 420 31836
rect 476 28420 532 38892
rect 700 38724 756 39116
rect 700 38658 756 38668
rect 700 34132 756 34142
rect 588 33012 644 33022
rect 588 30436 644 32956
rect 588 30370 644 30380
rect 700 29988 756 34076
rect 812 32340 868 53116
rect 924 32788 980 53564
rect 1036 52836 1092 52846
rect 1036 48692 1092 52780
rect 1148 52388 1204 53678
rect 1148 52322 1204 52332
rect 1260 53620 1316 55134
rect 1260 53058 1316 53564
rect 1260 53006 1262 53058
rect 1314 53006 1316 53058
rect 1260 52162 1316 53006
rect 1260 52110 1262 52162
rect 1314 52110 1316 52162
rect 1260 51378 1316 52110
rect 1372 52052 1428 55692
rect 1708 55636 1764 56924
rect 1484 55580 1764 55636
rect 1932 55858 1988 55870
rect 1932 55806 1934 55858
rect 1986 55806 1988 55858
rect 1484 54402 1540 55580
rect 1484 54350 1486 54402
rect 1538 54350 1540 54402
rect 1484 54338 1540 54350
rect 1708 55410 1764 55422
rect 1708 55358 1710 55410
rect 1762 55358 1764 55410
rect 1484 53842 1540 53854
rect 1484 53790 1486 53842
rect 1538 53790 1540 53842
rect 1484 52612 1540 53790
rect 1596 52836 1652 52846
rect 1596 52742 1652 52780
rect 1484 52546 1540 52556
rect 1596 52274 1652 52286
rect 1596 52222 1598 52274
rect 1650 52222 1652 52274
rect 1372 51996 1540 52052
rect 1260 51326 1262 51378
rect 1314 51326 1316 51378
rect 1260 51314 1316 51326
rect 1372 51378 1428 51390
rect 1372 51326 1374 51378
rect 1426 51326 1428 51378
rect 1260 51156 1316 51166
rect 1260 50482 1316 51100
rect 1260 50430 1262 50482
rect 1314 50430 1316 50482
rect 1260 49810 1316 50430
rect 1260 49758 1262 49810
rect 1314 49758 1316 49810
rect 1148 49252 1204 49262
rect 1148 49158 1204 49196
rect 1036 48626 1092 48636
rect 1148 48356 1204 48366
rect 1148 48262 1204 48300
rect 1260 47346 1316 49758
rect 1260 47294 1262 47346
rect 1314 47294 1316 47346
rect 1148 46788 1204 46798
rect 1036 45890 1092 45902
rect 1036 45838 1038 45890
rect 1090 45838 1092 45890
rect 1036 42868 1092 45838
rect 1148 45108 1204 46732
rect 1260 46786 1316 47294
rect 1372 47068 1428 51326
rect 1484 50820 1540 51996
rect 1484 50754 1540 50764
rect 1596 50706 1652 52222
rect 1708 51604 1764 55358
rect 1932 54740 1988 55806
rect 1932 54674 1988 54684
rect 1820 54292 1876 54302
rect 1820 54198 1876 54236
rect 1932 53732 1988 53742
rect 2044 53732 2100 57344
rect 2156 57204 2212 57214
rect 2156 54402 2212 57148
rect 2380 57204 2436 57214
rect 2380 56868 2436 57148
rect 2380 56802 2436 56812
rect 2380 56308 2436 56318
rect 2268 56196 2324 56206
rect 2268 55970 2324 56140
rect 2268 55918 2270 55970
rect 2322 55918 2324 55970
rect 2268 55906 2324 55918
rect 2156 54350 2158 54402
rect 2210 54350 2212 54402
rect 2156 54338 2212 54350
rect 2268 55524 2324 55534
rect 2156 53956 2212 53966
rect 2268 53956 2324 55468
rect 2156 53954 2324 53956
rect 2156 53902 2158 53954
rect 2210 53902 2324 53954
rect 2156 53900 2324 53902
rect 2156 53890 2212 53900
rect 2044 53676 2212 53732
rect 1932 53638 1988 53676
rect 2044 52276 2100 52286
rect 1708 51538 1764 51548
rect 1932 51940 1988 51950
rect 1820 51268 1876 51278
rect 1596 50654 1598 50706
rect 1650 50654 1652 50706
rect 1484 50596 1540 50606
rect 1484 49250 1540 50540
rect 1596 49924 1652 50654
rect 1596 49858 1652 49868
rect 1708 51212 1820 51268
rect 1596 49700 1652 49710
rect 1596 49606 1652 49644
rect 1484 49198 1486 49250
rect 1538 49198 1540 49250
rect 1484 49186 1540 49198
rect 1596 49364 1652 49374
rect 1484 48692 1540 48702
rect 1484 48020 1540 48636
rect 1596 48242 1652 49308
rect 1596 48190 1598 48242
rect 1650 48190 1652 48242
rect 1596 48178 1652 48190
rect 1596 48020 1652 48030
rect 1484 47964 1596 48020
rect 1596 47570 1652 47964
rect 1596 47518 1598 47570
rect 1650 47518 1652 47570
rect 1596 47506 1652 47518
rect 1708 47124 1764 51212
rect 1820 51174 1876 51212
rect 1820 50820 1876 50830
rect 1820 49250 1876 50764
rect 1932 49812 1988 51884
rect 1932 49746 1988 49756
rect 1820 49198 1822 49250
rect 1874 49198 1876 49250
rect 1820 49186 1876 49198
rect 1596 47068 1764 47124
rect 1820 48692 1876 48702
rect 1372 47012 1540 47068
rect 1260 46734 1262 46786
rect 1314 46734 1316 46786
rect 1260 45298 1316 46734
rect 1372 46116 1428 46126
rect 1372 46022 1428 46060
rect 1260 45242 1428 45298
rect 1260 45108 1316 45118
rect 1148 45106 1316 45108
rect 1148 45054 1262 45106
rect 1314 45054 1316 45106
rect 1148 45052 1316 45054
rect 1260 44996 1316 45052
rect 1260 44930 1316 44940
rect 1372 42980 1428 45242
rect 1036 42802 1092 42812
rect 1260 42924 1428 42980
rect 1484 44210 1540 47012
rect 1596 46564 1652 47068
rect 1596 46470 1652 46508
rect 1484 44158 1486 44210
rect 1538 44158 1540 44210
rect 1484 43538 1540 44158
rect 1484 43486 1486 43538
rect 1538 43486 1540 43538
rect 1260 42308 1316 42924
rect 1260 42242 1316 42252
rect 1372 42644 1428 42654
rect 1484 42644 1540 43486
rect 1708 45890 1764 45902
rect 1708 45838 1710 45890
rect 1762 45838 1764 45890
rect 1372 42642 1540 42644
rect 1372 42590 1374 42642
rect 1426 42590 1540 42642
rect 1372 42588 1540 42590
rect 1596 43428 1652 43438
rect 1260 41972 1316 41982
rect 1372 41972 1428 42588
rect 1260 41970 1428 41972
rect 1260 41918 1262 41970
rect 1314 41918 1428 41970
rect 1260 41916 1428 41918
rect 1484 42308 1540 42318
rect 1036 41524 1092 41534
rect 1036 39842 1092 41468
rect 1148 40962 1204 40974
rect 1148 40910 1150 40962
rect 1202 40910 1204 40962
rect 1148 40516 1204 40910
rect 1148 40450 1204 40460
rect 1148 40292 1204 40302
rect 1148 40198 1204 40236
rect 1260 40068 1316 41916
rect 1036 39790 1038 39842
rect 1090 39790 1092 39842
rect 1036 39778 1092 39790
rect 1148 40012 1316 40068
rect 1372 40068 1428 40078
rect 924 32722 980 32732
rect 1036 34356 1092 34366
rect 1036 32676 1092 34300
rect 1148 33572 1204 40012
rect 1372 39842 1428 40012
rect 1372 39790 1374 39842
rect 1426 39790 1428 39842
rect 1372 39778 1428 39790
rect 1260 38948 1316 38958
rect 1260 38854 1316 38892
rect 1260 38052 1316 38062
rect 1484 38052 1540 42252
rect 1596 41860 1652 43372
rect 1708 41972 1764 45838
rect 1820 44996 1876 48636
rect 1820 44930 1876 44940
rect 1932 48242 1988 48254
rect 1932 48190 1934 48242
rect 1986 48190 1988 48242
rect 1932 47124 1988 48190
rect 1932 44548 1988 47068
rect 2044 46340 2100 52220
rect 2156 51828 2212 53676
rect 2380 53396 2436 56252
rect 2492 54404 2548 57344
rect 2940 56084 2996 57344
rect 2940 56018 2996 56028
rect 3052 56868 3108 56878
rect 2604 55858 2660 55870
rect 2604 55806 2606 55858
rect 2658 55806 2660 55858
rect 2604 54628 2660 55806
rect 2940 55860 2996 55870
rect 3052 55860 3108 56812
rect 3388 56420 3444 57344
rect 3388 56354 3444 56364
rect 3612 56756 3668 56766
rect 3612 56196 3668 56700
rect 3836 56644 3892 57344
rect 4284 57204 4340 57344
rect 4284 57138 4340 57148
rect 3836 56588 4340 56644
rect 4284 56532 4340 56588
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4284 56466 4340 56476
rect 3804 56410 4068 56420
rect 4172 56420 4228 56430
rect 3612 56140 3780 56196
rect 2940 55858 3108 55860
rect 2940 55806 2942 55858
rect 2994 55806 3108 55858
rect 2940 55804 3108 55806
rect 3388 56082 3444 56094
rect 3388 56030 3390 56082
rect 3442 56030 3444 56082
rect 3388 55860 3444 56030
rect 3612 55972 3668 55982
rect 3724 55972 3780 56140
rect 3612 55970 3780 55972
rect 3612 55918 3614 55970
rect 3666 55918 3780 55970
rect 3612 55916 3780 55918
rect 3948 55972 4004 55982
rect 3612 55906 3668 55916
rect 3948 55878 4004 55916
rect 3500 55860 3556 55870
rect 3388 55804 3500 55860
rect 2940 55794 2996 55804
rect 3500 55794 3556 55804
rect 3388 55410 3444 55422
rect 3388 55358 3390 55410
rect 3442 55358 3444 55410
rect 3164 55300 3220 55310
rect 3052 55298 3220 55300
rect 3052 55246 3166 55298
rect 3218 55246 3220 55298
rect 3052 55244 3220 55246
rect 2604 54562 2660 54572
rect 2828 55074 2884 55086
rect 2828 55022 2830 55074
rect 2882 55022 2884 55074
rect 2716 54516 2772 54526
rect 2716 54422 2772 54460
rect 2492 54348 2660 54404
rect 2156 51762 2212 51772
rect 2268 53340 2436 53396
rect 2492 53842 2548 53854
rect 2492 53790 2494 53842
rect 2546 53790 2548 53842
rect 2156 49252 2212 49262
rect 2268 49252 2324 53340
rect 2156 49250 2324 49252
rect 2156 49198 2158 49250
rect 2210 49198 2324 49250
rect 2156 49196 2324 49198
rect 2492 49252 2548 53790
rect 2604 52052 2660 54348
rect 2716 53730 2772 53742
rect 2716 53678 2718 53730
rect 2770 53678 2772 53730
rect 2716 52276 2772 53678
rect 2828 53172 2884 55022
rect 2828 53106 2884 53116
rect 2940 54404 2996 54414
rect 2940 52948 2996 54348
rect 2940 52882 2996 52892
rect 2716 52210 2772 52220
rect 2828 52722 2884 52734
rect 2828 52670 2830 52722
rect 2882 52670 2884 52722
rect 2828 52164 2884 52670
rect 2940 52724 2996 52734
rect 2940 52276 2996 52668
rect 2940 52210 2996 52220
rect 2828 52098 2884 52108
rect 2604 51986 2660 51996
rect 2828 51938 2884 51950
rect 2828 51886 2830 51938
rect 2882 51886 2884 51938
rect 2828 50932 2884 51886
rect 2940 51156 2996 51166
rect 2940 51062 2996 51100
rect 2828 50866 2884 50876
rect 3052 50708 3108 55244
rect 3164 55234 3220 55244
rect 3276 55188 3332 55198
rect 3276 54516 3332 55132
rect 3388 55076 3444 55358
rect 3500 55412 3556 55422
rect 3500 55318 3556 55356
rect 4060 55188 4116 55198
rect 4060 55094 4116 55132
rect 3388 55010 3444 55020
rect 3804 54908 4068 54918
rect 3164 54404 3220 54414
rect 3164 54310 3220 54348
rect 3276 53956 3332 54460
rect 3164 53900 3332 53956
rect 3388 54852 3444 54862
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 3164 53844 3220 53900
rect 3388 53844 3444 54796
rect 4172 54292 4228 56364
rect 4732 56308 4788 57344
rect 4732 56242 4788 56252
rect 5068 56532 5124 56542
rect 4844 55970 4900 55982
rect 4844 55918 4846 55970
rect 4898 55918 4900 55970
rect 4284 55858 4340 55870
rect 4284 55806 4286 55858
rect 4338 55806 4340 55858
rect 4284 54852 4340 55806
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 4508 55524 4564 55534
rect 4508 55410 4564 55468
rect 4508 55358 4510 55410
rect 4562 55358 4564 55410
rect 4508 55300 4564 55358
rect 4508 55234 4564 55244
rect 4844 55076 4900 55918
rect 4956 55858 5012 55870
rect 4956 55806 4958 55858
rect 5010 55806 5012 55858
rect 4956 55636 5012 55806
rect 4956 55570 5012 55580
rect 4844 55010 4900 55020
rect 4956 55412 5012 55422
rect 4284 54786 4340 54796
rect 4284 54516 4340 54526
rect 4284 54422 4340 54460
rect 3164 53778 3220 53788
rect 3276 53788 3444 53844
rect 3500 54236 4228 54292
rect 3276 53508 3332 53788
rect 3164 53452 3332 53508
rect 3388 53618 3444 53630
rect 3388 53566 3390 53618
rect 3442 53566 3444 53618
rect 3388 53508 3444 53566
rect 3164 51940 3220 53452
rect 3388 53442 3444 53452
rect 3276 53172 3332 53182
rect 3276 52500 3332 53116
rect 3500 53060 3556 54236
rect 4464 54124 4728 54134
rect 3724 54068 3780 54078
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3612 53844 3668 53854
rect 3612 53172 3668 53788
rect 3724 53842 3780 54012
rect 4060 53956 4116 53966
rect 4116 53900 4228 53956
rect 4060 53890 4116 53900
rect 3724 53790 3726 53842
rect 3778 53790 3780 53842
rect 3724 53778 3780 53790
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 4172 53172 4228 53900
rect 4956 53732 5012 55356
rect 5068 55188 5124 56476
rect 5068 55122 5124 55132
rect 5068 54290 5124 54302
rect 5068 54238 5070 54290
rect 5122 54238 5124 54290
rect 5068 53956 5124 54238
rect 5068 53890 5124 53900
rect 5180 53844 5236 57344
rect 5628 56084 5684 57344
rect 5628 56018 5684 56028
rect 5740 57092 5796 57102
rect 5292 55858 5348 55870
rect 5292 55806 5294 55858
rect 5346 55806 5348 55858
rect 5292 55076 5348 55806
rect 5628 55860 5684 55870
rect 5740 55860 5796 57036
rect 6076 56308 6132 57344
rect 6076 56242 6132 56252
rect 6300 56084 6356 56094
rect 6300 55970 6356 56028
rect 6300 55918 6302 55970
rect 6354 55918 6356 55970
rect 6300 55906 6356 55918
rect 5964 55860 6020 55870
rect 5628 55858 5796 55860
rect 5628 55806 5630 55858
rect 5682 55806 5796 55858
rect 5628 55804 5796 55806
rect 5852 55858 6020 55860
rect 5852 55806 5966 55858
rect 6018 55806 6020 55858
rect 5852 55804 6020 55806
rect 5628 55794 5684 55804
rect 5628 55076 5684 55086
rect 5292 55010 5348 55020
rect 5516 55074 5684 55076
rect 5516 55022 5630 55074
rect 5682 55022 5684 55074
rect 5516 55020 5684 55022
rect 5404 54290 5460 54302
rect 5404 54238 5406 54290
rect 5458 54238 5460 54290
rect 5292 54180 5348 54190
rect 5292 53844 5348 54124
rect 5404 54068 5460 54238
rect 5404 54002 5460 54012
rect 5292 53788 5460 53844
rect 5180 53778 5236 53788
rect 4956 53676 5124 53732
rect 3612 53116 3892 53172
rect 3500 53004 3780 53060
rect 3724 52834 3780 53004
rect 3724 52782 3726 52834
rect 3778 52782 3780 52834
rect 3724 52770 3780 52782
rect 3388 52724 3444 52734
rect 3388 52630 3444 52668
rect 3276 52434 3332 52444
rect 3500 52612 3556 52622
rect 3500 52386 3556 52556
rect 3500 52334 3502 52386
rect 3554 52334 3556 52386
rect 3500 52322 3556 52334
rect 3612 52500 3668 52510
rect 3164 51874 3220 51884
rect 3612 51380 3668 52444
rect 3836 52386 3892 53116
rect 4060 53116 4228 53172
rect 4956 53506 5012 53518
rect 4956 53454 4958 53506
rect 5010 53454 5012 53506
rect 4060 52834 4116 53116
rect 4956 52948 5012 53454
rect 4956 52882 5012 52892
rect 4060 52782 4062 52834
rect 4114 52782 4116 52834
rect 4060 52770 4116 52782
rect 4172 52836 4228 52846
rect 3836 52334 3838 52386
rect 3890 52334 3892 52386
rect 3836 52322 3892 52334
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 3836 51604 3892 51614
rect 4172 51604 4228 52780
rect 4396 52724 4452 52762
rect 4396 52658 4452 52668
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4464 52490 4728 52500
rect 4732 52276 4788 52286
rect 4732 52182 4788 52220
rect 4284 52162 4340 52174
rect 4284 52110 4286 52162
rect 4338 52110 4340 52162
rect 4284 51940 4340 52110
rect 4284 51874 4340 51884
rect 4396 52052 4452 52062
rect 3836 51602 4228 51604
rect 3836 51550 3838 51602
rect 3890 51550 4228 51602
rect 3836 51548 4228 51550
rect 3836 51538 3892 51548
rect 4396 51490 4452 51996
rect 4396 51438 4398 51490
rect 4450 51438 4452 51490
rect 4396 51426 4452 51438
rect 4172 51380 4228 51390
rect 3612 51324 4004 51380
rect 3388 51266 3444 51278
rect 3388 51214 3390 51266
rect 3442 51214 3444 51266
rect 3388 51156 3444 51214
rect 3388 51090 3444 51100
rect 3500 51154 3556 51166
rect 3500 51102 3502 51154
rect 3554 51102 3556 51154
rect 3500 50932 3556 51102
rect 3500 50866 3556 50876
rect 2156 49186 2212 49196
rect 2492 49186 2548 49196
rect 2604 50652 3108 50708
rect 2268 49028 2324 49038
rect 2156 48580 2212 48590
rect 2156 48130 2212 48524
rect 2156 48078 2158 48130
rect 2210 48078 2212 48130
rect 2156 48066 2212 48078
rect 2044 46274 2100 46284
rect 2044 46004 2100 46014
rect 2044 45910 2100 45948
rect 2268 45444 2324 48972
rect 2492 48916 2548 48926
rect 2492 48822 2548 48860
rect 2492 46676 2548 46686
rect 2268 45378 2324 45388
rect 2380 45890 2436 45902
rect 2380 45838 2382 45890
rect 2434 45838 2436 45890
rect 2156 45108 2212 45118
rect 1932 44482 1988 44492
rect 2044 45106 2212 45108
rect 2044 45054 2158 45106
rect 2210 45054 2212 45106
rect 2044 45052 2212 45054
rect 1820 44436 1876 44474
rect 1820 44370 1876 44380
rect 2044 44324 2100 45052
rect 2156 45042 2212 45052
rect 2268 45108 2324 45118
rect 2044 44258 2100 44268
rect 2156 44548 2212 44558
rect 1820 44212 1876 44222
rect 1876 44156 1988 44212
rect 1820 44146 1876 44156
rect 1820 43428 1876 43438
rect 1820 42980 1876 43372
rect 1820 42886 1876 42924
rect 1932 42644 1988 44156
rect 1932 42578 1988 42588
rect 2044 43652 2100 43662
rect 2044 43314 2100 43596
rect 2044 43262 2046 43314
rect 2098 43262 2100 43314
rect 1708 41906 1764 41916
rect 1596 41766 1652 41804
rect 1708 41076 1764 41086
rect 1596 40404 1652 40414
rect 1596 40310 1652 40348
rect 1708 39842 1764 41020
rect 1932 40740 1988 40750
rect 1932 40404 1988 40684
rect 1708 39790 1710 39842
rect 1762 39790 1764 39842
rect 1708 39778 1764 39790
rect 1820 40402 1988 40404
rect 1820 40350 1934 40402
rect 1986 40350 1988 40402
rect 1820 40348 1988 40350
rect 1708 38724 1764 38762
rect 1708 38658 1764 38668
rect 1820 38500 1876 40348
rect 1932 40338 1988 40348
rect 2044 40180 2100 43262
rect 2156 40740 2212 44492
rect 2268 42980 2324 45052
rect 2268 42914 2324 42924
rect 2380 42420 2436 45838
rect 2380 42354 2436 42364
rect 2492 41860 2548 46620
rect 2604 45332 2660 50652
rect 3500 50594 3556 50606
rect 3500 50542 3502 50594
rect 3554 50542 3556 50594
rect 2828 50484 2884 50522
rect 2828 50418 2884 50428
rect 3052 50036 3108 50046
rect 3052 49812 3108 49980
rect 3500 49924 3556 50542
rect 3836 50594 3892 50606
rect 3836 50542 3838 50594
rect 3890 50542 3892 50594
rect 3612 50482 3668 50494
rect 3612 50430 3614 50482
rect 3666 50430 3668 50482
rect 3612 50036 3668 50430
rect 3836 50428 3892 50542
rect 3948 50594 4004 51324
rect 4172 51286 4228 51324
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 4732 50706 4788 50718
rect 4732 50654 4734 50706
rect 4786 50654 4788 50706
rect 3948 50542 3950 50594
rect 4002 50542 4004 50594
rect 3948 50530 4004 50542
rect 4508 50594 4564 50606
rect 4508 50542 4510 50594
rect 4562 50542 4564 50594
rect 4508 50484 4564 50542
rect 3836 50372 4228 50428
rect 4508 50418 4564 50428
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 3612 49980 3780 50036
rect 3500 49868 3668 49924
rect 3164 49812 3220 49822
rect 3052 49810 3220 49812
rect 3052 49758 3166 49810
rect 3218 49758 3220 49810
rect 3052 49756 3220 49758
rect 3164 49746 3220 49756
rect 3500 49700 3556 49710
rect 3500 49606 3556 49644
rect 2828 49586 2884 49598
rect 2828 49534 2830 49586
rect 2882 49534 2884 49586
rect 2828 49252 2884 49534
rect 3164 49588 3220 49598
rect 2828 49186 2884 49196
rect 2940 49364 2996 49374
rect 2940 49028 2996 49308
rect 2940 49026 3108 49028
rect 2940 48974 2942 49026
rect 2994 48974 3108 49026
rect 2940 48972 3108 48974
rect 2940 48962 2996 48972
rect 2940 48804 2996 48814
rect 2940 48356 2996 48748
rect 2716 48244 2772 48254
rect 2716 48150 2772 48188
rect 2828 47684 2884 47694
rect 2828 47590 2884 47628
rect 2828 46450 2884 46462
rect 2828 46398 2830 46450
rect 2882 46398 2884 46450
rect 2716 46002 2772 46014
rect 2716 45950 2718 46002
rect 2770 45950 2772 46002
rect 2716 45780 2772 45950
rect 2716 45714 2772 45724
rect 2828 45892 2884 46398
rect 2604 45266 2660 45276
rect 2716 45444 2772 45454
rect 2604 44996 2660 45006
rect 2604 43092 2660 44940
rect 2604 43026 2660 43036
rect 2716 42868 2772 45388
rect 2828 45106 2884 45836
rect 2828 45054 2830 45106
rect 2882 45054 2884 45106
rect 2828 45042 2884 45054
rect 2940 46004 2996 48300
rect 3052 48244 3108 48972
rect 3164 48468 3220 49532
rect 3388 49588 3444 49598
rect 3388 49494 3444 49532
rect 3500 49252 3556 49262
rect 3612 49252 3668 49868
rect 3500 49250 3668 49252
rect 3500 49198 3502 49250
rect 3554 49198 3668 49250
rect 3500 49196 3668 49198
rect 3500 49186 3556 49196
rect 3388 49026 3444 49038
rect 3388 48974 3390 49026
rect 3442 48974 3444 49026
rect 3388 48692 3444 48974
rect 3164 48412 3332 48468
rect 3052 47460 3108 48188
rect 3052 47394 3108 47404
rect 3164 48242 3220 48254
rect 3164 48190 3166 48242
rect 3218 48190 3220 48242
rect 3164 48020 3220 48190
rect 3052 47124 3108 47134
rect 3052 46228 3108 47068
rect 3164 46676 3220 47964
rect 3164 46610 3220 46620
rect 3276 46562 3332 48412
rect 3388 48356 3444 48636
rect 3388 48290 3444 48300
rect 3500 49028 3556 49038
rect 3388 47908 3444 47918
rect 3388 47682 3444 47852
rect 3388 47630 3390 47682
rect 3442 47630 3444 47682
rect 3388 47618 3444 47630
rect 3276 46510 3278 46562
rect 3330 46510 3332 46562
rect 3052 46162 3108 46172
rect 3164 46452 3220 46462
rect 3052 46004 3108 46014
rect 2940 46002 3108 46004
rect 2940 45950 3054 46002
rect 3106 45950 3108 46002
rect 2940 45948 3108 45950
rect 2940 43204 2996 45948
rect 3052 45938 3108 45948
rect 3164 45668 3220 46396
rect 3052 45612 3220 45668
rect 3052 44884 3108 45612
rect 3164 45444 3220 45454
rect 3164 44996 3220 45388
rect 3164 44930 3220 44940
rect 3052 44818 3108 44828
rect 2940 43138 2996 43148
rect 3052 44100 3108 44110
rect 3276 44100 3332 46510
rect 3388 46564 3444 46574
rect 3500 46564 3556 48972
rect 3724 48804 3780 49980
rect 3612 48748 3780 48804
rect 3836 49698 3892 49710
rect 3836 49646 3838 49698
rect 3890 49646 3892 49698
rect 3836 48804 3892 49646
rect 4172 49698 4228 50372
rect 4732 50260 4788 50654
rect 5068 50428 5124 53676
rect 5292 52836 5348 52846
rect 5292 52742 5348 52780
rect 5404 52500 5460 53788
rect 5516 52834 5572 55020
rect 5628 55010 5684 55020
rect 5852 54740 5908 55804
rect 5964 55794 6020 55804
rect 5740 54684 5908 54740
rect 5964 55524 6020 55534
rect 5628 53620 5684 53630
rect 5628 53526 5684 53564
rect 5740 53396 5796 54684
rect 5964 54628 6020 55468
rect 6524 55524 6580 57344
rect 6972 56196 7028 57344
rect 7420 56420 7476 57344
rect 7420 56354 7476 56364
rect 7868 56420 7924 57344
rect 7868 56354 7924 56364
rect 6860 56140 7028 56196
rect 8092 56194 8148 56206
rect 8092 56142 8094 56194
rect 8146 56142 8148 56194
rect 6748 56082 6804 56094
rect 6748 56030 6750 56082
rect 6802 56030 6804 56082
rect 6748 55636 6804 56030
rect 6748 55570 6804 55580
rect 6524 55458 6580 55468
rect 6188 55412 6244 55422
rect 6188 55410 6356 55412
rect 6188 55358 6190 55410
rect 6242 55358 6356 55410
rect 6188 55356 6356 55358
rect 6188 55346 6244 55356
rect 6076 55300 6132 55310
rect 6076 55206 6132 55244
rect 5964 54572 6132 54628
rect 5740 53330 5796 53340
rect 5852 54514 5908 54526
rect 5852 54462 5854 54514
rect 5906 54462 5908 54514
rect 5852 53060 5908 54462
rect 5964 54404 6020 54414
rect 5964 54310 6020 54348
rect 6076 53954 6132 54572
rect 6076 53902 6078 53954
rect 6130 53902 6132 53954
rect 6076 53890 6132 53902
rect 6188 54290 6244 54302
rect 6188 54238 6190 54290
rect 6242 54238 6244 54290
rect 6188 53284 6244 54238
rect 6076 53228 6244 53284
rect 5516 52782 5518 52834
rect 5570 52782 5572 52834
rect 5516 52612 5572 52782
rect 5740 53004 6020 53060
rect 5516 52546 5572 52556
rect 5628 52722 5684 52734
rect 5628 52670 5630 52722
rect 5682 52670 5684 52722
rect 5404 52434 5460 52444
rect 5628 51940 5684 52670
rect 5404 51884 5684 51940
rect 5404 51378 5460 51884
rect 5404 51326 5406 51378
rect 5458 51326 5460 51378
rect 5404 51314 5460 51326
rect 5516 51380 5572 51390
rect 5740 51380 5796 53004
rect 5516 51378 5796 51380
rect 5516 51326 5518 51378
rect 5570 51326 5796 51378
rect 5516 51324 5796 51326
rect 5852 52834 5908 52846
rect 5852 52782 5854 52834
rect 5906 52782 5908 52834
rect 5516 51314 5572 51324
rect 5628 51156 5684 51166
rect 5628 51062 5684 51100
rect 5740 51154 5796 51166
rect 5740 51102 5742 51154
rect 5794 51102 5796 51154
rect 5628 50708 5684 50718
rect 5292 50596 5348 50606
rect 5292 50594 5460 50596
rect 5292 50542 5294 50594
rect 5346 50542 5460 50594
rect 5292 50540 5460 50542
rect 5292 50530 5348 50540
rect 5068 50372 5348 50428
rect 4732 50194 4788 50204
rect 5068 50036 5124 50046
rect 4396 49812 4452 49822
rect 4396 49718 4452 49756
rect 4172 49646 4174 49698
rect 4226 49646 4228 49698
rect 4060 49586 4116 49598
rect 4060 49534 4062 49586
rect 4114 49534 4116 49586
rect 3948 49476 4004 49486
rect 3948 49138 4004 49420
rect 4060 49364 4116 49534
rect 4172 49588 4228 49646
rect 4172 49522 4228 49532
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 4060 49298 4116 49308
rect 3948 49086 3950 49138
rect 4002 49086 4004 49138
rect 3948 49028 4004 49086
rect 3948 48962 4004 48972
rect 4508 49026 4564 49038
rect 4508 48974 4510 49026
rect 4562 48974 4564 49026
rect 3612 46676 3668 48748
rect 3836 48738 3892 48748
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 4172 48580 4228 48590
rect 4172 48237 4228 48524
rect 4508 48468 4564 48974
rect 4508 48402 4564 48412
rect 4956 48468 5012 48478
rect 4956 48354 5012 48412
rect 4956 48302 4958 48354
rect 5010 48302 5012 48354
rect 4956 48290 5012 48302
rect 4172 48185 4174 48237
rect 4226 48185 4228 48237
rect 4172 48173 4228 48185
rect 5068 48020 5124 49980
rect 4172 47964 5012 48020
rect 4172 47908 4228 47964
rect 4956 47908 5012 47964
rect 5068 47954 5124 47964
rect 5180 49698 5236 49710
rect 5180 49646 5182 49698
rect 5234 49646 5236 49698
rect 4172 47842 4228 47852
rect 4464 47852 4728 47862
rect 4284 47796 4340 47806
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4956 47842 5012 47852
rect 4464 47786 4728 47796
rect 3724 47570 3780 47582
rect 3724 47518 3726 47570
rect 3778 47518 3780 47570
rect 3724 47236 3780 47518
rect 4060 47348 4116 47358
rect 4060 47346 4228 47348
rect 4060 47294 4062 47346
rect 4114 47294 4228 47346
rect 4060 47292 4228 47294
rect 4060 47282 4116 47292
rect 3724 47170 3780 47180
rect 4172 47124 4228 47292
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4172 47058 4228 47068
rect 3804 47002 4068 47012
rect 3836 46676 3892 46686
rect 3612 46674 3892 46676
rect 3612 46622 3838 46674
rect 3890 46622 3892 46674
rect 3612 46620 3892 46622
rect 3836 46610 3892 46620
rect 4284 46674 4340 47740
rect 4620 47684 4676 47694
rect 4396 47460 4452 47470
rect 4396 47366 4452 47404
rect 4620 47068 4676 47628
rect 5068 47572 5124 47582
rect 5068 47478 5124 47516
rect 4956 47458 5012 47470
rect 4956 47406 4958 47458
rect 5010 47406 5012 47458
rect 4956 47348 5012 47406
rect 5180 47460 5236 49646
rect 5292 48468 5348 50372
rect 5404 49476 5460 50540
rect 5628 49810 5684 50652
rect 5740 50428 5796 51102
rect 5852 51156 5908 52782
rect 5964 52386 6020 53004
rect 5964 52334 5966 52386
rect 6018 52334 6020 52386
rect 5964 52322 6020 52334
rect 5964 51380 6020 51390
rect 6076 51380 6132 53228
rect 6188 53060 6244 53070
rect 6188 52966 6244 53004
rect 6300 51828 6356 55356
rect 6412 55298 6468 55310
rect 6412 55246 6414 55298
rect 6466 55246 6468 55298
rect 6412 54964 6468 55246
rect 6412 54898 6468 54908
rect 6524 55300 6580 55310
rect 6300 51762 6356 51772
rect 6412 54514 6468 54526
rect 6412 54462 6414 54514
rect 6466 54462 6468 54514
rect 5964 51378 6132 51380
rect 5964 51326 5966 51378
rect 6018 51326 6132 51378
rect 5964 51324 6132 51326
rect 5964 51314 6020 51324
rect 6300 51266 6356 51278
rect 6300 51214 6302 51266
rect 6354 51214 6356 51266
rect 5852 51100 6244 51156
rect 6076 50594 6132 50606
rect 6076 50542 6078 50594
rect 6130 50542 6132 50594
rect 5740 50372 5908 50428
rect 5628 49758 5630 49810
rect 5682 49758 5684 49810
rect 5628 49746 5684 49758
rect 5404 49410 5460 49420
rect 5404 49252 5460 49262
rect 5404 48692 5460 49196
rect 5516 49026 5572 49038
rect 5516 48974 5518 49026
rect 5570 48974 5572 49026
rect 5516 48916 5572 48974
rect 5516 48850 5572 48860
rect 5628 49028 5684 49038
rect 5404 48636 5572 48692
rect 5292 48412 5460 48468
rect 5292 48244 5348 48254
rect 5292 48150 5348 48188
rect 5180 47394 5236 47404
rect 4956 47292 5124 47348
rect 4956 47124 5012 47134
rect 5068 47124 5124 47292
rect 5180 47124 5236 47134
rect 5068 47068 5180 47124
rect 4620 47012 4900 47068
rect 4284 46622 4286 46674
rect 4338 46622 4340 46674
rect 4284 46610 4340 46622
rect 3948 46564 4004 46574
rect 3500 46508 3780 46564
rect 3388 46470 3444 46508
rect 3388 45890 3444 45902
rect 3388 45838 3390 45890
rect 3442 45838 3444 45890
rect 3388 45668 3444 45838
rect 3724 45668 3780 46508
rect 3948 46470 4004 46508
rect 4060 46450 4116 46462
rect 4060 46398 4062 46450
rect 4114 46398 4116 46450
rect 4060 46340 4116 46398
rect 3836 46228 3892 46238
rect 4060 46228 4116 46284
rect 3836 45890 3892 46172
rect 3836 45838 3838 45890
rect 3890 45838 3892 45890
rect 3836 45826 3892 45838
rect 3948 46172 4116 46228
rect 4172 46450 4228 46462
rect 4172 46398 4174 46450
rect 4226 46398 4228 46450
rect 3388 45602 3444 45612
rect 3668 45612 3780 45668
rect 3948 45668 4004 46172
rect 4060 46004 4116 46014
rect 4060 45910 4116 45948
rect 3500 45332 3556 45342
rect 3668 45332 3724 45612
rect 3948 45602 4004 45612
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 4172 45444 4228 46398
rect 4284 46452 4340 46462
rect 4284 46116 4340 46396
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 4844 46116 4900 47012
rect 4284 46060 4564 46116
rect 4508 46002 4564 46060
rect 4508 45950 4510 46002
rect 4562 45950 4564 46002
rect 4508 45938 4564 45950
rect 4620 46060 4900 46116
rect 4620 45780 4676 46060
rect 4732 45892 4788 45902
rect 4732 45890 4900 45892
rect 4732 45838 4734 45890
rect 4786 45838 4900 45890
rect 4732 45836 4900 45838
rect 4732 45826 4788 45836
rect 4172 45378 4228 45388
rect 4284 45724 4676 45780
rect 3668 45276 3780 45332
rect 3500 45106 3556 45276
rect 3500 45054 3502 45106
rect 3554 45054 3556 45106
rect 3500 45042 3556 45054
rect 3388 44996 3444 45006
rect 3388 44902 3444 44940
rect 3052 44098 3332 44100
rect 3052 44046 3054 44098
rect 3106 44046 3332 44098
rect 3052 44044 3332 44046
rect 3500 44884 3556 44894
rect 2716 42802 2772 42812
rect 2940 42532 2996 42542
rect 2492 41794 2548 41804
rect 2604 42530 2996 42532
rect 2604 42478 2942 42530
rect 2994 42478 2996 42530
rect 2604 42476 2996 42478
rect 2268 41524 2324 41534
rect 2268 41410 2324 41468
rect 2268 41358 2270 41410
rect 2322 41358 2324 41410
rect 2268 41346 2324 41358
rect 2604 41188 2660 42476
rect 2940 42466 2996 42476
rect 3052 42308 3108 44044
rect 2940 42252 3108 42308
rect 3164 43652 3220 43662
rect 2156 40674 2212 40684
rect 2380 40964 2436 40974
rect 1708 38444 1876 38500
rect 1932 40124 2100 40180
rect 2156 40178 2212 40190
rect 2156 40126 2158 40178
rect 2210 40126 2212 40178
rect 1596 38164 1652 38174
rect 1596 38070 1652 38108
rect 1260 38050 1540 38052
rect 1260 37998 1262 38050
rect 1314 37998 1540 38050
rect 1260 37996 1540 37998
rect 1260 36482 1316 37996
rect 1372 37268 1428 37278
rect 1708 37268 1764 38444
rect 1932 38388 1988 40124
rect 2044 39844 2100 39854
rect 2044 39750 2100 39788
rect 2156 38836 2212 40126
rect 2380 39730 2436 40908
rect 2604 40402 2660 41132
rect 2716 41748 2772 41758
rect 2716 41186 2772 41692
rect 2716 41134 2718 41186
rect 2770 41134 2772 41186
rect 2716 41122 2772 41134
rect 2828 41746 2884 41758
rect 2828 41694 2830 41746
rect 2882 41694 2884 41746
rect 2604 40350 2606 40402
rect 2658 40350 2660 40402
rect 2604 39956 2660 40350
rect 2828 41076 2884 41694
rect 2828 40404 2884 41020
rect 2828 40338 2884 40348
rect 2604 39890 2660 39900
rect 2716 40180 2772 40190
rect 2940 40180 2996 42252
rect 3164 42084 3220 43596
rect 3388 43204 3444 43214
rect 3164 42018 3220 42028
rect 3276 42756 3332 42766
rect 3276 41970 3332 42700
rect 3388 42642 3444 43148
rect 3388 42590 3390 42642
rect 3442 42590 3444 42642
rect 3388 42532 3444 42590
rect 3388 42466 3444 42476
rect 3276 41918 3278 41970
rect 3330 41918 3332 41970
rect 3276 41906 3332 41918
rect 3500 41972 3556 44828
rect 3724 44322 3780 45276
rect 3948 45108 4004 45118
rect 3948 45014 4004 45052
rect 4284 44996 4340 45724
rect 4396 45332 4452 45342
rect 4396 45218 4452 45276
rect 4396 45166 4398 45218
rect 4450 45166 4452 45218
rect 4396 45154 4452 45166
rect 4620 45332 4676 45342
rect 4060 44940 4340 44996
rect 4060 44884 4116 44940
rect 4620 44884 4676 45276
rect 3724 44270 3726 44322
rect 3778 44270 3780 44322
rect 3724 44258 3780 44270
rect 3948 44828 4116 44884
rect 4284 44828 4676 44884
rect 3948 44322 4004 44828
rect 3948 44270 3950 44322
rect 4002 44270 4004 44322
rect 3948 44258 4004 44270
rect 4172 44772 4228 44782
rect 4060 44210 4116 44222
rect 4060 44158 4062 44210
rect 4114 44158 4116 44210
rect 4060 44100 4116 44158
rect 3612 44044 4116 44100
rect 3612 43538 3668 44044
rect 4172 43988 4228 44716
rect 4284 44660 4340 44828
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4284 44604 4396 44660
rect 4464 44650 4728 44660
rect 4340 44578 4396 44604
rect 4340 44522 4564 44578
rect 4508 44434 4564 44522
rect 4508 44382 4510 44434
rect 4562 44382 4564 44434
rect 4508 44370 4564 44382
rect 4284 44324 4340 44334
rect 4284 44322 4452 44324
rect 4284 44270 4286 44322
rect 4338 44270 4452 44322
rect 4284 44268 4452 44270
rect 4284 44258 4340 44268
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4172 43922 4228 43932
rect 3804 43866 4068 43876
rect 3612 43486 3614 43538
rect 3666 43486 3668 43538
rect 3612 43474 3668 43486
rect 4060 43540 4116 43550
rect 4060 43446 4116 43484
rect 4284 43540 4340 43550
rect 4284 43446 4340 43484
rect 3836 43316 3892 43326
rect 3164 41860 3220 41870
rect 2716 39842 2772 40124
rect 2716 39790 2718 39842
rect 2770 39790 2772 39842
rect 2716 39778 2772 39790
rect 2828 40124 2996 40180
rect 3052 41748 3108 41758
rect 2380 39678 2382 39730
rect 2434 39678 2436 39730
rect 2380 39666 2436 39678
rect 2492 39732 2548 39742
rect 2492 39730 2660 39732
rect 2492 39678 2494 39730
rect 2546 39678 2660 39730
rect 2492 39676 2660 39678
rect 2492 39666 2548 39676
rect 2604 39620 2660 39676
rect 2828 39620 2884 40124
rect 2604 39564 2884 39620
rect 2156 38770 2212 38780
rect 2380 39508 2436 39518
rect 2940 39508 2996 39518
rect 2380 38668 2436 39452
rect 1372 37266 1764 37268
rect 1372 37214 1374 37266
rect 1426 37214 1764 37266
rect 1372 37212 1764 37214
rect 1372 37202 1428 37212
rect 1596 36820 1652 36830
rect 1596 36594 1652 36764
rect 1596 36542 1598 36594
rect 1650 36542 1652 36594
rect 1596 36530 1652 36542
rect 1260 36430 1262 36482
rect 1314 36430 1316 36482
rect 1260 35308 1316 36430
rect 1484 36260 1540 36270
rect 1484 35693 1540 36204
rect 1484 35641 1486 35693
rect 1538 35641 1540 35693
rect 1260 35252 1428 35308
rect 1260 34804 1316 34814
rect 1372 34804 1428 35252
rect 1260 34802 1428 34804
rect 1260 34750 1262 34802
rect 1314 34750 1428 34802
rect 1260 34748 1428 34750
rect 1260 34132 1316 34748
rect 1260 34038 1316 34076
rect 1372 33572 1428 33582
rect 1148 33516 1316 33572
rect 1036 32610 1092 32620
rect 1148 33346 1204 33358
rect 1148 33294 1150 33346
rect 1202 33294 1204 33346
rect 812 32274 868 32284
rect 924 32564 980 32574
rect 812 32116 868 32126
rect 812 30100 868 32060
rect 924 31220 980 32508
rect 1148 32564 1204 33294
rect 1148 32498 1204 32508
rect 1260 32674 1316 33516
rect 1372 33478 1428 33516
rect 1484 33012 1540 35641
rect 1708 35364 1764 37212
rect 1708 35298 1764 35308
rect 1820 38332 1988 38388
rect 2268 38612 2436 38668
rect 2716 39506 2996 39508
rect 2716 39454 2942 39506
rect 2994 39454 2996 39506
rect 2716 39452 2996 39454
rect 1596 35026 1652 35038
rect 1596 34974 1598 35026
rect 1650 34974 1652 35026
rect 1596 34916 1652 34974
rect 1820 34916 1876 38332
rect 2156 37268 2212 37278
rect 1596 34860 1876 34916
rect 1708 33908 1764 33918
rect 1708 33814 1764 33852
rect 1820 33684 1876 34860
rect 1820 33618 1876 33628
rect 1932 37266 2212 37268
rect 1932 37214 2158 37266
rect 2210 37214 2212 37266
rect 1932 37212 2212 37214
rect 1820 33346 1876 33358
rect 1820 33294 1822 33346
rect 1874 33294 1876 33346
rect 1820 33124 1876 33294
rect 1820 33058 1876 33068
rect 1484 32946 1540 32956
rect 1260 32622 1262 32674
rect 1314 32622 1316 32674
rect 924 31154 980 31164
rect 1260 31778 1316 32622
rect 1484 32788 1540 32798
rect 1260 31726 1262 31778
rect 1314 31726 1316 31778
rect 1260 30210 1316 31726
rect 1372 32340 1428 32350
rect 1372 31332 1428 32284
rect 1484 31556 1540 32732
rect 1708 32452 1764 32462
rect 1708 32358 1764 32396
rect 1596 32340 1652 32350
rect 1596 31890 1652 32284
rect 1596 31838 1598 31890
rect 1650 31838 1652 31890
rect 1596 31826 1652 31838
rect 1484 31500 1652 31556
rect 1372 31276 1540 31332
rect 1260 30158 1262 30210
rect 1314 30158 1316 30210
rect 812 30044 980 30100
rect 700 29932 868 29988
rect 476 28354 532 28364
rect 700 29764 756 29774
rect 588 22932 644 22942
rect 364 18498 420 18508
rect 476 21588 532 21598
rect 476 16772 532 21532
rect 588 16884 644 22876
rect 700 22260 756 29708
rect 812 25732 868 29932
rect 812 25666 868 25676
rect 700 22194 756 22204
rect 812 25508 868 25518
rect 812 22036 868 25452
rect 924 23268 980 30044
rect 1260 29538 1316 30158
rect 1260 29486 1262 29538
rect 1314 29486 1316 29538
rect 1260 29474 1316 29486
rect 1372 30994 1428 31006
rect 1372 30942 1374 30994
rect 1426 30942 1428 30994
rect 1260 28532 1316 28542
rect 1148 28530 1316 28532
rect 1148 28478 1262 28530
rect 1314 28478 1316 28530
rect 1148 28476 1316 28478
rect 924 23202 980 23212
rect 1036 28420 1092 28430
rect 1036 27076 1092 28364
rect 1036 23156 1092 27020
rect 1148 27074 1204 28476
rect 1260 28466 1316 28476
rect 1372 27860 1428 30942
rect 1372 27766 1428 27804
rect 1484 27636 1540 31276
rect 1596 30322 1652 31500
rect 1596 30270 1598 30322
rect 1650 30270 1652 30322
rect 1596 29540 1652 30270
rect 1932 29540 1988 37212
rect 2156 37202 2212 37212
rect 2156 36820 2212 36830
rect 2044 33460 2100 33470
rect 2044 33366 2100 33404
rect 1596 29484 1764 29540
rect 1148 27022 1150 27074
rect 1202 27022 1204 27074
rect 1148 26908 1204 27022
rect 1372 27580 1540 27636
rect 1596 29316 1652 29326
rect 1596 28754 1652 29260
rect 1596 28702 1598 28754
rect 1650 28702 1652 28754
rect 1148 26852 1316 26908
rect 1260 26290 1316 26852
rect 1260 26238 1262 26290
rect 1314 26238 1316 26290
rect 1260 25508 1316 26238
rect 1372 26068 1428 27580
rect 1596 27524 1652 28702
rect 1596 27458 1652 27468
rect 1708 27298 1764 29484
rect 1932 29474 1988 29484
rect 2044 33012 2100 33022
rect 1708 27246 1710 27298
rect 1762 27246 1764 27298
rect 1708 27188 1764 27246
rect 1708 27122 1764 27132
rect 1372 26002 1428 26012
rect 1708 26068 1764 26078
rect 1260 25414 1316 25452
rect 1484 24722 1540 24734
rect 1484 24670 1486 24722
rect 1538 24670 1540 24722
rect 1148 24612 1204 24622
rect 1148 24518 1204 24556
rect 1260 23156 1316 23166
rect 1036 23154 1316 23156
rect 1036 23102 1262 23154
rect 1314 23102 1316 23154
rect 1036 23100 1316 23102
rect 700 21980 868 22036
rect 1148 22370 1204 22382
rect 1148 22318 1150 22370
rect 1202 22318 1204 22370
rect 700 18900 756 21980
rect 1036 21364 1092 21374
rect 1036 21270 1092 21308
rect 812 20916 868 20926
rect 812 19572 868 20860
rect 1148 20020 1204 22318
rect 1260 20802 1316 23100
rect 1372 22482 1428 22494
rect 1372 22430 1374 22482
rect 1426 22430 1428 22482
rect 1372 21700 1428 22430
rect 1372 21634 1428 21644
rect 1372 21476 1428 21486
rect 1372 21382 1428 21420
rect 1260 20750 1262 20802
rect 1314 20750 1316 20802
rect 1260 20244 1316 20750
rect 1260 20178 1316 20188
rect 1372 21140 1428 21150
rect 1148 19964 1316 20020
rect 1148 19796 1204 19806
rect 1148 19702 1204 19740
rect 812 19516 1092 19572
rect 700 18834 756 18844
rect 812 19124 868 19134
rect 588 16818 644 16828
rect 476 16706 532 16716
rect 588 16436 644 16446
rect 252 10210 308 10220
rect 364 14420 420 14430
rect 252 7364 308 7374
rect 140 7308 252 7364
rect 252 7298 308 7308
rect 364 7252 420 14364
rect 476 9268 532 9278
rect 476 8596 532 9212
rect 588 8708 644 16380
rect 700 14644 756 14654
rect 700 11172 756 14588
rect 700 11106 756 11116
rect 812 8932 868 19068
rect 1036 18338 1092 19516
rect 1260 18788 1316 19964
rect 1036 18286 1038 18338
rect 1090 18286 1092 18338
rect 1036 18274 1092 18286
rect 1148 18732 1316 18788
rect 924 18228 980 18238
rect 924 13636 980 18172
rect 1148 15538 1204 18732
rect 1372 18452 1428 21084
rect 1484 19796 1540 24670
rect 1708 24164 1764 26012
rect 1820 25732 1876 25742
rect 1820 25638 1876 25676
rect 1932 24724 1988 24734
rect 1820 24722 1988 24724
rect 1820 24670 1934 24722
rect 1986 24670 1988 24722
rect 1820 24668 1988 24670
rect 1820 24388 1876 24668
rect 1932 24658 1988 24668
rect 1820 24322 1876 24332
rect 1708 24108 1876 24164
rect 1708 23938 1764 23950
rect 1708 23886 1710 23938
rect 1762 23886 1764 23938
rect 1708 23828 1764 23886
rect 1708 23762 1764 23772
rect 1484 19730 1540 19740
rect 1596 23716 1652 23726
rect 1484 19348 1540 19358
rect 1484 19254 1540 19292
rect 1260 18396 1428 18452
rect 1260 16772 1316 18396
rect 1372 18228 1428 18266
rect 1372 18162 1428 18172
rect 1372 17666 1428 17678
rect 1372 17614 1374 17666
rect 1426 17614 1428 17666
rect 1372 17556 1428 17614
rect 1372 17490 1428 17500
rect 1260 16706 1316 16716
rect 1372 16324 1428 16334
rect 1260 16100 1316 16110
rect 1260 16006 1316 16044
rect 1148 15486 1150 15538
rect 1202 15486 1204 15538
rect 1148 15474 1204 15486
rect 1260 15764 1316 15774
rect 1148 14532 1204 14542
rect 1148 14438 1204 14476
rect 1036 14420 1092 14430
rect 1036 14326 1092 14364
rect 1260 13972 1316 15708
rect 1148 13916 1316 13972
rect 1036 13636 1092 13646
rect 924 13634 1092 13636
rect 924 13582 1038 13634
rect 1090 13582 1092 13634
rect 924 13580 1092 13582
rect 1036 13570 1092 13580
rect 1148 13186 1204 13916
rect 1372 13748 1428 16268
rect 1596 16210 1652 23660
rect 1820 22930 1876 24108
rect 1820 22878 1822 22930
rect 1874 22878 1876 22930
rect 1708 21476 1764 21486
rect 1708 21382 1764 21420
rect 1820 21364 1876 22878
rect 1932 22372 1988 22382
rect 1932 22278 1988 22316
rect 2044 21588 2100 32956
rect 2156 27860 2212 36764
rect 2156 27794 2212 27804
rect 2268 25172 2324 38612
rect 2380 38500 2436 38510
rect 2380 35698 2436 38444
rect 2492 38052 2548 38062
rect 2492 36260 2548 37996
rect 2716 37828 2772 39452
rect 2940 39442 2996 39452
rect 2828 38612 2884 38622
rect 2828 38610 2996 38612
rect 2828 38558 2830 38610
rect 2882 38558 2996 38610
rect 2828 38556 2996 38558
rect 2828 38546 2884 38556
rect 2716 36820 2772 37772
rect 2828 37826 2884 37838
rect 2828 37774 2830 37826
rect 2882 37774 2884 37826
rect 2828 37156 2884 37774
rect 2940 37266 2996 38556
rect 2940 37214 2942 37266
rect 2994 37214 2996 37266
rect 2940 37202 2996 37214
rect 3052 37268 3108 41692
rect 3164 40402 3220 41804
rect 3388 41860 3444 41870
rect 3388 41766 3444 41804
rect 3500 41636 3556 41916
rect 3612 43314 3892 43316
rect 3612 43262 3838 43314
rect 3890 43262 3892 43314
rect 3612 43260 3892 43262
rect 3612 41970 3668 43260
rect 3836 43250 3892 43260
rect 3948 43314 4004 43326
rect 4396 43316 4452 44268
rect 3948 43262 3950 43314
rect 4002 43262 4004 43314
rect 3724 43092 3780 43102
rect 3724 42754 3780 43036
rect 3724 42702 3726 42754
rect 3778 42702 3780 42754
rect 3724 42690 3780 42702
rect 3948 42532 4004 43262
rect 4284 43260 4452 43316
rect 4844 44322 4900 45836
rect 4956 45556 5012 47068
rect 5180 47058 5236 47068
rect 5068 46676 5124 46686
rect 5068 45890 5124 46620
rect 5068 45838 5070 45890
rect 5122 45838 5124 45890
rect 5068 45826 5124 45838
rect 5292 46674 5348 46686
rect 5292 46622 5294 46674
rect 5346 46622 5348 46674
rect 4956 45490 5012 45500
rect 5292 45556 5348 46622
rect 5292 45490 5348 45500
rect 5180 45444 5236 45454
rect 4956 44996 5012 45006
rect 4956 44902 5012 44940
rect 5068 44884 5124 44894
rect 5068 44790 5124 44828
rect 4844 44270 4846 44322
rect 4898 44270 4900 44322
rect 4284 42980 4340 43260
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 4396 42980 4452 42990
rect 4284 42978 4452 42980
rect 4284 42926 4398 42978
rect 4450 42926 4452 42978
rect 4284 42924 4452 42926
rect 4396 42914 4452 42924
rect 4844 42866 4900 44270
rect 4844 42814 4846 42866
rect 4898 42814 4900 42866
rect 4844 42802 4900 42814
rect 4956 44772 5012 44782
rect 4284 42756 4340 42766
rect 3948 42466 4004 42476
rect 4172 42700 4284 42756
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 3612 41918 3614 41970
rect 3666 41918 3668 41970
rect 3612 41906 3668 41918
rect 3724 41970 3780 41982
rect 3724 41918 3726 41970
rect 3778 41918 3780 41970
rect 3164 40350 3166 40402
rect 3218 40350 3220 40402
rect 3164 39508 3220 40350
rect 3276 41580 3556 41636
rect 3276 39956 3332 41580
rect 3276 39890 3332 39900
rect 3388 41076 3444 41086
rect 3388 39732 3444 41020
rect 3500 41074 3556 41086
rect 3500 41022 3502 41074
rect 3554 41022 3556 41074
rect 3500 40852 3556 41022
rect 3724 40964 3780 41918
rect 4060 41972 4116 41982
rect 4060 41878 4116 41916
rect 4060 41746 4116 41758
rect 4060 41694 4062 41746
rect 4114 41694 4116 41746
rect 3836 41186 3892 41198
rect 3836 41134 3838 41186
rect 3890 41134 3892 41186
rect 3836 41076 3892 41134
rect 4060 41076 4116 41694
rect 4172 41188 4228 42700
rect 4284 42662 4340 42700
rect 4284 42084 4340 42094
rect 4284 41970 4340 42028
rect 4284 41918 4286 41970
rect 4338 41918 4340 41970
rect 4284 41906 4340 41918
rect 4284 41692 4900 41748
rect 4284 41636 4340 41692
rect 4284 41570 4340 41580
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 4508 41300 4564 41310
rect 4508 41206 4564 41244
rect 4844 41300 4900 41692
rect 4844 41234 4900 41244
rect 4284 41188 4340 41198
rect 4172 41186 4340 41188
rect 4172 41134 4286 41186
rect 4338 41134 4340 41186
rect 4172 41132 4340 41134
rect 4284 41076 4340 41132
rect 4956 41076 5012 44716
rect 5180 44548 5236 45388
rect 5292 45220 5348 45230
rect 5292 45106 5348 45164
rect 5292 45054 5294 45106
rect 5346 45054 5348 45106
rect 5292 45042 5348 45054
rect 5068 44492 5236 44548
rect 5292 44660 5348 44670
rect 5068 41524 5124 44492
rect 5180 44324 5236 44334
rect 5180 43650 5236 44268
rect 5292 44322 5348 44604
rect 5404 44548 5460 48412
rect 5516 45106 5572 48636
rect 5628 48468 5684 48972
rect 5628 47458 5684 48412
rect 5740 48242 5796 48254
rect 5740 48190 5742 48242
rect 5794 48190 5796 48242
rect 5740 47796 5796 48190
rect 5740 47730 5796 47740
rect 5628 47406 5630 47458
rect 5682 47406 5684 47458
rect 5628 47394 5684 47406
rect 5516 45054 5518 45106
rect 5570 45054 5572 45106
rect 5516 45042 5572 45054
rect 5628 47236 5684 47246
rect 5516 44548 5572 44558
rect 5404 44546 5572 44548
rect 5404 44494 5518 44546
rect 5570 44494 5572 44546
rect 5404 44492 5572 44494
rect 5516 44482 5572 44492
rect 5292 44270 5294 44322
rect 5346 44270 5348 44322
rect 5292 44258 5348 44270
rect 5404 44212 5460 44222
rect 5180 43598 5182 43650
rect 5234 43598 5236 43650
rect 5180 43586 5236 43598
rect 5292 43876 5348 43886
rect 5292 43428 5348 43820
rect 5068 41458 5124 41468
rect 5180 43372 5348 43428
rect 4060 41020 4228 41076
rect 3836 41010 3892 41020
rect 3500 40786 3556 40796
rect 3612 40908 3780 40964
rect 3612 40628 3668 40908
rect 4172 40852 4228 41020
rect 4284 41010 4340 41020
rect 4396 41020 5012 41076
rect 4396 40852 4452 41020
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4172 40786 4228 40796
rect 4284 40796 4452 40852
rect 4732 40852 4788 40862
rect 4956 40852 5012 41020
rect 4788 40796 4900 40852
rect 3804 40730 4068 40740
rect 4284 40628 4340 40796
rect 4732 40786 4788 40796
rect 3612 40572 4004 40628
rect 3276 39676 3444 39732
rect 3500 40516 3556 40526
rect 3276 39620 3332 39676
rect 3276 39526 3332 39564
rect 3164 39442 3220 39452
rect 3388 39508 3444 39518
rect 3276 38948 3332 38958
rect 3276 38834 3332 38892
rect 3276 38782 3278 38834
rect 3330 38782 3332 38834
rect 3276 38770 3332 38782
rect 3388 38722 3444 39452
rect 3388 38670 3390 38722
rect 3442 38670 3444 38722
rect 3388 38658 3444 38670
rect 3500 37716 3556 40460
rect 3948 39842 4004 40572
rect 4172 40572 4340 40628
rect 4172 40402 4228 40572
rect 4172 40350 4174 40402
rect 4226 40350 4228 40402
rect 4172 40338 4228 40350
rect 4284 40404 4340 40414
rect 4844 40404 4900 40796
rect 4956 40786 5012 40796
rect 5068 41188 5124 41198
rect 4956 40404 5012 40414
rect 4844 40402 5012 40404
rect 4844 40350 4958 40402
rect 5010 40350 5012 40402
rect 4844 40348 5012 40350
rect 3948 39790 3950 39842
rect 4002 39790 4004 39842
rect 3948 39778 4004 39790
rect 4172 39956 4228 39966
rect 3724 39620 3780 39630
rect 3612 39618 3780 39620
rect 3612 39566 3726 39618
rect 3778 39566 3780 39618
rect 3612 39564 3780 39566
rect 3612 38836 3668 39564
rect 3724 39554 3780 39564
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 3836 38836 3892 38874
rect 3612 38780 3780 38836
rect 3612 38610 3668 38622
rect 3612 38558 3614 38610
rect 3666 38558 3668 38610
rect 3612 38388 3668 38558
rect 3612 38322 3668 38332
rect 3612 38052 3668 38062
rect 3612 37958 3668 37996
rect 3724 37828 3780 38780
rect 3836 38770 3892 38780
rect 4060 38836 4116 38846
rect 4060 38610 4116 38780
rect 4172 38834 4228 39900
rect 4172 38782 4174 38834
rect 4226 38782 4228 38834
rect 4172 38770 4228 38782
rect 4284 38836 4340 40348
rect 4956 40338 5012 40348
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 5068 39844 5124 41132
rect 5180 40290 5236 43372
rect 5404 42754 5460 44156
rect 5404 42702 5406 42754
rect 5458 42702 5460 42754
rect 5292 41860 5348 41870
rect 5292 41766 5348 41804
rect 5404 41188 5460 42702
rect 5516 43538 5572 43550
rect 5516 43486 5518 43538
rect 5570 43486 5572 43538
rect 5516 42196 5572 43486
rect 5628 42196 5684 47180
rect 5740 46452 5796 46462
rect 5740 46358 5796 46396
rect 5852 45556 5908 50372
rect 5964 49810 6020 49822
rect 5964 49758 5966 49810
rect 6018 49758 6020 49810
rect 5964 48804 6020 49758
rect 5964 48738 6020 48748
rect 6076 49700 6132 50542
rect 5964 48132 6020 48142
rect 5964 48038 6020 48076
rect 5964 47796 6020 47806
rect 5964 47236 6020 47740
rect 5964 47170 6020 47180
rect 5964 47012 6020 47022
rect 5964 46788 6020 46956
rect 5964 46722 6020 46732
rect 6076 46004 6132 49644
rect 6188 49698 6244 51100
rect 6300 50820 6356 51214
rect 6412 51268 6468 54462
rect 6524 53172 6580 55244
rect 6636 55298 6692 55310
rect 6636 55246 6638 55298
rect 6690 55246 6692 55298
rect 6636 54290 6692 55246
rect 6636 54238 6638 54290
rect 6690 54238 6692 54290
rect 6636 54180 6692 54238
rect 6636 54114 6692 54124
rect 6860 53284 6916 56140
rect 7420 56082 7476 56094
rect 7420 56030 7422 56082
rect 7474 56030 7476 56082
rect 6972 55860 7028 55870
rect 6972 55766 7028 55804
rect 7308 55636 7364 55646
rect 7308 55522 7364 55580
rect 7308 55470 7310 55522
rect 7362 55470 7364 55522
rect 7308 55458 7364 55470
rect 6972 55412 7028 55422
rect 6972 55318 7028 55356
rect 6860 53218 6916 53228
rect 6972 55188 7028 55198
rect 6524 53116 6692 53172
rect 6524 52948 6580 52958
rect 6524 52854 6580 52892
rect 6636 52724 6692 53116
rect 6412 51202 6468 51212
rect 6524 52668 6692 52724
rect 6748 52948 6804 52958
rect 6300 50754 6356 50764
rect 6188 49646 6190 49698
rect 6242 49646 6244 49698
rect 6188 49634 6244 49646
rect 6300 50148 6356 50158
rect 6188 47796 6244 47806
rect 6188 47458 6244 47740
rect 6188 47406 6190 47458
rect 6242 47406 6244 47458
rect 6188 47394 6244 47406
rect 6076 45938 6132 45948
rect 6188 47012 6244 47022
rect 6188 45890 6244 46956
rect 6188 45838 6190 45890
rect 6242 45838 6244 45890
rect 5852 45500 6132 45556
rect 5964 44994 6020 45006
rect 5964 44942 5966 44994
rect 6018 44942 6020 44994
rect 5852 44884 5908 44894
rect 5740 44882 5908 44884
rect 5740 44830 5854 44882
rect 5906 44830 5908 44882
rect 5740 44828 5908 44830
rect 5740 42420 5796 44828
rect 5852 44818 5908 44828
rect 5740 42354 5796 42364
rect 5852 44660 5908 44670
rect 5628 42140 5796 42196
rect 5516 42130 5572 42140
rect 5628 41972 5684 41982
rect 5628 41858 5684 41916
rect 5628 41806 5630 41858
rect 5682 41806 5684 41858
rect 5628 41794 5684 41806
rect 5628 41524 5684 41534
rect 5516 41188 5572 41198
rect 5404 41132 5516 41188
rect 5516 41094 5572 41132
rect 5404 40740 5460 40750
rect 5404 40514 5460 40684
rect 5404 40462 5406 40514
rect 5458 40462 5460 40514
rect 5404 40450 5460 40462
rect 5516 40404 5572 40414
rect 5516 40310 5572 40348
rect 5180 40238 5182 40290
rect 5234 40238 5236 40290
rect 5180 40226 5236 40238
rect 5404 40180 5460 40190
rect 5404 40086 5460 40124
rect 5628 40180 5684 41468
rect 5628 40114 5684 40124
rect 5740 39956 5796 42140
rect 5852 42194 5908 44604
rect 5964 43764 6020 44942
rect 5964 43698 6020 43708
rect 5852 42142 5854 42194
rect 5906 42142 5908 42194
rect 5852 42130 5908 42142
rect 5964 42756 6020 42766
rect 4620 39788 5124 39844
rect 5292 39900 5796 39956
rect 4620 39618 4676 39788
rect 4956 39620 5012 39630
rect 4620 39566 4622 39618
rect 4674 39566 4676 39618
rect 4620 39554 4676 39566
rect 4844 39618 5012 39620
rect 4844 39566 4958 39618
rect 5010 39566 5012 39618
rect 4844 39564 5012 39566
rect 4284 38770 4340 38780
rect 4396 39172 4452 39182
rect 4396 38834 4452 39116
rect 4396 38782 4398 38834
rect 4450 38782 4452 38834
rect 4396 38770 4452 38782
rect 4732 38724 4788 38734
rect 4844 38724 4900 39564
rect 4956 39554 5012 39564
rect 5180 39620 5236 39630
rect 5068 38836 5124 38846
rect 4788 38668 4900 38724
rect 4732 38658 4788 38668
rect 4060 38558 4062 38610
rect 4114 38558 4116 38610
rect 4060 38546 4116 38558
rect 4844 38500 4900 38668
rect 4956 38724 5012 38734
rect 4956 38630 5012 38668
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4844 38434 4900 38444
rect 4464 38378 4728 38388
rect 3948 38276 4004 38286
rect 5068 38276 5124 38780
rect 3948 38050 4004 38220
rect 4956 38220 5124 38276
rect 4620 38164 4676 38174
rect 4956 38164 5012 38220
rect 4620 38162 5012 38164
rect 4620 38110 4622 38162
rect 4674 38110 5012 38162
rect 4620 38108 5012 38110
rect 4620 38098 4676 38108
rect 3948 37998 3950 38050
rect 4002 37998 4004 38050
rect 3948 37986 4004 37998
rect 4508 38050 4564 38062
rect 4508 37998 4510 38050
rect 4562 37998 4564 38050
rect 4508 37940 4564 37998
rect 5068 38052 5124 38062
rect 4508 37884 5012 37940
rect 4396 37828 4452 37838
rect 3724 37772 4228 37828
rect 3500 37660 3668 37716
rect 3388 37604 3444 37614
rect 3444 37548 3556 37604
rect 3388 37538 3444 37548
rect 3052 37212 3444 37268
rect 2828 37090 2884 37100
rect 3388 37154 3444 37212
rect 3500 37266 3556 37548
rect 3500 37214 3502 37266
rect 3554 37214 3556 37266
rect 3500 37202 3556 37214
rect 3612 37268 3668 37660
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 3948 37268 4004 37278
rect 3612 37266 4004 37268
rect 3612 37214 3950 37266
rect 4002 37214 4004 37266
rect 3612 37212 4004 37214
rect 3948 37202 4004 37212
rect 3388 37102 3390 37154
rect 3442 37102 3444 37154
rect 3388 37090 3444 37102
rect 3668 37044 3724 37054
rect 3724 36988 3780 37044
rect 3668 36978 3780 36988
rect 2716 36754 2772 36764
rect 3724 36606 3780 36978
rect 4172 36708 4228 37772
rect 4452 37772 4676 37828
rect 4396 37762 4452 37772
rect 4396 37156 4452 37166
rect 4396 37062 4452 37100
rect 4620 37156 4676 37772
rect 4956 37716 5012 37884
rect 4956 37650 5012 37660
rect 5068 37558 5124 37996
rect 5180 38050 5236 39564
rect 5292 38834 5348 39900
rect 5292 38782 5294 38834
rect 5346 38782 5348 38834
rect 5292 38770 5348 38782
rect 5404 39172 5460 39182
rect 5180 37998 5182 38050
rect 5234 37998 5236 38050
rect 5180 37986 5236 37998
rect 4956 37502 5124 37558
rect 5180 37604 5236 37614
rect 4956 37156 5012 37502
rect 5068 37380 5124 37390
rect 5068 37266 5124 37324
rect 5068 37214 5070 37266
rect 5122 37214 5124 37266
rect 5068 37202 5124 37214
rect 4620 37090 4676 37100
rect 4900 37100 5012 37156
rect 4900 36932 4956 37100
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 4844 36876 4956 36932
rect 5068 37044 5124 37054
rect 3948 36652 4228 36708
rect 3724 36596 3836 36606
rect 3500 36594 3836 36596
rect 3500 36542 3782 36594
rect 3834 36542 3836 36594
rect 3500 36540 3836 36542
rect 2492 36194 2548 36204
rect 2828 36484 2884 36494
rect 2380 35646 2382 35698
rect 2434 35646 2436 35698
rect 2380 35634 2436 35646
rect 2828 35698 2884 36428
rect 2828 35646 2830 35698
rect 2882 35646 2884 35698
rect 2828 35634 2884 35646
rect 2940 36372 2996 36382
rect 2380 35476 2436 35486
rect 2380 33458 2436 35420
rect 2604 35252 2660 35262
rect 2604 34244 2660 35196
rect 2828 35028 2884 35038
rect 2828 34934 2884 34972
rect 2604 34178 2660 34188
rect 2716 34916 2772 34926
rect 2380 33406 2382 33458
rect 2434 33406 2436 33458
rect 2380 33394 2436 33406
rect 2492 33570 2548 33582
rect 2492 33518 2494 33570
rect 2546 33518 2548 33570
rect 2492 33460 2548 33518
rect 2716 33570 2772 34860
rect 2716 33518 2718 33570
rect 2770 33518 2772 33570
rect 2716 33506 2772 33518
rect 2828 33906 2884 33918
rect 2828 33854 2830 33906
rect 2882 33854 2884 33906
rect 2492 33394 2548 33404
rect 2828 33460 2884 33854
rect 2828 33394 2884 33404
rect 2940 33234 2996 36316
rect 3276 36372 3332 36382
rect 3276 36278 3332 36316
rect 3500 35924 3556 36540
rect 3780 36530 3836 36540
rect 3948 36372 4004 36652
rect 4284 36596 4340 36606
rect 4172 36594 4340 36596
rect 4172 36542 4286 36594
rect 4338 36542 4340 36594
rect 4172 36540 4340 36542
rect 3500 35858 3556 35868
rect 3612 36316 4004 36372
rect 4060 36482 4116 36494
rect 4060 36430 4062 36482
rect 4114 36430 4116 36482
rect 4060 36372 4116 36430
rect 3612 35698 3668 36316
rect 4060 36306 4116 36316
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 3612 35646 3614 35698
rect 3666 35646 3668 35698
rect 3388 35474 3444 35486
rect 3388 35422 3390 35474
rect 3442 35422 3444 35474
rect 3388 35308 3444 35422
rect 3388 35252 3556 35308
rect 3500 35140 3556 35252
rect 3612 35218 3668 35646
rect 3948 35924 4004 35934
rect 3948 35698 4004 35868
rect 3948 35646 3950 35698
rect 4002 35646 4004 35698
rect 3948 35634 4004 35646
rect 3836 35588 3892 35598
rect 3836 35364 3892 35532
rect 3724 35252 3780 35262
rect 3612 35196 3724 35218
rect 3612 35162 3780 35196
rect 3500 35074 3556 35084
rect 3388 35028 3444 35038
rect 3052 35026 3444 35028
rect 3052 34974 3390 35026
rect 3442 34974 3444 35026
rect 3052 34972 3444 34974
rect 3052 34132 3108 34972
rect 3388 34962 3444 34972
rect 3500 34916 3556 34954
rect 3500 34850 3556 34860
rect 3612 34914 3668 34926
rect 3612 34862 3614 34914
rect 3666 34862 3668 34914
rect 3612 34692 3668 34862
rect 3724 34916 3780 34926
rect 3724 34822 3780 34860
rect 3052 34066 3108 34076
rect 3500 34636 3668 34692
rect 3724 34692 3780 34702
rect 3836 34692 3892 35308
rect 3780 34636 3892 34692
rect 3948 34914 4004 34926
rect 3948 34862 3950 34914
rect 4002 34862 4004 34914
rect 3948 34692 4004 34862
rect 3276 34020 3332 34030
rect 3164 34018 3332 34020
rect 3164 33966 3278 34018
rect 3330 33966 3332 34018
rect 3164 33964 3332 33966
rect 3164 33572 3220 33964
rect 3276 33954 3332 33964
rect 3388 33906 3444 33918
rect 3388 33854 3390 33906
rect 3442 33854 3444 33906
rect 3388 33572 3444 33854
rect 3500 33796 3556 34636
rect 3724 34626 3780 34636
rect 3948 34626 4004 34636
rect 3804 34524 4068 34534
rect 3612 34468 3668 34478
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 3612 34356 3668 34412
rect 4172 34356 4228 36540
rect 4284 36530 4340 36540
rect 4732 36484 4788 36494
rect 4732 36390 4788 36428
rect 4508 36372 4564 36382
rect 4396 36148 4452 36158
rect 4284 35924 4340 35934
rect 4284 35140 4340 35868
rect 4396 35810 4452 36092
rect 4396 35758 4398 35810
rect 4450 35758 4452 35810
rect 4396 35746 4452 35758
rect 4508 36036 4564 36316
rect 4508 35588 4564 35980
rect 4508 35522 4564 35532
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4844 35308 4900 36876
rect 5068 36148 5124 36988
rect 5068 36082 5124 36092
rect 4956 35812 5012 35822
rect 4956 35718 5012 35756
rect 4844 35252 5012 35308
rect 4464 35242 4728 35252
rect 4844 35140 4900 35150
rect 4284 35084 4676 35140
rect 4620 34914 4676 35084
rect 4620 34862 4622 34914
rect 4674 34862 4676 34914
rect 4620 34850 4676 34862
rect 4284 34804 4340 34814
rect 4284 34802 4452 34804
rect 4284 34750 4286 34802
rect 4338 34750 4452 34802
rect 4284 34748 4452 34750
rect 4284 34738 4340 34748
rect 3612 34300 3780 34356
rect 3500 33730 3556 33740
rect 3612 33906 3668 33918
rect 3612 33854 3614 33906
rect 3666 33854 3668 33906
rect 3164 33506 3220 33516
rect 3276 33516 3444 33572
rect 2940 33182 2942 33234
rect 2994 33182 2996 33234
rect 2604 32788 2660 32798
rect 2380 30994 2436 31006
rect 2380 30942 2382 30994
rect 2434 30942 2436 30994
rect 2380 28084 2436 30942
rect 2604 29316 2660 32732
rect 2940 32564 2996 33182
rect 3276 33124 3332 33516
rect 3388 33348 3444 33358
rect 3388 33346 3556 33348
rect 3388 33294 3390 33346
rect 3442 33294 3556 33346
rect 3388 33292 3556 33294
rect 3388 33282 3444 33292
rect 3276 33068 3444 33124
rect 2716 32508 2996 32564
rect 2716 30324 2772 32508
rect 3276 32452 3332 32462
rect 3164 32450 3332 32452
rect 3164 32398 3278 32450
rect 3330 32398 3332 32450
rect 3164 32396 3332 32398
rect 2828 32340 2884 32350
rect 3164 32340 3220 32396
rect 3276 32386 3332 32396
rect 3388 32452 3444 33068
rect 3388 32358 3444 32396
rect 2828 32338 3220 32340
rect 2828 32286 2830 32338
rect 2882 32286 3220 32338
rect 2828 32284 3220 32286
rect 2828 32274 2884 32284
rect 2828 32116 2884 32126
rect 2828 32002 2884 32060
rect 2828 31950 2830 32002
rect 2882 31950 2884 32002
rect 2828 31938 2884 31950
rect 3164 31556 3220 32284
rect 3500 32116 3556 33292
rect 3612 32340 3668 33854
rect 3724 33346 3780 34300
rect 3836 34300 4228 34356
rect 4284 34580 4340 34590
rect 3836 34130 3892 34300
rect 3836 34078 3838 34130
rect 3890 34078 3892 34130
rect 3836 34066 3892 34078
rect 3948 34132 4004 34142
rect 3948 34038 4004 34076
rect 4172 34132 4228 34142
rect 4284 34132 4340 34524
rect 4396 34468 4452 34748
rect 4396 34402 4452 34412
rect 4172 34130 4340 34132
rect 4172 34078 4174 34130
rect 4226 34078 4340 34130
rect 4172 34076 4340 34078
rect 4844 34130 4900 35084
rect 4956 34468 5012 35252
rect 5068 35252 5124 35262
rect 5068 34914 5124 35196
rect 5068 34862 5070 34914
rect 5122 34862 5124 34914
rect 5068 34850 5124 34862
rect 4956 34402 5012 34412
rect 5068 34692 5124 34702
rect 5068 34242 5124 34636
rect 5068 34190 5070 34242
rect 5122 34190 5124 34242
rect 5068 34178 5124 34190
rect 4844 34078 4846 34130
rect 4898 34078 4900 34130
rect 4172 34066 4228 34076
rect 4844 34066 4900 34078
rect 4396 34020 4452 34030
rect 4396 33926 4452 33964
rect 3836 33908 3892 33918
rect 3892 33852 4116 33908
rect 3836 33842 3892 33852
rect 3948 33572 4004 33582
rect 4060 33572 4116 33852
rect 4464 33740 4728 33750
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4060 33516 4900 33572
rect 3948 33478 4004 33516
rect 3724 33294 3726 33346
rect 3778 33294 3780 33346
rect 3724 33282 3780 33294
rect 4396 33346 4452 33358
rect 4396 33294 4398 33346
rect 4450 33294 4452 33346
rect 4060 33124 4116 33134
rect 4116 33068 4340 33124
rect 4060 33058 4116 33068
rect 4284 33012 4340 33068
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4284 32946 4340 32956
rect 3804 32890 4068 32900
rect 4396 32900 4452 33294
rect 4732 33348 4788 33358
rect 4620 33012 4676 33022
rect 4732 33012 4788 33292
rect 4676 32956 4788 33012
rect 4844 33012 4900 33516
rect 5068 33346 5124 33358
rect 5068 33294 5070 33346
rect 5122 33294 5124 33346
rect 5068 33124 5124 33294
rect 5068 33058 5124 33068
rect 4620 32946 4676 32956
rect 4844 32946 4900 32956
rect 4396 32834 4452 32844
rect 3948 32676 4004 32686
rect 4172 32676 4228 32686
rect 4004 32620 4116 32676
rect 3948 32610 4004 32620
rect 3612 32274 3668 32284
rect 3836 32562 3892 32574
rect 3836 32510 3838 32562
rect 3890 32510 3892 32562
rect 3836 32228 3892 32510
rect 4060 32452 4116 32620
rect 4172 32582 4228 32620
rect 4620 32620 5012 32676
rect 4620 32564 4676 32620
rect 4620 32498 4676 32508
rect 4060 32386 4116 32396
rect 4956 32450 5012 32620
rect 4956 32398 4958 32450
rect 5010 32398 5012 32450
rect 4956 32386 5012 32398
rect 3836 32162 3892 32172
rect 3948 32338 4004 32350
rect 3948 32286 3950 32338
rect 4002 32286 4004 32338
rect 3388 31892 3444 31902
rect 3164 31490 3220 31500
rect 3276 31780 3332 31790
rect 3052 31332 3108 31342
rect 2940 30882 2996 30894
rect 2940 30830 2942 30882
rect 2994 30830 2996 30882
rect 2828 30436 2884 30446
rect 2940 30436 2996 30830
rect 2828 30434 2996 30436
rect 2828 30382 2830 30434
rect 2882 30382 2996 30434
rect 2828 30380 2996 30382
rect 2828 30370 2884 30380
rect 2716 30258 2772 30268
rect 2940 30212 2996 30380
rect 2940 30146 2996 30156
rect 2828 29428 2884 29438
rect 2828 29334 2884 29372
rect 2604 29250 2660 29260
rect 2380 27858 2436 28028
rect 2604 28980 2660 28990
rect 2380 27806 2382 27858
rect 2434 27806 2436 27858
rect 2380 27794 2436 27806
rect 2492 27972 2548 27982
rect 2492 27636 2548 27916
rect 2268 25106 2324 25116
rect 2380 27580 2548 27636
rect 2156 24724 2212 24734
rect 2156 24610 2212 24668
rect 2156 24558 2158 24610
rect 2210 24558 2212 24610
rect 2156 24546 2212 24558
rect 2268 22148 2324 22158
rect 1820 21298 1876 21308
rect 1932 21532 2100 21588
rect 2156 22146 2324 22148
rect 2156 22094 2270 22146
rect 2322 22094 2324 22146
rect 2156 22092 2324 22094
rect 1708 21028 1764 21038
rect 1708 20934 1764 20972
rect 1820 20356 1876 20366
rect 1708 18228 1764 18238
rect 1708 18134 1764 18172
rect 1820 18004 1876 20300
rect 1932 20132 1988 21532
rect 2044 21362 2100 21374
rect 2044 21310 2046 21362
rect 2098 21310 2100 21362
rect 2044 20580 2100 21310
rect 2044 20514 2100 20524
rect 1932 20066 1988 20076
rect 1596 16158 1598 16210
rect 1650 16158 1652 16210
rect 1596 16146 1652 16158
rect 1708 17948 1876 18004
rect 1932 19234 1988 19246
rect 1932 19182 1934 19234
rect 1986 19182 1988 19234
rect 1708 15540 1764 17948
rect 1820 16996 1876 17006
rect 1820 16100 1876 16940
rect 1820 16034 1876 16044
rect 1932 15764 1988 19182
rect 2156 19124 2212 22092
rect 2268 22082 2324 22092
rect 2156 19058 2212 19068
rect 2268 21364 2324 21374
rect 2268 19012 2324 21308
rect 2380 21028 2436 27580
rect 2604 27524 2660 28924
rect 2828 28868 2884 28878
rect 2828 28774 2884 28812
rect 2492 27468 2660 27524
rect 2716 27860 2772 27870
rect 2492 26180 2548 27468
rect 2716 27076 2772 27804
rect 2940 27748 2996 27758
rect 2828 27300 2884 27310
rect 2940 27300 2996 27692
rect 2828 27298 2996 27300
rect 2828 27246 2830 27298
rect 2882 27246 2996 27298
rect 2828 27244 2996 27246
rect 3052 27300 3108 31276
rect 3276 30996 3332 31724
rect 3388 31778 3444 31836
rect 3388 31726 3390 31778
rect 3442 31726 3444 31778
rect 3388 31714 3444 31726
rect 3276 30930 3332 30940
rect 3388 30770 3444 30782
rect 3388 30718 3390 30770
rect 3442 30718 3444 30770
rect 3388 30660 3444 30718
rect 3388 30594 3444 30604
rect 3500 30548 3556 32060
rect 3948 32116 4004 32286
rect 4172 32340 4228 32378
rect 4172 32274 4228 32284
rect 4284 32340 4340 32350
rect 4284 32338 4900 32340
rect 4284 32286 4286 32338
rect 4338 32286 4900 32338
rect 4284 32284 4900 32286
rect 4284 32274 4340 32284
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 3948 32050 4004 32060
rect 4844 32004 4900 32284
rect 4732 31948 4900 32004
rect 3612 31890 3668 31902
rect 3612 31838 3614 31890
rect 3666 31838 3668 31890
rect 3612 31780 3668 31838
rect 3612 31714 3668 31724
rect 4284 31780 4340 31790
rect 4284 31686 4340 31724
rect 3948 31666 4004 31678
rect 3948 31614 3950 31666
rect 4002 31614 4004 31666
rect 3948 31556 4004 31614
rect 3612 31500 4340 31556
rect 3612 31332 3668 31500
rect 4284 31444 4340 31500
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4284 31378 4340 31388
rect 4396 31500 4676 31556
rect 3804 31322 4068 31332
rect 3612 31266 3668 31276
rect 4396 31108 4452 31500
rect 4060 31052 4452 31108
rect 4508 31332 4564 31342
rect 4508 31108 4564 31276
rect 3612 30994 3668 31006
rect 3612 30942 3614 30994
rect 3666 30942 3668 30994
rect 3612 30772 3668 30942
rect 3612 30706 3668 30716
rect 3948 30996 4004 31006
rect 3948 30548 4004 30940
rect 4060 30660 4116 31052
rect 4508 31042 4564 31052
rect 4396 30884 4452 30894
rect 4060 30594 4116 30604
rect 4284 30882 4452 30884
rect 4284 30830 4398 30882
rect 4450 30830 4452 30882
rect 4284 30828 4452 30830
rect 3500 30492 4004 30548
rect 4172 30548 4228 30558
rect 4060 30212 4116 30222
rect 4060 30118 4116 30156
rect 3612 30098 3668 30110
rect 3612 30046 3614 30098
rect 3666 30046 3668 30098
rect 3612 29652 3668 30046
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 4060 29652 4116 29662
rect 3612 29596 4004 29652
rect 3276 29540 3332 29550
rect 3164 29316 3220 29326
rect 3164 27748 3220 29260
rect 3276 29314 3332 29484
rect 3836 29428 3892 29438
rect 3836 29334 3892 29372
rect 3276 29262 3278 29314
rect 3330 29262 3332 29314
rect 3276 28868 3332 29262
rect 3388 29202 3444 29214
rect 3388 29150 3390 29202
rect 3442 29150 3444 29202
rect 3388 28980 3444 29150
rect 3388 28914 3444 28924
rect 3276 28802 3332 28812
rect 3500 28754 3556 28766
rect 3500 28702 3502 28754
rect 3554 28702 3556 28754
rect 3276 28642 3332 28654
rect 3276 28590 3278 28642
rect 3330 28590 3332 28642
rect 3276 28420 3332 28590
rect 3276 28354 3332 28364
rect 3500 28084 3556 28702
rect 3612 28644 3668 28654
rect 3612 28550 3668 28588
rect 3948 28644 4004 29596
rect 4060 29426 4116 29596
rect 4172 29538 4228 30492
rect 4284 29764 4340 30828
rect 4396 30818 4452 30828
rect 4620 30772 4676 31500
rect 4732 31108 4788 31948
rect 4956 31890 5012 31902
rect 5180 31892 5236 37548
rect 5292 37380 5348 37390
rect 5292 37154 5348 37324
rect 5292 37102 5294 37154
rect 5346 37102 5348 37154
rect 5292 37090 5348 37102
rect 5292 35924 5348 35934
rect 5292 35698 5348 35868
rect 5292 35646 5294 35698
rect 5346 35646 5348 35698
rect 5292 35634 5348 35646
rect 5292 35028 5348 35038
rect 5292 34934 5348 34972
rect 5292 34580 5348 34590
rect 5292 34018 5348 34524
rect 5292 33966 5294 34018
rect 5346 33966 5348 34018
rect 5292 33684 5348 33966
rect 5292 33618 5348 33628
rect 5404 33572 5460 39116
rect 5628 38052 5684 38062
rect 5628 37958 5684 37996
rect 5964 37604 6020 42700
rect 6076 42532 6132 45500
rect 6188 45332 6244 45838
rect 6188 45266 6244 45276
rect 6188 45108 6244 45118
rect 6188 44322 6244 45052
rect 6188 44270 6190 44322
rect 6242 44270 6244 44322
rect 6188 44258 6244 44270
rect 6300 43876 6356 50092
rect 6412 48468 6468 48478
rect 6412 48242 6468 48412
rect 6412 48190 6414 48242
rect 6466 48190 6468 48242
rect 6412 48178 6468 48190
rect 6524 48244 6580 52668
rect 6636 52276 6692 52286
rect 6636 52162 6692 52220
rect 6636 52110 6638 52162
rect 6690 52110 6692 52162
rect 6636 51940 6692 52110
rect 6636 51874 6692 51884
rect 6748 52164 6804 52892
rect 6636 51604 6692 51614
rect 6636 50148 6692 51548
rect 6636 50082 6692 50092
rect 6748 51378 6804 52108
rect 6748 51326 6750 51378
rect 6802 51326 6804 51378
rect 6748 49810 6804 51326
rect 6860 51604 6916 51614
rect 6860 50708 6916 51548
rect 6972 50820 7028 55132
rect 7084 54516 7140 54526
rect 7084 54422 7140 54460
rect 7308 54290 7364 54302
rect 7308 54238 7310 54290
rect 7362 54238 7364 54290
rect 7308 53844 7364 54238
rect 7308 53778 7364 53788
rect 7420 53620 7476 56030
rect 7980 56084 8036 56094
rect 8092 56084 8148 56142
rect 7980 56082 8148 56084
rect 7980 56030 7982 56082
rect 8034 56030 8148 56082
rect 7980 56028 8148 56030
rect 7980 56018 8036 56028
rect 7644 55858 7700 55870
rect 7644 55806 7646 55858
rect 7698 55806 7700 55858
rect 7644 55636 7700 55806
rect 7644 55570 7700 55580
rect 7644 55300 7700 55310
rect 8092 55300 8148 56028
rect 8316 55636 8372 57344
rect 7644 55298 8036 55300
rect 7644 55246 7646 55298
rect 7698 55246 8036 55298
rect 7644 55244 8036 55246
rect 7644 55234 7700 55244
rect 7868 54516 7924 54526
rect 7756 54514 7924 54516
rect 7756 54462 7870 54514
rect 7922 54462 7924 54514
rect 7756 54460 7924 54462
rect 7420 53554 7476 53564
rect 7532 54404 7588 54414
rect 7196 53508 7252 53518
rect 7196 53414 7252 53452
rect 7532 53172 7588 54348
rect 7644 54292 7700 54302
rect 7644 54198 7700 54236
rect 7644 53620 7700 53630
rect 7756 53620 7812 54460
rect 7868 54450 7924 54460
rect 7980 53956 8036 55244
rect 8092 55206 8148 55244
rect 8204 55580 8372 55636
rect 8204 55076 8260 55580
rect 8764 55524 8820 57344
rect 9212 56980 9268 57344
rect 9212 56914 9268 56924
rect 9324 56420 9380 56430
rect 8764 55458 8820 55468
rect 9100 55858 9156 55870
rect 9100 55806 9102 55858
rect 9154 55806 9156 55858
rect 8316 55410 8372 55422
rect 8316 55358 8318 55410
rect 8370 55358 8372 55410
rect 8316 55188 8372 55358
rect 9100 55300 9156 55806
rect 9100 55206 9156 55244
rect 8316 55122 8372 55132
rect 7980 53890 8036 53900
rect 8092 55020 8260 55076
rect 7644 53618 7812 53620
rect 7644 53566 7646 53618
rect 7698 53566 7812 53618
rect 7644 53564 7812 53566
rect 7980 53618 8036 53630
rect 7980 53566 7982 53618
rect 8034 53566 8036 53618
rect 7644 53396 7700 53564
rect 7644 53330 7700 53340
rect 7868 53506 7924 53518
rect 7868 53454 7870 53506
rect 7922 53454 7924 53506
rect 7532 53116 7700 53172
rect 7084 52948 7140 52958
rect 7644 52948 7700 53116
rect 7084 52946 7476 52948
rect 7084 52894 7086 52946
rect 7138 52894 7476 52946
rect 7084 52892 7476 52894
rect 7084 52882 7140 52892
rect 7084 52724 7140 52734
rect 7084 52386 7140 52668
rect 7084 52334 7086 52386
rect 7138 52334 7140 52386
rect 7084 52322 7140 52334
rect 7196 52722 7252 52734
rect 7196 52670 7198 52722
rect 7250 52670 7252 52722
rect 7196 51492 7252 52670
rect 7196 51426 7252 51436
rect 7084 51378 7140 51390
rect 7084 51326 7086 51378
rect 7138 51326 7140 51378
rect 7084 51044 7140 51326
rect 7308 51268 7364 51278
rect 7308 51174 7364 51212
rect 7084 50978 7140 50988
rect 6972 50754 7028 50764
rect 6860 50614 6916 50652
rect 7196 50708 7252 50718
rect 6748 49758 6750 49810
rect 6802 49758 6804 49810
rect 6748 49746 6804 49758
rect 6860 50260 6916 50270
rect 6748 49140 6804 49150
rect 6524 48178 6580 48188
rect 6636 48914 6692 48926
rect 6636 48862 6638 48914
rect 6690 48862 6692 48914
rect 6300 43810 6356 43820
rect 6412 47460 6468 47470
rect 6188 43652 6244 43662
rect 6188 43538 6244 43596
rect 6188 43486 6190 43538
rect 6242 43486 6244 43538
rect 6188 43474 6244 43486
rect 6300 43426 6356 43438
rect 6300 43374 6302 43426
rect 6354 43374 6356 43426
rect 6300 43092 6356 43374
rect 6300 43026 6356 43036
rect 6412 42756 6468 47404
rect 6636 45668 6692 48862
rect 6748 48580 6804 49084
rect 6748 47012 6804 48524
rect 6748 46946 6804 46956
rect 6860 46788 6916 50204
rect 7196 50148 7252 50652
rect 7084 50092 7252 50148
rect 7308 50706 7364 50718
rect 7308 50654 7310 50706
rect 7362 50654 7364 50706
rect 6972 49924 7028 49934
rect 7084 49924 7140 50092
rect 7028 49868 7140 49924
rect 6972 49858 7028 49868
rect 7084 49250 7140 49868
rect 7196 49924 7252 49934
rect 7196 49810 7252 49868
rect 7196 49758 7198 49810
rect 7250 49758 7252 49810
rect 7196 49746 7252 49758
rect 7084 49198 7086 49250
rect 7138 49198 7140 49250
rect 7084 49186 7140 49198
rect 7196 48692 7252 48702
rect 6524 45612 6692 45668
rect 6748 46732 6916 46788
rect 6972 48242 7028 48254
rect 6972 48190 6974 48242
rect 7026 48190 7028 48242
rect 6524 45556 6580 45612
rect 6524 45218 6580 45500
rect 6524 45166 6526 45218
rect 6578 45166 6580 45218
rect 6524 45154 6580 45166
rect 6636 44436 6692 44446
rect 6636 44322 6692 44380
rect 6636 44270 6638 44322
rect 6690 44270 6692 44322
rect 6636 44258 6692 44270
rect 6412 42662 6468 42700
rect 6076 42476 6468 42532
rect 6300 42308 6356 42318
rect 6188 42196 6244 42206
rect 6188 42102 6244 42140
rect 6188 40852 6244 40862
rect 6188 40292 6244 40796
rect 6300 40516 6356 42252
rect 6300 40422 6356 40460
rect 6188 40236 6356 40292
rect 6076 39620 6132 39630
rect 6076 39618 6244 39620
rect 6076 39566 6078 39618
rect 6130 39566 6244 39618
rect 6076 39564 6244 39566
rect 6076 39554 6132 39564
rect 5964 37538 6020 37548
rect 6076 38834 6132 38846
rect 6076 38782 6078 38834
rect 6130 38782 6132 38834
rect 5852 37268 5908 37278
rect 6076 37268 6132 38782
rect 6188 38164 6244 39564
rect 6188 37828 6244 38108
rect 6188 37762 6244 37772
rect 5852 37266 6132 37268
rect 5852 37214 5854 37266
rect 5906 37214 6132 37266
rect 5852 37212 6132 37214
rect 5852 36708 5908 37212
rect 6188 37156 6244 37166
rect 6188 37062 6244 37100
rect 5628 36652 5908 36708
rect 5516 36482 5572 36494
rect 5516 36430 5518 36482
rect 5570 36430 5572 36482
rect 5516 35364 5572 36430
rect 5516 35298 5572 35308
rect 5292 32338 5348 32350
rect 5292 32286 5294 32338
rect 5346 32286 5348 32338
rect 5292 32116 5348 32286
rect 5404 32116 5460 33516
rect 5516 35140 5572 35150
rect 5516 34018 5572 35084
rect 5516 33966 5518 34018
rect 5570 33966 5572 34018
rect 5516 32564 5572 33966
rect 5516 32498 5572 32508
rect 5516 32340 5572 32350
rect 5516 32246 5572 32284
rect 5404 32060 5572 32116
rect 5292 32050 5348 32060
rect 4956 31838 4958 31890
rect 5010 31838 5012 31890
rect 4844 31780 4900 31790
rect 4844 31686 4900 31724
rect 4732 31042 4788 31052
rect 4956 30994 5012 31838
rect 5068 31836 5236 31892
rect 5068 31444 5124 31836
rect 5404 31780 5460 31790
rect 5292 31778 5460 31780
rect 5292 31726 5406 31778
rect 5458 31726 5460 31778
rect 5292 31724 5460 31726
rect 5068 31378 5124 31388
rect 5180 31556 5236 31566
rect 5068 31108 5124 31118
rect 5068 31014 5124 31052
rect 4956 30942 4958 30994
rect 5010 30942 5012 30994
rect 4956 30930 5012 30942
rect 5180 30994 5236 31500
rect 5180 30942 5182 30994
rect 5234 30942 5236 30994
rect 4620 30716 5012 30772
rect 4956 30660 5012 30716
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4956 30594 5012 30604
rect 4464 30538 4728 30548
rect 4844 30548 4900 30558
rect 4844 30436 4900 30492
rect 4732 30380 4900 30436
rect 4620 30322 4676 30334
rect 4620 30270 4622 30322
rect 4674 30270 4676 30322
rect 4508 30212 4564 30222
rect 4508 30118 4564 30156
rect 4396 30100 4452 30110
rect 4396 29876 4452 30044
rect 4396 29810 4452 29820
rect 4284 29698 4340 29708
rect 4172 29486 4174 29538
rect 4226 29486 4228 29538
rect 4172 29474 4228 29486
rect 4060 29374 4062 29426
rect 4114 29374 4116 29426
rect 4060 29362 4116 29374
rect 4396 29428 4452 29438
rect 4620 29428 4676 30270
rect 4396 29426 4676 29428
rect 4396 29374 4398 29426
rect 4450 29374 4676 29426
rect 4396 29372 4676 29374
rect 4396 29362 4452 29372
rect 4732 29204 4788 30380
rect 4172 29148 4788 29204
rect 4844 30212 4900 30222
rect 4172 29092 4228 29148
rect 4172 29026 4228 29036
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 3948 28550 4004 28588
rect 4396 28642 4452 28654
rect 4396 28590 4398 28642
rect 4450 28590 4452 28642
rect 4396 28420 4452 28590
rect 4844 28642 4900 30156
rect 5180 29652 5236 30942
rect 5292 30996 5348 31724
rect 5404 31714 5460 31724
rect 5516 31556 5572 32060
rect 5628 31892 5684 36652
rect 5852 36484 5908 36494
rect 6300 36484 6356 40236
rect 6412 38276 6468 42476
rect 6636 42084 6692 42094
rect 6524 41186 6580 41198
rect 6524 41134 6526 41186
rect 6578 41134 6580 41186
rect 6524 40852 6580 41134
rect 6524 40786 6580 40796
rect 6524 39844 6580 39854
rect 6636 39844 6692 42028
rect 6748 41188 6804 46732
rect 6860 46564 6916 46574
rect 6860 46470 6916 46508
rect 6860 44994 6916 45006
rect 6860 44942 6862 44994
rect 6914 44942 6916 44994
rect 6860 44100 6916 44942
rect 6972 44436 7028 48190
rect 7196 48242 7252 48636
rect 7196 48190 7198 48242
rect 7250 48190 7252 48242
rect 7196 48178 7252 48190
rect 7196 47572 7252 47582
rect 7084 47460 7140 47470
rect 7084 47366 7140 47404
rect 7084 45666 7140 45678
rect 7084 45614 7086 45666
rect 7138 45614 7140 45666
rect 7084 44660 7140 45614
rect 7084 44594 7140 44604
rect 6972 44370 7028 44380
rect 6860 44034 6916 44044
rect 6972 43988 7028 43998
rect 6972 43540 7028 43932
rect 6972 43538 7140 43540
rect 6972 43486 6974 43538
rect 7026 43486 7140 43538
rect 6972 43484 7140 43486
rect 6972 43474 7028 43484
rect 6860 42308 6916 42318
rect 6860 42082 6916 42252
rect 7084 42308 7140 43484
rect 7196 43428 7252 47516
rect 7308 43652 7364 50654
rect 7420 48468 7476 52892
rect 7644 52946 7812 52948
rect 7644 52894 7646 52946
rect 7698 52894 7812 52946
rect 7644 52892 7812 52894
rect 7644 52882 7700 52892
rect 7644 52612 7700 52622
rect 7532 50596 7588 50606
rect 7532 50502 7588 50540
rect 7420 48402 7476 48412
rect 7532 50260 7588 50270
rect 7532 49924 7588 50204
rect 7420 47796 7476 47806
rect 7420 45666 7476 47740
rect 7532 47236 7588 49868
rect 7644 49588 7700 52556
rect 7756 51604 7812 52892
rect 7756 51378 7812 51548
rect 7756 51326 7758 51378
rect 7810 51326 7812 51378
rect 7756 51314 7812 51326
rect 7868 49812 7924 53454
rect 7980 53172 8036 53566
rect 7980 53106 8036 53116
rect 7980 52164 8036 52174
rect 7980 50594 8036 52108
rect 8092 51044 8148 55020
rect 8988 54628 9044 54638
rect 8428 54514 8484 54526
rect 8428 54462 8430 54514
rect 8482 54462 8484 54514
rect 8316 53620 8372 53630
rect 8428 53620 8484 54462
rect 8988 54402 9044 54572
rect 8988 54350 8990 54402
rect 9042 54350 9044 54402
rect 8988 54338 9044 54350
rect 9212 54514 9268 54526
rect 9212 54462 9214 54514
rect 9266 54462 9268 54514
rect 8316 53618 8484 53620
rect 8316 53566 8318 53618
rect 8370 53566 8484 53618
rect 8316 53564 8484 53566
rect 8652 54290 8708 54302
rect 8652 54238 8654 54290
rect 8706 54238 8708 54290
rect 8316 53172 8372 53564
rect 8316 53116 8596 53172
rect 8316 52946 8372 52958
rect 8316 52894 8318 52946
rect 8370 52894 8372 52946
rect 8204 52164 8260 52174
rect 8204 52070 8260 52108
rect 8316 51716 8372 52894
rect 8092 50978 8148 50988
rect 8204 51660 8372 51716
rect 8428 52500 8484 52510
rect 8428 51716 8484 52444
rect 7980 50542 7982 50594
rect 8034 50542 8036 50594
rect 7980 50530 8036 50542
rect 8092 50820 8148 50830
rect 7868 49746 7924 49756
rect 7644 49532 7924 49588
rect 7756 47572 7812 47582
rect 7756 47478 7812 47516
rect 7532 47180 7700 47236
rect 7644 47068 7700 47180
rect 7420 45614 7422 45666
rect 7474 45614 7476 45666
rect 7420 45444 7476 45614
rect 7532 47012 7588 47022
rect 7644 47012 7812 47068
rect 7532 46674 7588 46956
rect 7532 46622 7534 46674
rect 7586 46622 7588 46674
rect 7532 45556 7588 46622
rect 7756 46788 7812 47012
rect 7756 46004 7812 46732
rect 7868 46676 7924 49532
rect 7980 48356 8036 48366
rect 7980 48242 8036 48300
rect 7980 48190 7982 48242
rect 8034 48190 8036 48242
rect 7980 48178 8036 48190
rect 7980 47460 8036 47498
rect 7980 47394 8036 47404
rect 7868 46610 7924 46620
rect 7980 47236 8036 47246
rect 7980 46788 8036 47180
rect 7980 46562 8036 46732
rect 7980 46510 7982 46562
rect 8034 46510 8036 46562
rect 7980 46498 8036 46510
rect 7980 46004 8036 46014
rect 7756 46002 8036 46004
rect 7756 45950 7982 46002
rect 8034 45950 8036 46002
rect 7756 45948 8036 45950
rect 7532 45490 7588 45500
rect 7420 45378 7476 45388
rect 7756 45108 7812 45118
rect 7532 44322 7588 44334
rect 7532 44270 7534 44322
rect 7586 44270 7588 44322
rect 7532 44100 7588 44270
rect 7532 44034 7588 44044
rect 7308 43596 7700 43652
rect 7420 43428 7476 43438
rect 7196 43372 7364 43428
rect 7196 43204 7252 43214
rect 7196 42866 7252 43148
rect 7196 42814 7198 42866
rect 7250 42814 7252 42866
rect 7196 42802 7252 42814
rect 7308 42644 7364 43372
rect 7084 42242 7140 42252
rect 7196 42588 7364 42644
rect 6860 42030 6862 42082
rect 6914 42030 6916 42082
rect 6860 42018 6916 42030
rect 6972 42084 7028 42094
rect 6748 41122 6804 41132
rect 6860 41636 6916 41646
rect 6860 40852 6916 41580
rect 6524 39842 6692 39844
rect 6524 39790 6526 39842
rect 6578 39790 6692 39842
rect 6524 39788 6692 39790
rect 6748 40796 6916 40852
rect 6748 40178 6804 40796
rect 6748 40126 6750 40178
rect 6802 40126 6804 40178
rect 6524 39778 6580 39788
rect 6636 39620 6692 39630
rect 6636 38722 6692 39564
rect 6748 39172 6804 40126
rect 6860 40068 6916 40078
rect 6860 39842 6916 40012
rect 6860 39790 6862 39842
rect 6914 39790 6916 39842
rect 6860 39778 6916 39790
rect 6748 39106 6804 39116
rect 6972 38948 7028 42028
rect 7084 41524 7140 41534
rect 7084 41410 7140 41468
rect 7084 41358 7086 41410
rect 7138 41358 7140 41410
rect 7084 41346 7140 41358
rect 7196 39730 7252 42588
rect 7420 42084 7476 43372
rect 7532 42866 7588 42878
rect 7532 42814 7534 42866
rect 7586 42814 7588 42866
rect 7532 42532 7588 42814
rect 7532 42466 7588 42476
rect 7420 42018 7476 42028
rect 7420 41860 7476 41870
rect 7308 41804 7420 41860
rect 7308 41746 7364 41804
rect 7420 41794 7476 41804
rect 7308 41694 7310 41746
rect 7362 41694 7364 41746
rect 7308 41682 7364 41694
rect 7308 41188 7364 41198
rect 7308 41094 7364 41132
rect 7420 40180 7476 40190
rect 7308 39956 7364 39966
rect 7308 39842 7364 39900
rect 7308 39790 7310 39842
rect 7362 39790 7364 39842
rect 7308 39778 7364 39790
rect 7196 39678 7198 39730
rect 7250 39678 7252 39730
rect 7196 39666 7252 39678
rect 7308 39396 7364 39406
rect 7420 39396 7476 40124
rect 7308 39394 7476 39396
rect 7308 39342 7310 39394
rect 7362 39342 7476 39394
rect 7308 39340 7476 39342
rect 7308 39330 7364 39340
rect 7644 39284 7700 43596
rect 7756 41524 7812 45052
rect 7868 43540 7924 43550
rect 7868 42754 7924 43484
rect 7868 42702 7870 42754
rect 7922 42702 7924 42754
rect 7868 42690 7924 42702
rect 7756 41458 7812 41468
rect 7756 41186 7812 41198
rect 7756 41134 7758 41186
rect 7810 41134 7812 41186
rect 7756 40964 7812 41134
rect 7756 40898 7812 40908
rect 7980 40628 8036 45948
rect 8092 45108 8148 50764
rect 8204 50036 8260 51660
rect 8428 51650 8484 51660
rect 8428 51380 8484 51390
rect 8428 51286 8484 51324
rect 8316 50596 8372 50606
rect 8316 50502 8372 50540
rect 8540 50428 8596 53116
rect 8652 52500 8708 54238
rect 8988 53620 9044 53630
rect 9212 53620 9268 54462
rect 8988 53618 9268 53620
rect 8988 53566 8990 53618
rect 9042 53566 9268 53618
rect 8988 53564 9268 53566
rect 8652 52434 8708 52444
rect 8876 53508 8932 53518
rect 8876 52274 8932 53452
rect 8988 52724 9044 53564
rect 9324 53284 9380 56364
rect 9436 56196 9492 56206
rect 9436 55410 9492 56140
rect 9660 55524 9716 57344
rect 10108 57316 10164 57344
rect 10108 57250 10164 57260
rect 10108 56420 10164 56430
rect 9660 55458 9716 55468
rect 9884 56082 9940 56094
rect 9884 56030 9886 56082
rect 9938 56030 9940 56082
rect 9436 55358 9438 55410
rect 9490 55358 9492 55410
rect 9436 55346 9492 55358
rect 9548 55412 9604 55422
rect 9548 53396 9604 55356
rect 9772 55410 9828 55422
rect 9772 55358 9774 55410
rect 9826 55358 9828 55410
rect 9772 54516 9828 55358
rect 9884 55412 9940 56030
rect 10108 55970 10164 56364
rect 10108 55918 10110 55970
rect 10162 55918 10164 55970
rect 10108 55906 10164 55918
rect 10444 55858 10500 55870
rect 10444 55806 10446 55858
rect 10498 55806 10500 55858
rect 10444 55524 10500 55806
rect 10444 55458 10500 55468
rect 9884 55346 9940 55356
rect 9772 54450 9828 54460
rect 9996 55298 10052 55310
rect 9996 55246 9998 55298
rect 10050 55246 10052 55298
rect 9772 54292 9828 54302
rect 9996 54292 10052 55246
rect 10444 55300 10500 55310
rect 10444 55206 10500 55244
rect 9828 54236 10052 54292
rect 10220 54964 10276 54974
rect 9772 54198 9828 54236
rect 9884 53956 9940 53966
rect 9660 53842 9716 53854
rect 9660 53790 9662 53842
rect 9714 53790 9716 53842
rect 9660 53620 9716 53790
rect 9660 53554 9716 53564
rect 9772 53508 9828 53518
rect 9548 53340 9716 53396
rect 9324 53218 9380 53228
rect 9324 52946 9380 52958
rect 9324 52894 9326 52946
rect 9378 52894 9380 52946
rect 9324 52836 9380 52894
rect 9324 52770 9380 52780
rect 8988 52668 9268 52724
rect 8988 52388 9044 52398
rect 8988 52294 9044 52332
rect 8876 52222 8878 52274
rect 8930 52222 8932 52274
rect 8876 52210 8932 52222
rect 9100 52276 9156 52286
rect 8876 51828 8932 51838
rect 8764 51604 8820 51614
rect 8764 50484 8820 51548
rect 8540 50372 8708 50428
rect 8764 50418 8820 50428
rect 8204 49970 8260 49980
rect 8316 49924 8372 49934
rect 8316 49810 8372 49868
rect 8316 49758 8318 49810
rect 8370 49758 8372 49810
rect 8316 49746 8372 49758
rect 8428 49588 8484 49598
rect 8316 49140 8372 49150
rect 8204 49028 8260 49038
rect 8204 48934 8260 48972
rect 8316 47570 8372 49084
rect 8316 47518 8318 47570
rect 8370 47518 8372 47570
rect 8316 47506 8372 47518
rect 8204 47346 8260 47358
rect 8204 47294 8206 47346
rect 8258 47294 8260 47346
rect 8204 47124 8260 47294
rect 8204 47058 8260 47068
rect 8204 45890 8260 45902
rect 8204 45838 8206 45890
rect 8258 45838 8260 45890
rect 8204 45556 8260 45838
rect 8204 45490 8260 45500
rect 8092 45042 8148 45052
rect 8092 44882 8148 44894
rect 8092 44830 8094 44882
rect 8146 44830 8148 44882
rect 8092 44772 8148 44830
rect 8092 44706 8148 44716
rect 8204 44436 8260 44446
rect 8204 44342 8260 44380
rect 8092 44324 8148 44334
rect 8092 44230 8148 44268
rect 8204 44100 8260 44110
rect 8204 44006 8260 44044
rect 8428 43988 8484 49532
rect 8652 48356 8708 50372
rect 8652 48290 8708 48300
rect 8764 49588 8820 49598
rect 8652 48130 8708 48142
rect 8652 48078 8654 48130
rect 8706 48078 8708 48130
rect 8540 48018 8596 48030
rect 8540 47966 8542 48018
rect 8594 47966 8596 48018
rect 8540 47572 8596 47966
rect 8540 47506 8596 47516
rect 8652 46564 8708 48078
rect 8652 45108 8708 46508
rect 8764 46340 8820 49532
rect 8876 48804 8932 51772
rect 9100 50594 9156 52220
rect 9100 50542 9102 50594
rect 9154 50542 9156 50594
rect 9100 50428 9156 50542
rect 8988 50372 9156 50428
rect 9212 50428 9268 52668
rect 9324 52388 9380 52398
rect 9324 51378 9380 52332
rect 9548 52050 9604 52062
rect 9548 51998 9550 52050
rect 9602 51998 9604 52050
rect 9548 51940 9604 51998
rect 9548 51874 9604 51884
rect 9324 51326 9326 51378
rect 9378 51326 9380 51378
rect 9324 51314 9380 51326
rect 9548 51604 9604 51614
rect 9548 51268 9604 51548
rect 9548 50818 9604 51212
rect 9548 50766 9550 50818
rect 9602 50766 9604 50818
rect 9548 50754 9604 50766
rect 9212 50372 9604 50428
rect 8988 49140 9044 50372
rect 9324 50260 9380 50270
rect 9324 50036 9380 50204
rect 9212 49810 9268 49822
rect 9212 49758 9214 49810
rect 9266 49758 9268 49810
rect 9212 49476 9268 49758
rect 9212 49410 9268 49420
rect 8988 49084 9268 49140
rect 8876 48710 8932 48748
rect 8988 48914 9044 48926
rect 8988 48862 8990 48914
rect 9042 48862 9044 48914
rect 8988 48356 9044 48862
rect 8876 48300 9044 48356
rect 9100 48916 9156 48926
rect 8876 47460 8932 48300
rect 8988 48130 9044 48142
rect 8988 48078 8990 48130
rect 9042 48078 9044 48130
rect 8988 47684 9044 48078
rect 8988 47618 9044 47628
rect 9100 47570 9156 48860
rect 9212 48692 9268 49084
rect 9324 49138 9380 49980
rect 9324 49086 9326 49138
rect 9378 49086 9380 49138
rect 9324 49074 9380 49086
rect 9436 49028 9492 49038
rect 9212 48636 9380 48692
rect 9100 47518 9102 47570
rect 9154 47518 9156 47570
rect 9100 47506 9156 47518
rect 8988 47460 9044 47470
rect 8876 47404 8988 47460
rect 8988 46452 9044 47404
rect 9212 47236 9268 47246
rect 9100 46452 9156 46462
rect 8988 46450 9156 46452
rect 8988 46398 9102 46450
rect 9154 46398 9156 46450
rect 8988 46396 9156 46398
rect 8764 46274 8820 46284
rect 8988 45668 9044 45678
rect 8988 45574 9044 45612
rect 8652 45042 8708 45052
rect 8764 45332 8820 45342
rect 9100 45332 9156 46396
rect 9212 46116 9268 47180
rect 9324 47012 9380 48636
rect 9436 48242 9492 48972
rect 9436 48190 9438 48242
rect 9490 48190 9492 48242
rect 9436 47458 9492 48190
rect 9436 47406 9438 47458
rect 9490 47406 9492 47458
rect 9436 47394 9492 47406
rect 9324 46946 9380 46956
rect 9212 46050 9268 46060
rect 9212 45892 9268 45902
rect 9212 45444 9268 45836
rect 9212 45378 9268 45388
rect 9324 45666 9380 45678
rect 9324 45614 9326 45666
rect 9378 45614 9380 45666
rect 8540 44994 8596 45006
rect 8540 44942 8542 44994
rect 8594 44942 8596 44994
rect 8540 44660 8596 44942
rect 8764 44994 8820 45276
rect 8988 45276 9156 45332
rect 8764 44942 8766 44994
rect 8818 44942 8820 44994
rect 8764 44930 8820 44942
rect 8876 45218 8932 45230
rect 8876 45166 8878 45218
rect 8930 45166 8932 45218
rect 8540 44594 8596 44604
rect 8428 43922 8484 43932
rect 8764 43428 8820 43438
rect 8540 43314 8596 43326
rect 8540 43262 8542 43314
rect 8594 43262 8596 43314
rect 8428 43204 8484 43214
rect 8204 43092 8260 43102
rect 8204 42978 8260 43036
rect 8204 42926 8206 42978
rect 8258 42926 8260 42978
rect 8204 42914 8260 42926
rect 8092 42644 8148 42654
rect 8092 42084 8148 42588
rect 8428 42308 8484 43148
rect 8428 42242 8484 42252
rect 8092 42028 8372 42084
rect 8092 41412 8148 41422
rect 8092 41318 8148 41356
rect 8316 40852 8372 42028
rect 8316 40786 8372 40796
rect 8428 41746 8484 41758
rect 8428 41694 8430 41746
rect 8482 41694 8484 41746
rect 7980 40572 8372 40628
rect 8316 40514 8372 40572
rect 8316 40462 8318 40514
rect 8370 40462 8372 40514
rect 8316 40450 8372 40462
rect 8204 40404 8260 40414
rect 6636 38670 6638 38722
rect 6690 38670 6692 38722
rect 6636 38658 6692 38670
rect 6748 38892 7028 38948
rect 7420 39228 7700 39284
rect 7868 40178 7924 40190
rect 7868 40126 7870 40178
rect 7922 40126 7924 40178
rect 7868 39618 7924 40126
rect 8204 39732 8260 40348
rect 8428 39844 8484 41694
rect 8540 41300 8596 43262
rect 8764 41972 8820 43372
rect 8876 42756 8932 45166
rect 8988 43316 9044 45276
rect 9324 45220 9380 45614
rect 9212 45164 9380 45220
rect 8988 43250 9044 43260
rect 9100 44210 9156 44222
rect 9100 44158 9102 44210
rect 9154 44158 9156 44210
rect 9100 43538 9156 44158
rect 9100 43486 9102 43538
rect 9154 43486 9156 43538
rect 8988 42756 9044 42766
rect 8876 42754 9044 42756
rect 8876 42702 8990 42754
rect 9042 42702 9044 42754
rect 8876 42700 9044 42702
rect 8988 42690 9044 42700
rect 8876 42308 8932 42318
rect 8876 41972 8932 42252
rect 9100 42308 9156 43486
rect 9212 43092 9268 45164
rect 9212 43026 9268 43036
rect 9324 44994 9380 45006
rect 9324 44942 9326 44994
rect 9378 44942 9380 44994
rect 9324 43652 9380 44942
rect 9100 42242 9156 42252
rect 9212 42530 9268 42542
rect 9212 42478 9214 42530
rect 9266 42478 9268 42530
rect 8988 42196 9044 42206
rect 8988 42102 9044 42140
rect 9212 42082 9268 42478
rect 9324 42196 9380 43596
rect 9324 42130 9380 42140
rect 9436 44772 9492 44782
rect 9212 42030 9214 42082
rect 9266 42030 9268 42082
rect 9212 42018 9268 42030
rect 9324 41972 9380 41982
rect 8876 41916 9156 41972
rect 8764 41906 8820 41916
rect 8540 41234 8596 41244
rect 8764 41188 8820 41198
rect 8764 40404 8820 41132
rect 8652 40402 8820 40404
rect 8652 40350 8766 40402
rect 8818 40350 8820 40402
rect 8652 40348 8820 40350
rect 8428 39788 8596 39844
rect 8204 39676 8372 39732
rect 7868 39566 7870 39618
rect 7922 39566 7924 39618
rect 6412 38210 6468 38220
rect 6636 38052 6692 38062
rect 5740 35812 5796 35822
rect 5740 35698 5796 35756
rect 5740 35646 5742 35698
rect 5794 35646 5796 35698
rect 5740 35634 5796 35646
rect 5852 35588 5908 36428
rect 5740 35252 5796 35262
rect 5740 33796 5796 35196
rect 5852 34914 5908 35532
rect 6076 36482 6356 36484
rect 6076 36430 6302 36482
rect 6354 36430 6356 36482
rect 6076 36428 6356 36430
rect 5964 35476 6020 35486
rect 5964 35382 6020 35420
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34850 5908 34862
rect 5740 33730 5796 33740
rect 5852 34580 5908 34590
rect 5852 33348 5908 34524
rect 6076 34580 6132 36428
rect 6300 36418 6356 36428
rect 6412 38050 6692 38052
rect 6412 37998 6638 38050
rect 6690 37998 6692 38050
rect 6412 37996 6692 37998
rect 6412 36260 6468 37996
rect 6636 37986 6692 37996
rect 6300 36204 6468 36260
rect 6524 37604 6580 37614
rect 6076 34514 6132 34524
rect 6188 36148 6244 36158
rect 6076 34132 6132 34142
rect 6076 34038 6132 34076
rect 5964 33348 6020 33358
rect 5852 33346 6020 33348
rect 5852 33294 5966 33346
rect 6018 33294 6020 33346
rect 5852 33292 6020 33294
rect 5852 32450 5908 32462
rect 5852 32398 5854 32450
rect 5906 32398 5908 32450
rect 5740 32338 5796 32350
rect 5740 32286 5742 32338
rect 5794 32286 5796 32338
rect 5740 32004 5796 32286
rect 5740 31938 5796 31948
rect 5628 31826 5684 31836
rect 5516 31490 5572 31500
rect 5852 30996 5908 32398
rect 5964 32452 6020 33292
rect 5964 32386 6020 32396
rect 6188 32004 6244 36092
rect 6300 34914 6356 36204
rect 6412 35588 6468 35598
rect 6412 35494 6468 35532
rect 6300 34862 6302 34914
rect 6354 34862 6356 34914
rect 6300 34132 6356 34862
rect 6300 34066 6356 34076
rect 6188 31778 6244 31948
rect 6188 31726 6190 31778
rect 6242 31726 6244 31778
rect 6188 31444 6244 31726
rect 6188 31378 6244 31388
rect 6412 34020 6468 34030
rect 6412 32562 6468 33964
rect 6524 34018 6580 37548
rect 6524 33966 6526 34018
rect 6578 33966 6580 34018
rect 6524 33954 6580 33966
rect 6636 34804 6692 34814
rect 6524 33684 6580 33694
rect 6524 33570 6580 33628
rect 6524 33518 6526 33570
rect 6578 33518 6580 33570
rect 6524 33506 6580 33518
rect 6636 33460 6692 34748
rect 6636 33366 6692 33404
rect 6636 33012 6692 33022
rect 6412 32510 6414 32562
rect 6466 32510 6468 32562
rect 6188 31108 6244 31118
rect 6188 31014 6244 31052
rect 6412 31108 6468 32510
rect 5852 30940 6020 30996
rect 5292 30210 5348 30940
rect 5516 30884 5572 30894
rect 5516 30882 5908 30884
rect 5516 30830 5518 30882
rect 5570 30830 5908 30882
rect 5516 30828 5908 30830
rect 5516 30818 5572 30828
rect 5292 30158 5294 30210
rect 5346 30158 5348 30210
rect 5292 30146 5348 30158
rect 5628 30212 5684 30222
rect 5628 30118 5684 30156
rect 5180 29586 5236 29596
rect 5852 29650 5908 30828
rect 5964 30660 6020 30940
rect 5964 30594 6020 30604
rect 5852 29598 5854 29650
rect 5906 29598 5908 29650
rect 5852 29586 5908 29598
rect 6076 30212 6132 30222
rect 5404 29540 5460 29550
rect 5180 29426 5236 29438
rect 5180 29374 5182 29426
rect 5234 29374 5236 29426
rect 4956 29316 5012 29326
rect 4956 29222 5012 29260
rect 5068 29202 5124 29214
rect 5068 29150 5070 29202
rect 5122 29150 5124 29202
rect 4956 28756 5012 28766
rect 4956 28662 5012 28700
rect 4844 28590 4846 28642
rect 4898 28590 4900 28642
rect 4844 28578 4900 28590
rect 4452 28364 4564 28420
rect 4396 28354 4452 28364
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 4172 28196 4228 28206
rect 3500 28028 3668 28084
rect 3500 27860 3556 27870
rect 3500 27766 3556 27804
rect 3388 27748 3444 27758
rect 3164 27746 3444 27748
rect 3164 27694 3390 27746
rect 3442 27694 3444 27746
rect 3164 27692 3444 27694
rect 3388 27682 3444 27692
rect 3612 27412 3668 28028
rect 3500 27356 3668 27412
rect 3724 27860 3780 27870
rect 3948 27860 4004 27870
rect 3724 27412 3780 27804
rect 3500 27300 3556 27356
rect 3724 27346 3780 27356
rect 3836 27804 3948 27860
rect 2828 27234 2884 27244
rect 3052 27234 3108 27244
rect 3276 27298 3556 27300
rect 3276 27246 3502 27298
rect 3554 27246 3556 27298
rect 3276 27244 3556 27246
rect 3164 27188 3220 27198
rect 2716 27020 2996 27076
rect 2828 26852 2884 26862
rect 2828 26514 2884 26796
rect 2828 26462 2830 26514
rect 2882 26462 2884 26514
rect 2828 26450 2884 26462
rect 2492 26114 2548 26124
rect 2940 25956 2996 27020
rect 2716 25900 2996 25956
rect 3052 25956 3108 25966
rect 2492 24612 2548 24622
rect 2492 22596 2548 24556
rect 2492 22530 2548 22540
rect 2604 23938 2660 23950
rect 2604 23886 2606 23938
rect 2658 23886 2660 23938
rect 2604 22372 2660 23886
rect 2716 22708 2772 25900
rect 2940 25732 2996 25742
rect 3052 25732 3108 25900
rect 2940 25730 3108 25732
rect 2940 25678 2942 25730
rect 2994 25678 3108 25730
rect 2940 25676 3108 25678
rect 2940 25666 2996 25676
rect 2828 24722 2884 24734
rect 2828 24670 2830 24722
rect 2882 24670 2884 24722
rect 2828 23380 2884 24670
rect 3164 24612 3220 27132
rect 3276 26402 3332 27244
rect 3500 27234 3556 27244
rect 3612 27188 3668 27198
rect 3612 27094 3668 27132
rect 3500 26852 3556 26862
rect 3836 26852 3892 27804
rect 3948 27766 4004 27804
rect 3948 27300 4004 27310
rect 3948 27186 4004 27244
rect 3948 27134 3950 27186
rect 4002 27134 4004 27186
rect 3948 26964 4004 27134
rect 3948 26898 4004 26908
rect 3500 26850 3668 26852
rect 3500 26798 3502 26850
rect 3554 26798 3668 26850
rect 3500 26796 3668 26798
rect 3500 26786 3556 26796
rect 3276 26350 3278 26402
rect 3330 26350 3332 26402
rect 3276 25956 3332 26350
rect 3500 26628 3556 26638
rect 3276 25890 3332 25900
rect 3388 26066 3444 26078
rect 3388 26014 3390 26066
rect 3442 26014 3444 26066
rect 3388 25508 3444 26014
rect 3500 25678 3556 26572
rect 3612 26292 3668 26796
rect 3836 26786 3892 26796
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 3948 26292 4004 26302
rect 3612 26290 4004 26292
rect 3612 26238 3950 26290
rect 4002 26238 4004 26290
rect 3612 26236 4004 26238
rect 3948 26226 4004 26236
rect 4172 26290 4228 28140
rect 4396 28084 4452 28094
rect 4396 27970 4452 28028
rect 4396 27918 4398 27970
rect 4450 27918 4452 27970
rect 4396 27906 4452 27918
rect 4396 27748 4452 27758
rect 4508 27748 4564 28364
rect 4452 27692 4564 27748
rect 4732 28196 4788 28206
rect 4396 27682 4452 27692
rect 4732 27636 4788 28140
rect 4956 27746 5012 27758
rect 4956 27694 4958 27746
rect 5010 27694 5012 27746
rect 4732 27580 4844 27636
rect 4464 27468 4728 27478
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4788 27300 4844 27580
rect 4956 27524 5012 27694
rect 4956 27458 5012 27468
rect 4732 27244 4844 27300
rect 4396 27076 4452 27086
rect 4620 27076 4676 27086
rect 4396 27074 4620 27076
rect 4396 27022 4398 27074
rect 4450 27022 4620 27074
rect 4396 27020 4620 27022
rect 4396 27010 4452 27020
rect 4620 27010 4676 27020
rect 4732 27074 4788 27244
rect 4956 27188 5012 27198
rect 4956 27094 5012 27132
rect 4732 27022 4734 27074
rect 4786 27022 4788 27074
rect 4732 27010 4788 27022
rect 4956 26964 5012 26974
rect 4396 26628 4452 26638
rect 4396 26516 4452 26572
rect 4172 26238 4174 26290
rect 4226 26238 4228 26290
rect 4172 26226 4228 26238
rect 4284 26460 4452 26516
rect 3836 26066 3892 26078
rect 3836 26014 3838 26066
rect 3890 26014 3892 26066
rect 3836 25844 3892 26014
rect 4060 26068 4116 26078
rect 4284 26068 4340 26460
rect 4956 26404 5012 26908
rect 4956 26338 5012 26348
rect 4396 26292 4452 26302
rect 4396 26198 4452 26236
rect 5068 26292 5124 29150
rect 5068 26226 5124 26236
rect 4060 26066 4340 26068
rect 4060 26014 4062 26066
rect 4114 26014 4340 26066
rect 4060 26012 4340 26014
rect 5068 26066 5124 26078
rect 5068 26014 5070 26066
rect 5122 26014 5124 26066
rect 4060 26002 4116 26012
rect 4464 25900 4728 25910
rect 3836 25778 3892 25788
rect 4284 25844 4340 25854
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 4844 25844 4900 25854
rect 4284 25732 4340 25788
rect 4396 25732 4452 25742
rect 4284 25730 4452 25732
rect 4284 25678 4398 25730
rect 4450 25678 4452 25730
rect 3500 25622 4116 25678
rect 4284 25676 4452 25678
rect 4396 25666 4452 25676
rect 4060 25618 4116 25622
rect 4620 25620 4676 25630
rect 4060 25566 4062 25618
rect 4114 25566 4116 25618
rect 4060 25554 4116 25566
rect 4508 25564 4620 25620
rect 3388 25442 3444 25452
rect 4172 25508 4228 25518
rect 4396 25508 4452 25518
rect 4508 25508 4564 25564
rect 4620 25554 4676 25564
rect 4228 25506 4564 25508
rect 4228 25454 4398 25506
rect 4450 25454 4564 25506
rect 4228 25452 4564 25454
rect 4732 25508 4788 25518
rect 4844 25508 4900 25788
rect 4732 25506 4900 25508
rect 4732 25454 4734 25506
rect 4786 25454 4900 25506
rect 4732 25452 4900 25454
rect 4172 25442 4228 25452
rect 4396 25442 4452 25452
rect 4732 25442 4788 25452
rect 3612 25396 3668 25406
rect 3388 25172 3444 25182
rect 3276 24724 3332 24734
rect 3276 24630 3332 24668
rect 3052 23938 3108 23950
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 2940 23380 2996 23390
rect 2828 23378 2996 23380
rect 2828 23326 2942 23378
rect 2994 23326 2996 23378
rect 2828 23324 2996 23326
rect 2940 23314 2996 23324
rect 2716 22642 2772 22652
rect 2828 23156 2884 23166
rect 2492 22316 2660 22372
rect 2492 21140 2548 22316
rect 2716 22260 2772 22270
rect 2716 22166 2772 22204
rect 2828 22148 2884 23100
rect 3052 22596 3108 23886
rect 2828 22082 2884 22092
rect 2940 22540 3108 22596
rect 2716 21700 2772 21710
rect 2716 21606 2772 21644
rect 2940 21140 2996 22540
rect 2492 21084 2772 21140
rect 2380 20972 2660 21028
rect 2380 20692 2436 20702
rect 2380 19906 2436 20636
rect 2380 19854 2382 19906
rect 2434 19854 2436 19906
rect 2380 19842 2436 19854
rect 2492 19346 2548 19358
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2380 19236 2436 19246
rect 2380 19142 2436 19180
rect 2268 18956 2436 19012
rect 2044 18900 2100 18910
rect 2044 18450 2100 18844
rect 2044 18398 2046 18450
rect 2098 18398 2100 18450
rect 2044 18386 2100 18398
rect 2156 17668 2212 17678
rect 2156 17574 2212 17612
rect 2268 16772 2324 16782
rect 2268 16678 2324 16716
rect 1932 15698 1988 15708
rect 2156 16660 2212 16670
rect 1708 15484 2100 15540
rect 1932 15316 1988 15326
rect 1484 15204 1540 15214
rect 1484 14418 1540 15148
rect 1596 14642 1652 14654
rect 1596 14590 1598 14642
rect 1650 14590 1652 14642
rect 1596 14532 1652 14590
rect 1820 14644 1876 14654
rect 1820 14550 1876 14588
rect 1596 14466 1652 14476
rect 1484 14366 1486 14418
rect 1538 14366 1540 14418
rect 1484 14354 1540 14366
rect 1148 13134 1150 13186
rect 1202 13134 1204 13186
rect 1148 13122 1204 13134
rect 1260 13692 1428 13748
rect 1708 13860 1764 13870
rect 1148 12292 1204 12302
rect 1148 12198 1204 12236
rect 1148 11956 1204 11966
rect 1036 8932 1092 8942
rect 812 8930 1092 8932
rect 812 8878 1038 8930
rect 1090 8878 1092 8930
rect 812 8876 1092 8878
rect 1036 8866 1092 8876
rect 588 8652 1092 8708
rect 476 8540 980 8596
rect 812 8372 868 8382
rect 364 7186 420 7196
rect 476 7588 532 7598
rect 252 6244 308 6254
rect 28 6188 252 6244
rect 252 6178 308 6188
rect 476 3668 532 7532
rect 700 7028 756 7038
rect 476 3612 644 3668
rect 476 3444 532 3454
rect 476 2660 532 3388
rect 588 2660 644 3612
rect 700 2884 756 6972
rect 812 3668 868 8316
rect 812 3602 868 3612
rect 924 3388 980 8540
rect 1036 5346 1092 8652
rect 1148 7476 1204 11900
rect 1260 11844 1316 13692
rect 1372 13524 1428 13534
rect 1708 13524 1764 13804
rect 1372 13522 1764 13524
rect 1372 13470 1374 13522
rect 1426 13470 1764 13522
rect 1372 13468 1764 13470
rect 1372 13458 1428 13468
rect 1932 12628 1988 15260
rect 1820 12572 1988 12628
rect 1260 11778 1316 11788
rect 1484 12178 1540 12190
rect 1484 12126 1486 12178
rect 1538 12126 1540 12178
rect 1260 11620 1316 11630
rect 1260 11394 1316 11564
rect 1260 11342 1262 11394
rect 1314 11342 1316 11394
rect 1260 11330 1316 11342
rect 1372 10948 1428 10958
rect 1372 10610 1428 10892
rect 1372 10558 1374 10610
rect 1426 10558 1428 10610
rect 1372 10546 1428 10558
rect 1260 9044 1316 9054
rect 1260 8950 1316 8988
rect 1148 7420 1428 7476
rect 1260 7252 1316 7262
rect 1036 5294 1038 5346
rect 1090 5294 1092 5346
rect 1036 5282 1092 5294
rect 1148 6916 1204 6926
rect 924 3332 1092 3388
rect 700 2818 756 2828
rect 1036 2772 1092 3332
rect 1148 2994 1204 6860
rect 1260 6130 1316 7196
rect 1372 6356 1428 7420
rect 1484 6916 1540 12126
rect 1820 11620 1876 12572
rect 1932 12180 1988 12190
rect 1932 12086 1988 12124
rect 1820 11554 1876 11564
rect 1596 11508 1652 11518
rect 1596 11414 1652 11452
rect 1596 11172 1652 11182
rect 1596 8372 1652 11116
rect 2044 10612 2100 15484
rect 2156 14530 2212 16604
rect 2268 15764 2324 15774
rect 2268 14644 2324 15708
rect 2380 15202 2436 18956
rect 2492 18900 2548 19294
rect 2492 18834 2548 18844
rect 2492 18676 2548 18686
rect 2492 15316 2548 18620
rect 2492 15250 2548 15260
rect 2380 15150 2382 15202
rect 2434 15150 2436 15202
rect 2380 15138 2436 15150
rect 2380 14756 2436 14766
rect 2380 14662 2436 14700
rect 2268 14578 2324 14588
rect 2492 14644 2548 14654
rect 2492 14550 2548 14588
rect 2156 14478 2158 14530
rect 2210 14478 2212 14530
rect 2156 14420 2212 14478
rect 2156 14354 2212 14364
rect 2156 14084 2212 14094
rect 2604 14084 2660 20972
rect 2716 20356 2772 21084
rect 2828 21084 2996 21140
rect 3052 22370 3108 22382
rect 3052 22318 3054 22370
rect 3106 22318 3108 22370
rect 2828 21026 2884 21084
rect 2828 20974 2830 21026
rect 2882 20974 2884 21026
rect 2828 20962 2884 20974
rect 3052 20916 3108 22318
rect 3052 20850 3108 20860
rect 3164 21362 3220 24556
rect 3388 23548 3444 25116
rect 3612 23604 3668 25340
rect 5068 25172 5124 26014
rect 5180 25678 5236 29374
rect 5404 29426 5460 29484
rect 5404 29374 5406 29426
rect 5458 29374 5460 29426
rect 5404 29362 5460 29374
rect 5964 29428 6020 29438
rect 5964 29334 6020 29372
rect 5852 28980 5908 28990
rect 5404 28644 5460 28654
rect 5292 28642 5460 28644
rect 5292 28590 5406 28642
rect 5458 28590 5460 28642
rect 5292 28588 5460 28590
rect 5292 27860 5348 28588
rect 5404 28578 5460 28588
rect 5292 27188 5348 27804
rect 5852 27858 5908 28924
rect 6076 28756 6132 30156
rect 6300 30100 6356 30110
rect 6300 29650 6356 30044
rect 6412 29876 6468 31052
rect 6412 29810 6468 29820
rect 6524 32564 6580 32574
rect 6300 29598 6302 29650
rect 6354 29598 6356 29650
rect 6300 29586 6356 29598
rect 6412 29540 6468 29550
rect 6524 29540 6580 32508
rect 6636 30770 6692 32956
rect 6748 32450 6804 38892
rect 7308 38612 7364 38622
rect 6860 38500 6916 38510
rect 6860 37156 6916 38444
rect 7084 38276 7140 38286
rect 7084 38182 7140 38220
rect 7308 38274 7364 38556
rect 7308 38222 7310 38274
rect 7362 38222 7364 38274
rect 6860 37090 6916 37100
rect 6860 36708 6916 36718
rect 6860 36614 6916 36652
rect 7196 36708 7252 36718
rect 7196 36614 7252 36652
rect 7308 36596 7364 38222
rect 7420 38162 7476 39228
rect 7420 38110 7422 38162
rect 7474 38110 7476 38162
rect 7420 38098 7476 38110
rect 7532 38836 7588 38846
rect 7308 36530 7364 36540
rect 7420 37042 7476 37054
rect 7420 36990 7422 37042
rect 7474 36990 7476 37042
rect 6972 36148 7028 36158
rect 6972 35698 7028 36092
rect 7420 36148 7476 36990
rect 7532 36706 7588 38780
rect 7868 38724 7924 39566
rect 7980 39618 8036 39630
rect 7980 39566 7982 39618
rect 8034 39566 8036 39618
rect 7980 39508 8036 39566
rect 7980 39060 8036 39452
rect 8204 39508 8260 39518
rect 8204 39414 8260 39452
rect 7980 38994 8036 39004
rect 8204 38836 8260 38846
rect 8204 38742 8260 38780
rect 7868 38658 7924 38668
rect 7756 38610 7812 38622
rect 7756 38558 7758 38610
rect 7810 38558 7812 38610
rect 7756 38388 7812 38558
rect 7756 38332 7924 38388
rect 7756 38164 7812 38174
rect 7756 38070 7812 38108
rect 7868 36932 7924 38332
rect 8316 38162 8372 39676
rect 8428 39618 8484 39630
rect 8428 39566 8430 39618
rect 8482 39566 8484 39618
rect 8428 38724 8484 39566
rect 8428 38658 8484 38668
rect 8540 39172 8596 39788
rect 8316 38110 8318 38162
rect 8370 38110 8372 38162
rect 8316 38098 8372 38110
rect 8092 38050 8148 38062
rect 8092 37998 8094 38050
rect 8146 37998 8148 38050
rect 8092 37828 8148 37998
rect 8204 38052 8260 38062
rect 8204 37958 8260 37996
rect 8540 37828 8596 39116
rect 8652 38834 8708 40348
rect 8764 40338 8820 40348
rect 8876 41074 8932 41086
rect 8876 41022 8878 41074
rect 8930 41022 8932 41074
rect 8876 40068 8932 41022
rect 9100 40964 9156 41916
rect 9324 41878 9380 41916
rect 9324 41188 9380 41226
rect 9436 41188 9492 44716
rect 9548 44660 9604 50372
rect 9660 47460 9716 53340
rect 9772 52724 9828 53452
rect 9884 53170 9940 53900
rect 9996 53732 10052 53742
rect 9996 53638 10052 53676
rect 9884 53118 9886 53170
rect 9938 53118 9940 53170
rect 9884 53106 9940 53118
rect 9996 52834 10052 52846
rect 9996 52782 9998 52834
rect 10050 52782 10052 52834
rect 9884 52724 9940 52734
rect 9772 52722 9940 52724
rect 9772 52670 9886 52722
rect 9938 52670 9940 52722
rect 9772 52668 9940 52670
rect 9772 51828 9828 52668
rect 9884 52658 9940 52668
rect 9996 52500 10052 52782
rect 9772 51762 9828 51772
rect 9884 52444 10052 52500
rect 10108 52612 10164 52622
rect 9884 50820 9940 52444
rect 10108 52388 10164 52556
rect 9996 52332 10164 52388
rect 9996 52274 10052 52332
rect 9996 52222 9998 52274
rect 10050 52222 10052 52274
rect 9996 52052 10052 52222
rect 9996 51986 10052 51996
rect 10108 51940 10164 51950
rect 10108 51490 10164 51884
rect 10108 51438 10110 51490
rect 10162 51438 10164 51490
rect 10108 51426 10164 51438
rect 9884 50754 9940 50764
rect 9772 49812 9828 49822
rect 9772 49252 9828 49756
rect 10108 49810 10164 49822
rect 10108 49758 10110 49810
rect 10162 49758 10164 49810
rect 10108 49476 10164 49758
rect 9772 49186 9828 49196
rect 9884 49420 10164 49476
rect 9772 49028 9828 49038
rect 9772 48934 9828 48972
rect 9884 48804 9940 49420
rect 10108 49252 10164 49262
rect 10108 49026 10164 49196
rect 10108 48974 10110 49026
rect 10162 48974 10164 49026
rect 10108 48962 10164 48974
rect 9884 48748 10164 48804
rect 10108 48692 10164 48748
rect 10108 48626 10164 48636
rect 9884 48580 9940 48590
rect 9660 47394 9716 47404
rect 9772 48468 9828 48478
rect 9772 48242 9828 48412
rect 9772 48190 9774 48242
rect 9826 48190 9828 48242
rect 9772 45892 9828 48190
rect 9884 47908 9940 48524
rect 10108 48244 10164 48254
rect 9996 48132 10052 48142
rect 10108 48132 10164 48188
rect 9996 48130 10164 48132
rect 9996 48078 9998 48130
rect 10050 48078 10164 48130
rect 9996 48076 10164 48078
rect 9996 48066 10052 48076
rect 9884 47458 9940 47852
rect 10108 47572 10164 47582
rect 10108 47478 10164 47516
rect 9884 47406 9886 47458
rect 9938 47406 9940 47458
rect 9884 47394 9940 47406
rect 9884 47124 9940 47134
rect 9884 46674 9940 47068
rect 9884 46622 9886 46674
rect 9938 46622 9940 46674
rect 9884 46610 9940 46622
rect 10108 46676 10164 46686
rect 10220 46676 10276 54908
rect 10332 54740 10388 54750
rect 10332 54402 10388 54684
rect 10332 54350 10334 54402
rect 10386 54350 10388 54402
rect 10332 54338 10388 54350
rect 10556 54292 10612 57344
rect 11004 56644 11060 57344
rect 11452 56868 11508 57344
rect 11452 56802 11508 56812
rect 11900 56868 11956 57344
rect 11900 56802 11956 56812
rect 10892 56588 11060 56644
rect 11676 56644 11732 56654
rect 11900 56644 11956 56654
rect 11732 56588 11844 56644
rect 10780 56532 10836 56542
rect 10780 55970 10836 56476
rect 10780 55918 10782 55970
rect 10834 55918 10836 55970
rect 10780 55906 10836 55918
rect 10668 55748 10724 55758
rect 10668 54628 10724 55692
rect 10668 54562 10724 54572
rect 10780 55410 10836 55422
rect 10780 55358 10782 55410
rect 10834 55358 10836 55410
rect 10556 54226 10612 54236
rect 10668 54290 10724 54302
rect 10668 54238 10670 54290
rect 10722 54238 10724 54290
rect 10332 53618 10388 53630
rect 10332 53566 10334 53618
rect 10386 53566 10388 53618
rect 10332 53508 10388 53566
rect 10332 53442 10388 53452
rect 10668 53508 10724 54238
rect 10668 53442 10724 53452
rect 10780 53396 10836 55358
rect 10892 54516 10948 56588
rect 11676 56578 11732 56588
rect 11004 55972 11060 55982
rect 11004 55412 11060 55916
rect 11116 55860 11172 55870
rect 11564 55860 11620 55870
rect 11116 55858 11284 55860
rect 11116 55806 11118 55858
rect 11170 55806 11284 55858
rect 11116 55804 11284 55806
rect 11116 55794 11172 55804
rect 11116 55412 11172 55422
rect 11004 55410 11172 55412
rect 11004 55358 11118 55410
rect 11170 55358 11172 55410
rect 11004 55356 11172 55358
rect 11116 55346 11172 55356
rect 11228 55300 11284 55804
rect 11564 55766 11620 55804
rect 11788 55748 11844 56588
rect 11900 55970 11956 56588
rect 12348 56308 12404 57344
rect 12348 56242 12404 56252
rect 12796 56084 12852 57344
rect 13244 56756 13300 57344
rect 13244 56690 13300 56700
rect 13468 56756 13524 56766
rect 11900 55918 11902 55970
rect 11954 55918 11956 55970
rect 11900 55906 11956 55918
rect 12012 56028 12852 56084
rect 13244 56308 13300 56318
rect 13244 56082 13300 56252
rect 13244 56030 13246 56082
rect 13298 56030 13300 56082
rect 11788 55682 11844 55692
rect 11452 55300 11508 55310
rect 11228 55298 11508 55300
rect 11228 55246 11454 55298
rect 11506 55246 11508 55298
rect 11228 55244 11508 55246
rect 11452 54740 11508 55244
rect 11900 55300 11956 55310
rect 11900 55206 11956 55244
rect 11452 54674 11508 54684
rect 10892 54450 10948 54460
rect 11004 54628 11060 54638
rect 11004 54402 11060 54572
rect 11900 54628 11956 54638
rect 11900 54514 11956 54572
rect 11900 54462 11902 54514
rect 11954 54462 11956 54514
rect 11676 54404 11732 54414
rect 11004 54350 11006 54402
rect 11058 54350 11060 54402
rect 11004 54338 11060 54350
rect 11452 54402 11732 54404
rect 11452 54350 11678 54402
rect 11730 54350 11732 54402
rect 11452 54348 11732 54350
rect 11340 54290 11396 54302
rect 11340 54238 11342 54290
rect 11394 54238 11396 54290
rect 11004 53620 11060 53630
rect 11004 53526 11060 53564
rect 11340 53620 11396 54238
rect 11340 53554 11396 53564
rect 10780 53330 10836 53340
rect 10444 53284 10500 53294
rect 10332 49140 10388 49150
rect 10332 49046 10388 49084
rect 10332 48692 10388 48702
rect 10332 47012 10388 48636
rect 10332 46946 10388 46956
rect 10108 46674 10276 46676
rect 10108 46622 10110 46674
rect 10162 46622 10276 46674
rect 10108 46620 10276 46622
rect 10108 46610 10164 46620
rect 10220 46450 10276 46462
rect 10220 46398 10222 46450
rect 10274 46398 10276 46450
rect 9772 45826 9828 45836
rect 9884 46002 9940 46014
rect 9884 45950 9886 46002
rect 9938 45950 9940 46002
rect 9884 45668 9940 45950
rect 9884 45220 9940 45612
rect 9548 44594 9604 44604
rect 9660 45164 9940 45220
rect 9996 45890 10052 45902
rect 9996 45838 9998 45890
rect 10050 45838 10052 45890
rect 9996 45332 10052 45838
rect 9548 44434 9604 44446
rect 9548 44382 9550 44434
rect 9602 44382 9604 44434
rect 9548 43876 9604 44382
rect 9548 43810 9604 43820
rect 9548 43652 9604 43662
rect 9548 42866 9604 43596
rect 9660 43540 9716 45164
rect 9884 44996 9940 45006
rect 9884 44436 9940 44940
rect 9660 43474 9716 43484
rect 9772 44100 9828 44110
rect 9660 43314 9716 43326
rect 9660 43262 9662 43314
rect 9714 43262 9716 43314
rect 9660 43092 9716 43262
rect 9660 43026 9716 43036
rect 9548 42814 9550 42866
rect 9602 42814 9604 42866
rect 9548 42802 9604 42814
rect 9660 42868 9716 42878
rect 9660 42530 9716 42812
rect 9772 42866 9828 44044
rect 9884 43652 9940 44380
rect 9996 43988 10052 45276
rect 10220 45332 10276 46398
rect 10220 45266 10276 45276
rect 10332 46450 10388 46462
rect 10332 46398 10334 46450
rect 10386 46398 10388 46450
rect 9996 43922 10052 43932
rect 10108 45106 10164 45118
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 9884 43586 9940 43596
rect 9772 42814 9774 42866
rect 9826 42814 9828 42866
rect 9772 42802 9828 42814
rect 9996 43092 10052 43102
rect 9660 42478 9662 42530
rect 9714 42478 9716 42530
rect 9660 42466 9716 42478
rect 9100 40402 9156 40908
rect 9100 40350 9102 40402
rect 9154 40350 9156 40402
rect 9100 40338 9156 40350
rect 9212 41132 9324 41188
rect 9380 41132 9492 41188
rect 9548 42196 9604 42206
rect 8652 38782 8654 38834
rect 8706 38782 8708 38834
rect 8652 38770 8708 38782
rect 8764 40012 8932 40068
rect 7980 37772 8596 37828
rect 7980 37156 8036 37772
rect 8316 37604 8372 37614
rect 8092 37380 8148 37390
rect 8092 37378 8260 37380
rect 8092 37326 8094 37378
rect 8146 37326 8260 37378
rect 8092 37324 8260 37326
rect 8092 37314 8148 37324
rect 8204 37268 8260 37324
rect 8204 37202 8260 37212
rect 8316 37156 8372 37548
rect 8540 37604 8596 37614
rect 8428 37156 8484 37166
rect 7980 37100 8148 37156
rect 8316 37154 8484 37156
rect 8316 37102 8430 37154
rect 8482 37102 8484 37154
rect 8316 37100 8484 37102
rect 7868 36866 7924 36876
rect 7532 36654 7534 36706
rect 7586 36654 7588 36706
rect 7532 36642 7588 36654
rect 7756 36820 7812 36830
rect 7420 36082 7476 36092
rect 7756 36036 7812 36764
rect 8092 36820 8148 37100
rect 8428 37090 8484 37100
rect 8092 36754 8148 36764
rect 8204 37044 8260 37054
rect 7868 36596 7924 36606
rect 8204 36596 8260 36988
rect 7868 36594 8260 36596
rect 7868 36542 7870 36594
rect 7922 36542 8260 36594
rect 7868 36540 8260 36542
rect 8316 36596 8372 36606
rect 7868 36530 7924 36540
rect 8316 36502 8372 36540
rect 8204 36372 8260 36382
rect 8204 36278 8260 36316
rect 7756 35980 8372 36036
rect 7980 35700 8036 35710
rect 6972 35646 6974 35698
rect 7026 35646 7028 35698
rect 6972 35634 7028 35646
rect 7756 35698 8036 35700
rect 7756 35646 7982 35698
rect 8034 35646 8036 35698
rect 7756 35644 8036 35646
rect 7756 35588 7812 35644
rect 7980 35634 8036 35644
rect 7308 35532 7812 35588
rect 7196 35364 7252 35374
rect 7308 35308 7364 35532
rect 7868 35476 7924 35486
rect 7196 35252 7364 35308
rect 7420 35364 7476 35374
rect 7084 33348 7140 33358
rect 7084 33254 7140 33292
rect 6748 32398 6750 32450
rect 6802 32398 6804 32450
rect 6748 32386 6804 32398
rect 6860 32900 6916 32910
rect 6636 30718 6638 30770
rect 6690 30718 6692 30770
rect 6636 30660 6692 30718
rect 6636 30594 6692 30604
rect 6636 30212 6692 30222
rect 6636 30118 6692 30156
rect 6412 29538 6580 29540
rect 6412 29486 6414 29538
rect 6466 29486 6580 29538
rect 6412 29484 6580 29486
rect 6412 29474 6468 29484
rect 6076 28642 6132 28700
rect 6076 28590 6078 28642
rect 6130 28590 6132 28642
rect 6076 28578 6132 28590
rect 6636 28868 6692 28878
rect 5852 27806 5854 27858
rect 5906 27806 5908 27858
rect 5516 27636 5572 27646
rect 5404 27188 5460 27198
rect 5292 27186 5460 27188
rect 5292 27134 5406 27186
rect 5458 27134 5460 27186
rect 5292 27132 5460 27134
rect 5404 27122 5460 27132
rect 5404 25844 5460 25854
rect 5516 25844 5572 27580
rect 5740 27524 5796 27534
rect 5460 25788 5572 25844
rect 5628 25844 5684 25854
rect 5404 25778 5460 25788
rect 5180 25622 5348 25678
rect 5292 25620 5348 25622
rect 5292 25554 5348 25564
rect 3804 25116 4068 25126
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 3804 25050 4068 25060
rect 4284 25116 5124 25172
rect 5180 25508 5236 25518
rect 4172 24722 4228 24734
rect 4172 24670 4174 24722
rect 4226 24670 4228 24722
rect 3948 24612 4004 24622
rect 3948 24276 4004 24556
rect 3948 24210 4004 24220
rect 3724 24164 3780 24174
rect 3724 24070 3780 24108
rect 3836 23940 3892 23950
rect 3836 23846 3892 23884
rect 3164 21310 3166 21362
rect 3218 21310 3220 21362
rect 2716 20290 2772 20300
rect 2828 20804 2884 20814
rect 2716 20132 2772 20142
rect 2716 18788 2772 20076
rect 2716 18722 2772 18732
rect 2716 18450 2772 18462
rect 2716 18398 2718 18450
rect 2770 18398 2772 18450
rect 2716 16996 2772 18398
rect 2716 15428 2772 16940
rect 2828 16322 2884 20748
rect 3164 20692 3220 21310
rect 3276 23492 3332 23502
rect 3388 23492 3556 23548
rect 3612 23538 3668 23548
rect 3804 23548 4068 23558
rect 3276 20914 3332 23436
rect 3388 22932 3444 22942
rect 3388 22838 3444 22876
rect 3388 22596 3444 22606
rect 3388 21924 3444 22540
rect 3388 21858 3444 21868
rect 3500 21140 3556 23492
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4172 23548 4228 24670
rect 4284 23938 4340 25116
rect 5068 24948 5124 24958
rect 5180 24948 5236 25452
rect 5404 25396 5460 25406
rect 5068 24946 5236 24948
rect 5068 24894 5070 24946
rect 5122 24894 5236 24946
rect 5068 24892 5236 24894
rect 5292 25394 5460 25396
rect 5292 25342 5406 25394
rect 5458 25342 5460 25394
rect 5292 25340 5460 25342
rect 5292 25060 5348 25340
rect 5404 25330 5460 25340
rect 5628 25396 5684 25788
rect 5628 25330 5684 25340
rect 5068 24882 5124 24892
rect 4956 24610 5012 24622
rect 4956 24558 4958 24610
rect 5010 24558 5012 24610
rect 4844 24388 4900 24398
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23874 4340 23886
rect 4732 23826 4788 23838
rect 4732 23774 4734 23826
rect 4786 23774 4788 23826
rect 4172 23492 4676 23548
rect 3804 23482 4068 23492
rect 3612 23380 3668 23390
rect 3612 22370 3668 23324
rect 4060 23268 4116 23278
rect 4060 23174 4116 23212
rect 3724 22932 3780 22942
rect 4172 22932 4228 22942
rect 3724 22930 4004 22932
rect 3724 22878 3726 22930
rect 3778 22878 4004 22930
rect 3724 22876 4004 22878
rect 3724 22866 3780 22876
rect 3612 22318 3614 22370
rect 3666 22318 3668 22370
rect 3612 22306 3668 22318
rect 3724 22482 3780 22494
rect 3724 22430 3726 22482
rect 3778 22430 3780 22482
rect 3724 22372 3780 22430
rect 3724 22306 3780 22316
rect 3948 22372 4004 22876
rect 4620 22932 4676 23492
rect 4732 23492 4788 23774
rect 4732 23426 4788 23436
rect 4844 23156 4900 24332
rect 4956 23548 5012 24558
rect 5068 24164 5124 24174
rect 5068 24050 5124 24108
rect 5292 24052 5348 25004
rect 5516 25284 5572 25294
rect 5516 24946 5572 25228
rect 5516 24894 5518 24946
rect 5570 24894 5572 24946
rect 5516 24882 5572 24894
rect 5628 24836 5684 24846
rect 5404 24610 5460 24622
rect 5404 24558 5406 24610
rect 5458 24558 5460 24610
rect 5404 24164 5460 24558
rect 5516 24612 5572 24622
rect 5516 24518 5572 24556
rect 5628 24388 5684 24780
rect 5404 24098 5460 24108
rect 5516 24332 5684 24388
rect 5068 23998 5070 24050
rect 5122 23998 5124 24050
rect 5068 23828 5124 23998
rect 5068 23762 5124 23772
rect 5180 23996 5348 24052
rect 4956 23492 5124 23548
rect 4844 23090 4900 23100
rect 4620 22876 4900 22932
rect 4172 22838 4228 22876
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4844 22708 4900 22876
rect 4844 22642 4900 22652
rect 3948 22306 4004 22316
rect 4172 22370 4228 22382
rect 4172 22318 4174 22370
rect 4226 22318 4228 22370
rect 4172 22148 4228 22318
rect 3500 21074 3556 21084
rect 3612 22092 4228 22148
rect 4956 22372 5012 22382
rect 3276 20862 3278 20914
rect 3330 20862 3332 20914
rect 3276 20850 3332 20862
rect 3612 20804 3668 22092
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 4172 21812 4228 21822
rect 3164 20626 3220 20636
rect 3500 20802 3668 20804
rect 3500 20750 3614 20802
rect 3666 20750 3668 20802
rect 3500 20748 3668 20750
rect 4060 21140 4116 21150
rect 4060 20804 4116 21084
rect 4172 21028 4228 21756
rect 4284 21700 4340 21710
rect 4956 21700 5012 22316
rect 5068 21924 5124 23492
rect 5068 21858 5124 21868
rect 5180 23156 5236 23996
rect 5404 23938 5460 23950
rect 5404 23886 5406 23938
rect 5458 23886 5460 23938
rect 4956 21644 5124 21700
rect 4284 21606 4340 21644
rect 4956 21364 5012 21374
rect 4844 21362 5012 21364
rect 4844 21310 4958 21362
rect 5010 21310 5012 21362
rect 4844 21308 5012 21310
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4464 21130 4728 21140
rect 4284 21028 4340 21038
rect 4172 21026 4340 21028
rect 4172 20974 4286 21026
rect 4338 20974 4340 21026
rect 4172 20972 4340 20974
rect 4284 20962 4340 20972
rect 4732 20916 4788 20926
rect 4732 20822 4788 20860
rect 4172 20804 4228 20814
rect 4060 20802 4228 20804
rect 4060 20750 4174 20802
rect 4226 20750 4228 20802
rect 4060 20748 4228 20750
rect 3276 20468 3332 20478
rect 3276 19906 3332 20412
rect 3276 19854 3278 19906
rect 3330 19854 3332 19906
rect 3276 19842 3332 19854
rect 3164 19236 3220 19246
rect 3164 19234 3332 19236
rect 3164 19182 3166 19234
rect 3218 19182 3332 19234
rect 3164 19180 3332 19182
rect 3164 19170 3220 19180
rect 3164 18340 3220 18350
rect 3164 18246 3220 18284
rect 2828 16270 2830 16322
rect 2882 16270 2884 16322
rect 2828 16258 2884 16270
rect 2940 17666 2996 17678
rect 2940 17614 2942 17666
rect 2994 17614 2996 17666
rect 2716 15334 2772 15372
rect 2828 15876 2884 15886
rect 2156 13858 2212 14028
rect 2156 13806 2158 13858
rect 2210 13806 2212 13858
rect 2156 13794 2212 13806
rect 2492 14028 2660 14084
rect 2716 14084 2772 14094
rect 2380 13300 2436 13310
rect 2268 13188 2324 13198
rect 2268 13094 2324 13132
rect 2268 12628 2324 12638
rect 2156 12404 2212 12414
rect 2156 12066 2212 12348
rect 2156 12014 2158 12066
rect 2210 12014 2212 12066
rect 2156 12002 2212 12014
rect 2156 10612 2212 10622
rect 2044 10610 2212 10612
rect 2044 10558 2158 10610
rect 2210 10558 2212 10610
rect 2044 10556 2212 10558
rect 2156 10546 2212 10556
rect 1932 10500 1988 10510
rect 1820 10276 1876 10286
rect 1708 9826 1764 9838
rect 1708 9774 1710 9826
rect 1762 9774 1764 9826
rect 1708 9156 1764 9774
rect 1708 9090 1764 9100
rect 1708 8932 1764 8942
rect 1820 8932 1876 10220
rect 1932 9042 1988 10444
rect 2268 10052 2324 12572
rect 2380 10276 2436 13244
rect 2492 12964 2548 14028
rect 2604 13524 2660 13534
rect 2604 13430 2660 13468
rect 2492 12898 2548 12908
rect 2716 12962 2772 14028
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2604 12066 2660 12078
rect 2604 12014 2606 12066
rect 2658 12014 2660 12066
rect 2380 10210 2436 10220
rect 2492 11396 2548 11406
rect 2492 10052 2548 11340
rect 1932 8990 1934 9042
rect 1986 8990 1988 9042
rect 1932 8978 1988 8990
rect 2044 9996 2324 10052
rect 2380 9996 2548 10052
rect 1708 8930 1876 8932
rect 1708 8878 1710 8930
rect 1762 8878 1876 8930
rect 1708 8876 1876 8878
rect 1708 8866 1764 8876
rect 2044 8708 2100 9996
rect 1596 8306 1652 8316
rect 1932 8652 2100 8708
rect 2156 9828 2212 9838
rect 1484 6850 1540 6860
rect 1596 8146 1652 8158
rect 1596 8094 1598 8146
rect 1650 8094 1652 8146
rect 1596 8036 1652 8094
rect 1596 7586 1652 7980
rect 1596 7534 1598 7586
rect 1650 7534 1652 7586
rect 1484 6692 1540 6702
rect 1596 6692 1652 7534
rect 1484 6690 1652 6692
rect 1484 6638 1486 6690
rect 1538 6638 1652 6690
rect 1484 6636 1652 6638
rect 1484 6626 1540 6636
rect 1372 6290 1428 6300
rect 1260 6078 1262 6130
rect 1314 6078 1316 6130
rect 1260 6066 1316 6078
rect 1372 6132 1428 6142
rect 1372 5346 1428 6076
rect 1596 6020 1652 6636
rect 1596 5954 1652 5964
rect 1708 8148 1764 8158
rect 1372 5294 1374 5346
rect 1426 5294 1428 5346
rect 1372 5282 1428 5294
rect 1708 5236 1764 8092
rect 1708 5170 1764 5180
rect 1820 8036 1876 8046
rect 1820 4452 1876 7980
rect 1932 7028 1988 8652
rect 2044 8484 2100 8494
rect 2044 8390 2100 8428
rect 2044 8260 2100 8270
rect 2044 7362 2100 8204
rect 2044 7310 2046 7362
rect 2098 7310 2100 7362
rect 2044 7298 2100 7310
rect 1932 6972 2100 7028
rect 1932 6804 1988 6814
rect 1932 6710 1988 6748
rect 1932 5236 1988 5246
rect 2044 5236 2100 6972
rect 1932 5234 2100 5236
rect 1932 5182 1934 5234
rect 1986 5182 2100 5234
rect 1932 5180 2100 5182
rect 1932 5170 1988 5180
rect 1820 4396 1988 4452
rect 1372 4338 1428 4350
rect 1372 4286 1374 4338
rect 1426 4286 1428 4338
rect 1372 4116 1428 4286
rect 1820 4228 1876 4238
rect 1820 4134 1876 4172
rect 1372 4050 1428 4060
rect 1372 3780 1428 3790
rect 1372 3686 1428 3724
rect 1596 3556 1652 3566
rect 1596 3462 1652 3500
rect 1932 3388 1988 4396
rect 2044 3780 2100 3790
rect 2156 3780 2212 9772
rect 2268 7476 2324 7486
rect 2268 4228 2324 7420
rect 2380 6468 2436 9996
rect 2492 9828 2548 9838
rect 2492 9734 2548 9772
rect 2380 6402 2436 6412
rect 2492 9604 2548 9614
rect 2380 5908 2436 5918
rect 2380 5794 2436 5852
rect 2380 5742 2382 5794
rect 2434 5742 2436 5794
rect 2380 5730 2436 5742
rect 2492 5348 2548 9548
rect 2492 5282 2548 5292
rect 2380 5124 2436 5134
rect 2380 5122 2548 5124
rect 2380 5070 2382 5122
rect 2434 5070 2548 5122
rect 2380 5068 2548 5070
rect 2380 5058 2436 5068
rect 2268 4162 2324 4172
rect 2380 4900 2436 4910
rect 2380 4116 2436 4844
rect 2380 4050 2436 4060
rect 2044 3778 2212 3780
rect 2044 3726 2046 3778
rect 2098 3726 2212 3778
rect 2044 3724 2212 3726
rect 2044 3714 2100 3724
rect 2380 3556 2436 3566
rect 2380 3462 2436 3500
rect 1932 3332 2212 3388
rect 1148 2942 1150 2994
rect 1202 2942 1204 2994
rect 1148 2930 1204 2942
rect 1036 2716 1652 2772
rect 588 2604 756 2660
rect 476 2594 532 2604
rect 700 112 756 2604
rect 1596 2210 1652 2716
rect 1596 2158 1598 2210
rect 1650 2158 1652 2210
rect 1596 2146 1652 2158
rect 2156 2212 2212 3332
rect 2268 2772 2324 2782
rect 2268 2658 2324 2716
rect 2268 2606 2270 2658
rect 2322 2606 2324 2658
rect 2268 2594 2324 2606
rect 2268 2212 2324 2222
rect 2156 2210 2324 2212
rect 2156 2158 2270 2210
rect 2322 2158 2324 2210
rect 2156 2156 2324 2158
rect 2268 2146 2324 2156
rect 1932 1986 1988 1998
rect 1932 1934 1934 1986
rect 1986 1934 1988 1986
rect 1372 1874 1428 1886
rect 1372 1822 1374 1874
rect 1426 1822 1428 1874
rect 1372 1764 1428 1822
rect 1372 1698 1428 1708
rect 1932 1764 1988 1934
rect 1932 1698 1988 1708
rect 2044 1988 2100 1998
rect 1148 1540 1204 1550
rect 1036 1204 1092 1214
rect 1036 1110 1092 1148
rect 1148 112 1204 1484
rect 1596 1540 1652 1550
rect 1372 1092 1428 1102
rect 1372 998 1428 1036
rect 1596 112 1652 1484
rect 1820 1204 1876 1214
rect 1820 1110 1876 1148
rect 2044 1090 2100 1932
rect 2492 1426 2548 5068
rect 2604 4564 2660 12014
rect 2716 9604 2772 12910
rect 2828 12068 2884 15820
rect 2828 12002 2884 12012
rect 2828 11620 2884 11630
rect 2940 11620 2996 17614
rect 3164 16548 3220 16558
rect 3052 15428 3108 15438
rect 3052 14530 3108 15372
rect 3052 14478 3054 14530
rect 3106 14478 3108 14530
rect 3052 14084 3108 14478
rect 3052 14018 3108 14028
rect 3164 15316 3220 16492
rect 3276 16212 3332 19180
rect 3388 18564 3444 18574
rect 3388 17890 3444 18508
rect 3388 17838 3390 17890
rect 3442 17838 3444 17890
rect 3388 17826 3444 17838
rect 3388 17108 3444 17118
rect 3500 17108 3556 20748
rect 3612 20738 3668 20748
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 3612 20132 3668 20142
rect 3612 20018 3668 20076
rect 3612 19966 3614 20018
rect 3666 19966 3668 20018
rect 3612 19954 3668 19966
rect 3948 20020 4004 20030
rect 3948 19906 4004 19964
rect 3948 19854 3950 19906
rect 4002 19854 4004 19906
rect 3948 19842 4004 19854
rect 3612 19234 3668 19246
rect 3612 19182 3614 19234
rect 3666 19182 3668 19234
rect 3612 17892 3668 19182
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 4172 18564 4228 20748
rect 4396 20020 4452 20030
rect 4284 19794 4340 19806
rect 4284 19742 4286 19794
rect 4338 19742 4340 19794
rect 4284 18900 4340 19742
rect 4396 19796 4452 19964
rect 4844 20020 4900 21308
rect 4956 21298 5012 21308
rect 4956 20468 5012 20478
rect 4956 20130 5012 20412
rect 4956 20078 4958 20130
rect 5010 20078 5012 20130
rect 4956 20066 5012 20078
rect 4844 19954 4900 19964
rect 4396 19730 4452 19740
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 5068 19346 5124 21644
rect 5180 21588 5236 23100
rect 5292 23828 5348 23838
rect 5292 21588 5348 23772
rect 5404 21812 5460 23886
rect 5516 23042 5572 24332
rect 5516 22990 5518 23042
rect 5570 22990 5572 23042
rect 5516 22978 5572 22990
rect 5628 23940 5684 23950
rect 5404 21746 5460 21756
rect 5292 21532 5460 21588
rect 5180 21522 5236 21532
rect 5292 21362 5348 21374
rect 5292 21310 5294 21362
rect 5346 21310 5348 21362
rect 5068 19294 5070 19346
rect 5122 19294 5124 19346
rect 5068 19282 5124 19294
rect 5180 21140 5236 21150
rect 4284 18834 4340 18844
rect 4620 19234 4676 19246
rect 4620 19182 4622 19234
rect 4674 19182 4676 19234
rect 4620 18788 4676 19182
rect 4620 18722 4676 18732
rect 4172 18498 4228 18508
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 5068 18340 5124 18350
rect 5180 18340 5236 21084
rect 5292 21028 5348 21310
rect 5292 20962 5348 20972
rect 5404 20638 5460 21532
rect 5516 20804 5572 20814
rect 5516 20710 5572 20748
rect 5404 20582 5572 20638
rect 5068 18338 5236 18340
rect 5068 18286 5070 18338
rect 5122 18286 5236 18338
rect 5068 18284 5236 18286
rect 5068 18274 5124 18284
rect 4464 18060 4728 18070
rect 3612 17826 3668 17836
rect 4284 18004 4340 18014
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 5068 18004 5124 18014
rect 3612 17666 3668 17678
rect 3612 17614 3614 17666
rect 3666 17614 3668 17666
rect 3612 17556 3668 17614
rect 3948 17668 4004 17678
rect 3948 17574 4004 17612
rect 3612 17490 3668 17500
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 4284 17220 4340 17948
rect 5068 17666 5124 17948
rect 5068 17614 5070 17666
rect 5122 17614 5124 17666
rect 4396 17554 4452 17566
rect 4396 17502 4398 17554
rect 4450 17502 4452 17554
rect 4396 17444 4452 17502
rect 4396 17378 4452 17388
rect 4732 17554 4788 17566
rect 4732 17502 4734 17554
rect 4786 17502 4788 17554
rect 4732 17444 4788 17502
rect 4732 17378 4788 17388
rect 4284 17154 4340 17164
rect 3388 17106 3556 17108
rect 3388 17054 3390 17106
rect 3442 17054 3556 17106
rect 3388 17052 3556 17054
rect 3388 17042 3444 17052
rect 3724 16882 3780 16894
rect 4284 16884 4340 16894
rect 3724 16830 3726 16882
rect 3778 16830 3780 16882
rect 3388 16772 3444 16782
rect 3388 16436 3444 16716
rect 3724 16548 3780 16830
rect 3724 16482 3780 16492
rect 4060 16882 4340 16884
rect 4060 16830 4286 16882
rect 4338 16830 4340 16882
rect 4060 16828 4340 16830
rect 4060 16548 4116 16828
rect 4284 16818 4340 16828
rect 4172 16660 4228 16670
rect 4172 16566 4228 16604
rect 4396 16660 4452 16670
rect 4396 16658 4900 16660
rect 4396 16606 4398 16658
rect 4450 16606 4900 16658
rect 4396 16604 4900 16606
rect 4396 16594 4452 16604
rect 4060 16482 4116 16492
rect 4464 16492 4728 16502
rect 3612 16436 3668 16446
rect 3388 16370 3444 16380
rect 3500 16380 3612 16436
rect 3276 16156 3444 16212
rect 3276 15986 3332 15998
rect 3276 15934 3278 15986
rect 3330 15934 3332 15986
rect 3276 15876 3332 15934
rect 3276 15810 3332 15820
rect 2828 11618 2996 11620
rect 2828 11566 2830 11618
rect 2882 11566 2996 11618
rect 2828 11564 2996 11566
rect 3052 13524 3108 13534
rect 2828 11554 2884 11564
rect 2940 11060 2996 11070
rect 2940 10610 2996 11004
rect 2940 10558 2942 10610
rect 2994 10558 2996 10610
rect 2940 10546 2996 10558
rect 3052 10164 3108 13468
rect 2716 9538 2772 9548
rect 2828 10108 3108 10164
rect 2716 9042 2772 9054
rect 2716 8990 2718 9042
rect 2770 8990 2772 9042
rect 2716 8596 2772 8990
rect 2716 8530 2772 8540
rect 2828 7700 2884 10108
rect 3052 9828 3108 9838
rect 2828 7634 2884 7644
rect 2940 9826 3108 9828
rect 2940 9774 3054 9826
rect 3106 9774 3108 9826
rect 2940 9772 3108 9774
rect 2828 6020 2884 6030
rect 2828 5926 2884 5964
rect 2940 5796 2996 9772
rect 3052 9762 3108 9772
rect 3052 8932 3108 8942
rect 3052 8484 3108 8876
rect 3052 8418 3108 8428
rect 3164 8260 3220 15260
rect 3276 15314 3332 15326
rect 3276 15262 3278 15314
rect 3330 15262 3332 15314
rect 3276 14756 3332 15262
rect 3276 14690 3332 14700
rect 3388 13636 3444 16156
rect 3500 15764 3556 16380
rect 3612 16370 3668 16380
rect 4172 16436 4228 16446
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4228 16380 4340 16436
rect 4464 16426 4728 16436
rect 4172 16370 4228 16380
rect 4284 16322 4340 16380
rect 4284 16270 4286 16322
rect 4338 16270 4340 16322
rect 4284 16258 4340 16270
rect 3500 15698 3556 15708
rect 3612 16098 3668 16110
rect 3612 16046 3614 16098
rect 3666 16046 3668 16098
rect 3612 15652 3668 16046
rect 4060 16100 4116 16110
rect 4060 16006 4116 16044
rect 3804 15708 4068 15718
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 3612 15586 3668 15596
rect 4172 15540 4228 15550
rect 3724 15426 3780 15438
rect 3724 15374 3726 15426
rect 3778 15374 3780 15426
rect 3500 15314 3556 15326
rect 3500 15262 3502 15314
rect 3554 15262 3556 15314
rect 3500 14868 3556 15262
rect 3612 15316 3668 15326
rect 3724 15316 3780 15374
rect 3668 15260 3780 15316
rect 4172 15314 4228 15484
rect 4172 15262 4174 15314
rect 4226 15262 4228 15314
rect 3612 15250 3668 15260
rect 4172 15250 4228 15262
rect 3948 15204 4004 15242
rect 3948 15138 4004 15148
rect 4060 15090 4116 15102
rect 4060 15038 4062 15090
rect 4114 15038 4116 15090
rect 4060 14980 4116 15038
rect 4060 14914 4116 14924
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 3500 14812 3668 14868
rect 4464 14858 4728 14868
rect 3500 14642 3556 14654
rect 3500 14590 3502 14642
rect 3554 14590 3556 14642
rect 3500 13972 3556 14590
rect 3612 14308 3668 14812
rect 4620 14756 4676 14766
rect 4620 14662 4676 14700
rect 4844 14532 4900 16604
rect 4956 16100 5012 16138
rect 4956 16034 5012 16044
rect 4956 15876 5012 15886
rect 4956 15314 5012 15820
rect 4956 15262 4958 15314
rect 5010 15262 5012 15314
rect 4956 15250 5012 15262
rect 5068 15148 5124 17614
rect 5180 15316 5236 18284
rect 5404 20018 5460 20030
rect 5404 19966 5406 20018
rect 5458 19966 5460 20018
rect 5404 19234 5460 19966
rect 5404 19182 5406 19234
rect 5458 19182 5460 19234
rect 5404 18450 5460 19182
rect 5404 18398 5406 18450
rect 5458 18398 5460 18450
rect 5404 18004 5460 18398
rect 5404 17938 5460 17948
rect 5516 17666 5572 20582
rect 5628 18116 5684 23884
rect 5740 23548 5796 27468
rect 5852 27412 5908 27806
rect 6076 28196 6132 28206
rect 5964 27636 6020 27646
rect 5964 27542 6020 27580
rect 5852 27356 6020 27412
rect 5852 26292 5908 26302
rect 5852 25618 5908 26236
rect 5852 25566 5854 25618
rect 5906 25566 5908 25618
rect 5852 25172 5908 25566
rect 5852 25106 5908 25116
rect 5964 24388 6020 27356
rect 6076 27074 6132 28140
rect 6412 27746 6468 27758
rect 6412 27694 6414 27746
rect 6466 27694 6468 27746
rect 6076 27022 6078 27074
rect 6130 27022 6132 27074
rect 6076 25956 6132 27022
rect 6188 27636 6244 27646
rect 6188 26404 6244 27580
rect 6188 26338 6244 26348
rect 6300 27188 6356 27198
rect 6300 26178 6356 27132
rect 6412 27076 6468 27694
rect 6412 27010 6468 27020
rect 6636 26852 6692 28812
rect 6636 26402 6692 26796
rect 6636 26350 6638 26402
rect 6690 26350 6692 26402
rect 6636 26338 6692 26350
rect 6748 28644 6804 28654
rect 6300 26126 6302 26178
rect 6354 26126 6356 26178
rect 6300 26114 6356 26126
rect 6076 25890 6132 25900
rect 6188 26066 6244 26078
rect 6188 26014 6190 26066
rect 6242 26014 6244 26066
rect 6076 25396 6132 25406
rect 6076 24610 6132 25340
rect 6188 24836 6244 26014
rect 6188 24770 6244 24780
rect 6300 25620 6356 25630
rect 6300 24722 6356 25564
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 6300 24658 6356 24670
rect 6412 25060 6468 25070
rect 6412 24834 6468 25004
rect 6412 24782 6414 24834
rect 6466 24782 6468 24834
rect 6076 24558 6078 24610
rect 6130 24558 6132 24610
rect 6076 24546 6132 24558
rect 5964 24332 6244 24388
rect 6076 24164 6132 24174
rect 6076 24070 6132 24108
rect 5964 23938 6020 23950
rect 5964 23886 5966 23938
rect 6018 23886 6020 23938
rect 5964 23828 6020 23886
rect 5740 23492 5908 23548
rect 5852 22370 5908 23492
rect 5852 22318 5854 22370
rect 5906 22318 5908 22370
rect 5852 21476 5908 22318
rect 5852 21410 5908 21420
rect 5964 20468 6020 23772
rect 6188 21588 6244 24332
rect 6412 23268 6468 24782
rect 6748 24836 6804 28588
rect 6860 27860 6916 32844
rect 7084 31780 7140 31790
rect 7196 31780 7252 35252
rect 7308 34914 7364 34926
rect 7308 34862 7310 34914
rect 7362 34862 7364 34914
rect 7308 32116 7364 34862
rect 7420 33346 7476 35308
rect 7756 34916 7812 34926
rect 7756 34822 7812 34860
rect 7644 33906 7700 33918
rect 7644 33854 7646 33906
rect 7698 33854 7700 33906
rect 7420 33294 7422 33346
rect 7474 33294 7476 33346
rect 7420 33282 7476 33294
rect 7532 33460 7588 33470
rect 7308 32060 7476 32116
rect 6860 27794 6916 27804
rect 6972 31778 7252 31780
rect 6972 31726 7086 31778
rect 7138 31726 7252 31778
rect 6972 31724 7252 31726
rect 7308 31892 7364 31902
rect 6860 27300 6916 27310
rect 6860 26740 6916 27244
rect 6972 27076 7028 31724
rect 7084 31714 7140 31724
rect 7196 30996 7252 31006
rect 6972 26982 7028 27020
rect 7084 30212 7140 30222
rect 7084 28642 7140 30156
rect 7084 28590 7086 28642
rect 7138 28590 7140 28642
rect 6860 26674 6916 26684
rect 7084 26516 7140 28590
rect 7196 27858 7252 30940
rect 7196 27806 7198 27858
rect 7250 27806 7252 27858
rect 7196 27412 7252 27806
rect 7196 27346 7252 27356
rect 7308 26740 7364 31836
rect 7420 30212 7476 32060
rect 7532 31890 7588 33404
rect 7644 32228 7700 33854
rect 7756 33796 7812 33806
rect 7756 32340 7812 33740
rect 7756 32274 7812 32284
rect 7644 32162 7700 32172
rect 7868 32116 7924 35420
rect 7980 35026 8036 35038
rect 7980 34974 7982 35026
rect 8034 34974 8036 35026
rect 7980 34804 8036 34974
rect 8092 35028 8148 35038
rect 8092 34934 8148 34972
rect 7980 34738 8036 34748
rect 8092 34132 8148 34142
rect 8092 33458 8148 34076
rect 8092 33406 8094 33458
rect 8146 33406 8148 33458
rect 8092 33394 8148 33406
rect 8204 33906 8260 33918
rect 8204 33854 8206 33906
rect 8258 33854 8260 33906
rect 8204 33346 8260 33854
rect 8316 33684 8372 35980
rect 8428 34580 8484 34590
rect 8428 34020 8484 34524
rect 8428 33954 8484 33964
rect 8316 33628 8484 33684
rect 8204 33294 8206 33346
rect 8258 33294 8260 33346
rect 8204 33282 8260 33294
rect 8428 33124 8484 33628
rect 8428 33058 8484 33068
rect 7980 32788 8036 32798
rect 7980 32694 8036 32732
rect 8428 32676 8484 32686
rect 8316 32674 8484 32676
rect 8316 32622 8430 32674
rect 8482 32622 8484 32674
rect 8316 32620 8484 32622
rect 8204 32340 8260 32350
rect 8316 32340 8372 32620
rect 8428 32610 8484 32620
rect 8260 32284 8372 32340
rect 8428 32452 8484 32462
rect 8204 32274 8260 32284
rect 7868 32050 7924 32060
rect 7532 31838 7534 31890
rect 7586 31838 7588 31890
rect 7532 31826 7588 31838
rect 7644 31892 7700 31902
rect 7980 31892 8036 31902
rect 8204 31892 8260 31902
rect 7644 31890 7812 31892
rect 7644 31838 7646 31890
rect 7698 31838 7812 31890
rect 7644 31836 7812 31838
rect 7644 31826 7700 31836
rect 7420 30146 7476 30156
rect 7644 31556 7700 31566
rect 7420 29876 7476 29886
rect 7420 29426 7476 29820
rect 7420 29374 7422 29426
rect 7474 29374 7476 29426
rect 7420 28980 7476 29374
rect 7644 29316 7700 31500
rect 7756 30770 7812 31836
rect 7756 30718 7758 30770
rect 7810 30718 7812 30770
rect 7756 30212 7812 30718
rect 7868 31778 7924 31790
rect 7868 31726 7870 31778
rect 7922 31726 7924 31778
rect 7868 30436 7924 31726
rect 7980 30660 8036 31836
rect 7980 30594 8036 30604
rect 8092 31890 8260 31892
rect 8092 31838 8206 31890
rect 8258 31838 8260 31890
rect 8092 31836 8260 31838
rect 7868 30370 7924 30380
rect 7756 30118 7812 30156
rect 7868 29986 7924 29998
rect 7868 29934 7870 29986
rect 7922 29934 7924 29986
rect 7868 29876 7924 29934
rect 7868 29810 7924 29820
rect 8092 29876 8148 31836
rect 8204 31826 8260 31836
rect 8316 31780 8372 31790
rect 8428 31780 8484 32396
rect 8316 31778 8484 31780
rect 8316 31726 8318 31778
rect 8370 31726 8484 31778
rect 8316 31724 8484 31726
rect 8316 31714 8372 31724
rect 8204 31554 8260 31566
rect 8204 31502 8206 31554
rect 8258 31502 8260 31554
rect 8204 31444 8260 31502
rect 8204 31378 8260 31388
rect 8316 31556 8372 31566
rect 8204 31108 8260 31118
rect 8316 31108 8372 31500
rect 8540 31332 8596 37548
rect 8652 35924 8708 35934
rect 8652 33796 8708 35868
rect 8652 33730 8708 33740
rect 8764 34468 8820 40012
rect 8876 39844 8932 39854
rect 8876 39730 8932 39788
rect 8876 39678 8878 39730
rect 8930 39678 8932 39730
rect 8876 39666 8932 39678
rect 9212 39618 9268 41132
rect 9324 41122 9380 41132
rect 9548 41076 9604 42140
rect 9996 41858 10052 43036
rect 10108 42532 10164 45054
rect 10332 44884 10388 46398
rect 10444 45220 10500 53228
rect 10668 53284 10724 53294
rect 10556 53060 10612 53070
rect 10668 53060 10724 53228
rect 10556 53058 10724 53060
rect 10556 53006 10558 53058
rect 10610 53006 10724 53058
rect 10556 53004 10724 53006
rect 10556 52994 10612 53004
rect 10892 52836 10948 52846
rect 10668 52834 10948 52836
rect 10668 52782 10894 52834
rect 10946 52782 10948 52834
rect 10668 52780 10948 52782
rect 10556 52724 10612 52734
rect 10556 51604 10612 52668
rect 10556 51538 10612 51548
rect 10556 51268 10612 51278
rect 10668 51268 10724 52780
rect 10892 52770 10948 52780
rect 11004 52836 11060 52846
rect 10556 51266 10668 51268
rect 10556 51214 10558 51266
rect 10610 51214 10668 51266
rect 10556 51212 10668 51214
rect 10556 51202 10612 51212
rect 10668 51174 10724 51212
rect 10668 50370 10724 50382
rect 10668 50318 10670 50370
rect 10722 50318 10724 50370
rect 10556 49810 10612 49822
rect 10556 49758 10558 49810
rect 10610 49758 10612 49810
rect 10556 49028 10612 49758
rect 10668 49812 10724 50318
rect 10668 49028 10724 49756
rect 11004 49700 11060 52780
rect 11452 52500 11508 54348
rect 11676 54338 11732 54348
rect 11900 54404 11956 54462
rect 11900 54338 11956 54348
rect 12012 54068 12068 56028
rect 13244 56018 13300 56030
rect 13468 55970 13524 56700
rect 13468 55918 13470 55970
rect 13522 55918 13524 55970
rect 13468 55906 13524 55918
rect 12460 55860 12516 55870
rect 12460 55858 12628 55860
rect 12460 55806 12462 55858
rect 12514 55806 12628 55858
rect 12460 55804 12628 55806
rect 12460 55794 12516 55804
rect 12124 55410 12180 55422
rect 12124 55358 12126 55410
rect 12178 55358 12180 55410
rect 12124 54964 12180 55358
rect 12460 55410 12516 55422
rect 12460 55358 12462 55410
rect 12514 55358 12516 55410
rect 12460 55076 12516 55358
rect 12572 55300 12628 55804
rect 13132 55468 13524 55524
rect 12796 55300 12852 55310
rect 13020 55300 13076 55310
rect 12572 55298 12852 55300
rect 12572 55246 12798 55298
rect 12850 55246 12852 55298
rect 12572 55244 12852 55246
rect 12460 55010 12516 55020
rect 12796 55076 12852 55244
rect 12796 55010 12852 55020
rect 12908 55298 13076 55300
rect 12908 55246 13022 55298
rect 13074 55246 13076 55298
rect 12908 55244 13076 55246
rect 12124 54898 12180 54908
rect 12124 54628 12180 54638
rect 12124 54626 12404 54628
rect 12124 54574 12126 54626
rect 12178 54574 12404 54626
rect 12124 54572 12404 54574
rect 12124 54562 12180 54572
rect 12348 54516 12404 54572
rect 12796 54516 12852 54526
rect 12348 54514 12852 54516
rect 12348 54462 12798 54514
rect 12850 54462 12852 54514
rect 12348 54460 12852 54462
rect 12796 54450 12852 54460
rect 11788 54012 12068 54068
rect 12236 54402 12292 54414
rect 12236 54350 12238 54402
rect 12290 54350 12292 54402
rect 11676 53730 11732 53742
rect 11676 53678 11678 53730
rect 11730 53678 11732 53730
rect 11676 52836 11732 53678
rect 11788 53060 11844 54012
rect 11788 52994 11844 53004
rect 12012 53732 12068 53742
rect 11676 52770 11732 52780
rect 11116 52444 11508 52500
rect 11116 52386 11172 52444
rect 11116 52334 11118 52386
rect 11170 52334 11172 52386
rect 11116 52322 11172 52334
rect 11004 49634 11060 49644
rect 11116 52052 11172 52062
rect 10780 49028 10836 49038
rect 10668 49026 10836 49028
rect 10668 48974 10782 49026
rect 10834 48974 10836 49026
rect 10668 48972 10836 48974
rect 10556 48962 10612 48972
rect 10556 48244 10612 48254
rect 10780 48244 10836 48972
rect 11116 48692 11172 51996
rect 11452 51492 11508 52444
rect 12012 52388 12068 53676
rect 12236 53172 12292 54350
rect 12684 54180 12740 54190
rect 12460 53732 12516 53742
rect 12460 53638 12516 53676
rect 12684 53732 12740 54124
rect 12684 53666 12740 53676
rect 12236 53116 12516 53172
rect 12124 52948 12180 52958
rect 12348 52948 12404 52958
rect 12124 52946 12348 52948
rect 12124 52894 12126 52946
rect 12178 52894 12348 52946
rect 12124 52892 12348 52894
rect 12124 52882 12180 52892
rect 12348 52882 12404 52892
rect 12460 52388 12516 53116
rect 11900 52332 12068 52388
rect 12348 52332 12516 52388
rect 12572 52388 12628 52398
rect 12908 52388 12964 55244
rect 13020 55234 13076 55244
rect 13020 54740 13076 54750
rect 13020 54514 13076 54684
rect 13132 54628 13188 55468
rect 13468 55410 13524 55468
rect 13468 55358 13470 55410
rect 13522 55358 13524 55410
rect 13468 55346 13524 55358
rect 13580 55298 13636 55310
rect 13580 55246 13582 55298
rect 13634 55246 13636 55298
rect 13132 54562 13188 54572
rect 13244 55186 13300 55198
rect 13244 55134 13246 55186
rect 13298 55134 13300 55186
rect 13020 54462 13022 54514
rect 13074 54462 13076 54514
rect 13020 54450 13076 54462
rect 13244 54516 13300 55134
rect 13356 54516 13412 54526
rect 13244 54514 13412 54516
rect 13244 54462 13358 54514
rect 13410 54462 13412 54514
rect 13244 54460 13412 54462
rect 13356 54450 13412 54460
rect 13132 54290 13188 54302
rect 13132 54238 13134 54290
rect 13186 54238 13188 54290
rect 12572 52386 12964 52388
rect 12572 52334 12574 52386
rect 12626 52334 12964 52386
rect 12572 52332 12964 52334
rect 13020 53730 13076 53742
rect 13020 53678 13022 53730
rect 13074 53678 13076 53730
rect 11788 52164 11844 52174
rect 11452 51426 11508 51436
rect 11564 52050 11620 52062
rect 11564 51998 11566 52050
rect 11618 51998 11620 52050
rect 11340 50596 11396 50606
rect 11340 50502 11396 50540
rect 11340 50372 11396 50382
rect 11340 49810 11396 50316
rect 11340 49758 11342 49810
rect 11394 49758 11396 49810
rect 11116 48626 11172 48636
rect 11228 49586 11284 49598
rect 11228 49534 11230 49586
rect 11282 49534 11284 49586
rect 11228 48468 11284 49534
rect 11340 49588 11396 49758
rect 11340 49522 11396 49532
rect 10556 48242 10836 48244
rect 10556 48190 10558 48242
rect 10610 48190 10836 48242
rect 10556 48188 10836 48190
rect 10892 48412 11284 48468
rect 11340 49026 11396 49038
rect 11340 48974 11342 49026
rect 11394 48974 11396 49026
rect 10556 47570 10612 48188
rect 10556 47518 10558 47570
rect 10610 47518 10612 47570
rect 10556 47506 10612 47518
rect 10668 48020 10724 48030
rect 10556 46564 10612 46574
rect 10556 46470 10612 46508
rect 10668 46452 10724 47964
rect 10668 46386 10724 46396
rect 10892 45780 10948 48412
rect 11004 48244 11060 48254
rect 11004 46562 11060 48188
rect 11228 48244 11284 48254
rect 11228 48150 11284 48188
rect 11340 47908 11396 48974
rect 11564 48580 11620 51998
rect 11676 52052 11732 52062
rect 11676 51602 11732 51996
rect 11676 51550 11678 51602
rect 11730 51550 11732 51602
rect 11676 51538 11732 51550
rect 11564 48514 11620 48524
rect 11676 50932 11732 50942
rect 11116 47852 11396 47908
rect 11116 47796 11172 47852
rect 11116 47730 11172 47740
rect 11228 47684 11284 47694
rect 11228 47068 11284 47628
rect 11452 47684 11508 47694
rect 11340 47460 11396 47470
rect 11452 47460 11508 47628
rect 11676 47572 11732 50876
rect 11788 50594 11844 52108
rect 11788 50542 11790 50594
rect 11842 50542 11844 50594
rect 11788 50530 11844 50542
rect 11788 49812 11844 49822
rect 11788 49718 11844 49756
rect 11340 47458 11508 47460
rect 11340 47406 11342 47458
rect 11394 47406 11508 47458
rect 11340 47404 11508 47406
rect 11564 47516 11732 47572
rect 11340 47394 11396 47404
rect 11228 47012 11508 47068
rect 11004 46510 11006 46562
rect 11058 46510 11060 46562
rect 11004 46452 11060 46510
rect 11004 46386 11060 46396
rect 11116 46674 11172 46686
rect 11116 46622 11118 46674
rect 11170 46622 11172 46674
rect 11004 45892 11060 45902
rect 11004 45798 11060 45836
rect 10780 45724 10948 45780
rect 10668 45668 10724 45678
rect 10668 45574 10724 45612
rect 10444 45164 10724 45220
rect 10332 44818 10388 44828
rect 10444 44882 10500 44894
rect 10444 44830 10446 44882
rect 10498 44830 10500 44882
rect 10332 44100 10388 44110
rect 10108 42466 10164 42476
rect 10220 43316 10276 43326
rect 9996 41806 9998 41858
rect 10050 41806 10052 41858
rect 9996 41794 10052 41806
rect 9660 41748 9716 41758
rect 9660 41654 9716 41692
rect 9436 41020 9604 41076
rect 9660 41300 9716 41310
rect 9324 40404 9380 40414
rect 9324 40290 9380 40348
rect 9324 40238 9326 40290
rect 9378 40238 9380 40290
rect 9324 40226 9380 40238
rect 9212 39566 9214 39618
rect 9266 39566 9268 39618
rect 9212 39554 9268 39566
rect 9100 38834 9156 38846
rect 9100 38782 9102 38834
rect 9154 38782 9156 38834
rect 8988 38612 9044 38622
rect 8876 38164 8932 38174
rect 8876 38070 8932 38108
rect 8988 38162 9044 38556
rect 8988 38110 8990 38162
rect 9042 38110 9044 38162
rect 8988 38098 9044 38110
rect 8876 37604 8932 37614
rect 9100 37604 9156 38782
rect 9212 38724 9268 38762
rect 9212 38658 9268 38668
rect 8932 37548 9156 37604
rect 9212 38164 9268 38174
rect 8876 37538 8932 37548
rect 9212 37492 9268 38108
rect 9324 38052 9380 38062
rect 9324 37958 9380 37996
rect 8988 37436 9268 37492
rect 8876 36594 8932 36606
rect 8876 36542 8878 36594
rect 8930 36542 8932 36594
rect 8876 36372 8932 36542
rect 8876 36306 8932 36316
rect 8988 36036 9044 37436
rect 9436 37380 9492 41020
rect 9660 40404 9716 41244
rect 9884 41300 9940 41310
rect 9884 41298 10052 41300
rect 9884 41246 9886 41298
rect 9938 41246 10052 41298
rect 9884 41244 10052 41246
rect 9884 41234 9940 41244
rect 9772 41188 9828 41198
rect 9772 41094 9828 41132
rect 9772 40404 9828 40414
rect 9660 40402 9828 40404
rect 9660 40350 9774 40402
rect 9826 40350 9828 40402
rect 9660 40348 9828 40350
rect 9660 38834 9716 40348
rect 9772 40338 9828 40348
rect 9772 39732 9828 39742
rect 9772 39618 9828 39676
rect 9772 39566 9774 39618
rect 9826 39566 9828 39618
rect 9772 39554 9828 39566
rect 9884 39730 9940 39742
rect 9884 39678 9886 39730
rect 9938 39678 9940 39730
rect 9884 38948 9940 39678
rect 9884 38882 9940 38892
rect 9660 38782 9662 38834
rect 9714 38782 9716 38834
rect 9660 38770 9716 38782
rect 9772 38724 9828 38734
rect 9772 38612 9940 38668
rect 9548 38500 9604 38510
rect 9548 38274 9604 38444
rect 9548 38222 9550 38274
rect 9602 38222 9604 38274
rect 9548 38210 9604 38222
rect 9772 38050 9828 38062
rect 9772 37998 9774 38050
rect 9826 37998 9828 38050
rect 9660 37938 9716 37950
rect 9660 37886 9662 37938
rect 9714 37886 9716 37938
rect 9660 37604 9716 37886
rect 9660 37538 9716 37548
rect 8988 35812 9044 35980
rect 8876 35756 9044 35812
rect 9100 37324 9492 37380
rect 8876 35308 8932 35756
rect 8988 35588 9044 35598
rect 8988 35494 9044 35532
rect 8876 35252 9044 35308
rect 8764 33236 8820 34412
rect 8876 33236 8932 33246
rect 8764 33234 8932 33236
rect 8764 33182 8878 33234
rect 8930 33182 8932 33234
rect 8764 33180 8932 33182
rect 8876 32900 8932 33180
rect 8876 32834 8932 32844
rect 8764 32562 8820 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 32228 8820 32510
rect 8988 32564 9044 35252
rect 8988 32498 9044 32508
rect 8764 32162 8820 32172
rect 8876 31666 8932 31678
rect 8876 31614 8878 31666
rect 8930 31614 8932 31666
rect 8876 31332 8932 31614
rect 8596 31276 8820 31332
rect 8540 31266 8596 31276
rect 8204 31106 8372 31108
rect 8204 31054 8206 31106
rect 8258 31054 8372 31106
rect 8204 31052 8372 31054
rect 8204 31042 8260 31052
rect 8540 30996 8596 31006
rect 8540 30902 8596 30940
rect 8764 30996 8820 31276
rect 8876 31266 8932 31276
rect 8988 30996 9044 31006
rect 8764 30994 9044 30996
rect 8764 30942 8990 30994
rect 9042 30942 9044 30994
rect 8764 30940 9044 30942
rect 8428 30660 8484 30670
rect 8204 30100 8260 30110
rect 8204 30006 8260 30044
rect 8316 29988 8372 29998
rect 8316 29894 8372 29932
rect 8092 29810 8148 29820
rect 7756 29316 7812 29326
rect 7644 29314 7812 29316
rect 7644 29262 7758 29314
rect 7810 29262 7812 29314
rect 7644 29260 7812 29262
rect 7756 29250 7812 29260
rect 7420 28914 7476 28924
rect 7532 28754 7588 28766
rect 7532 28702 7534 28754
rect 7586 28702 7588 28754
rect 7532 28532 7588 28702
rect 7756 28644 7812 28654
rect 7532 28466 7588 28476
rect 7644 28642 7812 28644
rect 7644 28590 7758 28642
rect 7810 28590 7812 28642
rect 7644 28588 7812 28590
rect 7644 26908 7700 28588
rect 7756 28578 7812 28588
rect 8204 28644 8260 28654
rect 8204 28550 8260 28588
rect 8316 28420 8372 28430
rect 8204 28418 8372 28420
rect 8204 28366 8318 28418
rect 8370 28366 8372 28418
rect 8204 28364 8372 28366
rect 7980 28196 8036 28206
rect 7868 27972 7924 27982
rect 7756 27860 7812 27870
rect 7756 27298 7812 27804
rect 7756 27246 7758 27298
rect 7810 27246 7812 27298
rect 7756 27234 7812 27246
rect 7868 27298 7924 27916
rect 7980 27858 8036 28140
rect 7980 27806 7982 27858
rect 8034 27806 8036 27858
rect 7980 27524 8036 27806
rect 7980 27458 8036 27468
rect 7868 27246 7870 27298
rect 7922 27246 7924 27298
rect 7868 27234 7924 27246
rect 7980 27188 8036 27198
rect 7980 27094 8036 27132
rect 7868 27076 7924 27086
rect 7868 26964 7924 27020
rect 7868 26908 8036 26964
rect 7644 26852 7812 26908
rect 7308 26674 7364 26684
rect 7644 26740 7700 26750
rect 7084 26460 7364 26516
rect 7196 26180 7252 26190
rect 7084 25956 7140 25966
rect 6972 25620 7028 25630
rect 6972 25526 7028 25564
rect 6860 24836 6916 24846
rect 6748 24780 6860 24836
rect 6860 24742 6916 24780
rect 6524 24498 6580 24510
rect 6524 24446 6526 24498
rect 6578 24446 6580 24498
rect 6524 24164 6580 24446
rect 6524 24098 6580 24108
rect 6748 23938 6804 23950
rect 6748 23886 6750 23938
rect 6802 23886 6804 23938
rect 6748 23716 6804 23886
rect 6748 23650 6804 23660
rect 7084 23938 7140 25900
rect 7084 23886 7086 23938
rect 7138 23886 7140 23938
rect 6860 23604 6916 23614
rect 6748 23380 6804 23390
rect 6860 23380 6916 23548
rect 6748 23378 6916 23380
rect 6748 23326 6750 23378
rect 6802 23326 6916 23378
rect 6748 23324 6916 23326
rect 6748 23314 6804 23324
rect 6412 23202 6468 23212
rect 6972 23268 7028 23278
rect 6188 21522 6244 21532
rect 6524 23156 6580 23166
rect 6524 22258 6580 23100
rect 6524 22206 6526 22258
rect 6578 22206 6580 22258
rect 6524 21252 6580 22206
rect 6972 22482 7028 23212
rect 6972 22430 6974 22482
rect 7026 22430 7028 22482
rect 6748 21476 6804 21486
rect 6748 21382 6804 21420
rect 6972 21364 7028 22430
rect 7084 22260 7140 23886
rect 7196 22820 7252 26124
rect 7308 25844 7364 26460
rect 7644 26402 7700 26684
rect 7644 26350 7646 26402
rect 7698 26350 7700 26402
rect 7644 26338 7700 26350
rect 7420 26180 7476 26190
rect 7420 25844 7476 26124
rect 7364 25788 7476 25844
rect 7756 25844 7812 26796
rect 7868 26516 7924 26526
rect 7868 25844 7924 26460
rect 7980 25956 8036 26908
rect 8204 26404 8260 28364
rect 8316 28354 8372 28364
rect 8428 27636 8484 30604
rect 8764 30660 8820 30940
rect 8988 30930 9044 30940
rect 9100 30772 9156 37324
rect 9772 37268 9828 37998
rect 9884 38050 9940 38612
rect 9884 37998 9886 38050
rect 9938 37998 9940 38050
rect 9884 37986 9940 37998
rect 9436 37212 9828 37268
rect 9884 37268 9940 37278
rect 9324 36932 9380 36942
rect 9212 36708 9268 36718
rect 9212 36614 9268 36652
rect 9324 35698 9380 36876
rect 9436 36706 9492 37212
rect 9660 37044 9716 37054
rect 9660 36950 9716 36988
rect 9772 36932 9828 36942
rect 9436 36654 9438 36706
rect 9490 36654 9492 36706
rect 9436 36642 9492 36654
rect 9660 36820 9716 36830
rect 9660 36706 9716 36764
rect 9660 36654 9662 36706
rect 9714 36654 9716 36706
rect 9660 36642 9716 36654
rect 9772 36594 9828 36876
rect 9772 36542 9774 36594
rect 9826 36542 9828 36594
rect 9772 36530 9828 36542
rect 9436 36484 9492 36494
rect 9436 35924 9492 36428
rect 9436 35858 9492 35868
rect 9548 36372 9604 36382
rect 9324 35646 9326 35698
rect 9378 35646 9380 35698
rect 9324 35634 9380 35646
rect 9324 34804 9380 34814
rect 9324 33906 9380 34748
rect 9324 33854 9326 33906
rect 9378 33854 9380 33906
rect 9212 33346 9268 33358
rect 9212 33294 9214 33346
rect 9266 33294 9268 33346
rect 9212 32788 9268 33294
rect 9212 32722 9268 32732
rect 9212 32564 9268 32574
rect 9212 32470 9268 32508
rect 9212 32228 9268 32238
rect 9212 31778 9268 32172
rect 9324 31892 9380 33854
rect 9436 32452 9492 32462
rect 9436 32358 9492 32396
rect 9324 31826 9380 31836
rect 9212 31726 9214 31778
rect 9266 31726 9268 31778
rect 9212 30996 9268 31726
rect 9548 31668 9604 36316
rect 9772 35698 9828 35710
rect 9772 35646 9774 35698
rect 9826 35646 9828 35698
rect 9772 34244 9828 35646
rect 9772 34178 9828 34188
rect 9884 34130 9940 37212
rect 9996 36932 10052 41244
rect 10220 40516 10276 43260
rect 10332 41860 10388 44044
rect 10444 43428 10500 44830
rect 10668 44436 10724 45164
rect 10668 44370 10724 44380
rect 10668 44098 10724 44110
rect 10668 44046 10670 44098
rect 10722 44046 10724 44098
rect 10668 43988 10724 44046
rect 10780 44100 10836 45724
rect 10780 44034 10836 44044
rect 10892 45556 10948 45566
rect 10668 43922 10724 43932
rect 10892 43708 10948 45500
rect 11004 45332 11060 45342
rect 11116 45332 11172 46622
rect 11452 46116 11508 47012
rect 11564 46228 11620 47516
rect 11788 46674 11844 46686
rect 11788 46622 11790 46674
rect 11842 46622 11844 46674
rect 11788 46452 11844 46622
rect 11788 46386 11844 46396
rect 11564 46172 11844 46228
rect 11452 46060 11620 46116
rect 11564 46002 11620 46060
rect 11564 45950 11566 46002
rect 11618 45950 11620 46002
rect 11564 45938 11620 45950
rect 11452 45890 11508 45902
rect 11452 45838 11454 45890
rect 11506 45838 11508 45890
rect 11004 45330 11284 45332
rect 11004 45278 11006 45330
rect 11058 45278 11284 45330
rect 11004 45276 11284 45278
rect 11004 45266 11060 45276
rect 11228 44324 11284 45276
rect 11340 45106 11396 45118
rect 11340 45054 11342 45106
rect 11394 45054 11396 45106
rect 11340 44772 11396 45054
rect 11340 44706 11396 44716
rect 11340 44324 11396 44334
rect 11228 44322 11396 44324
rect 11228 44270 11342 44322
rect 11394 44270 11396 44322
rect 11228 44268 11396 44270
rect 11340 44258 11396 44268
rect 11116 44154 11172 44166
rect 11116 44102 11118 44154
rect 11170 44102 11172 44154
rect 11116 43988 11172 44102
rect 11116 43922 11172 43932
rect 10780 43652 10836 43662
rect 10892 43652 11060 43708
rect 10780 43558 10836 43596
rect 11004 43586 11060 43596
rect 11340 43652 11396 43662
rect 11340 43558 11396 43596
rect 10444 43362 10500 43372
rect 10556 43540 10612 43550
rect 10444 42980 10500 42990
rect 10556 42980 10612 43484
rect 11452 43540 11508 45838
rect 11676 45220 11732 45230
rect 11564 44996 11620 45006
rect 11564 44902 11620 44940
rect 11564 44772 11620 44782
rect 11564 43876 11620 44716
rect 11676 44324 11732 45164
rect 11788 44996 11844 46172
rect 11900 45220 11956 52332
rect 12012 52162 12068 52174
rect 12012 52110 12014 52162
rect 12066 52110 12068 52162
rect 12012 52052 12068 52110
rect 12012 51986 12068 51996
rect 12124 51492 12180 51502
rect 12124 51398 12180 51436
rect 12348 51380 12404 52332
rect 12572 52322 12628 52332
rect 12460 52164 12516 52174
rect 12460 52070 12516 52108
rect 12908 52164 12964 52174
rect 12684 51716 12740 51726
rect 12348 51314 12404 51324
rect 12460 51660 12684 51716
rect 12460 51268 12516 51660
rect 12684 51650 12740 51660
rect 12460 51202 12516 51212
rect 12796 51268 12852 51278
rect 12796 51174 12852 51212
rect 12236 51156 12292 51166
rect 12236 51062 12292 51100
rect 12684 51044 12740 51054
rect 12460 50932 12516 50942
rect 12348 50820 12404 50830
rect 12348 50726 12404 50764
rect 12012 50708 12068 50718
rect 12012 49588 12068 50652
rect 12236 50594 12292 50606
rect 12236 50542 12238 50594
rect 12290 50542 12292 50594
rect 12236 50036 12292 50542
rect 12236 49970 12292 49980
rect 12460 50596 12516 50876
rect 12684 50708 12740 50988
rect 12236 49700 12292 49710
rect 12236 49606 12292 49644
rect 12012 49522 12068 49532
rect 12460 49026 12516 50540
rect 12460 48974 12462 49026
rect 12514 48974 12516 49026
rect 12124 48244 12180 48254
rect 12124 48242 12404 48244
rect 12124 48190 12126 48242
rect 12178 48190 12404 48242
rect 12124 48188 12404 48190
rect 12124 48178 12180 48188
rect 11900 45154 11956 45164
rect 12012 47460 12068 47470
rect 11788 44940 11956 44996
rect 11676 44258 11732 44268
rect 11676 44100 11732 44110
rect 11676 44098 11844 44100
rect 11676 44046 11678 44098
rect 11730 44046 11844 44098
rect 11676 44044 11844 44046
rect 11676 44034 11732 44044
rect 11564 43820 11732 43876
rect 11452 43474 11508 43484
rect 11228 43428 11284 43438
rect 11228 43334 11284 43372
rect 11564 43426 11620 43438
rect 11564 43374 11566 43426
rect 11618 43374 11620 43426
rect 10444 42978 10612 42980
rect 10444 42926 10446 42978
rect 10498 42926 10612 42978
rect 10444 42924 10612 42926
rect 11564 43316 11620 43374
rect 10444 42914 10500 42924
rect 11004 42866 11060 42878
rect 11004 42814 11006 42866
rect 11058 42814 11060 42866
rect 10556 42532 10612 42542
rect 10780 42532 10836 42542
rect 10612 42530 10836 42532
rect 10612 42478 10782 42530
rect 10834 42478 10836 42530
rect 10612 42476 10836 42478
rect 10444 42084 10500 42094
rect 10444 41970 10500 42028
rect 10444 41918 10446 41970
rect 10498 41918 10500 41970
rect 10444 41906 10500 41918
rect 10332 41794 10388 41804
rect 10332 41300 10388 41338
rect 10332 41234 10388 41244
rect 10444 41186 10500 41198
rect 10444 41134 10446 41186
rect 10498 41134 10500 41186
rect 10220 40450 10276 40460
rect 10332 41076 10388 41086
rect 10332 40402 10388 41020
rect 10332 40350 10334 40402
rect 10386 40350 10388 40402
rect 10332 40338 10388 40350
rect 9996 36866 10052 36876
rect 10108 39844 10164 39854
rect 10108 36820 10164 39788
rect 10444 39618 10500 41134
rect 10444 39566 10446 39618
rect 10498 39566 10500 39618
rect 10444 39554 10500 39566
rect 10332 38836 10388 38874
rect 10332 38770 10388 38780
rect 10556 38668 10612 42476
rect 10780 42466 10836 42476
rect 10892 42308 10948 42318
rect 10892 41858 10948 42252
rect 11004 41972 11060 42814
rect 11452 42866 11508 42878
rect 11452 42814 11454 42866
rect 11506 42814 11508 42866
rect 11452 42532 11508 42814
rect 11564 42754 11620 43260
rect 11564 42702 11566 42754
rect 11618 42702 11620 42754
rect 11564 42690 11620 42702
rect 11676 42532 11732 43820
rect 11788 43538 11844 44044
rect 11788 43486 11790 43538
rect 11842 43486 11844 43538
rect 11788 43474 11844 43486
rect 11452 42476 11732 42532
rect 11788 42644 11844 42654
rect 11004 41906 11060 41916
rect 11116 42308 11172 42318
rect 10892 41806 10894 41858
rect 10946 41806 10948 41858
rect 10892 41794 10948 41806
rect 11004 41746 11060 41758
rect 11004 41694 11006 41746
rect 11058 41694 11060 41746
rect 10668 41300 10724 41310
rect 10668 39732 10724 41244
rect 10668 39666 10724 39676
rect 10892 40180 10948 40190
rect 10892 39618 10948 40124
rect 10892 39566 10894 39618
rect 10946 39566 10948 39618
rect 10108 36754 10164 36764
rect 10220 38612 10612 38668
rect 10780 38724 10836 38734
rect 10108 36372 10164 36382
rect 10108 36278 10164 36316
rect 9996 35588 10052 35598
rect 10220 35588 10276 38612
rect 10556 38052 10612 38062
rect 10556 37958 10612 37996
rect 10332 37268 10388 37278
rect 10332 37174 10388 37212
rect 10780 37154 10836 38668
rect 10780 37102 10782 37154
rect 10834 37102 10836 37154
rect 10780 37090 10836 37102
rect 10444 37044 10500 37054
rect 10444 36484 10500 36988
rect 9996 35586 10276 35588
rect 9996 35534 9998 35586
rect 10050 35534 10276 35586
rect 9996 35532 10276 35534
rect 10332 36482 10500 36484
rect 10332 36430 10446 36482
rect 10498 36430 10500 36482
rect 10332 36428 10500 36430
rect 9996 35522 10052 35532
rect 10332 34914 10388 36428
rect 10444 36418 10500 36428
rect 10444 36148 10500 36158
rect 10444 35698 10500 36092
rect 10444 35646 10446 35698
rect 10498 35646 10500 35698
rect 10444 35634 10500 35646
rect 10556 35812 10612 35822
rect 10332 34862 10334 34914
rect 10386 34862 10388 34914
rect 10332 34850 10388 34862
rect 9884 34078 9886 34130
rect 9938 34078 9940 34130
rect 9884 33796 9940 34078
rect 9884 33730 9940 33740
rect 9996 34804 10052 34814
rect 9996 33908 10052 34748
rect 10556 34244 10612 35756
rect 10892 35308 10948 39566
rect 11004 38724 11060 41694
rect 11116 41186 11172 42252
rect 11788 42084 11844 42588
rect 11116 41134 11118 41186
rect 11170 41134 11172 41186
rect 11116 41122 11172 41134
rect 11340 41636 11396 41646
rect 11340 40964 11396 41580
rect 11340 40402 11396 40908
rect 11340 40350 11342 40402
rect 11394 40350 11396 40402
rect 11340 40338 11396 40350
rect 11788 39284 11844 42028
rect 11900 40290 11956 44940
rect 12012 42084 12068 47404
rect 12124 47458 12180 47470
rect 12124 47406 12126 47458
rect 12178 47406 12180 47458
rect 12124 47348 12180 47406
rect 12124 47282 12180 47292
rect 12124 46450 12180 46462
rect 12124 46398 12126 46450
rect 12178 46398 12180 46450
rect 12124 46340 12180 46398
rect 12124 46274 12180 46284
rect 12348 46116 12404 48188
rect 12460 46452 12516 48974
rect 12460 46386 12516 46396
rect 12572 50652 12740 50708
rect 12348 46060 12516 46116
rect 12460 46002 12516 46060
rect 12460 45950 12462 46002
rect 12514 45950 12516 46002
rect 12348 45890 12404 45902
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 12124 44996 12180 45006
rect 12124 44902 12180 44940
rect 12348 44772 12404 45838
rect 12460 45892 12516 45950
rect 12460 45826 12516 45836
rect 12348 44706 12404 44716
rect 12236 44212 12292 44222
rect 12236 44210 12404 44212
rect 12236 44158 12238 44210
rect 12290 44158 12404 44210
rect 12236 44156 12404 44158
rect 12236 44146 12292 44156
rect 12236 43988 12292 43998
rect 12236 43650 12292 43932
rect 12236 43598 12238 43650
rect 12290 43598 12292 43650
rect 12236 43586 12292 43598
rect 12236 43428 12292 43438
rect 12348 43428 12404 44156
rect 12292 43372 12404 43428
rect 12124 43316 12180 43326
rect 12124 43222 12180 43260
rect 12124 42756 12180 42766
rect 12124 42532 12180 42700
rect 12236 42644 12292 43372
rect 12236 42550 12292 42588
rect 12124 42308 12180 42476
rect 12124 42252 12404 42308
rect 12012 42018 12068 42028
rect 12348 42084 12404 42252
rect 12348 42018 12404 42028
rect 12124 41972 12180 41982
rect 12124 41878 12180 41916
rect 12012 41636 12068 41646
rect 12012 41186 12068 41580
rect 12460 41412 12516 41422
rect 12572 41412 12628 50652
rect 12908 50484 12964 52108
rect 13020 52052 13076 53678
rect 13132 53172 13188 54238
rect 13244 54290 13300 54302
rect 13244 54238 13246 54290
rect 13298 54238 13300 54290
rect 13244 53956 13300 54238
rect 13244 53890 13300 53900
rect 13132 53116 13300 53172
rect 13244 53060 13300 53116
rect 13356 53060 13412 53070
rect 13244 53004 13356 53060
rect 13020 51380 13076 51996
rect 13132 52946 13188 52958
rect 13132 52894 13134 52946
rect 13186 52894 13188 52946
rect 13132 52388 13188 52894
rect 13132 51604 13188 52332
rect 13244 52276 13300 52286
rect 13244 52162 13300 52220
rect 13244 52110 13246 52162
rect 13298 52110 13300 52162
rect 13244 51940 13300 52110
rect 13244 51874 13300 51884
rect 13132 51548 13300 51604
rect 13132 51380 13188 51390
rect 13020 51378 13188 51380
rect 13020 51326 13134 51378
rect 13186 51326 13188 51378
rect 13020 51324 13188 51326
rect 13020 50594 13076 51324
rect 13132 51314 13188 51324
rect 13020 50542 13022 50594
rect 13074 50542 13076 50594
rect 13020 50530 13076 50542
rect 12684 50428 12964 50484
rect 12684 48468 12740 50428
rect 13132 49924 13188 49934
rect 13244 49924 13300 51548
rect 13132 49922 13300 49924
rect 13132 49870 13134 49922
rect 13186 49870 13300 49922
rect 13132 49868 13300 49870
rect 13132 49858 13188 49868
rect 13244 49026 13300 49868
rect 13356 49140 13412 53004
rect 13580 52948 13636 55246
rect 13692 54852 13748 57344
rect 14140 57092 14196 57344
rect 14140 57026 14196 57036
rect 14028 56082 14084 56094
rect 14028 56030 14030 56082
rect 14082 56030 14084 56082
rect 13692 54786 13748 54796
rect 13804 55300 13860 55310
rect 13804 54402 13860 55244
rect 13804 54350 13806 54402
rect 13858 54350 13860 54402
rect 13804 54338 13860 54350
rect 13692 53842 13748 53854
rect 13692 53790 13694 53842
rect 13746 53790 13748 53842
rect 13692 53620 13748 53790
rect 13692 53554 13748 53564
rect 13916 53730 13972 53742
rect 13916 53678 13918 53730
rect 13970 53678 13972 53730
rect 13916 53172 13972 53678
rect 14028 53396 14084 56030
rect 14588 56084 14644 57344
rect 14588 56018 14644 56028
rect 14364 55970 14420 55982
rect 14364 55918 14366 55970
rect 14418 55918 14420 55970
rect 14140 54292 14196 54302
rect 14140 54198 14196 54236
rect 14028 53330 14084 53340
rect 14252 53730 14308 53742
rect 14252 53678 14254 53730
rect 14306 53678 14308 53730
rect 13916 53106 13972 53116
rect 13468 52892 13636 52948
rect 13468 51156 13524 52892
rect 13580 52724 13636 52734
rect 13580 52630 13636 52668
rect 14140 52724 14196 52734
rect 13692 52162 13748 52174
rect 13692 52110 13694 52162
rect 13746 52110 13748 52162
rect 13580 51378 13636 51390
rect 13580 51326 13582 51378
rect 13634 51326 13636 51378
rect 13580 51268 13636 51326
rect 13580 51202 13636 51212
rect 13468 51090 13524 51100
rect 13468 50594 13524 50606
rect 13468 50542 13470 50594
rect 13522 50542 13524 50594
rect 13468 49700 13524 50542
rect 13468 49634 13524 49644
rect 13580 49588 13636 49598
rect 13580 49494 13636 49532
rect 13356 49084 13524 49140
rect 13244 48974 13246 49026
rect 13298 48974 13300 49026
rect 12684 48402 12740 48412
rect 12796 48804 12852 48814
rect 12684 47572 12740 47582
rect 12684 45106 12740 47516
rect 12796 47236 12852 48748
rect 13244 48354 13300 48974
rect 13468 48692 13524 49084
rect 13244 48302 13246 48354
rect 13298 48302 13300 48354
rect 13020 47460 13076 47470
rect 13020 47366 13076 47404
rect 12796 47180 13076 47236
rect 12908 46564 12964 46574
rect 12908 45218 12964 46508
rect 12908 45166 12910 45218
rect 12962 45166 12964 45218
rect 12908 45154 12964 45166
rect 12684 45054 12686 45106
rect 12738 45054 12740 45106
rect 12684 45042 12740 45054
rect 13020 45106 13076 47180
rect 13244 47068 13300 48302
rect 13356 48636 13524 48692
rect 13356 47572 13412 48636
rect 13692 48244 13748 52110
rect 13804 51380 13860 51390
rect 13804 51266 13860 51324
rect 13804 51214 13806 51266
rect 13858 51214 13860 51266
rect 13804 51202 13860 51214
rect 14140 50820 14196 52668
rect 14252 51940 14308 53678
rect 14364 52612 14420 55918
rect 15036 55972 15092 57344
rect 15484 56420 15540 57344
rect 15036 55906 15092 55916
rect 15372 56364 15540 56420
rect 14476 55412 14532 55422
rect 14476 55318 14532 55356
rect 14700 55298 14756 55310
rect 14700 55246 14702 55298
rect 14754 55246 14756 55298
rect 14476 54292 14532 54302
rect 14700 54292 14756 55246
rect 15148 55298 15204 55310
rect 15148 55246 15150 55298
rect 15202 55246 15204 55298
rect 14924 54628 14980 54638
rect 14924 54404 14980 54572
rect 14924 54338 14980 54348
rect 14476 54290 14756 54292
rect 14476 54238 14478 54290
rect 14530 54238 14756 54290
rect 14476 54236 14756 54238
rect 15148 54292 15204 55246
rect 15372 55300 15428 56364
rect 15596 55858 15652 55870
rect 15596 55806 15598 55858
rect 15650 55806 15652 55858
rect 15372 55234 15428 55244
rect 15484 55410 15540 55422
rect 15484 55358 15486 55410
rect 15538 55358 15540 55410
rect 15484 54628 15540 55358
rect 15484 54562 15540 54572
rect 15596 55076 15652 55806
rect 15820 55412 15876 55422
rect 15820 55318 15876 55356
rect 14476 54180 14532 54236
rect 15148 54198 15204 54236
rect 14476 54114 14532 54124
rect 15148 53842 15204 53854
rect 15148 53790 15150 53842
rect 15202 53790 15204 53842
rect 15036 53732 15092 53742
rect 14700 53620 14756 53630
rect 14364 52546 14420 52556
rect 14588 53618 14868 53620
rect 14588 53566 14702 53618
rect 14754 53566 14868 53618
rect 14588 53564 14868 53566
rect 14252 51378 14308 51884
rect 14252 51326 14254 51378
rect 14306 51326 14308 51378
rect 14252 51314 14308 51326
rect 14476 52276 14532 52286
rect 14140 50764 14308 50820
rect 13804 50708 13860 50718
rect 13804 49364 13860 50652
rect 14140 50596 14196 50606
rect 14140 49924 14196 50540
rect 14252 50428 14308 50764
rect 14476 50596 14532 52220
rect 14588 50708 14644 53564
rect 14700 53554 14756 53564
rect 14812 53508 14868 53564
rect 15036 53508 15092 53676
rect 14812 53452 15092 53508
rect 15148 53060 15204 53790
rect 15148 52994 15204 53004
rect 15484 53730 15540 53742
rect 15484 53678 15486 53730
rect 15538 53678 15540 53730
rect 14700 52724 14756 52734
rect 14700 52722 14980 52724
rect 14700 52670 14702 52722
rect 14754 52670 14980 52722
rect 14700 52668 14980 52670
rect 14700 52658 14756 52668
rect 14700 52162 14756 52174
rect 14700 52110 14702 52162
rect 14754 52110 14756 52162
rect 14700 51716 14756 52110
rect 14700 51650 14756 51660
rect 14924 51156 14980 52668
rect 15148 52722 15204 52734
rect 15148 52670 15150 52722
rect 15202 52670 15204 52722
rect 15148 52612 15204 52670
rect 15148 52546 15204 52556
rect 15260 52724 15316 52734
rect 15260 52386 15316 52668
rect 15484 52612 15540 53678
rect 15484 52546 15540 52556
rect 15260 52334 15262 52386
rect 15314 52334 15316 52386
rect 15260 52322 15316 52334
rect 15596 52274 15652 55020
rect 15932 54964 15988 57344
rect 16156 55300 16212 55310
rect 16156 55298 16324 55300
rect 16156 55246 16158 55298
rect 16210 55246 16324 55298
rect 16156 55244 16324 55246
rect 16156 55234 16212 55244
rect 15932 54908 16212 54964
rect 16044 54628 16100 54638
rect 16044 54514 16100 54572
rect 16044 54462 16046 54514
rect 16098 54462 16100 54514
rect 16044 54450 16100 54462
rect 15820 54292 15876 54302
rect 15820 54198 15876 54236
rect 15932 53956 15988 53966
rect 15708 53732 15764 53742
rect 15708 53060 15764 53676
rect 15820 53730 15876 53742
rect 15820 53678 15822 53730
rect 15874 53678 15876 53730
rect 15820 53508 15876 53678
rect 15820 53442 15876 53452
rect 15708 52966 15764 53004
rect 15932 52836 15988 53900
rect 16156 53954 16212 54908
rect 16268 54292 16324 55244
rect 16380 54964 16436 57344
rect 16828 56420 16884 57344
rect 16828 56354 16884 56364
rect 16828 55972 16884 55982
rect 16828 55878 16884 55916
rect 16380 54898 16436 54908
rect 16492 55858 16548 55870
rect 16492 55806 16494 55858
rect 16546 55806 16548 55858
rect 16492 54852 16548 55806
rect 17164 55860 17220 55870
rect 17164 55766 17220 55804
rect 16716 55186 16772 55198
rect 16716 55134 16718 55186
rect 16770 55134 16772 55186
rect 16716 55076 16772 55134
rect 17164 55186 17220 55198
rect 17164 55134 17166 55186
rect 17218 55134 17220 55186
rect 16716 55010 16772 55020
rect 16828 55074 16884 55086
rect 16828 55022 16830 55074
rect 16882 55022 16884 55074
rect 16828 54964 16884 55022
rect 17164 55076 17220 55134
rect 17164 55010 17220 55020
rect 16828 54898 16884 54908
rect 16492 54786 16548 54796
rect 16380 54628 16436 54638
rect 16380 54402 16436 54572
rect 17276 54628 17332 57344
rect 17724 56532 17780 57344
rect 18172 56644 18228 57344
rect 18620 56756 18676 57344
rect 18620 56690 18676 56700
rect 18844 56756 18900 56766
rect 18172 56578 18228 56588
rect 17724 56466 17780 56476
rect 18620 56532 18676 56542
rect 17612 56420 17668 56430
rect 17388 56082 17444 56094
rect 17388 56030 17390 56082
rect 17442 56030 17444 56082
rect 17388 55076 17444 56030
rect 17500 55412 17556 55422
rect 17500 55318 17556 55356
rect 17612 55300 17668 56364
rect 17948 56082 18004 56094
rect 17948 56030 17950 56082
rect 18002 56030 18004 56082
rect 17948 55524 18004 56030
rect 18172 56084 18228 56094
rect 18172 55970 18228 56028
rect 18172 55918 18174 55970
rect 18226 55918 18228 55970
rect 18172 55906 18228 55918
rect 18508 55858 18564 55870
rect 18508 55806 18510 55858
rect 18562 55806 18564 55858
rect 18508 55636 18564 55806
rect 17948 55458 18004 55468
rect 18396 55580 18564 55636
rect 17612 55234 17668 55244
rect 17836 55410 17892 55422
rect 17836 55358 17838 55410
rect 17890 55358 17892 55410
rect 17836 55300 17892 55358
rect 17836 55234 17892 55244
rect 18284 55298 18340 55310
rect 18284 55246 18286 55298
rect 18338 55246 18340 55298
rect 17388 55010 17444 55020
rect 17276 54562 17332 54572
rect 18284 54516 18340 55246
rect 18396 55188 18452 55580
rect 18508 55412 18564 55422
rect 18620 55412 18676 56476
rect 18508 55410 18676 55412
rect 18508 55358 18510 55410
rect 18562 55358 18676 55410
rect 18508 55356 18676 55358
rect 18732 56308 18788 56318
rect 18508 55346 18564 55356
rect 18396 55132 18564 55188
rect 18508 55076 18564 55132
rect 18508 55010 18564 55020
rect 18284 54450 18340 54460
rect 16380 54350 16382 54402
rect 16434 54350 16436 54402
rect 16380 54338 16436 54350
rect 18508 54404 18564 54414
rect 18508 54310 18564 54348
rect 16268 54226 16324 54236
rect 17276 54290 17332 54302
rect 17276 54238 17278 54290
rect 17330 54238 17332 54290
rect 16156 53902 16158 53954
rect 16210 53902 16212 53954
rect 16156 53890 16212 53902
rect 16940 53618 16996 53630
rect 16940 53566 16942 53618
rect 16994 53566 16996 53618
rect 16940 53508 16996 53566
rect 16996 53452 17108 53508
rect 16940 53442 16996 53452
rect 16492 53172 16548 53182
rect 16044 52948 16100 52958
rect 16100 52892 16212 52948
rect 16044 52854 16100 52892
rect 15932 52770 15988 52780
rect 15596 52222 15598 52274
rect 15650 52222 15652 52274
rect 15596 52210 15652 52222
rect 15148 52164 15204 52174
rect 15148 52070 15204 52108
rect 15932 52164 15988 52174
rect 15932 52070 15988 52108
rect 16044 52050 16100 52062
rect 16044 51998 16046 52050
rect 16098 51998 16100 52050
rect 15708 51492 15764 51502
rect 15036 51380 15092 51390
rect 15036 51286 15092 51324
rect 15708 51380 15764 51436
rect 15820 51380 15876 51390
rect 15708 51378 15876 51380
rect 15708 51326 15822 51378
rect 15874 51326 15876 51378
rect 15708 51324 15876 51326
rect 15148 51156 15204 51166
rect 14924 51100 15092 51156
rect 14588 50642 14644 50652
rect 14924 50706 14980 50718
rect 14924 50654 14926 50706
rect 14978 50654 14980 50706
rect 14476 50530 14532 50540
rect 14924 50428 14980 50654
rect 14252 50372 14532 50428
rect 14140 49858 14196 49868
rect 13804 49308 14196 49364
rect 13692 48178 13748 48188
rect 13804 49138 13860 49150
rect 13804 49086 13806 49138
rect 13858 49086 13860 49138
rect 13692 48020 13748 48030
rect 13692 47926 13748 47964
rect 13356 47506 13412 47516
rect 13468 47908 13524 47918
rect 13468 47348 13524 47852
rect 13468 47282 13524 47292
rect 13692 47124 13748 47134
rect 13244 47012 13412 47068
rect 13132 46674 13188 46686
rect 13132 46622 13134 46674
rect 13186 46622 13188 46674
rect 13132 45892 13188 46622
rect 13132 45826 13188 45836
rect 13132 45668 13188 45678
rect 13132 45574 13188 45612
rect 13020 45054 13022 45106
rect 13074 45054 13076 45106
rect 13020 45042 13076 45054
rect 13244 45108 13300 45118
rect 13244 45014 13300 45052
rect 12796 44772 12852 44782
rect 12684 44434 12740 44446
rect 12684 44382 12686 44434
rect 12738 44382 12740 44434
rect 12684 43764 12740 44382
rect 12684 43698 12740 43708
rect 12684 43316 12740 43326
rect 12684 42978 12740 43260
rect 12684 42926 12686 42978
rect 12738 42926 12740 42978
rect 12684 42914 12740 42926
rect 12796 42756 12852 44716
rect 13356 44772 13412 47012
rect 13580 46564 13636 46574
rect 13580 46470 13636 46508
rect 13692 46340 13748 47068
rect 13580 46284 13748 46340
rect 13804 46788 13860 49086
rect 14028 47908 14084 47918
rect 13916 47796 13972 47806
rect 13916 47458 13972 47740
rect 13916 47406 13918 47458
rect 13970 47406 13972 47458
rect 13916 47394 13972 47406
rect 14028 46900 14084 47852
rect 13804 46340 13860 46732
rect 13356 44706 13412 44716
rect 13468 45666 13524 45678
rect 13468 45614 13470 45666
rect 13522 45614 13524 45666
rect 12460 41410 12628 41412
rect 12460 41358 12462 41410
rect 12514 41358 12628 41410
rect 12460 41356 12628 41358
rect 12684 42700 12852 42756
rect 13132 44436 13188 44446
rect 12460 41346 12516 41356
rect 12684 41188 12740 42700
rect 12796 42196 12852 42206
rect 12796 41970 12852 42140
rect 12796 41918 12798 41970
rect 12850 41918 12852 41970
rect 12796 41906 12852 41918
rect 12908 42084 12964 42094
rect 12908 41970 12964 42028
rect 12908 41918 12910 41970
rect 12962 41918 12964 41970
rect 12908 41906 12964 41918
rect 13020 41860 13076 41870
rect 12796 41524 12852 41534
rect 12796 41410 12852 41468
rect 12796 41358 12798 41410
rect 12850 41358 12852 41410
rect 12796 41346 12852 41358
rect 12012 41134 12014 41186
rect 12066 41134 12068 41186
rect 12012 41122 12068 41134
rect 12348 41132 12740 41188
rect 12796 41188 12852 41198
rect 11900 40238 11902 40290
rect 11954 40238 11956 40290
rect 11900 40226 11956 40238
rect 12236 40740 12292 40750
rect 12236 40402 12292 40684
rect 12236 40350 12238 40402
rect 12290 40350 12292 40402
rect 11900 39732 11956 39742
rect 11900 39618 11956 39676
rect 11900 39566 11902 39618
rect 11954 39566 11956 39618
rect 11900 39554 11956 39566
rect 11788 39218 11844 39228
rect 11900 39172 11956 39182
rect 11788 39060 11844 39070
rect 11788 38966 11844 39004
rect 11900 38946 11956 39116
rect 11900 38894 11902 38946
rect 11954 38894 11956 38946
rect 11900 38882 11956 38894
rect 11004 38658 11060 38668
rect 11340 38834 11396 38846
rect 11340 38782 11342 38834
rect 11394 38782 11396 38834
rect 11004 38164 11060 38174
rect 11004 38070 11060 38108
rect 11340 37828 11396 38782
rect 12124 38276 12180 38286
rect 12124 38182 12180 38220
rect 11564 38164 11620 38174
rect 11396 37772 11508 37828
rect 11340 37762 11396 37772
rect 11228 37604 11284 37614
rect 11116 36594 11172 36606
rect 11116 36542 11118 36594
rect 11170 36542 11172 36594
rect 11004 36484 11060 36494
rect 11004 36390 11060 36428
rect 10556 34150 10612 34188
rect 10668 35252 10948 35308
rect 11116 35364 11172 36542
rect 11228 35698 11284 37548
rect 11228 35646 11230 35698
rect 11282 35646 11284 35698
rect 11228 35634 11284 35646
rect 11340 36820 11396 36830
rect 11116 35298 11172 35308
rect 9884 33460 9940 33470
rect 9884 33366 9940 33404
rect 9772 33346 9828 33358
rect 9772 33294 9774 33346
rect 9826 33294 9828 33346
rect 9772 33236 9828 33294
rect 9996 33236 10052 33852
rect 9772 33180 10052 33236
rect 10332 33346 10388 33358
rect 10332 33294 10334 33346
rect 10386 33294 10388 33346
rect 9772 32452 9828 33180
rect 9884 32788 9940 32798
rect 9884 32564 9940 32732
rect 9884 32562 10052 32564
rect 9884 32510 9886 32562
rect 9938 32510 10052 32562
rect 9884 32508 10052 32510
rect 9884 32498 9940 32508
rect 9772 32386 9828 32396
rect 9996 32004 10052 32508
rect 10332 32116 10388 33294
rect 10556 33012 10612 33022
rect 10556 32340 10612 32956
rect 10332 32050 10388 32060
rect 10444 32284 10612 32340
rect 10668 32562 10724 35252
rect 11004 35026 11060 35038
rect 11004 34974 11006 35026
rect 11058 34974 11060 35026
rect 10892 34914 10948 34926
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10780 33572 10836 33582
rect 10892 33572 10948 34862
rect 11004 34132 11060 34974
rect 11004 34066 11060 34076
rect 11004 33908 11060 33918
rect 11004 33814 11060 33852
rect 10892 33516 11172 33572
rect 10780 33348 10836 33516
rect 10892 33348 10948 33358
rect 10780 33346 10948 33348
rect 10780 33294 10894 33346
rect 10946 33294 10948 33346
rect 10780 33292 10948 33294
rect 10668 32510 10670 32562
rect 10722 32510 10724 32562
rect 9996 31948 10276 32004
rect 9660 31892 9716 31902
rect 9660 31780 9716 31836
rect 9884 31892 9940 31902
rect 10220 31892 10276 31948
rect 10332 31892 10388 31902
rect 9884 31890 10164 31892
rect 9884 31838 9886 31890
rect 9938 31838 10164 31890
rect 9884 31836 10164 31838
rect 9884 31826 9940 31836
rect 9772 31780 9828 31790
rect 9660 31778 9828 31780
rect 9660 31726 9774 31778
rect 9826 31726 9828 31778
rect 9660 31724 9828 31726
rect 9772 31714 9828 31724
rect 9548 31612 9716 31668
rect 9212 30930 9268 30940
rect 9548 31444 9604 31454
rect 8764 30594 8820 30604
rect 8876 30716 9156 30772
rect 9212 30770 9268 30782
rect 9212 30718 9214 30770
rect 9266 30718 9268 30770
rect 8764 29764 8820 29774
rect 8764 28756 8820 29708
rect 8876 29204 8932 30716
rect 9100 30210 9156 30222
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 8988 30100 9044 30110
rect 8988 29650 9044 30044
rect 8988 29598 8990 29650
rect 9042 29598 9044 29650
rect 8988 29428 9044 29598
rect 8988 29362 9044 29372
rect 9100 29204 9156 30158
rect 9212 29428 9268 30718
rect 9436 30548 9492 30558
rect 9324 30436 9380 30446
rect 9324 30342 9380 30380
rect 9436 30210 9492 30492
rect 9548 30434 9604 31388
rect 9660 30772 9716 31612
rect 9996 31444 10052 31454
rect 9884 30996 9940 31006
rect 9884 30902 9940 30940
rect 9660 30716 9940 30772
rect 9548 30382 9550 30434
rect 9602 30382 9604 30434
rect 9548 30370 9604 30382
rect 9436 30158 9438 30210
rect 9490 30158 9492 30210
rect 9436 30146 9492 30158
rect 9772 30212 9828 30222
rect 9772 30118 9828 30156
rect 9884 29988 9940 30716
rect 9772 29932 9940 29988
rect 9660 29876 9716 29886
rect 9324 29428 9380 29438
rect 9212 29426 9380 29428
rect 9212 29374 9326 29426
rect 9378 29374 9380 29426
rect 9212 29372 9380 29374
rect 9324 29362 9380 29372
rect 9660 29426 9716 29820
rect 9660 29374 9662 29426
rect 9714 29374 9716 29426
rect 9660 29362 9716 29374
rect 9548 29204 9604 29214
rect 8876 29148 9044 29204
rect 9100 29202 9604 29204
rect 9100 29150 9550 29202
rect 9602 29150 9604 29202
rect 9100 29148 9604 29150
rect 8764 28690 8820 28700
rect 8876 28642 8932 28654
rect 8876 28590 8878 28642
rect 8930 28590 8932 28642
rect 8876 27972 8932 28590
rect 8988 28530 9044 29148
rect 9548 29138 9604 29148
rect 9772 28980 9828 29932
rect 9884 29428 9940 29438
rect 9884 29334 9940 29372
rect 9436 28924 9828 28980
rect 9324 28754 9380 28766
rect 9324 28702 9326 28754
rect 9378 28702 9380 28754
rect 9100 28644 9156 28654
rect 9100 28642 9268 28644
rect 9100 28590 9102 28642
rect 9154 28590 9268 28642
rect 9100 28588 9268 28590
rect 9100 28578 9156 28588
rect 8988 28478 8990 28530
rect 9042 28478 9044 28530
rect 8988 28466 9044 28478
rect 8876 27906 8932 27916
rect 9100 28308 9156 28318
rect 8540 27748 8596 27758
rect 8540 27654 8596 27692
rect 8876 27748 8932 27758
rect 8876 27654 8932 27692
rect 8428 27570 8484 27580
rect 8764 27634 8820 27646
rect 8764 27582 8766 27634
rect 8818 27582 8820 27634
rect 8764 27524 8820 27582
rect 8764 27468 9044 27524
rect 8988 27188 9044 27468
rect 8428 27074 8484 27086
rect 8428 27022 8430 27074
rect 8482 27022 8484 27074
rect 8428 26516 8484 27022
rect 8428 26450 8484 26460
rect 8988 26850 9044 27132
rect 8988 26798 8990 26850
rect 9042 26798 9044 26850
rect 8204 26348 8372 26404
rect 8092 26292 8148 26302
rect 8092 26180 8148 26236
rect 8316 26292 8372 26348
rect 8316 26226 8372 26236
rect 8764 26180 8820 26190
rect 8092 26178 8260 26180
rect 8092 26126 8094 26178
rect 8146 26126 8260 26178
rect 8092 26124 8260 26126
rect 8092 26114 8148 26124
rect 8204 25956 8260 26124
rect 7980 25900 8148 25956
rect 7868 25788 8036 25844
rect 7308 25778 7364 25788
rect 7756 25778 7812 25788
rect 7644 25618 7700 25630
rect 7644 25566 7646 25618
rect 7698 25566 7700 25618
rect 7420 25508 7476 25518
rect 7420 25414 7476 25452
rect 7532 25396 7588 25406
rect 7532 25302 7588 25340
rect 7644 24948 7700 25566
rect 7756 25618 7812 25630
rect 7756 25566 7758 25618
rect 7810 25566 7812 25618
rect 7756 25284 7812 25566
rect 7868 25620 7924 25630
rect 7868 25526 7924 25564
rect 7756 25218 7812 25228
rect 7644 24892 7812 24948
rect 7308 24722 7364 24734
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 23716 7364 24670
rect 7644 24724 7700 24734
rect 7644 24630 7700 24668
rect 7756 24612 7812 24892
rect 7308 23650 7364 23660
rect 7420 23940 7476 23950
rect 7420 23156 7476 23884
rect 7756 23604 7812 24556
rect 7868 24498 7924 24510
rect 7868 24446 7870 24498
rect 7922 24446 7924 24498
rect 7868 23940 7924 24446
rect 7868 23874 7924 23884
rect 7756 23538 7812 23548
rect 7868 23716 7924 23726
rect 7420 23090 7476 23100
rect 7868 23154 7924 23660
rect 7868 23102 7870 23154
rect 7922 23102 7924 23154
rect 7196 22754 7252 22764
rect 7532 23042 7588 23054
rect 7532 22990 7534 23042
rect 7586 22990 7588 23042
rect 7532 22596 7588 22990
rect 7868 22932 7924 23102
rect 7980 23156 8036 25788
rect 7980 23090 8036 23100
rect 8092 23938 8148 25900
rect 8204 25890 8260 25900
rect 8764 25508 8820 26124
rect 8988 26180 9044 26798
rect 8988 26114 9044 26124
rect 8764 25442 8820 25452
rect 8428 25284 8484 25294
rect 8092 23886 8094 23938
rect 8146 23886 8148 23938
rect 7868 22876 8036 22932
rect 7084 22204 7252 22260
rect 6972 21298 7028 21308
rect 7084 22036 7140 22046
rect 6524 21196 6804 21252
rect 5964 20402 6020 20412
rect 6300 20802 6356 20814
rect 6524 20804 6580 20814
rect 6300 20750 6302 20802
rect 6354 20750 6356 20802
rect 6300 20468 6356 20750
rect 6300 20402 6356 20412
rect 6412 20748 6524 20804
rect 6188 20244 6244 20254
rect 5740 20020 5796 20030
rect 5740 19926 5796 19964
rect 5964 19794 6020 19806
rect 5964 19742 5966 19794
rect 6018 19742 6020 19794
rect 5852 19684 5908 19694
rect 5852 19460 5908 19628
rect 5852 19234 5908 19404
rect 5964 19348 6020 19742
rect 5964 19282 6020 19292
rect 6076 19346 6132 19358
rect 6076 19294 6078 19346
rect 6130 19294 6132 19346
rect 5852 19182 5854 19234
rect 5906 19182 5908 19234
rect 5852 19170 5908 19182
rect 6076 19236 6132 19294
rect 6076 19170 6132 19180
rect 6188 19012 6244 20188
rect 5964 18956 6244 19012
rect 6300 20020 6356 20030
rect 5852 18564 5908 18574
rect 5852 18450 5908 18508
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5852 18386 5908 18398
rect 5628 18050 5684 18060
rect 5740 17892 5796 17930
rect 5740 17826 5796 17836
rect 5516 17614 5518 17666
rect 5570 17614 5572 17666
rect 5404 16996 5460 17006
rect 5404 16902 5460 16940
rect 5516 16436 5572 17614
rect 5628 17780 5684 17790
rect 5628 16770 5684 17724
rect 5628 16718 5630 16770
rect 5682 16718 5684 16770
rect 5628 16706 5684 16718
rect 5852 17668 5908 17678
rect 5516 16370 5572 16380
rect 5516 16098 5572 16110
rect 5516 16046 5518 16098
rect 5570 16046 5572 16098
rect 5516 15428 5572 16046
rect 5516 15362 5572 15372
rect 5740 15652 5796 15662
rect 5740 15426 5796 15596
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 15362 5796 15374
rect 5180 15250 5236 15260
rect 5292 15204 5348 15242
rect 5068 15092 5236 15148
rect 5292 15138 5348 15148
rect 5180 14756 5236 15092
rect 5180 14690 5236 14700
rect 5292 14980 5348 14990
rect 5292 14644 5348 14924
rect 5852 14756 5908 17612
rect 5964 16996 6020 18956
rect 6076 18788 6132 18798
rect 6076 18338 6132 18732
rect 6076 18286 6078 18338
rect 6130 18286 6132 18338
rect 6076 18274 6132 18286
rect 6188 18452 6244 18462
rect 6188 17778 6244 18396
rect 6188 17726 6190 17778
rect 6242 17726 6244 17778
rect 6188 17714 6244 17726
rect 6300 17556 6356 19964
rect 5964 16882 6020 16940
rect 5964 16830 5966 16882
rect 6018 16830 6020 16882
rect 5964 16818 6020 16830
rect 6188 17500 6356 17556
rect 6412 18564 6468 20748
rect 6524 20738 6580 20748
rect 5740 14700 5908 14756
rect 5964 16660 6020 16670
rect 5964 15652 6020 16604
rect 5292 14588 5404 14644
rect 5348 14542 5404 14588
rect 4284 14476 4900 14532
rect 4956 14532 5012 14542
rect 3836 14308 3892 14318
rect 3612 14252 3836 14308
rect 3836 14242 3892 14252
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 4172 14084 4228 14094
rect 3500 13906 3556 13916
rect 3388 13580 3556 13636
rect 3500 13412 3556 13580
rect 3724 13522 3780 13534
rect 3724 13470 3726 13522
rect 3778 13470 3780 13522
rect 3724 13412 3780 13470
rect 3500 13356 3780 13412
rect 3948 13188 4004 13198
rect 3500 13132 3948 13188
rect 3500 13076 3556 13132
rect 3948 13122 4004 13132
rect 3500 12982 3556 13020
rect 3836 12964 3892 12974
rect 3612 12962 3892 12964
rect 3612 12910 3838 12962
rect 3890 12910 3892 12962
rect 3612 12908 3892 12910
rect 3388 12516 3444 12526
rect 3276 12292 3332 12302
rect 3276 12178 3332 12236
rect 3276 12126 3278 12178
rect 3330 12126 3332 12178
rect 3276 12114 3332 12126
rect 3052 8204 3220 8260
rect 3276 11956 3332 11966
rect 3052 6690 3108 8204
rect 3164 8036 3220 8046
rect 3276 8036 3332 11900
rect 3388 11618 3444 12460
rect 3612 11956 3668 12908
rect 3836 12852 3892 12908
rect 4172 12852 4228 14028
rect 4284 13188 4340 14476
rect 4844 14308 4900 14318
rect 4732 14196 4788 14206
rect 4732 13636 4788 14140
rect 4844 13972 4900 14252
rect 4956 14196 5012 14476
rect 5348 14530 5460 14542
rect 5348 14478 5406 14530
rect 5458 14478 5460 14530
rect 5348 14466 5460 14478
rect 5628 14532 5684 14542
rect 5068 14420 5124 14430
rect 5348 14420 5404 14466
rect 5068 14418 5236 14420
rect 5068 14366 5070 14418
rect 5122 14366 5236 14418
rect 5068 14364 5236 14366
rect 5068 14354 5124 14364
rect 5180 14308 5236 14364
rect 5180 14242 5236 14252
rect 5292 14364 5404 14420
rect 4956 14140 5124 14196
rect 4956 13972 5012 13982
rect 4844 13970 5012 13972
rect 4844 13918 4958 13970
rect 5010 13918 5012 13970
rect 4844 13916 5012 13918
rect 4956 13906 5012 13916
rect 4732 13570 4788 13580
rect 5068 13634 5124 14140
rect 5180 14084 5236 14094
rect 5292 14084 5348 14364
rect 5236 14028 5348 14084
rect 5404 14084 5460 14094
rect 5180 14018 5236 14028
rect 5068 13582 5070 13634
rect 5122 13582 5124 13634
rect 5068 13570 5124 13582
rect 5292 13634 5348 13646
rect 5292 13582 5294 13634
rect 5346 13582 5348 13634
rect 5292 13524 5348 13582
rect 5292 13458 5348 13468
rect 5068 13412 5124 13422
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4508 13188 4564 13198
rect 4284 13186 4564 13188
rect 4284 13134 4510 13186
rect 4562 13134 4564 13186
rect 4284 13132 4564 13134
rect 4508 13122 4564 13132
rect 4620 13076 4676 13086
rect 4396 12964 4452 12974
rect 4620 12964 4676 13020
rect 4396 12962 4676 12964
rect 4396 12910 4398 12962
rect 4450 12910 4676 12962
rect 4396 12908 4676 12910
rect 5068 12962 5124 13356
rect 5068 12910 5070 12962
rect 5122 12910 5124 12962
rect 4396 12898 4452 12908
rect 5068 12898 5124 12910
rect 5404 12852 5460 14028
rect 3836 12796 4228 12852
rect 5180 12796 5460 12852
rect 4508 12628 4564 12638
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4396 12516 4452 12526
rect 3804 12506 4068 12516
rect 4284 12460 4396 12516
rect 3612 11890 3668 11900
rect 3724 12180 3780 12190
rect 3388 11566 3390 11618
rect 3442 11566 3444 11618
rect 3388 11554 3444 11566
rect 3500 11844 3556 11854
rect 3388 10388 3444 10398
rect 3500 10388 3556 11788
rect 3724 11284 3780 12124
rect 3724 11218 3780 11228
rect 4172 12178 4228 12190
rect 4172 12126 4174 12178
rect 4226 12126 4228 12178
rect 4172 12068 4228 12126
rect 4172 11284 4228 12012
rect 4284 11620 4340 12460
rect 4396 12450 4452 12460
rect 4508 12292 4564 12572
rect 4508 12226 4564 12236
rect 4956 12292 5012 12302
rect 4956 12198 5012 12236
rect 5180 12180 5236 12796
rect 5628 12404 5684 14476
rect 5740 12964 5796 14700
rect 5852 14532 5908 14542
rect 5852 14438 5908 14476
rect 5964 13858 6020 15596
rect 6076 16100 6132 16110
rect 6076 15314 6132 16044
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 6076 14980 6132 15262
rect 6076 14914 6132 14924
rect 6076 14644 6132 14654
rect 6076 14550 6132 14588
rect 5964 13806 5966 13858
rect 6018 13806 6020 13858
rect 5964 13794 6020 13806
rect 6076 14308 6132 14318
rect 5740 12962 5908 12964
rect 5740 12910 5742 12962
rect 5794 12910 5908 12962
rect 5740 12908 5908 12910
rect 5740 12898 5796 12908
rect 5516 12348 5684 12404
rect 5740 12516 5796 12526
rect 5404 12292 5460 12302
rect 5516 12292 5572 12348
rect 5404 12290 5572 12292
rect 5404 12238 5406 12290
rect 5458 12238 5572 12290
rect 5404 12236 5572 12238
rect 5404 12226 5460 12236
rect 5180 12114 5236 12124
rect 5628 12180 5684 12190
rect 4844 12068 4900 12078
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4508 11620 4564 11630
rect 4284 11618 4564 11620
rect 4284 11566 4510 11618
rect 4562 11566 4564 11618
rect 4284 11564 4564 11566
rect 4508 11554 4564 11564
rect 4172 11218 4228 11228
rect 4396 11060 4452 11070
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 4172 10948 4228 10958
rect 4172 10836 4228 10892
rect 4060 10780 4228 10836
rect 3612 10612 3668 10622
rect 3612 10518 3668 10556
rect 4060 10610 4116 10780
rect 4396 10722 4452 11004
rect 4396 10670 4398 10722
rect 4450 10670 4452 10722
rect 4396 10658 4452 10670
rect 4060 10558 4062 10610
rect 4114 10558 4116 10610
rect 4060 10546 4116 10558
rect 3500 10332 3668 10388
rect 3388 10294 3444 10332
rect 3612 10052 3668 10332
rect 3500 9996 3668 10052
rect 4172 10276 4228 10286
rect 3164 8034 3332 8036
rect 3164 7982 3166 8034
rect 3218 7982 3332 8034
rect 3164 7980 3332 7982
rect 3388 9940 3444 9950
rect 3388 8036 3444 9884
rect 3500 8932 3556 9996
rect 3724 9940 3780 9950
rect 3500 8866 3556 8876
rect 3612 9938 3780 9940
rect 3612 9886 3726 9938
rect 3778 9886 3780 9938
rect 3612 9884 3780 9886
rect 3612 8820 3668 9884
rect 3724 9874 3780 9884
rect 3948 9828 4004 9838
rect 3948 9734 4004 9772
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 3612 8754 3668 8764
rect 3948 8932 4004 8942
rect 3948 8482 4004 8876
rect 3948 8430 3950 8482
rect 4002 8430 4004 8482
rect 3948 8418 4004 8430
rect 3612 8372 3668 8382
rect 4172 8372 4228 10220
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4732 9940 4788 9950
rect 4732 9846 4788 9884
rect 4396 9826 4452 9838
rect 4396 9774 4398 9826
rect 4450 9774 4452 9826
rect 4284 9604 4340 9614
rect 4284 9266 4340 9548
rect 4396 9380 4452 9774
rect 4396 9314 4452 9324
rect 4284 9214 4286 9266
rect 4338 9214 4340 9266
rect 4284 9202 4340 9214
rect 4284 8932 4340 8942
rect 4284 8596 4340 8876
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 4284 8530 4340 8540
rect 4284 8372 4340 8382
rect 4172 8370 4340 8372
rect 4172 8318 4286 8370
rect 4338 8318 4340 8370
rect 4172 8316 4340 8318
rect 3612 8278 3668 8316
rect 4284 8306 4340 8316
rect 4508 8260 4564 8270
rect 4508 8166 4564 8204
rect 3164 7970 3220 7980
rect 3388 7970 3444 7980
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3164 7700 3220 7710
rect 4844 7700 4900 12012
rect 5068 11956 5124 11966
rect 5068 11954 5460 11956
rect 5068 11902 5070 11954
rect 5122 11902 5460 11954
rect 5068 11900 5460 11902
rect 5068 11890 5124 11900
rect 4956 11620 5012 11630
rect 5180 11620 5236 11630
rect 4956 11394 5012 11564
rect 4956 11342 4958 11394
rect 5010 11342 5012 11394
rect 4956 11330 5012 11342
rect 5068 11564 5180 11620
rect 5068 10612 5124 11564
rect 5180 11554 5236 11564
rect 5068 10546 5124 10556
rect 5180 11396 5236 11406
rect 3164 7606 3220 7644
rect 3836 7644 4900 7700
rect 4956 10498 5012 10510
rect 4956 10446 4958 10498
rect 5010 10446 5012 10498
rect 4956 7698 5012 10446
rect 5068 10388 5124 10398
rect 5068 10294 5124 10332
rect 5180 10164 5236 11340
rect 5404 11394 5460 11900
rect 5628 11732 5684 12124
rect 5740 12178 5796 12460
rect 5740 12126 5742 12178
rect 5794 12126 5796 12178
rect 5740 12114 5796 12126
rect 5852 12068 5908 12908
rect 6076 12180 6132 14252
rect 6188 13524 6244 17500
rect 6300 16436 6356 16446
rect 6300 16100 6356 16380
rect 6300 16006 6356 16044
rect 6188 13458 6244 13468
rect 6300 13746 6356 13758
rect 6300 13694 6302 13746
rect 6354 13694 6356 13746
rect 6188 13076 6244 13086
rect 6188 12292 6244 13020
rect 6300 12516 6356 13694
rect 6412 12964 6468 18508
rect 6524 20018 6580 20030
rect 6524 19966 6526 20018
rect 6578 19966 6580 20018
rect 6524 19234 6580 19966
rect 6524 19182 6526 19234
rect 6578 19182 6580 19234
rect 6524 18452 6580 19182
rect 6524 18358 6580 18396
rect 6636 20020 6692 20030
rect 6636 18228 6692 19964
rect 6636 18162 6692 18172
rect 6524 17220 6580 17230
rect 6524 15428 6580 17164
rect 6748 16100 6804 21196
rect 7084 19234 7140 21980
rect 7196 21924 7252 22204
rect 7532 22036 7588 22540
rect 7980 22148 8036 22876
rect 8092 22708 8148 23886
rect 8316 25228 8428 25284
rect 8316 23154 8372 25228
rect 8428 25218 8484 25228
rect 8316 23102 8318 23154
rect 8370 23102 8372 23154
rect 8316 23090 8372 23102
rect 8428 24722 8484 24734
rect 8428 24670 8430 24722
rect 8482 24670 8484 24722
rect 8428 23268 8484 24670
rect 9100 24722 9156 28252
rect 9212 27858 9268 28588
rect 9324 27970 9380 28702
rect 9324 27918 9326 27970
rect 9378 27918 9380 27970
rect 9324 27906 9380 27918
rect 9212 27806 9214 27858
rect 9266 27806 9268 27858
rect 9212 26514 9268 27806
rect 9212 26462 9214 26514
rect 9266 26462 9268 26514
rect 9212 26450 9268 26462
rect 9100 24670 9102 24722
rect 9154 24670 9156 24722
rect 9100 24658 9156 24670
rect 9212 25394 9268 25406
rect 9212 25342 9214 25394
rect 9266 25342 9268 25394
rect 9212 25284 9268 25342
rect 8988 24164 9044 24174
rect 8988 24070 9044 24108
rect 9212 23716 9268 25228
rect 9324 23940 9380 23950
rect 9324 23846 9380 23884
rect 9100 23660 9268 23716
rect 9324 23716 9380 23726
rect 8428 23212 9044 23268
rect 8092 22642 8148 22652
rect 8092 22148 8148 22158
rect 7980 22146 8148 22148
rect 7980 22094 8094 22146
rect 8146 22094 8148 22146
rect 7980 22092 8148 22094
rect 7532 21980 7924 22036
rect 7196 21868 7700 21924
rect 7196 21586 7252 21598
rect 7196 21534 7198 21586
rect 7250 21534 7252 21586
rect 7196 21364 7252 21534
rect 7196 21298 7252 21308
rect 7532 21588 7588 21598
rect 7196 20018 7252 20030
rect 7196 19966 7198 20018
rect 7250 19966 7252 20018
rect 7196 19796 7252 19966
rect 7196 19730 7252 19740
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 7084 19170 7140 19182
rect 7196 19236 7252 19246
rect 6972 17668 7028 17678
rect 6972 17574 7028 17612
rect 6972 17332 7028 17342
rect 6972 16994 7028 17276
rect 6972 16942 6974 16994
rect 7026 16942 7028 16994
rect 6972 16930 7028 16942
rect 7084 17108 7140 17118
rect 6860 16324 6916 16334
rect 6860 16230 6916 16268
rect 7084 16322 7140 17052
rect 7196 16436 7252 19180
rect 7308 18452 7364 18462
rect 7308 18358 7364 18396
rect 7532 17668 7588 21532
rect 7644 20020 7700 21868
rect 7756 21812 7812 21822
rect 7756 21474 7812 21756
rect 7756 21422 7758 21474
rect 7810 21422 7812 21474
rect 7756 21410 7812 21422
rect 7868 21476 7924 21980
rect 7868 21410 7924 21420
rect 8092 21364 8148 22092
rect 8316 21924 8372 21934
rect 8204 21700 8260 21710
rect 8204 21586 8260 21644
rect 8204 21534 8206 21586
rect 8258 21534 8260 21586
rect 8204 21522 8260 21534
rect 8092 21298 8148 21308
rect 8092 20692 8148 20702
rect 7980 20020 8036 20030
rect 7644 20018 8036 20020
rect 7644 19966 7982 20018
rect 8034 19966 8036 20018
rect 7644 19964 8036 19966
rect 7756 19796 7812 19806
rect 7532 17602 7588 17612
rect 7644 19124 7700 19134
rect 7532 16772 7588 16782
rect 7420 16660 7476 16670
rect 7420 16566 7476 16604
rect 7196 16380 7364 16436
rect 7084 16270 7086 16322
rect 7138 16270 7140 16322
rect 7084 16258 7140 16270
rect 7308 16100 7364 16380
rect 7420 16324 7476 16334
rect 7532 16324 7588 16716
rect 7476 16268 7588 16324
rect 7644 16324 7700 19068
rect 7756 16884 7812 19740
rect 7756 16818 7812 16828
rect 7868 18116 7924 18126
rect 7868 17666 7924 18060
rect 7868 17614 7870 17666
rect 7922 17614 7924 17666
rect 7756 16324 7812 16334
rect 7644 16322 7812 16324
rect 7644 16270 7758 16322
rect 7810 16270 7812 16322
rect 7644 16268 7812 16270
rect 7420 16230 7476 16268
rect 7756 16258 7812 16268
rect 6748 16044 6916 16100
rect 6524 13300 6580 15372
rect 6636 15316 6692 15326
rect 6636 14868 6692 15260
rect 6748 15092 6804 15102
rect 6748 14998 6804 15036
rect 6860 14980 6916 16044
rect 7196 15202 7252 15214
rect 7196 15150 7198 15202
rect 7250 15150 7252 15202
rect 6860 14914 6916 14924
rect 7084 14980 7140 14990
rect 6636 14812 6804 14868
rect 6636 14644 6692 14654
rect 6636 14530 6692 14588
rect 6636 14478 6638 14530
rect 6690 14478 6692 14530
rect 6636 13636 6692 14478
rect 6748 14532 6804 14812
rect 6748 14476 6916 14532
rect 6636 13570 6692 13580
rect 6748 13748 6804 13758
rect 6748 13412 6804 13692
rect 6860 13746 6916 14476
rect 7084 14308 7140 14924
rect 7196 14644 7252 15150
rect 7196 14578 7252 14588
rect 7084 14242 7140 14252
rect 7308 14530 7364 16044
rect 7868 14644 7924 17614
rect 7980 17220 8036 19964
rect 8092 18564 8148 20636
rect 8204 19236 8260 19246
rect 8204 19142 8260 19180
rect 8204 18564 8260 18574
rect 8092 18508 8204 18564
rect 8204 18450 8260 18508
rect 8204 18398 8206 18450
rect 8258 18398 8260 18450
rect 8204 18386 8260 18398
rect 7980 17154 8036 17164
rect 7868 14578 7924 14588
rect 7980 16996 8036 17006
rect 7980 15314 8036 16940
rect 8092 16210 8148 16222
rect 8092 16158 8094 16210
rect 8146 16158 8148 16210
rect 8092 15652 8148 16158
rect 8092 15586 8148 15596
rect 7980 15262 7982 15314
rect 8034 15262 8036 15314
rect 7308 14478 7310 14530
rect 7362 14478 7364 14530
rect 6860 13694 6862 13746
rect 6914 13694 6916 13746
rect 6860 13682 6916 13694
rect 7084 13748 7140 13758
rect 6748 13346 6804 13356
rect 6972 13522 7028 13534
rect 6972 13470 6974 13522
rect 7026 13470 7028 13522
rect 6636 13300 6692 13310
rect 6524 13244 6636 13300
rect 6636 13234 6692 13244
rect 6972 13188 7028 13470
rect 6972 13122 7028 13132
rect 6636 12964 6692 12974
rect 6412 12962 6692 12964
rect 6412 12910 6638 12962
rect 6690 12910 6692 12962
rect 6412 12908 6692 12910
rect 6300 12450 6356 12460
rect 6188 12236 6356 12292
rect 6076 12124 6244 12180
rect 5852 12002 5908 12012
rect 5964 11732 6020 11742
rect 5404 11342 5406 11394
rect 5458 11342 5460 11394
rect 5404 11330 5460 11342
rect 5516 11676 5684 11732
rect 5740 11676 5964 11732
rect 5516 11396 5572 11676
rect 5628 11396 5684 11406
rect 5516 11394 5684 11396
rect 5516 11342 5630 11394
rect 5682 11342 5684 11394
rect 5516 11340 5684 11342
rect 5628 11330 5684 11340
rect 5292 11284 5348 11294
rect 5292 10612 5348 11228
rect 5740 11172 5796 11676
rect 5964 11666 6020 11676
rect 5852 11508 5908 11546
rect 6188 11458 6244 12124
rect 6300 12178 6356 12236
rect 6300 12126 6302 12178
rect 6354 12126 6356 12178
rect 6300 12114 6356 12126
rect 6524 12068 6580 12078
rect 6412 12012 6524 12068
rect 5852 11442 5908 11452
rect 5964 11394 6020 11406
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11284 6020 11342
rect 5628 11116 5796 11172
rect 5852 11228 6020 11284
rect 6132 11402 6244 11458
rect 6300 11956 6356 11966
rect 6300 11508 6356 11900
rect 6412 11954 6468 12012
rect 6524 12002 6580 12012
rect 6412 11902 6414 11954
rect 6466 11902 6468 11954
rect 6412 11890 6468 11902
rect 6636 11844 6692 12908
rect 6524 11788 6692 11844
rect 6748 12964 6804 12974
rect 5628 11060 5684 11116
rect 5628 10994 5684 11004
rect 5628 10836 5684 10846
rect 5292 10546 5348 10556
rect 5516 10612 5572 10622
rect 5516 10518 5572 10556
rect 5292 10388 5348 10426
rect 5292 10322 5348 10332
rect 5068 10108 5236 10164
rect 5292 10164 5348 10174
rect 5068 8260 5124 10108
rect 5292 10052 5348 10108
rect 5180 9996 5348 10052
rect 5180 9154 5236 9996
rect 5292 9828 5348 9838
rect 5292 9734 5348 9772
rect 5180 9102 5182 9154
rect 5234 9102 5236 9154
rect 5180 8932 5236 9102
rect 5180 8866 5236 8876
rect 5628 8930 5684 10780
rect 5628 8878 5630 8930
rect 5682 8878 5684 8930
rect 5292 8708 5348 8718
rect 5348 8652 5460 8708
rect 5292 8642 5348 8652
rect 5292 8372 5348 8382
rect 5180 8260 5236 8270
rect 5068 8204 5180 8260
rect 5180 8166 5236 8204
rect 4956 7646 4958 7698
rect 5010 7646 5012 7698
rect 3612 7364 3668 7374
rect 3612 7270 3668 7308
rect 3388 7028 3444 7038
rect 3388 6804 3444 6972
rect 3836 6914 3892 7644
rect 4956 7634 5012 7646
rect 5292 7588 5348 8316
rect 5068 7532 5348 7588
rect 3948 7476 4004 7486
rect 3948 7382 4004 7420
rect 5068 7474 5124 7532
rect 5068 7422 5070 7474
rect 5122 7422 5124 7474
rect 5068 7410 5124 7422
rect 3836 6862 3838 6914
rect 3890 6862 3892 6914
rect 3836 6850 3892 6862
rect 4172 7364 4228 7374
rect 4172 6916 4228 7308
rect 4284 7362 4340 7374
rect 4284 7310 4286 7362
rect 4338 7310 4340 7362
rect 4284 7140 4340 7310
rect 4396 7364 4452 7374
rect 5404 7364 5460 8652
rect 5628 8484 5684 8878
rect 5852 8932 5908 11228
rect 6132 11172 6188 11402
rect 6076 11116 6188 11172
rect 5964 10612 6020 10622
rect 5964 10518 6020 10556
rect 6076 10500 6132 11116
rect 6300 11060 6356 11452
rect 6076 10434 6132 10444
rect 6188 11004 6356 11060
rect 6412 11732 6580 11788
rect 5852 8866 5908 8876
rect 6076 10276 6132 10286
rect 6188 10276 6244 11004
rect 6300 10836 6356 10846
rect 6300 10610 6356 10780
rect 6300 10558 6302 10610
rect 6354 10558 6356 10610
rect 6300 10546 6356 10558
rect 6132 10220 6244 10276
rect 6300 10276 6356 10286
rect 5628 8418 5684 8428
rect 5740 8820 5796 8830
rect 4396 7270 4452 7308
rect 5180 7308 5460 7364
rect 5516 8260 5572 8270
rect 4844 7252 4900 7262
rect 5180 7252 5236 7308
rect 4284 7074 4340 7084
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4172 6860 4452 6916
rect 3388 6748 3556 6804
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6626 3108 6638
rect 3500 6690 3556 6748
rect 4396 6802 4452 6860
rect 4396 6750 4398 6802
rect 4450 6750 4452 6802
rect 4396 6738 4452 6750
rect 3500 6638 3502 6690
rect 3554 6638 3556 6690
rect 3500 6626 3556 6638
rect 4284 6690 4340 6702
rect 4284 6638 4286 6690
rect 4338 6638 4340 6690
rect 4172 6468 4228 6478
rect 2828 5740 2996 5796
rect 3388 6356 3444 6366
rect 2716 5124 2772 5134
rect 2716 5030 2772 5068
rect 2828 4900 2884 5740
rect 2940 5234 2996 5246
rect 2940 5182 2942 5234
rect 2994 5182 2996 5234
rect 2940 5012 2996 5182
rect 2940 4946 2996 4956
rect 2604 4498 2660 4508
rect 2716 4844 2884 4900
rect 2716 4452 2772 4844
rect 2940 4564 2996 4602
rect 2940 4498 2996 4508
rect 2716 4396 2884 4452
rect 2716 4116 2772 4126
rect 2716 2882 2772 4060
rect 2828 3778 2884 4396
rect 2828 3726 2830 3778
rect 2882 3726 2884 3778
rect 2828 3714 2884 3726
rect 3276 4340 3332 4350
rect 3276 3332 3332 4284
rect 3388 4226 3444 6300
rect 3804 6300 4068 6310
rect 3500 6244 3556 6254
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3500 5794 3556 6188
rect 3500 5742 3502 5794
rect 3554 5742 3556 5794
rect 3500 5730 3556 5742
rect 4060 5908 4116 5918
rect 3836 5684 3892 5694
rect 3836 5590 3892 5628
rect 3612 5124 3668 5134
rect 3612 5030 3668 5068
rect 4060 5122 4116 5852
rect 4060 5070 4062 5122
rect 4114 5070 4116 5122
rect 4060 5058 4116 5070
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 3948 4564 4004 4574
rect 3724 4340 3780 4350
rect 3724 4246 3780 4284
rect 3388 4174 3390 4226
rect 3442 4174 3444 4226
rect 3388 4162 3444 4174
rect 3500 4004 3556 4014
rect 3500 3444 3556 3948
rect 3948 3778 4004 4508
rect 4060 4228 4116 4238
rect 4172 4228 4228 6412
rect 4284 6356 4340 6638
rect 4620 6692 4676 6702
rect 4620 6598 4676 6636
rect 4844 6690 4900 7196
rect 5068 7196 5236 7252
rect 4844 6638 4846 6690
rect 4898 6638 4900 6690
rect 4844 6626 4900 6638
rect 4956 7140 5012 7150
rect 4284 6290 4340 6300
rect 4844 6020 4900 6030
rect 4464 5516 4728 5526
rect 4284 5460 4340 5470
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4284 4900 4340 5404
rect 4284 4844 4676 4900
rect 4396 4676 4452 4686
rect 4396 4338 4452 4620
rect 4620 4452 4676 4844
rect 4620 4386 4676 4396
rect 4396 4286 4398 4338
rect 4450 4286 4452 4338
rect 4396 4274 4452 4286
rect 4508 4340 4564 4350
rect 4060 4226 4228 4228
rect 4060 4174 4062 4226
rect 4114 4174 4228 4226
rect 4060 4172 4228 4174
rect 4060 4162 4116 4172
rect 4508 4116 4564 4284
rect 4284 4060 4564 4116
rect 4844 4116 4900 5964
rect 4956 5122 5012 7084
rect 4956 5070 4958 5122
rect 5010 5070 5012 5122
rect 4956 5058 5012 5070
rect 5068 4338 5124 7196
rect 5404 7140 5460 7150
rect 5516 7140 5572 8204
rect 5628 7476 5684 7486
rect 5628 7382 5684 7420
rect 5460 7084 5572 7140
rect 5628 7140 5684 7150
rect 5404 7074 5460 7084
rect 5292 7028 5348 7038
rect 5292 6690 5348 6972
rect 5292 6638 5294 6690
rect 5346 6638 5348 6690
rect 5292 6626 5348 6638
rect 5516 6580 5572 6590
rect 5180 6468 5236 6478
rect 5180 6018 5236 6412
rect 5180 5966 5182 6018
rect 5234 5966 5236 6018
rect 5180 5954 5236 5966
rect 5292 6356 5348 6366
rect 5180 5796 5236 5806
rect 5180 5572 5236 5740
rect 5180 5506 5236 5516
rect 5292 4340 5348 6300
rect 5516 5794 5572 6524
rect 5628 6356 5684 7084
rect 5628 6290 5684 6300
rect 5516 5742 5518 5794
rect 5570 5742 5572 5794
rect 5516 5730 5572 5742
rect 5628 5348 5684 5358
rect 5740 5348 5796 8764
rect 6076 8820 6132 10220
rect 6300 9828 6356 10220
rect 6076 8754 6132 8764
rect 6188 9826 6356 9828
rect 6188 9774 6302 9826
rect 6354 9774 6356 9826
rect 6188 9772 6356 9774
rect 5964 8260 6020 8270
rect 5852 6468 5908 6478
rect 5852 5796 5908 6412
rect 5964 5908 6020 8204
rect 6188 6690 6244 9772
rect 6300 9762 6356 9772
rect 6412 9828 6468 11732
rect 6636 11620 6692 11630
rect 6636 11394 6692 11564
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11330 6692 11342
rect 6636 10500 6692 10510
rect 6412 9762 6468 9772
rect 6524 10386 6580 10398
rect 6524 10334 6526 10386
rect 6578 10334 6580 10386
rect 6300 8484 6356 8494
rect 6300 8258 6356 8428
rect 6524 8372 6580 10334
rect 6636 9156 6692 10444
rect 6748 9828 6804 12908
rect 6972 12962 7028 12974
rect 6972 12910 6974 12962
rect 7026 12910 7028 12962
rect 6972 12180 7028 12910
rect 6972 12114 7028 12124
rect 7084 12178 7140 13692
rect 7084 12126 7086 12178
rect 7138 12126 7140 12178
rect 7084 12114 7140 12126
rect 7196 12516 7252 12526
rect 6748 9762 6804 9772
rect 6860 12066 6916 12078
rect 6860 12014 6862 12066
rect 6914 12014 6916 12066
rect 6860 10612 6916 12014
rect 6972 11508 7028 11518
rect 6972 11414 7028 11452
rect 6860 9938 6916 10556
rect 7084 10836 7140 10846
rect 6860 9886 6862 9938
rect 6914 9886 6916 9938
rect 6748 9268 6804 9278
rect 6860 9268 6916 9886
rect 6972 10498 7028 10510
rect 6972 10446 6974 10498
rect 7026 10446 7028 10498
rect 6972 9604 7028 10446
rect 6972 9538 7028 9548
rect 6748 9266 6916 9268
rect 6748 9214 6750 9266
rect 6802 9214 6916 9266
rect 6748 9212 6916 9214
rect 6972 9268 7028 9278
rect 6748 9202 6804 9212
rect 6636 8484 6692 9100
rect 6636 8418 6692 8428
rect 6748 8932 6804 8942
rect 6524 8306 6580 8316
rect 6300 8206 6302 8258
rect 6354 8206 6356 8258
rect 6300 8194 6356 8206
rect 6188 6638 6190 6690
rect 6242 6638 6244 6690
rect 6188 6626 6244 6638
rect 6300 7700 6356 7710
rect 5964 5842 6020 5852
rect 6188 6356 6244 6366
rect 5852 5730 5908 5740
rect 5628 5346 5796 5348
rect 5628 5294 5630 5346
rect 5682 5294 5796 5346
rect 5628 5292 5796 5294
rect 5628 5282 5684 5292
rect 5068 4286 5070 4338
rect 5122 4286 5124 4338
rect 5068 4274 5124 4286
rect 5180 4284 5348 4340
rect 5516 5124 5572 5134
rect 4844 4060 5124 4116
rect 3948 3726 3950 3778
rect 4002 3726 4004 3778
rect 3948 3714 4004 3726
rect 4172 4004 4228 4014
rect 3276 3266 3332 3276
rect 3388 3332 3556 3388
rect 3388 3108 3444 3332
rect 2716 2830 2718 2882
rect 2770 2830 2772 2882
rect 2716 2436 2772 2830
rect 3276 3052 3444 3108
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3276 2436 3332 3052
rect 3388 2884 3444 2894
rect 3388 2658 3444 2828
rect 3724 2772 3780 2782
rect 3724 2678 3780 2716
rect 3388 2606 3390 2658
rect 3442 2606 3444 2658
rect 3388 2594 3444 2606
rect 4060 2546 4116 2558
rect 4060 2494 4062 2546
rect 4114 2494 4116 2546
rect 3276 2380 3388 2436
rect 2716 2370 2772 2380
rect 3332 2324 3388 2380
rect 4060 2324 4116 2494
rect 3332 2268 3556 2324
rect 3164 2212 3220 2222
rect 2492 1374 2494 1426
rect 2546 1374 2548 1426
rect 2492 1362 2548 1374
rect 2604 2098 2660 2110
rect 2604 2046 2606 2098
rect 2658 2046 2660 2098
rect 2604 1316 2660 2046
rect 3164 1986 3220 2156
rect 3164 1934 3166 1986
rect 3218 1934 3220 1986
rect 3164 1922 3220 1934
rect 3276 2100 3332 2110
rect 2604 1250 2660 1260
rect 2940 1428 2996 1438
rect 2044 1038 2046 1090
rect 2098 1038 2100 1090
rect 2044 1026 2100 1038
rect 2044 644 2100 654
rect 2044 112 2100 588
rect 2492 644 2548 654
rect 2492 112 2548 588
rect 2940 112 2996 1372
rect 3276 532 3332 2044
rect 3500 2098 3556 2268
rect 4060 2258 4116 2268
rect 3500 2046 3502 2098
rect 3554 2046 3556 2098
rect 3500 2034 3556 2046
rect 3612 1876 3668 1886
rect 3388 1652 3444 1662
rect 3444 1596 3556 1652
rect 3388 1586 3444 1596
rect 3276 466 3332 476
rect 3388 1204 3444 1214
rect 3388 112 3444 1148
rect 3500 980 3556 1596
rect 3612 1090 3668 1820
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 4172 1428 4228 3948
rect 4284 2770 4340 4060
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 5068 3780 5124 4060
rect 5180 3892 5236 4284
rect 5292 4116 5348 4126
rect 5292 4114 5460 4116
rect 5292 4062 5294 4114
rect 5346 4062 5460 4114
rect 5292 4060 5460 4062
rect 5292 4050 5348 4060
rect 5180 3836 5348 3892
rect 5068 3724 5236 3780
rect 5180 3554 5236 3724
rect 5180 3502 5182 3554
rect 5234 3502 5236 3554
rect 4284 2718 4286 2770
rect 4338 2718 4340 2770
rect 4284 2706 4340 2718
rect 4396 3442 4452 3454
rect 4396 3390 4398 3442
rect 4450 3390 4452 3442
rect 4396 2548 4452 3390
rect 5068 3444 5124 3454
rect 4508 2996 4564 3006
rect 4508 2772 4564 2940
rect 4508 2706 4564 2716
rect 5068 2772 5124 3388
rect 5068 2706 5124 2716
rect 4284 2492 4452 2548
rect 4284 2436 4340 2492
rect 4284 2212 4340 2380
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 5068 2324 5124 2334
rect 4284 2156 4452 2212
rect 3612 1038 3614 1090
rect 3666 1038 3668 1090
rect 3612 1026 3668 1038
rect 3836 1372 4228 1428
rect 4396 1540 4452 2156
rect 4732 2100 4788 2110
rect 4732 2006 4788 2044
rect 3500 914 3556 924
rect 3836 112 3892 1372
rect 4172 1204 4228 1214
rect 4396 1204 4452 1484
rect 4172 1202 4452 1204
rect 4172 1150 4174 1202
rect 4226 1150 4452 1202
rect 4172 1148 4452 1150
rect 4508 1876 4564 1886
rect 4172 1138 4228 1148
rect 4508 980 4564 1820
rect 4844 1204 4900 1214
rect 4844 1110 4900 1148
rect 4284 924 4564 980
rect 4284 112 4340 924
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 5068 644 5124 2268
rect 5180 2212 5236 3502
rect 5180 2146 5236 2156
rect 5292 2210 5348 3836
rect 5292 2158 5294 2210
rect 5346 2158 5348 2210
rect 5292 2146 5348 2158
rect 5180 980 5236 990
rect 5180 886 5236 924
rect 4732 588 5124 644
rect 5180 756 5236 766
rect 4732 112 4788 588
rect 5180 112 5236 700
rect 5404 420 5460 4060
rect 5516 1428 5572 5068
rect 5740 5124 5796 5134
rect 5628 4788 5684 4798
rect 5628 4338 5684 4732
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 5628 4274 5684 4286
rect 5628 3892 5684 3902
rect 5628 3778 5684 3836
rect 5628 3726 5630 3778
rect 5682 3726 5684 3778
rect 5628 3714 5684 3726
rect 5628 2996 5684 3006
rect 5740 2996 5796 5068
rect 5964 4114 6020 4126
rect 5964 4062 5966 4114
rect 6018 4062 6020 4114
rect 5964 3108 6020 4062
rect 5964 3042 6020 3052
rect 5628 2994 5796 2996
rect 5628 2942 5630 2994
rect 5682 2942 5796 2994
rect 5628 2940 5796 2942
rect 5628 2930 5684 2940
rect 6188 2100 6244 6300
rect 6300 4900 6356 7644
rect 6412 7588 6468 7598
rect 6412 7474 6468 7532
rect 6412 7422 6414 7474
rect 6466 7422 6468 7474
rect 6412 7410 6468 7422
rect 6412 6916 6468 6926
rect 6412 6468 6468 6860
rect 6412 6402 6468 6412
rect 6636 6690 6692 6702
rect 6636 6638 6638 6690
rect 6690 6638 6692 6690
rect 6636 6580 6692 6638
rect 6636 6356 6692 6524
rect 6636 6290 6692 6300
rect 6412 6132 6468 6142
rect 6412 5796 6468 6076
rect 6748 6130 6804 8876
rect 6748 6078 6750 6130
rect 6802 6078 6804 6130
rect 6748 6066 6804 6078
rect 6860 8258 6916 8270
rect 6860 8206 6862 8258
rect 6914 8206 6916 8258
rect 6412 5740 6580 5796
rect 6300 4834 6356 4844
rect 6524 4338 6580 5740
rect 6748 5572 6804 5582
rect 6636 5460 6692 5470
rect 6636 5012 6692 5404
rect 6748 5346 6804 5516
rect 6860 5460 6916 8206
rect 6972 8260 7028 9212
rect 7084 8596 7140 10780
rect 7196 10610 7252 12460
rect 7308 12180 7364 14478
rect 7868 13972 7924 13982
rect 7420 13748 7476 13758
rect 7420 13654 7476 13692
rect 7756 13188 7812 13198
rect 7868 13188 7924 13916
rect 7980 13746 8036 15262
rect 8092 14868 8148 14878
rect 8092 14530 8148 14812
rect 8092 14478 8094 14530
rect 8146 14478 8148 14530
rect 8092 14466 8148 14478
rect 8316 14084 8372 21868
rect 8428 21586 8484 23212
rect 8988 23154 9044 23212
rect 8988 23102 8990 23154
rect 9042 23102 9044 23154
rect 8988 23090 9044 23102
rect 8540 23044 8596 23054
rect 8540 22950 8596 22988
rect 9100 22820 9156 23660
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 8428 21522 8484 21534
rect 8652 22764 9156 22820
rect 9212 23492 9268 23502
rect 8540 17108 8596 17118
rect 8540 17014 8596 17052
rect 8316 14018 8372 14028
rect 8428 14644 8484 14654
rect 7980 13694 7982 13746
rect 8034 13694 8036 13746
rect 7980 13682 8036 13694
rect 8204 13748 8260 13758
rect 8204 13654 8260 13692
rect 8428 13524 8484 14588
rect 8316 13300 8372 13310
rect 7980 13188 8036 13198
rect 7868 13186 8036 13188
rect 7868 13134 7982 13186
rect 8034 13134 8036 13186
rect 7868 13132 8036 13134
rect 7420 12962 7476 12974
rect 7420 12910 7422 12962
rect 7474 12910 7476 12962
rect 7420 12404 7476 12910
rect 7532 12964 7588 12974
rect 7532 12870 7588 12908
rect 7644 12962 7700 12974
rect 7644 12910 7646 12962
rect 7698 12910 7700 12962
rect 7420 12338 7476 12348
rect 7420 12180 7476 12190
rect 7308 12178 7476 12180
rect 7308 12126 7422 12178
rect 7474 12126 7476 12178
rect 7308 12124 7476 12126
rect 7420 12114 7476 12124
rect 7644 12068 7700 12910
rect 7644 12002 7700 12012
rect 7196 10558 7198 10610
rect 7250 10558 7252 10610
rect 7196 10546 7252 10558
rect 7644 10612 7700 10622
rect 7644 10518 7700 10556
rect 7644 10388 7700 10398
rect 7308 9938 7364 9950
rect 7308 9886 7310 9938
rect 7362 9886 7364 9938
rect 7308 9268 7364 9886
rect 7420 9828 7476 9838
rect 7420 9380 7476 9772
rect 7420 9324 7588 9380
rect 7196 9212 7364 9268
rect 7196 8930 7252 9212
rect 7308 9044 7364 9082
rect 7308 8978 7364 8988
rect 7196 8878 7198 8930
rect 7250 8878 7252 8930
rect 7196 8866 7252 8878
rect 7420 8820 7476 8830
rect 7420 8726 7476 8764
rect 7084 8540 7476 8596
rect 6972 8194 7028 8204
rect 7308 8370 7364 8382
rect 7308 8318 7310 8370
rect 7362 8318 7364 8370
rect 6972 7474 7028 7486
rect 6972 7422 6974 7474
rect 7026 7422 7028 7474
rect 6972 6580 7028 7422
rect 7196 7028 7252 7038
rect 7308 7028 7364 8318
rect 7420 8258 7476 8540
rect 7420 8206 7422 8258
rect 7474 8206 7476 8258
rect 7420 8194 7476 8206
rect 7308 6972 7476 7028
rect 6972 6514 7028 6524
rect 7084 6804 7140 6814
rect 7196 6804 7252 6972
rect 7308 6804 7364 6814
rect 7196 6802 7364 6804
rect 7196 6750 7310 6802
rect 7362 6750 7364 6802
rect 7196 6748 7364 6750
rect 6860 5394 6916 5404
rect 6972 6356 7028 6366
rect 6748 5294 6750 5346
rect 6802 5294 6804 5346
rect 6748 5282 6804 5294
rect 6636 4956 6804 5012
rect 6524 4286 6526 4338
rect 6578 4286 6580 4338
rect 6524 4274 6580 4286
rect 6300 4228 6356 4238
rect 6300 4134 6356 4172
rect 6524 4004 6580 4014
rect 6412 2212 6468 2222
rect 6412 2118 6468 2156
rect 6188 2034 6244 2044
rect 6076 1652 6132 1662
rect 5628 1428 5684 1438
rect 5516 1426 5684 1428
rect 5516 1374 5630 1426
rect 5682 1374 5684 1426
rect 5516 1372 5684 1374
rect 5628 1362 5684 1372
rect 5404 354 5460 364
rect 5628 1204 5684 1214
rect 5628 112 5684 1148
rect 6076 112 6132 1596
rect 6524 112 6580 3948
rect 6748 3778 6804 4956
rect 6972 4676 7028 6300
rect 7084 5906 7140 6748
rect 7308 6738 7364 6748
rect 7084 5854 7086 5906
rect 7138 5854 7140 5906
rect 7084 5842 7140 5854
rect 7308 6468 7364 6478
rect 7420 6468 7476 6972
rect 7532 6690 7588 9324
rect 7644 9042 7700 10332
rect 7756 9380 7812 13132
rect 7980 13122 8036 13132
rect 8092 13076 8148 13086
rect 8092 10276 8148 13020
rect 8204 12962 8260 12974
rect 8204 12910 8206 12962
rect 8258 12910 8260 12962
rect 8204 11844 8260 12910
rect 8204 11778 8260 11788
rect 8204 11620 8260 11630
rect 8204 11526 8260 11564
rect 8204 11284 8260 11294
rect 8204 10276 8260 11228
rect 8316 10612 8372 13244
rect 8428 11284 8484 13468
rect 8652 12852 8708 22764
rect 8764 21588 8820 21598
rect 8764 20804 8820 21532
rect 9212 21364 9268 23436
rect 9212 21298 9268 21308
rect 9324 20998 9380 23660
rect 9436 22036 9492 28924
rect 9884 28532 9940 28542
rect 9884 27970 9940 28476
rect 9996 28308 10052 31388
rect 10108 30210 10164 31836
rect 10220 31890 10388 31892
rect 10220 31838 10334 31890
rect 10386 31838 10388 31890
rect 10220 31836 10388 31838
rect 10220 30996 10276 31836
rect 10332 31826 10388 31836
rect 10220 30930 10276 30940
rect 10332 31668 10388 31678
rect 10332 30994 10388 31612
rect 10332 30942 10334 30994
rect 10386 30942 10388 30994
rect 10332 30436 10388 30942
rect 10332 30370 10388 30380
rect 10108 30158 10110 30210
rect 10162 30158 10164 30210
rect 10108 30146 10164 30158
rect 10220 30212 10276 30222
rect 10220 30118 10276 30156
rect 10332 30210 10388 30222
rect 10332 30158 10334 30210
rect 10386 30158 10388 30210
rect 10332 30100 10388 30158
rect 10332 30034 10388 30044
rect 10332 28532 10388 28542
rect 10332 28438 10388 28476
rect 9996 28242 10052 28252
rect 10108 28420 10164 28430
rect 10108 28084 10164 28364
rect 9884 27918 9886 27970
rect 9938 27918 9940 27970
rect 9660 27524 9716 27534
rect 9548 27076 9604 27086
rect 9548 26740 9604 27020
rect 9548 26674 9604 26684
rect 9660 26516 9716 27468
rect 9548 26460 9716 26516
rect 9772 26516 9828 26526
rect 9548 25396 9604 26460
rect 9772 26422 9828 26460
rect 9660 26292 9716 26302
rect 9660 26198 9716 26236
rect 9772 26180 9828 26190
rect 9772 26086 9828 26124
rect 9660 25620 9716 25630
rect 9660 25618 9828 25620
rect 9660 25566 9662 25618
rect 9714 25566 9828 25618
rect 9660 25564 9828 25566
rect 9660 25554 9716 25564
rect 9548 25340 9716 25396
rect 9548 24050 9604 24062
rect 9548 23998 9550 24050
rect 9602 23998 9604 24050
rect 9548 23604 9604 23998
rect 9548 23538 9604 23548
rect 9660 22932 9716 25340
rect 9772 24836 9828 25564
rect 9884 25284 9940 27918
rect 9884 25218 9940 25228
rect 9996 28028 10164 28084
rect 9996 25508 10052 28028
rect 10220 27746 10276 27758
rect 10220 27694 10222 27746
rect 10274 27694 10276 27746
rect 10108 27300 10164 27310
rect 10108 27206 10164 27244
rect 10220 27118 10276 27694
rect 9772 24276 9828 24780
rect 9996 24722 10052 25452
rect 9996 24670 9998 24722
rect 10050 24670 10052 24722
rect 9996 24658 10052 24670
rect 10108 27062 10276 27118
rect 10332 27748 10388 27758
rect 10108 25956 10164 27062
rect 10332 26514 10388 27692
rect 10332 26462 10334 26514
rect 10386 26462 10388 26514
rect 10332 26450 10388 26462
rect 9772 24210 9828 24220
rect 9884 24050 9940 24062
rect 9884 23998 9886 24050
rect 9938 23998 9940 24050
rect 9772 23156 9828 23166
rect 9772 23062 9828 23100
rect 9884 23044 9940 23998
rect 9884 22978 9940 22988
rect 9996 23716 10052 23726
rect 9436 21970 9492 21980
rect 9548 22876 9716 22932
rect 9548 21588 9604 22876
rect 9548 21140 9604 21532
rect 9548 21074 9604 21084
rect 9660 22708 9716 22718
rect 8764 20738 8820 20748
rect 9212 20942 9380 20998
rect 9100 20690 9156 20702
rect 9100 20638 9102 20690
rect 9154 20638 9156 20690
rect 8764 20020 8820 20030
rect 9100 20020 9156 20638
rect 9212 20692 9268 20942
rect 9436 20914 9492 20926
rect 9436 20862 9438 20914
rect 9490 20862 9492 20914
rect 9212 20626 9268 20636
rect 9324 20804 9380 20814
rect 8764 20018 9156 20020
rect 8764 19966 8766 20018
rect 8818 19966 9156 20018
rect 8764 19964 9156 19966
rect 8764 19954 8820 19964
rect 8876 19234 8932 19246
rect 8876 19182 8878 19234
rect 8930 19182 8932 19234
rect 8876 17892 8932 19182
rect 8988 18338 9044 18350
rect 8988 18286 8990 18338
rect 9042 18286 9044 18338
rect 8988 18116 9044 18286
rect 8988 18050 9044 18060
rect 8876 17826 8932 17836
rect 8652 12786 8708 12796
rect 8764 17668 8820 17678
rect 8764 17332 8820 17612
rect 9100 17668 9156 19964
rect 9212 20132 9268 20142
rect 9212 19906 9268 20076
rect 9212 19854 9214 19906
rect 9266 19854 9268 19906
rect 9212 19842 9268 19854
rect 9212 19460 9268 19470
rect 9212 19366 9268 19404
rect 9324 19458 9380 20748
rect 9436 20020 9492 20862
rect 9660 20916 9716 22652
rect 9996 22484 10052 23660
rect 10108 23548 10164 25900
rect 10220 26178 10276 26190
rect 10220 26126 10222 26178
rect 10274 26126 10276 26178
rect 10220 25060 10276 26126
rect 10332 26180 10388 26190
rect 10332 26086 10388 26124
rect 10220 24994 10276 25004
rect 10444 23828 10500 32284
rect 10556 30210 10612 30222
rect 10556 30158 10558 30210
rect 10610 30158 10612 30210
rect 10556 29988 10612 30158
rect 10668 30100 10724 32510
rect 10892 32116 10948 33292
rect 10892 32050 10948 32060
rect 11004 33124 11060 33134
rect 10780 32004 10836 32014
rect 10780 31780 10836 31948
rect 10892 31780 10948 31790
rect 10780 31778 10948 31780
rect 10780 31726 10894 31778
rect 10946 31726 10948 31778
rect 10780 31724 10948 31726
rect 10892 31714 10948 31724
rect 10668 30034 10724 30044
rect 10780 31332 10836 31342
rect 10556 29922 10612 29932
rect 10780 28980 10836 31276
rect 10892 30436 10948 30446
rect 10892 29876 10948 30380
rect 10892 29810 10948 29820
rect 10780 28914 10836 28924
rect 10892 28868 10948 28878
rect 10780 28754 10836 28766
rect 10780 28702 10782 28754
rect 10834 28702 10836 28754
rect 10668 28308 10724 28318
rect 10668 27076 10724 28252
rect 10668 26982 10724 27020
rect 10780 27300 10836 28702
rect 10892 28308 10948 28812
rect 10892 28242 10948 28252
rect 10780 26964 10836 27244
rect 10780 26898 10836 26908
rect 10892 27636 10948 27646
rect 10108 23492 10388 23548
rect 10220 22708 10276 22718
rect 10220 22594 10276 22652
rect 10220 22542 10222 22594
rect 10274 22542 10276 22594
rect 10220 22530 10276 22542
rect 9772 22428 10164 22484
rect 9772 22370 9828 22428
rect 9772 22318 9774 22370
rect 9826 22318 9828 22370
rect 9772 22306 9828 22318
rect 9884 22148 9940 22158
rect 9772 21588 9828 21598
rect 9772 21494 9828 21532
rect 9660 20850 9716 20860
rect 9436 19954 9492 19964
rect 9772 20692 9828 20702
rect 9324 19406 9326 19458
rect 9378 19406 9380 19458
rect 9324 19394 9380 19406
rect 9772 19796 9828 20636
rect 9884 19908 9940 22092
rect 9884 19842 9940 19852
rect 9996 22036 10052 22046
rect 9772 19346 9828 19740
rect 9772 19294 9774 19346
rect 9826 19294 9828 19346
rect 9436 19234 9492 19246
rect 9436 19182 9438 19234
rect 9490 19182 9492 19234
rect 9324 18452 9380 18462
rect 9324 18358 9380 18396
rect 9100 17574 9156 17612
rect 8540 12740 8596 12750
rect 8540 12178 8596 12684
rect 8540 12126 8542 12178
rect 8594 12126 8596 12178
rect 8540 12114 8596 12126
rect 8652 12516 8708 12526
rect 8428 11218 8484 11228
rect 8316 10546 8372 10556
rect 8428 10948 8484 10958
rect 8204 10220 8372 10276
rect 8092 10210 8148 10220
rect 8204 10052 8260 10062
rect 7868 9826 7924 9838
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9604 7924 9774
rect 7868 9538 7924 9548
rect 7756 9324 8148 9380
rect 7644 8990 7646 9042
rect 7698 8990 7700 9042
rect 7644 8978 7700 8990
rect 7756 9156 7812 9166
rect 7756 8484 7812 9100
rect 7868 9042 7924 9054
rect 7868 8990 7870 9042
rect 7922 8990 7924 9042
rect 7868 8932 7924 8990
rect 7868 8866 7924 8876
rect 7756 8428 8036 8484
rect 7868 8258 7924 8270
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7756 7924 7812 7934
rect 7756 7474 7812 7868
rect 7756 7422 7758 7474
rect 7810 7422 7812 7474
rect 7756 7410 7812 7422
rect 7644 7252 7700 7262
rect 7644 7158 7700 7196
rect 7532 6638 7534 6690
rect 7586 6638 7588 6690
rect 7532 6626 7588 6638
rect 7868 6580 7924 8206
rect 7980 6916 8036 8428
rect 8092 8428 8148 9324
rect 8204 8932 8260 9996
rect 8316 9938 8372 10220
rect 8316 9886 8318 9938
rect 8370 9886 8372 9938
rect 8316 9604 8372 9886
rect 8316 9538 8372 9548
rect 8316 8932 8372 8942
rect 8204 8930 8372 8932
rect 8204 8878 8318 8930
rect 8370 8878 8372 8930
rect 8204 8876 8372 8878
rect 8316 8866 8372 8876
rect 8428 8820 8484 10892
rect 8540 10612 8596 10650
rect 8540 10546 8596 10556
rect 8652 9940 8708 12460
rect 8652 9874 8708 9884
rect 8652 8932 8708 8942
rect 8652 8838 8708 8876
rect 8428 8754 8484 8764
rect 8092 8372 8260 8428
rect 8316 8372 8372 8382
rect 8204 8370 8372 8372
rect 8204 8318 8318 8370
rect 8370 8318 8372 8370
rect 8204 8316 8372 8318
rect 8316 8306 8372 8316
rect 8652 8260 8708 8270
rect 8428 7700 8484 7710
rect 8204 7476 8260 7486
rect 7980 6850 8036 6860
rect 8092 7474 8260 7476
rect 8092 7422 8206 7474
rect 8258 7422 8260 7474
rect 8092 7420 8260 7422
rect 7980 6692 8036 6702
rect 8092 6692 8148 7420
rect 8204 7410 8260 7420
rect 8316 7252 8372 7262
rect 7980 6690 8148 6692
rect 7980 6638 7982 6690
rect 8034 6638 8148 6690
rect 7980 6636 8148 6638
rect 7980 6626 8036 6636
rect 7868 6514 7924 6524
rect 7420 6412 7812 6468
rect 7196 5796 7252 5806
rect 6748 3726 6750 3778
rect 6802 3726 6804 3778
rect 6748 3714 6804 3726
rect 6860 4620 7028 4676
rect 7084 5236 7140 5246
rect 6860 3388 6916 4620
rect 6972 4228 7028 4238
rect 6972 4134 7028 4172
rect 7084 3892 7140 5180
rect 7196 5010 7252 5740
rect 7308 5794 7364 6412
rect 7756 6020 7812 6412
rect 7756 5964 7924 6020
rect 7308 5742 7310 5794
rect 7362 5742 7364 5794
rect 7308 5124 7364 5742
rect 7420 5796 7476 5806
rect 7756 5796 7812 5806
rect 7420 5702 7476 5740
rect 7532 5794 7812 5796
rect 7532 5742 7758 5794
rect 7810 5742 7812 5794
rect 7532 5740 7812 5742
rect 7308 5058 7364 5068
rect 7196 4958 7198 5010
rect 7250 4958 7252 5010
rect 7196 4946 7252 4958
rect 7308 4788 7364 4798
rect 7308 4338 7364 4732
rect 7532 4564 7588 5740
rect 7756 5730 7812 5740
rect 7644 5572 7700 5582
rect 7644 4900 7700 5516
rect 7756 5236 7812 5246
rect 7868 5236 7924 5964
rect 8092 5906 8148 6636
rect 8092 5854 8094 5906
rect 8146 5854 8148 5906
rect 8092 5460 8148 5854
rect 8092 5394 8148 5404
rect 8204 6916 8260 6926
rect 7980 5348 8036 5386
rect 7980 5282 8036 5292
rect 7756 5234 7924 5236
rect 7756 5182 7758 5234
rect 7810 5182 7924 5234
rect 7756 5180 7924 5182
rect 7756 5170 7812 5180
rect 7980 5124 8036 5134
rect 7980 5030 8036 5068
rect 8204 5122 8260 6860
rect 8316 6802 8372 7196
rect 8316 6750 8318 6802
rect 8370 6750 8372 6802
rect 8316 6738 8372 6750
rect 8204 5070 8206 5122
rect 8258 5070 8260 5122
rect 8204 5058 8260 5070
rect 7644 4844 8036 4900
rect 7308 4286 7310 4338
rect 7362 4286 7364 4338
rect 7308 4228 7364 4286
rect 7308 4162 7364 4172
rect 7420 4508 7588 4564
rect 7756 4676 7812 4686
rect 7084 3836 7364 3892
rect 7308 3778 7364 3836
rect 7308 3726 7310 3778
rect 7362 3726 7364 3778
rect 7308 3714 7364 3726
rect 7196 3556 7252 3566
rect 7252 3500 7364 3556
rect 7196 3490 7252 3500
rect 6860 3332 7252 3388
rect 6636 2772 6692 2782
rect 6636 2100 6692 2716
rect 7196 2770 7252 3332
rect 7196 2718 7198 2770
rect 7250 2718 7252 2770
rect 6860 2660 6916 2670
rect 6860 2566 6916 2604
rect 6636 2034 6692 2044
rect 6972 1988 7028 1998
rect 7196 1988 7252 2718
rect 7308 2660 7364 3500
rect 7308 2594 7364 2604
rect 6972 1986 7252 1988
rect 6972 1934 6974 1986
rect 7026 1934 7252 1986
rect 6972 1932 7252 1934
rect 7308 2212 7364 2222
rect 6972 1922 7028 1932
rect 7196 1652 7252 1662
rect 6972 1540 7028 1550
rect 6860 1204 6916 1214
rect 6860 1090 6916 1148
rect 6860 1038 6862 1090
rect 6914 1038 6916 1090
rect 6860 1026 6916 1038
rect 6972 112 7028 1484
rect 7196 1202 7252 1596
rect 7196 1150 7198 1202
rect 7250 1150 7252 1202
rect 7196 196 7252 1150
rect 7308 308 7364 2156
rect 7420 1652 7476 4508
rect 7532 4228 7588 4266
rect 7532 4162 7588 4172
rect 7420 1586 7476 1596
rect 7532 4004 7588 4014
rect 7532 756 7588 3948
rect 7644 3668 7700 3678
rect 7644 3574 7700 3612
rect 7756 3444 7812 4620
rect 7868 4114 7924 4126
rect 7868 4062 7870 4114
rect 7922 4062 7924 4114
rect 7868 3780 7924 4062
rect 7868 3714 7924 3724
rect 7980 3778 8036 4844
rect 8092 4338 8148 4350
rect 8092 4286 8094 4338
rect 8146 4286 8148 4338
rect 8092 4228 8148 4286
rect 8092 4162 8148 4172
rect 8316 4116 8372 4126
rect 7980 3726 7982 3778
rect 8034 3726 8036 3778
rect 7980 3714 8036 3726
rect 8092 4004 8148 4014
rect 7644 3388 7812 3444
rect 8092 3388 8148 3948
rect 8316 3778 8372 4060
rect 8316 3726 8318 3778
rect 8370 3726 8372 3778
rect 8316 3714 8372 3726
rect 7644 2882 7700 3388
rect 7644 2830 7646 2882
rect 7698 2830 7700 2882
rect 7644 2818 7700 2830
rect 7868 3332 8148 3388
rect 7532 690 7588 700
rect 7756 978 7812 990
rect 7756 926 7758 978
rect 7810 926 7812 978
rect 7756 308 7812 926
rect 7308 242 7364 252
rect 7420 252 7700 308
rect 7196 130 7252 140
rect 7420 112 7476 252
rect 672 0 784 112
rect 1120 0 1232 112
rect 1568 0 1680 112
rect 2016 0 2128 112
rect 2464 0 2576 112
rect 2912 0 3024 112
rect 3360 0 3472 112
rect 3808 0 3920 112
rect 4256 0 4368 112
rect 4704 0 4816 112
rect 5152 0 5264 112
rect 5600 0 5712 112
rect 6048 0 6160 112
rect 6496 0 6608 112
rect 6944 0 7056 112
rect 7392 0 7504 112
rect 7644 84 7700 252
rect 7756 242 7812 252
rect 7868 112 7924 3332
rect 7980 3220 8036 3230
rect 7980 2210 8036 3164
rect 8092 2772 8148 2782
rect 8092 2678 8148 2716
rect 8428 2658 8484 7644
rect 8652 7588 8708 8204
rect 8652 7494 8708 7532
rect 8764 6020 8820 17276
rect 9324 17444 9380 17454
rect 8988 16996 9044 17006
rect 8988 16902 9044 16940
rect 8876 16884 8932 16894
rect 8876 16210 8932 16828
rect 9324 16882 9380 17388
rect 9324 16830 9326 16882
rect 9378 16830 9380 16882
rect 9324 16818 9380 16830
rect 8988 16436 9044 16446
rect 8988 16322 9044 16380
rect 8988 16270 8990 16322
rect 9042 16270 9044 16322
rect 8988 16258 9044 16270
rect 9436 16324 9492 19182
rect 9660 18788 9716 18798
rect 9436 16258 9492 16268
rect 9548 18116 9604 18126
rect 9548 17778 9604 18060
rect 9660 18004 9716 18732
rect 9772 18228 9828 19294
rect 9772 18162 9828 18172
rect 9884 19348 9940 19358
rect 9884 18450 9940 19292
rect 9996 18788 10052 21980
rect 9996 18722 10052 18732
rect 10108 18676 10164 22428
rect 10332 22372 10388 23492
rect 10220 22316 10388 22372
rect 10220 19572 10276 22316
rect 10444 20244 10500 23772
rect 10556 26740 10612 26750
rect 10556 22036 10612 26684
rect 10556 21970 10612 21980
rect 10668 26516 10724 26526
rect 10668 23154 10724 26460
rect 10780 25956 10836 25966
rect 10780 25730 10836 25900
rect 10780 25678 10782 25730
rect 10834 25678 10836 25730
rect 10780 25666 10836 25678
rect 10668 23102 10670 23154
rect 10722 23102 10724 23154
rect 10556 21700 10612 21710
rect 10556 21606 10612 21644
rect 10668 21252 10724 23102
rect 10556 21196 10724 21252
rect 10780 23156 10836 23166
rect 10556 20468 10612 21196
rect 10668 20916 10724 20926
rect 10668 20822 10724 20860
rect 10556 20402 10612 20412
rect 10780 20468 10836 23100
rect 10892 22708 10948 27580
rect 10892 22642 10948 22652
rect 11004 22372 11060 33068
rect 11116 25620 11172 33516
rect 11340 33012 11396 36764
rect 11340 32946 11396 32956
rect 11452 34916 11508 37772
rect 11452 32788 11508 34860
rect 11340 32732 11508 32788
rect 11340 30994 11396 32732
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 30930 11396 30942
rect 11452 32564 11508 32574
rect 11228 29428 11284 29438
rect 11228 29314 11284 29372
rect 11228 29262 11230 29314
rect 11282 29262 11284 29314
rect 11228 28084 11284 29262
rect 11340 29202 11396 29214
rect 11340 29150 11342 29202
rect 11394 29150 11396 29202
rect 11340 28308 11396 29150
rect 11452 28980 11508 32508
rect 11452 28914 11508 28924
rect 11340 28242 11396 28252
rect 11452 28084 11508 28094
rect 11228 28082 11508 28084
rect 11228 28030 11454 28082
rect 11506 28030 11508 28082
rect 11228 28028 11508 28030
rect 11452 28018 11508 28028
rect 11452 27076 11508 27086
rect 11228 25620 11284 25630
rect 11116 25618 11284 25620
rect 11116 25566 11230 25618
rect 11282 25566 11284 25618
rect 11116 25564 11284 25566
rect 11004 22306 11060 22316
rect 11116 23940 11172 23950
rect 11116 21812 11172 23884
rect 11228 23044 11284 25564
rect 11340 25284 11396 25294
rect 11340 23938 11396 25228
rect 11340 23886 11342 23938
rect 11394 23886 11396 23938
rect 11340 23874 11396 23886
rect 11228 22978 11284 22988
rect 11340 22372 11396 22382
rect 11340 22278 11396 22316
rect 11116 21746 11172 21756
rect 10780 20402 10836 20412
rect 10892 21588 10948 21598
rect 10892 21474 10948 21532
rect 10892 21422 10894 21474
rect 10946 21422 10948 21474
rect 10444 20188 10612 20244
rect 10332 19796 10388 19806
rect 10332 19702 10388 19740
rect 10220 19516 10388 19572
rect 10220 19234 10276 19246
rect 10220 19182 10222 19234
rect 10274 19182 10276 19234
rect 10220 19124 10276 19182
rect 10220 19058 10276 19068
rect 10108 18620 10276 18676
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9660 17948 9828 18004
rect 9548 17726 9550 17778
rect 9602 17726 9604 17778
rect 8876 16158 8878 16210
rect 8930 16158 8932 16210
rect 8876 16146 8932 16158
rect 9212 15988 9268 15998
rect 9100 15652 9156 15662
rect 8876 15316 8932 15326
rect 8988 15316 9044 15326
rect 8876 15314 8988 15316
rect 8876 15262 8878 15314
rect 8930 15262 8988 15314
rect 8876 15260 8988 15262
rect 8876 15250 8932 15260
rect 8876 14756 8932 14766
rect 8876 14662 8932 14700
rect 8988 13748 9044 15260
rect 9100 14530 9156 15596
rect 9212 15204 9268 15932
rect 9324 15986 9380 15998
rect 9324 15934 9326 15986
rect 9378 15934 9380 15986
rect 9324 15540 9380 15934
rect 9324 15474 9380 15484
rect 9324 15204 9380 15214
rect 9212 15202 9380 15204
rect 9212 15150 9326 15202
rect 9378 15150 9380 15202
rect 9212 15148 9380 15150
rect 9324 15138 9380 15148
rect 9100 14478 9102 14530
rect 9154 14478 9156 14530
rect 9100 14466 9156 14478
rect 9436 15092 9492 15102
rect 8876 13746 9044 13748
rect 8876 13694 8990 13746
rect 9042 13694 9044 13746
rect 8876 13692 9044 13694
rect 8876 12292 8932 13692
rect 8988 13682 9044 13692
rect 9436 13300 9492 15036
rect 9548 14980 9604 17726
rect 9660 16996 9716 17006
rect 9660 16098 9716 16940
rect 9772 16882 9828 17948
rect 9772 16830 9774 16882
rect 9826 16830 9828 16882
rect 9772 16324 9828 16830
rect 9884 16548 9940 18398
rect 9996 18340 10052 18350
rect 9996 18246 10052 18284
rect 9996 16884 10052 16894
rect 9996 16770 10052 16828
rect 9996 16718 9998 16770
rect 10050 16718 10052 16770
rect 9996 16706 10052 16718
rect 9996 16548 10052 16558
rect 9884 16492 9996 16548
rect 9996 16482 10052 16492
rect 9772 16268 10052 16324
rect 9660 16046 9662 16098
rect 9714 16046 9716 16098
rect 9660 16034 9716 16046
rect 9996 15428 10052 16268
rect 10108 16100 10164 16110
rect 10108 16006 10164 16044
rect 9660 15204 9716 15242
rect 9660 15138 9716 15148
rect 9772 15092 9828 15102
rect 9548 14924 9716 14980
rect 9548 14420 9604 14430
rect 9548 13634 9604 14364
rect 9548 13582 9550 13634
rect 9602 13582 9604 13634
rect 9548 13570 9604 13582
rect 9436 13234 9492 13244
rect 8988 13076 9044 13086
rect 8988 12982 9044 13020
rect 9548 13074 9604 13086
rect 9548 13022 9550 13074
rect 9602 13022 9604 13074
rect 9100 12964 9156 12974
rect 9100 12870 9156 12908
rect 8988 12738 9044 12750
rect 9436 12740 9492 12750
rect 8988 12686 8990 12738
rect 9042 12686 9044 12738
rect 8988 12516 9044 12686
rect 8988 12450 9044 12460
rect 9100 12738 9492 12740
rect 9100 12686 9438 12738
rect 9490 12686 9492 12738
rect 9100 12684 9492 12686
rect 8988 12292 9044 12302
rect 8876 12290 9044 12292
rect 8876 12238 8990 12290
rect 9042 12238 9044 12290
rect 8876 12236 9044 12238
rect 8988 12226 9044 12236
rect 8876 11396 8932 11406
rect 9100 11396 9156 12684
rect 9436 12674 9492 12684
rect 9324 12178 9380 12190
rect 9324 12126 9326 12178
rect 9378 12126 9380 12178
rect 9324 11620 9380 12126
rect 9548 11844 9604 13022
rect 9548 11778 9604 11788
rect 9324 11554 9380 11564
rect 9660 11620 9716 14924
rect 9772 13746 9828 15036
rect 9884 14644 9940 14654
rect 9884 14550 9940 14588
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 13682 9828 13694
rect 9772 12738 9828 12750
rect 9772 12686 9774 12738
rect 9826 12686 9828 12738
rect 9772 11956 9828 12686
rect 9884 12180 9940 12190
rect 9996 12180 10052 15372
rect 9884 12178 10052 12180
rect 9884 12126 9886 12178
rect 9938 12126 10052 12178
rect 9884 12124 10052 12126
rect 10108 15540 10164 15550
rect 10108 12850 10164 15484
rect 10220 15428 10276 18620
rect 10332 17220 10388 19516
rect 10556 19222 10612 20188
rect 10780 19908 10836 19918
rect 10780 19814 10836 19852
rect 10780 19348 10836 19358
rect 10780 19254 10836 19292
rect 10556 19170 10558 19222
rect 10610 19170 10612 19222
rect 10556 19158 10612 19170
rect 10668 19124 10724 19134
rect 10332 17154 10388 17164
rect 10556 18452 10612 18462
rect 10556 16996 10612 18396
rect 10668 18450 10724 19068
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 17444 10724 18398
rect 10892 18116 10948 21422
rect 11452 21252 11508 27020
rect 11564 24052 11620 38108
rect 11900 37042 11956 37054
rect 11900 36990 11902 37042
rect 11954 36990 11956 37042
rect 11676 36484 11732 36494
rect 11900 36484 11956 36990
rect 12124 36484 12180 36494
rect 11676 36482 11956 36484
rect 11676 36430 11678 36482
rect 11730 36430 11956 36482
rect 11676 36428 11956 36430
rect 12012 36482 12180 36484
rect 12012 36430 12126 36482
rect 12178 36430 12180 36482
rect 12012 36428 12180 36430
rect 11676 34914 11732 36428
rect 12012 36372 12068 36428
rect 12124 36418 12180 36428
rect 11676 34862 11678 34914
rect 11730 34862 11732 34914
rect 11676 34850 11732 34862
rect 11788 36316 12068 36372
rect 11788 29652 11844 36316
rect 11900 35812 11956 35822
rect 11900 32564 11956 35756
rect 12124 35812 12180 35822
rect 12236 35812 12292 40350
rect 12348 37044 12404 41132
rect 12460 40740 12516 40750
rect 12460 39172 12516 40684
rect 12684 40516 12740 40526
rect 12460 39106 12516 39116
rect 12572 39284 12628 39294
rect 12348 36978 12404 36988
rect 12460 38948 12516 38958
rect 12348 36484 12404 36494
rect 12460 36484 12516 38892
rect 12572 37940 12628 39228
rect 12684 39060 12740 40460
rect 12796 40290 12852 41132
rect 12796 40238 12798 40290
rect 12850 40238 12852 40290
rect 12796 40226 12852 40238
rect 12908 39618 12964 39630
rect 12908 39566 12910 39618
rect 12962 39566 12964 39618
rect 12684 39004 12852 39060
rect 12684 38836 12740 38846
rect 12684 38742 12740 38780
rect 12796 38612 12852 39004
rect 12908 38836 12964 39566
rect 12908 38770 12964 38780
rect 13020 38834 13076 41804
rect 13132 41410 13188 44380
rect 13356 44324 13412 44334
rect 13244 43540 13300 43578
rect 13244 43474 13300 43484
rect 13132 41358 13134 41410
rect 13186 41358 13188 41410
rect 13132 41346 13188 41358
rect 13244 43316 13300 43326
rect 13020 38782 13022 38834
rect 13074 38782 13076 38834
rect 13020 38770 13076 38782
rect 13132 40178 13188 40190
rect 13132 40126 13134 40178
rect 13186 40126 13188 40178
rect 13132 38668 13188 40126
rect 13244 40068 13300 43260
rect 13356 41970 13412 44268
rect 13468 42084 13524 45614
rect 13468 42018 13524 42028
rect 13356 41918 13358 41970
rect 13410 41918 13412 41970
rect 13356 41906 13412 41918
rect 13468 41860 13524 41870
rect 13356 41186 13412 41198
rect 13356 41134 13358 41186
rect 13410 41134 13412 41186
rect 13356 40740 13412 41134
rect 13356 40674 13412 40684
rect 13468 40404 13524 41804
rect 13580 40516 13636 46284
rect 13804 46274 13860 46284
rect 13916 46844 14084 46900
rect 13804 44100 13860 44110
rect 13804 44006 13860 44044
rect 13580 40450 13636 40460
rect 13692 43426 13748 43438
rect 13692 43374 13694 43426
rect 13746 43374 13748 43426
rect 13692 41076 13748 43374
rect 13916 43428 13972 46844
rect 14028 45892 14084 45902
rect 14028 45798 14084 45836
rect 14028 45332 14084 45342
rect 14028 45218 14084 45276
rect 14028 45166 14030 45218
rect 14082 45166 14084 45218
rect 14028 45154 14084 45166
rect 14140 44996 14196 49308
rect 14476 48580 14532 50372
rect 14476 48514 14532 48524
rect 14588 50372 14980 50428
rect 13916 43362 13972 43372
rect 14028 44940 14196 44996
rect 14252 48020 14308 48030
rect 14252 44996 14308 47964
rect 13468 40338 13524 40348
rect 13580 40292 13636 40302
rect 13580 40198 13636 40236
rect 13244 40012 13524 40068
rect 13356 39844 13412 39854
rect 12908 38612 12964 38622
rect 12796 38610 12964 38612
rect 12796 38558 12910 38610
rect 12962 38558 12964 38610
rect 12796 38556 12964 38558
rect 12908 38546 12964 38556
rect 13020 38612 13188 38668
rect 13244 39172 13300 39182
rect 12796 37940 12852 37950
rect 12572 37938 12852 37940
rect 12572 37886 12798 37938
rect 12850 37886 12852 37938
rect 12572 37884 12852 37886
rect 12684 37044 12740 37054
rect 12348 36482 12516 36484
rect 12348 36430 12350 36482
rect 12402 36430 12516 36482
rect 12348 36428 12516 36430
rect 12572 36820 12628 36830
rect 12348 36418 12404 36428
rect 12180 35756 12292 35812
rect 12348 36148 12404 36158
rect 12124 35698 12180 35756
rect 12124 35646 12126 35698
rect 12178 35646 12180 35698
rect 12124 35634 12180 35646
rect 12348 35028 12404 36092
rect 12572 35308 12628 36764
rect 12348 34962 12404 34972
rect 12460 35252 12628 35308
rect 12012 34914 12068 34926
rect 12012 34862 12014 34914
rect 12066 34862 12068 34914
rect 12012 34580 12068 34862
rect 12012 33348 12068 34524
rect 12124 33906 12180 33918
rect 12124 33854 12126 33906
rect 12178 33854 12180 33906
rect 12124 33572 12180 33854
rect 12124 33506 12180 33516
rect 12012 33346 12180 33348
rect 12012 33294 12014 33346
rect 12066 33294 12180 33346
rect 12012 33292 12180 33294
rect 12012 33282 12068 33292
rect 11900 32498 11956 32508
rect 12012 32900 12068 32910
rect 11900 32004 11956 32014
rect 11900 31778 11956 31948
rect 11900 31726 11902 31778
rect 11954 31726 11956 31778
rect 11900 31714 11956 31726
rect 12012 31780 12068 32844
rect 12012 31714 12068 31724
rect 12124 31444 12180 33292
rect 12236 32452 12292 32462
rect 12236 31668 12292 32396
rect 12236 31602 12292 31612
rect 12348 31780 12404 31790
rect 12124 31378 12180 31388
rect 12236 30324 12292 30334
rect 12236 30210 12292 30268
rect 12236 30158 12238 30210
rect 12290 30158 12292 30210
rect 12236 30146 12292 30158
rect 11788 29586 11844 29596
rect 11676 29428 11732 29438
rect 11676 29334 11732 29372
rect 11900 29314 11956 29326
rect 11900 29262 11902 29314
rect 11954 29262 11956 29314
rect 11900 28868 11956 29262
rect 12236 29316 12292 29326
rect 12236 29222 12292 29260
rect 11788 28866 11956 28868
rect 11788 28814 11902 28866
rect 11954 28814 11956 28866
rect 11788 28812 11956 28814
rect 11676 27524 11732 27534
rect 11676 26852 11732 27468
rect 11788 27188 11844 28812
rect 11900 28802 11956 28812
rect 12124 29202 12180 29214
rect 12124 29150 12126 29202
rect 12178 29150 12180 29202
rect 12124 27972 12180 29150
rect 12348 29204 12404 31724
rect 12460 29652 12516 35252
rect 12572 32004 12628 32014
rect 12572 31556 12628 31948
rect 12572 31490 12628 31500
rect 12684 31444 12740 36988
rect 12796 35700 12852 37884
rect 12796 35634 12852 35644
rect 13020 35252 13076 38612
rect 13244 38274 13300 39116
rect 13244 38222 13246 38274
rect 13298 38222 13300 38274
rect 13244 38210 13300 38222
rect 13244 37156 13300 37166
rect 13020 35186 13076 35196
rect 13132 36482 13188 36494
rect 13132 36430 13134 36482
rect 13186 36430 13188 36482
rect 13020 34916 13076 34926
rect 13020 34822 13076 34860
rect 12908 33234 12964 33246
rect 12908 33182 12910 33234
rect 12962 33182 12964 33234
rect 12908 33124 12964 33182
rect 12908 33058 12964 33068
rect 13132 31780 13188 36430
rect 13244 35476 13300 37100
rect 13356 36708 13412 39788
rect 13468 39842 13524 40012
rect 13468 39790 13470 39842
rect 13522 39790 13524 39842
rect 13468 39508 13524 39790
rect 13468 39442 13524 39452
rect 13356 36642 13412 36652
rect 13580 38500 13636 38510
rect 13580 36596 13636 38444
rect 13692 38164 13748 41020
rect 13804 42530 13860 42542
rect 13804 42478 13806 42530
rect 13858 42478 13860 42530
rect 13804 40404 13860 42478
rect 13916 41748 13972 41758
rect 13916 40740 13972 41692
rect 13916 40674 13972 40684
rect 13916 40404 13972 40414
rect 13804 40402 13972 40404
rect 13804 40350 13918 40402
rect 13970 40350 13972 40402
rect 13804 40348 13972 40350
rect 13916 40338 13972 40348
rect 13916 40180 13972 40190
rect 13692 38098 13748 38108
rect 13804 38388 13860 38398
rect 13804 37268 13860 38332
rect 13804 37202 13860 37212
rect 13580 36530 13636 36540
rect 13244 35410 13300 35420
rect 13468 36372 13524 36382
rect 13468 34692 13524 36316
rect 13916 35924 13972 40124
rect 13468 34626 13524 34636
rect 13580 35868 13972 35924
rect 13244 33572 13300 33582
rect 13244 33346 13300 33516
rect 13244 33294 13246 33346
rect 13298 33294 13300 33346
rect 13244 33282 13300 33294
rect 13132 31714 13188 31724
rect 13244 33124 13300 33134
rect 12684 31378 12740 31388
rect 13020 31332 13076 31342
rect 12684 30324 12740 30334
rect 12684 30230 12740 30268
rect 12460 29586 12516 29596
rect 12908 29652 12964 29662
rect 12908 29558 12964 29596
rect 13020 29428 13076 31276
rect 13132 30884 13188 30894
rect 13132 30790 13188 30828
rect 12348 29138 12404 29148
rect 12908 29372 13076 29428
rect 12348 28644 12404 28654
rect 12348 28196 12404 28588
rect 12572 28644 12628 28654
rect 12572 28550 12628 28588
rect 12348 28130 12404 28140
rect 12796 28308 12852 28318
rect 12124 27916 12740 27972
rect 12124 27748 12180 27758
rect 11900 27634 11956 27646
rect 11900 27582 11902 27634
rect 11954 27582 11956 27634
rect 11900 27412 11956 27582
rect 11900 27346 11956 27356
rect 12012 27300 12068 27310
rect 12124 27300 12180 27692
rect 12012 27298 12180 27300
rect 12012 27246 12014 27298
rect 12066 27246 12180 27298
rect 12012 27244 12180 27246
rect 12236 27746 12292 27758
rect 12236 27694 12238 27746
rect 12290 27694 12292 27746
rect 12236 27300 12292 27694
rect 12684 27636 12740 27916
rect 12796 27858 12852 28252
rect 12796 27806 12798 27858
rect 12850 27806 12852 27858
rect 12796 27794 12852 27806
rect 12684 27580 12852 27636
rect 12012 27234 12068 27244
rect 12236 27234 12292 27244
rect 11900 27188 11956 27198
rect 11788 27132 11900 27188
rect 11900 27094 11956 27132
rect 12460 27188 12516 27198
rect 12460 27094 12516 27132
rect 12348 27074 12404 27086
rect 12348 27022 12350 27074
rect 12402 27022 12404 27074
rect 11676 26786 11732 26796
rect 12124 26852 12180 26862
rect 11676 25956 11732 25966
rect 11676 25506 11732 25900
rect 11900 25844 11956 25854
rect 11676 25454 11678 25506
rect 11730 25454 11732 25506
rect 11676 25442 11732 25454
rect 11788 25508 11844 25518
rect 11788 24836 11844 25452
rect 11788 24770 11844 24780
rect 11676 24052 11732 24062
rect 11564 23996 11676 24052
rect 11676 23958 11732 23996
rect 11452 21186 11508 21196
rect 11788 22596 11844 22606
rect 11788 22482 11844 22540
rect 11788 22430 11790 22482
rect 11842 22430 11844 22482
rect 11340 20916 11396 20926
rect 11116 20804 11172 20814
rect 11116 20710 11172 20748
rect 11228 20692 11284 20702
rect 11228 20598 11284 20636
rect 11116 19908 11172 19918
rect 11116 19814 11172 19852
rect 11340 19906 11396 20860
rect 11564 20914 11620 20926
rect 11564 20862 11566 20914
rect 11618 20862 11620 20914
rect 11340 19854 11342 19906
rect 11394 19854 11396 19906
rect 11340 19842 11396 19854
rect 11452 20468 11508 20478
rect 11004 19796 11060 19806
rect 11004 19460 11060 19740
rect 11004 19236 11060 19404
rect 11004 19180 11172 19236
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 18340 11060 18398
rect 11004 18274 11060 18284
rect 10892 18050 10948 18060
rect 11116 17892 11172 19180
rect 11228 19234 11284 19246
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 11228 18452 11284 19182
rect 11228 18386 11284 18396
rect 11340 18564 11396 18574
rect 11228 17892 11284 17902
rect 11116 17890 11284 17892
rect 11116 17838 11230 17890
rect 11282 17838 11284 17890
rect 11116 17836 11284 17838
rect 11228 17826 11284 17836
rect 11116 17668 11172 17678
rect 11004 17666 11172 17668
rect 11004 17614 11118 17666
rect 11170 17614 11172 17666
rect 11004 17612 11172 17614
rect 10724 17388 10836 17444
rect 10668 17350 10724 17388
rect 10556 16882 10612 16940
rect 10556 16830 10558 16882
rect 10610 16830 10612 16882
rect 10556 16818 10612 16830
rect 10668 16548 10724 16558
rect 10332 16324 10388 16334
rect 10332 16230 10388 16268
rect 10556 16324 10612 16334
rect 10556 15876 10612 16268
rect 10556 15810 10612 15820
rect 10220 15362 10276 15372
rect 10556 15428 10612 15438
rect 10332 14530 10388 14542
rect 10332 14478 10334 14530
rect 10386 14478 10388 14530
rect 10108 12798 10110 12850
rect 10162 12798 10164 12850
rect 9884 12114 9940 12124
rect 9996 11956 10052 11966
rect 9772 11954 10052 11956
rect 9772 11902 9998 11954
rect 10050 11902 10052 11954
rect 9772 11900 10052 11902
rect 9996 11890 10052 11900
rect 9660 11554 9716 11564
rect 8876 11394 9156 11396
rect 8876 11342 8878 11394
rect 8930 11342 9156 11394
rect 8876 11340 9156 11342
rect 9212 11508 9268 11518
rect 8876 11330 8932 11340
rect 9100 11172 9156 11182
rect 9100 11078 9156 11116
rect 9100 10948 9156 10958
rect 8876 10724 8932 10734
rect 8876 10050 8932 10668
rect 8876 9998 8878 10050
rect 8930 9998 8932 10050
rect 8876 9986 8932 9998
rect 9100 9268 9156 10892
rect 9212 10610 9268 11452
rect 9548 11394 9604 11406
rect 9548 11342 9550 11394
rect 9602 11342 9604 11394
rect 9212 10558 9214 10610
rect 9266 10558 9268 10610
rect 9212 10052 9268 10558
rect 9212 9986 9268 9996
rect 9324 11282 9380 11294
rect 9324 11230 9326 11282
rect 9378 11230 9380 11282
rect 9324 9940 9380 11230
rect 9548 10164 9604 11342
rect 9772 11394 9828 11406
rect 9772 11342 9774 11394
rect 9826 11342 9828 11394
rect 9660 11282 9716 11294
rect 9660 11230 9662 11282
rect 9714 11230 9716 11282
rect 9660 10276 9716 11230
rect 9772 10724 9828 11342
rect 9772 10658 9828 10668
rect 10108 10500 10164 12798
rect 10220 13188 10276 13198
rect 10220 11506 10276 13132
rect 10220 11454 10222 11506
rect 10274 11454 10276 11506
rect 10220 11442 10276 11454
rect 10332 11508 10388 14478
rect 10556 13858 10612 15372
rect 10556 13806 10558 13858
rect 10610 13806 10612 13858
rect 10556 13794 10612 13806
rect 10668 14530 10724 16492
rect 10780 16210 10836 17388
rect 11004 16436 11060 17612
rect 11116 17602 11172 17612
rect 11228 17332 11284 17342
rect 11228 16882 11284 17276
rect 11228 16830 11230 16882
rect 11282 16830 11284 16882
rect 11228 16818 11284 16830
rect 11004 16370 11060 16380
rect 10780 16158 10782 16210
rect 10834 16158 10836 16210
rect 10780 16146 10836 16158
rect 11116 16212 11172 16222
rect 10892 15204 10948 15242
rect 10892 15138 10948 15148
rect 10892 14644 10948 14654
rect 10668 14478 10670 14530
rect 10722 14478 10724 14530
rect 10332 11442 10388 11452
rect 10444 13748 10500 13758
rect 10332 10612 10388 10622
rect 10444 10612 10500 13692
rect 10556 13188 10612 13198
rect 10556 12962 10612 13132
rect 10556 12910 10558 12962
rect 10610 12910 10612 12962
rect 10556 12178 10612 12910
rect 10556 12126 10558 12178
rect 10610 12126 10612 12178
rect 10556 11394 10612 12126
rect 10556 11342 10558 11394
rect 10610 11342 10612 11394
rect 10556 10836 10612 11342
rect 10556 10770 10612 10780
rect 10444 10556 10612 10612
rect 10332 10500 10388 10556
rect 10108 10444 10276 10500
rect 10332 10444 10500 10500
rect 9772 10388 9828 10398
rect 9996 10388 10052 10398
rect 9772 10294 9828 10332
rect 9884 10332 9996 10388
rect 9660 10210 9716 10220
rect 9548 10098 9604 10108
rect 9324 9874 9380 9884
rect 9884 9940 9940 10332
rect 9996 10322 10052 10332
rect 9884 9846 9940 9884
rect 9212 9826 9268 9838
rect 9212 9774 9214 9826
rect 9266 9774 9268 9826
rect 9212 9716 9268 9774
rect 9436 9716 9492 9726
rect 9212 9714 9492 9716
rect 9212 9662 9438 9714
rect 9490 9662 9492 9714
rect 9212 9660 9492 9662
rect 9100 9202 9156 9212
rect 9324 8708 9380 9660
rect 9436 9650 9492 9660
rect 9660 9380 9716 9390
rect 9548 9268 9604 9278
rect 9436 9156 9492 9166
rect 9548 9156 9604 9212
rect 9436 9154 9604 9156
rect 9436 9102 9438 9154
rect 9490 9102 9604 9154
rect 9436 9100 9604 9102
rect 9436 9090 9492 9100
rect 9324 8642 9380 8652
rect 9548 8260 9604 8270
rect 9548 8166 9604 8204
rect 8988 8146 9044 8158
rect 8988 8094 8990 8146
rect 9042 8094 9044 8146
rect 8876 8034 8932 8046
rect 8876 7982 8878 8034
rect 8930 7982 8932 8034
rect 8876 6916 8932 7982
rect 8988 7252 9044 8094
rect 9100 7924 9156 7934
rect 9100 7474 9156 7868
rect 9100 7422 9102 7474
rect 9154 7422 9156 7474
rect 9100 7410 9156 7422
rect 8988 7186 9044 7196
rect 9324 7252 9380 7262
rect 8876 6850 8932 6860
rect 9324 6914 9380 7196
rect 9324 6862 9326 6914
rect 9378 6862 9380 6914
rect 9324 6850 9380 6862
rect 9100 6804 9156 6814
rect 9100 6710 9156 6748
rect 8876 6692 8932 6702
rect 8876 6598 8932 6636
rect 9212 6692 9268 6702
rect 9212 6598 9268 6636
rect 9436 6690 9492 6702
rect 9436 6638 9438 6690
rect 9490 6638 9492 6690
rect 8652 5964 8820 6020
rect 9100 6580 9156 6590
rect 8540 5908 8596 5918
rect 8540 5814 8596 5852
rect 8428 2606 8430 2658
rect 8482 2606 8484 2658
rect 8428 2594 8484 2606
rect 8540 5124 8596 5134
rect 8540 2324 8596 5068
rect 8652 2772 8708 5964
rect 9100 5908 9156 6524
rect 9212 5908 9268 5918
rect 9100 5906 9268 5908
rect 9100 5854 9214 5906
rect 9266 5854 9268 5906
rect 9100 5852 9268 5854
rect 9212 5842 9268 5852
rect 8764 5796 8820 5806
rect 8764 5702 8820 5740
rect 9212 5460 9268 5470
rect 9212 5346 9268 5404
rect 9212 5294 9214 5346
rect 9266 5294 9268 5346
rect 9212 5282 9268 5294
rect 9436 5348 9492 6638
rect 9660 5796 9716 9324
rect 9884 9268 9940 9278
rect 9884 8930 9940 9212
rect 9884 8878 9886 8930
rect 9938 8878 9940 8930
rect 9884 8148 9940 8878
rect 9884 8082 9940 8092
rect 10108 9268 10164 9278
rect 10108 7812 10164 9212
rect 9660 5730 9716 5740
rect 9772 7756 10164 7812
rect 9436 5282 9492 5292
rect 8876 5234 8932 5246
rect 8876 5182 8878 5234
rect 8930 5182 8932 5234
rect 8876 4900 8932 5182
rect 9548 5234 9604 5246
rect 9548 5182 9550 5234
rect 9602 5182 9604 5234
rect 8988 5012 9044 5022
rect 9044 4956 9156 5012
rect 8988 4946 9044 4956
rect 8876 4834 8932 4844
rect 8876 4564 8932 4574
rect 8876 4450 8932 4508
rect 8876 4398 8878 4450
rect 8930 4398 8932 4450
rect 8876 4386 8932 4398
rect 9100 3778 9156 4956
rect 9548 4340 9604 5182
rect 9772 5124 9828 7756
rect 10108 7588 10164 7598
rect 9996 7476 10052 7486
rect 9996 7382 10052 7420
rect 10108 6802 10164 7532
rect 10108 6750 10110 6802
rect 10162 6750 10164 6802
rect 10108 6738 10164 6750
rect 9996 6690 10052 6702
rect 9996 6638 9998 6690
rect 10050 6638 10052 6690
rect 9884 6356 9940 6366
rect 9884 5906 9940 6300
rect 9884 5854 9886 5906
rect 9938 5854 9940 5906
rect 9884 5842 9940 5854
rect 9996 5236 10052 6638
rect 10108 5236 10164 5246
rect 9996 5180 10108 5236
rect 10108 5170 10164 5180
rect 9772 5058 9828 5068
rect 9884 5122 9940 5134
rect 9884 5070 9886 5122
rect 9938 5070 9940 5122
rect 9548 4274 9604 4284
rect 9100 3726 9102 3778
rect 9154 3726 9156 3778
rect 9100 3714 9156 3726
rect 9212 4226 9268 4238
rect 9212 4174 9214 4226
rect 9266 4174 9268 4226
rect 9212 3444 9268 4174
rect 9772 3780 9828 3790
rect 9772 3686 9828 3724
rect 9436 3668 9492 3678
rect 9436 3666 9716 3668
rect 9436 3614 9438 3666
rect 9490 3614 9716 3666
rect 9436 3612 9716 3614
rect 9436 3602 9492 3612
rect 9212 3378 9268 3388
rect 9324 3220 9380 3230
rect 8652 2706 8708 2716
rect 8876 2772 8932 2782
rect 8932 2716 9156 2772
rect 8876 2678 8932 2716
rect 8540 2258 8596 2268
rect 7980 2158 7982 2210
rect 8034 2158 8036 2210
rect 7980 2146 8036 2158
rect 8540 2100 8596 2110
rect 8204 1988 8260 1998
rect 8204 1894 8260 1932
rect 7980 1652 8036 1662
rect 7980 308 8036 1596
rect 8316 1652 8372 1662
rect 8092 980 8148 990
rect 8092 886 8148 924
rect 7980 242 8036 252
rect 8316 112 8372 1596
rect 8540 1204 8596 2044
rect 9100 1986 9156 2716
rect 9100 1934 9102 1986
rect 9154 1934 9156 1986
rect 9100 1922 9156 1934
rect 9324 2658 9380 3164
rect 9324 2606 9326 2658
rect 9378 2606 9380 2658
rect 9324 1988 9380 2606
rect 9660 2660 9716 3612
rect 9884 3388 9940 5070
rect 10108 3666 10164 3678
rect 10108 3614 10110 3666
rect 10162 3614 10164 3666
rect 10108 3556 10164 3614
rect 10108 3490 10164 3500
rect 10220 3388 10276 10444
rect 10332 8260 10388 8270
rect 10332 8166 10388 8204
rect 10332 6580 10388 6590
rect 10332 6486 10388 6524
rect 9884 3332 10052 3388
rect 9660 2594 9716 2604
rect 9660 2212 9716 2222
rect 9660 2118 9716 2156
rect 9324 1922 9380 1932
rect 9660 1988 9716 1998
rect 9212 1652 9268 1662
rect 8764 1540 8820 1550
rect 8764 1426 8820 1484
rect 8764 1374 8766 1426
rect 8818 1374 8820 1426
rect 8764 1362 8820 1374
rect 8540 1138 8596 1148
rect 8764 1204 8820 1214
rect 8764 112 8820 1148
rect 9212 112 9268 1596
rect 9660 112 9716 1932
rect 9884 1316 9940 1326
rect 9884 1090 9940 1260
rect 9884 1038 9886 1090
rect 9938 1038 9940 1090
rect 9884 1026 9940 1038
rect 9996 980 10052 3332
rect 9996 914 10052 924
rect 10108 3332 10276 3388
rect 10332 5796 10388 5806
rect 10332 3388 10388 5740
rect 10444 5122 10500 10444
rect 10556 7924 10612 10556
rect 10668 8148 10724 14478
rect 10780 14642 10948 14644
rect 10780 14590 10894 14642
rect 10946 14590 10948 14642
rect 10780 14588 10948 14590
rect 10780 9940 10836 14588
rect 10892 14578 10948 14588
rect 11004 13748 11060 13758
rect 11004 13634 11060 13692
rect 11004 13582 11006 13634
rect 11058 13582 11060 13634
rect 11004 13570 11060 13582
rect 11116 13524 11172 16156
rect 11340 16098 11396 18508
rect 11452 18116 11508 20412
rect 11564 20130 11620 20862
rect 11788 20692 11844 22430
rect 11900 21476 11956 25788
rect 12012 25508 12068 25518
rect 12012 25414 12068 25452
rect 12124 22596 12180 26796
rect 12236 25732 12292 25742
rect 12348 25732 12404 27022
rect 12684 27074 12740 27086
rect 12684 27022 12686 27074
rect 12738 27022 12740 27074
rect 12684 26292 12740 27022
rect 12684 26226 12740 26236
rect 12796 26290 12852 27580
rect 12908 27186 12964 29372
rect 13020 28644 13076 28654
rect 13020 28642 13188 28644
rect 13020 28590 13022 28642
rect 13074 28590 13188 28642
rect 13020 28588 13188 28590
rect 13020 28578 13076 28588
rect 13020 28308 13076 28318
rect 13020 28084 13076 28252
rect 13020 28018 13076 28028
rect 13132 27860 13188 28588
rect 13244 28532 13300 33068
rect 13468 32562 13524 32574
rect 13468 32510 13470 32562
rect 13522 32510 13524 32562
rect 13468 32452 13524 32510
rect 13468 32386 13524 32396
rect 13468 30994 13524 31006
rect 13468 30942 13470 30994
rect 13522 30942 13524 30994
rect 13244 28466 13300 28476
rect 13356 30884 13412 30894
rect 13356 28642 13412 30828
rect 13468 29652 13524 30942
rect 13580 29988 13636 35868
rect 13916 35700 13972 35710
rect 13916 35308 13972 35644
rect 13804 35252 13972 35308
rect 13692 34692 13748 34702
rect 13692 34598 13748 34636
rect 13804 33684 13860 35252
rect 13916 34692 13972 34702
rect 13916 34020 13972 34636
rect 14028 34242 14084 44940
rect 14252 44930 14308 44940
rect 14364 47348 14420 47358
rect 14364 44772 14420 47292
rect 14588 47124 14644 50372
rect 14812 49924 14868 49934
rect 14700 49812 14756 49822
rect 14700 49718 14756 49756
rect 14812 49588 14868 49868
rect 15036 49924 15092 51100
rect 15148 50428 15204 51100
rect 15260 50596 15316 50634
rect 15260 50530 15316 50540
rect 15596 50594 15652 50606
rect 15596 50542 15598 50594
rect 15650 50542 15652 50594
rect 15596 50428 15652 50542
rect 15708 50596 15764 51324
rect 15820 51314 15876 51324
rect 16044 51380 16100 51998
rect 16156 51492 16212 52892
rect 16492 52946 16548 53116
rect 16492 52894 16494 52946
rect 16546 52894 16548 52946
rect 16492 52882 16548 52894
rect 16716 52724 16772 52734
rect 16268 52722 16772 52724
rect 16268 52670 16718 52722
rect 16770 52670 16772 52722
rect 16268 52668 16772 52670
rect 16268 52162 16324 52668
rect 16716 52658 16772 52668
rect 16268 52110 16270 52162
rect 16322 52110 16324 52162
rect 16268 52098 16324 52110
rect 16828 52276 16884 52286
rect 16828 52162 16884 52220
rect 16828 52110 16830 52162
rect 16882 52110 16884 52162
rect 16828 52098 16884 52110
rect 16156 51426 16212 51436
rect 16940 52052 16996 52062
rect 16044 51314 16100 51324
rect 16492 51266 16548 51278
rect 16492 51214 16494 51266
rect 16546 51214 16548 51266
rect 16380 51154 16436 51166
rect 16380 51102 16382 51154
rect 16434 51102 16436 51154
rect 16268 50708 16324 50718
rect 15708 50530 15764 50540
rect 15820 50594 15876 50606
rect 15820 50542 15822 50594
rect 15874 50542 15876 50594
rect 15148 50372 15316 50428
rect 15036 49858 15092 49868
rect 14700 49532 14868 49588
rect 15148 49700 15204 49710
rect 14700 47460 14756 49532
rect 15148 49476 15204 49644
rect 15148 49410 15204 49420
rect 14924 48916 14980 48926
rect 14924 48822 14980 48860
rect 15260 48356 15316 50372
rect 15260 48262 15316 48300
rect 15372 50372 15652 50428
rect 15820 50372 15876 50542
rect 16156 50594 16212 50606
rect 16156 50542 16158 50594
rect 16210 50542 16212 50594
rect 14812 48018 14868 48030
rect 14812 47966 14814 48018
rect 14866 47966 14868 48018
rect 14812 47908 14868 47966
rect 14812 47842 14868 47852
rect 15148 47572 15204 47582
rect 14700 47366 14756 47404
rect 14924 47570 15204 47572
rect 14924 47518 15150 47570
rect 15202 47518 15204 47570
rect 14924 47516 15204 47518
rect 14588 47058 14644 47068
rect 14588 46788 14644 46798
rect 14588 46002 14644 46732
rect 14588 45950 14590 46002
rect 14642 45950 14644 46002
rect 14476 45220 14532 45230
rect 14476 45106 14532 45164
rect 14476 45054 14478 45106
rect 14530 45054 14532 45106
rect 14476 45042 14532 45054
rect 14252 44716 14420 44772
rect 14252 41970 14308 44716
rect 14252 41918 14254 41970
rect 14306 41918 14308 41970
rect 14140 40740 14196 40750
rect 14140 39732 14196 40684
rect 14252 40292 14308 41918
rect 14252 40226 14308 40236
rect 14364 44322 14420 44334
rect 14364 44270 14366 44322
rect 14418 44270 14420 44322
rect 14364 42754 14420 44270
rect 14364 42702 14366 42754
rect 14418 42702 14420 42754
rect 14364 41186 14420 42702
rect 14588 42644 14644 45950
rect 14700 46450 14756 46462
rect 14700 46398 14702 46450
rect 14754 46398 14756 46450
rect 14700 45220 14756 46398
rect 14700 45154 14756 45164
rect 14812 45109 14868 45146
rect 14812 45108 14814 45109
rect 14866 45108 14868 45109
rect 14812 45042 14868 45052
rect 14924 44660 14980 47516
rect 15148 47506 15204 47516
rect 15260 47458 15316 47470
rect 15260 47406 15262 47458
rect 15314 47406 15316 47458
rect 15260 47348 15316 47406
rect 15260 47282 15316 47292
rect 15036 46788 15092 46798
rect 15148 46788 15204 46798
rect 15092 46786 15204 46788
rect 15092 46734 15150 46786
rect 15202 46734 15204 46786
rect 15092 46732 15204 46734
rect 15036 46722 15092 46732
rect 15148 46722 15204 46732
rect 15260 46676 15316 46686
rect 15036 44884 15092 44894
rect 15036 44790 15092 44828
rect 14924 44604 15092 44660
rect 14588 42578 14644 42588
rect 14812 44434 14868 44446
rect 14812 44382 14814 44434
rect 14866 44382 14868 44434
rect 14812 42196 14868 44382
rect 15036 43708 15092 44604
rect 15148 44324 15204 44334
rect 15148 43876 15204 44268
rect 15148 43810 15204 43820
rect 15036 43652 15204 43708
rect 15148 43540 15204 43652
rect 15148 43474 15204 43484
rect 14924 43316 14980 43326
rect 14924 43314 15204 43316
rect 14924 43262 14926 43314
rect 14978 43262 15204 43314
rect 14924 43260 15204 43262
rect 14924 43250 14980 43260
rect 14924 42866 14980 42878
rect 14924 42814 14926 42866
rect 14978 42814 14980 42866
rect 14924 42644 14980 42814
rect 14924 42578 14980 42588
rect 14700 42140 14868 42196
rect 14924 42420 14980 42430
rect 14700 41860 14756 42140
rect 14924 42084 14980 42364
rect 14924 42018 14980 42028
rect 14812 41972 14868 41982
rect 14812 41878 14868 41916
rect 14700 41794 14756 41804
rect 14812 41300 14868 41310
rect 14812 41206 14868 41244
rect 14364 41134 14366 41186
rect 14418 41134 14420 41186
rect 14364 40180 14420 41134
rect 14588 40516 14644 40526
rect 14476 40404 14532 40414
rect 14476 40310 14532 40348
rect 14588 40292 14644 40460
rect 15148 40402 15204 43260
rect 15260 41300 15316 46620
rect 15372 43876 15428 50372
rect 15820 50306 15876 50316
rect 16044 50482 16100 50494
rect 16044 50430 16046 50482
rect 16098 50430 16100 50482
rect 15708 50036 15764 50046
rect 15484 49812 15540 49822
rect 15708 49812 15764 49980
rect 15540 49756 15652 49812
rect 15484 49718 15540 49756
rect 15484 49026 15540 49038
rect 15484 48974 15486 49026
rect 15538 48974 15540 49026
rect 15484 46900 15540 48974
rect 15596 48242 15652 49756
rect 15708 49746 15764 49756
rect 15932 49812 15988 49822
rect 15932 49718 15988 49756
rect 16044 49250 16100 50430
rect 16156 49698 16212 50542
rect 16156 49646 16158 49698
rect 16210 49646 16212 49698
rect 16156 49634 16212 49646
rect 16044 49198 16046 49250
rect 16098 49198 16100 49250
rect 16044 49186 16100 49198
rect 15596 48190 15598 48242
rect 15650 48190 15652 48242
rect 15596 47460 15652 48190
rect 15708 49026 15764 49038
rect 15708 48974 15710 49026
rect 15762 48974 15764 49026
rect 15708 47908 15764 48974
rect 15932 49026 15988 49038
rect 15932 48974 15934 49026
rect 15986 48974 15988 49026
rect 15932 48804 15988 48974
rect 16044 49028 16100 49038
rect 16044 48914 16100 48972
rect 16044 48862 16046 48914
rect 16098 48862 16100 48914
rect 16044 48850 16100 48862
rect 15932 48738 15988 48748
rect 16044 48468 16100 48478
rect 15708 47842 15764 47852
rect 15820 48356 15876 48366
rect 15708 47460 15764 47470
rect 15596 47458 15764 47460
rect 15596 47406 15710 47458
rect 15762 47406 15764 47458
rect 15596 47404 15764 47406
rect 15484 46844 15652 46900
rect 15484 46676 15540 46686
rect 15484 46582 15540 46620
rect 15372 43810 15428 43820
rect 15484 45780 15540 45790
rect 15372 43540 15428 43550
rect 15372 43446 15428 43484
rect 15484 42868 15540 45724
rect 15596 43650 15652 46844
rect 15708 46676 15764 47404
rect 15708 46610 15764 46620
rect 15820 46900 15876 48300
rect 16044 48242 16100 48412
rect 16268 48244 16324 50652
rect 16380 48356 16436 51102
rect 16492 50372 16548 51214
rect 16828 51266 16884 51278
rect 16828 51214 16830 51266
rect 16882 51214 16884 51266
rect 16828 51156 16884 51214
rect 16940 51268 16996 51996
rect 16940 51202 16996 51212
rect 17052 51156 17108 53452
rect 17276 52164 17332 54238
rect 18396 54180 18452 54190
rect 17388 53842 17444 53854
rect 17388 53790 17390 53842
rect 17442 53790 17444 53842
rect 17388 53396 17444 53790
rect 18396 53844 18452 54124
rect 18732 54180 18788 56252
rect 18844 55970 18900 56700
rect 18844 55918 18846 55970
rect 18898 55918 18900 55970
rect 18844 55906 18900 55918
rect 19068 55972 19124 57344
rect 19292 56196 19348 56206
rect 19292 56082 19348 56140
rect 19516 56084 19572 57344
rect 19292 56030 19294 56082
rect 19346 56030 19348 56082
rect 19292 56018 19348 56030
rect 19404 56028 19572 56084
rect 19068 55906 19124 55916
rect 19180 55636 19236 55646
rect 19180 55410 19236 55580
rect 19180 55358 19182 55410
rect 19234 55358 19236 55410
rect 19180 55346 19236 55358
rect 18956 55298 19012 55310
rect 18956 55246 18958 55298
rect 19010 55246 19012 55298
rect 18732 54114 18788 54124
rect 18844 54514 18900 54526
rect 18844 54462 18846 54514
rect 18898 54462 18900 54514
rect 18396 53778 18452 53788
rect 18620 53844 18676 53854
rect 17388 53330 17444 53340
rect 18508 53506 18564 53518
rect 18508 53454 18510 53506
rect 18562 53454 18564 53506
rect 18508 53172 18564 53454
rect 17612 53116 18564 53172
rect 17388 52948 17444 52958
rect 17612 52948 17668 53116
rect 17388 52946 17668 52948
rect 17388 52894 17390 52946
rect 17442 52894 17668 52946
rect 17388 52892 17668 52894
rect 17724 52948 17780 52958
rect 17388 52882 17444 52892
rect 17724 52854 17780 52892
rect 17948 52948 18004 52958
rect 17948 52724 18004 52892
rect 17948 52658 18004 52668
rect 17276 52098 17332 52108
rect 17948 52162 18004 52174
rect 17948 52110 17950 52162
rect 18002 52110 18004 52162
rect 17164 51492 17220 51502
rect 17164 51380 17220 51436
rect 17164 51378 17444 51380
rect 17164 51326 17166 51378
rect 17218 51326 17444 51378
rect 17164 51324 17444 51326
rect 17164 51314 17220 51324
rect 17052 51100 17332 51156
rect 16828 51090 16884 51100
rect 17164 50820 17220 50830
rect 16492 50306 16548 50316
rect 16940 50484 16996 50494
rect 17052 50484 17108 50494
rect 16996 50482 17108 50484
rect 16996 50430 17054 50482
rect 17106 50430 17108 50482
rect 16996 50428 17108 50430
rect 16940 50036 16996 50428
rect 17052 50418 17108 50428
rect 16940 49970 16996 49980
rect 17052 50260 17108 50270
rect 16828 49924 16884 49934
rect 16716 49868 16828 49924
rect 16716 49810 16772 49868
rect 16716 49758 16718 49810
rect 16770 49758 16772 49810
rect 16716 49746 16772 49758
rect 16380 48290 16436 48300
rect 16492 49700 16548 49710
rect 16044 48190 16046 48242
rect 16098 48190 16100 48242
rect 16044 48178 16100 48190
rect 16156 48188 16324 48244
rect 16156 48020 16212 48188
rect 16044 47964 16212 48020
rect 16268 48018 16324 48030
rect 16268 47966 16270 48018
rect 16322 47966 16324 48018
rect 15932 47908 15988 47918
rect 15932 47124 15988 47852
rect 15932 47058 15988 47068
rect 16044 47068 16100 47964
rect 16268 47908 16324 47966
rect 16492 47908 16548 49644
rect 16828 49588 16884 49868
rect 16716 49532 16884 49588
rect 16716 48244 16772 49532
rect 17052 48916 17108 50204
rect 17164 49252 17220 50764
rect 17276 49252 17332 51100
rect 17388 50594 17444 51324
rect 17612 51378 17668 51390
rect 17612 51326 17614 51378
rect 17666 51326 17668 51378
rect 17612 51268 17668 51326
rect 17612 51202 17668 51212
rect 17836 51268 17892 51278
rect 17836 51174 17892 51212
rect 17388 50542 17390 50594
rect 17442 50542 17444 50594
rect 17388 50530 17444 50542
rect 17500 50932 17556 50942
rect 17500 50596 17556 50876
rect 17500 50530 17556 50540
rect 17724 50932 17780 50942
rect 17388 49812 17444 49822
rect 17388 49810 17556 49812
rect 17388 49758 17390 49810
rect 17442 49758 17556 49810
rect 17388 49756 17556 49758
rect 17388 49746 17444 49756
rect 17276 49196 17444 49252
rect 17164 49186 17220 49196
rect 17276 49028 17332 49038
rect 17276 48934 17332 48972
rect 16940 48802 16996 48814
rect 16940 48750 16942 48802
rect 16994 48750 16996 48802
rect 16828 48244 16884 48254
rect 16716 48242 16884 48244
rect 16716 48190 16830 48242
rect 16882 48190 16884 48242
rect 16716 48188 16884 48190
rect 16828 48178 16884 48188
rect 16828 48020 16884 48030
rect 16940 48020 16996 48750
rect 16884 47964 16996 48020
rect 16828 47954 16884 47964
rect 16268 47842 16324 47852
rect 16380 47852 16548 47908
rect 16716 47908 16772 47918
rect 17052 47908 17108 48860
rect 16156 47348 16212 47358
rect 16156 47254 16212 47292
rect 16044 47012 16324 47068
rect 15820 46844 16100 46900
rect 15708 45666 15764 45678
rect 15708 45614 15710 45666
rect 15762 45614 15764 45666
rect 15708 45106 15764 45614
rect 15708 45054 15710 45106
rect 15762 45054 15764 45106
rect 15708 45042 15764 45054
rect 15596 43598 15598 43650
rect 15650 43598 15652 43650
rect 15596 43586 15652 43598
rect 15820 43538 15876 46844
rect 15932 46674 15988 46686
rect 15932 46622 15934 46674
rect 15986 46622 15988 46674
rect 15932 46452 15988 46622
rect 16044 46564 16100 46844
rect 16044 46498 16100 46508
rect 15932 46386 15988 46396
rect 16156 46450 16212 46462
rect 16156 46398 16158 46450
rect 16210 46398 16212 46450
rect 16156 45444 16212 46398
rect 16156 45378 16212 45388
rect 16044 45108 16100 45118
rect 16044 45014 16100 45052
rect 16268 44324 16324 47012
rect 15820 43486 15822 43538
rect 15874 43486 15876 43538
rect 15820 43474 15876 43486
rect 15932 44268 16324 44324
rect 15484 42802 15540 42812
rect 15820 42196 15876 42206
rect 15484 41972 15540 41982
rect 15484 41858 15540 41916
rect 15484 41806 15486 41858
rect 15538 41806 15540 41858
rect 15484 41794 15540 41806
rect 15708 41970 15764 41982
rect 15708 41918 15710 41970
rect 15762 41918 15764 41970
rect 15260 41234 15316 41244
rect 15596 41300 15652 41310
rect 15148 40350 15150 40402
rect 15202 40350 15204 40402
rect 15148 40338 15204 40350
rect 15596 40402 15652 41244
rect 15596 40350 15598 40402
rect 15650 40350 15652 40402
rect 15596 40338 15652 40350
rect 15708 40404 15764 41918
rect 15708 40338 15764 40348
rect 14588 40290 14756 40292
rect 14588 40238 14590 40290
rect 14642 40238 14756 40290
rect 14588 40236 14756 40238
rect 14588 40226 14644 40236
rect 14364 40124 14532 40180
rect 14140 39666 14196 39676
rect 14252 39620 14308 39630
rect 14140 39508 14196 39518
rect 14140 38052 14196 39452
rect 14252 38948 14308 39564
rect 14364 38948 14420 38958
rect 14252 38946 14420 38948
rect 14252 38894 14366 38946
rect 14418 38894 14420 38946
rect 14252 38892 14420 38894
rect 14252 38500 14308 38892
rect 14364 38882 14420 38892
rect 14252 38434 14308 38444
rect 14476 38388 14532 40124
rect 14588 39394 14644 39406
rect 14588 39342 14590 39394
rect 14642 39342 14644 39394
rect 14588 38836 14644 39342
rect 14588 38770 14644 38780
rect 14476 38322 14532 38332
rect 14140 37996 14644 38052
rect 14364 37826 14420 37838
rect 14364 37774 14366 37826
rect 14418 37774 14420 37826
rect 14364 35924 14420 37774
rect 14476 37604 14532 37614
rect 14476 37156 14532 37548
rect 14476 37062 14532 37100
rect 14476 36820 14532 36830
rect 14476 36482 14532 36764
rect 14476 36430 14478 36482
rect 14530 36430 14532 36482
rect 14476 36418 14532 36430
rect 14364 35868 14532 35924
rect 14364 35588 14420 35598
rect 14364 35494 14420 35532
rect 14028 34190 14030 34242
rect 14082 34190 14084 34242
rect 14028 34178 14084 34190
rect 14140 34692 14196 34702
rect 14140 34244 14196 34636
rect 14140 34178 14196 34188
rect 14476 34130 14532 35868
rect 14588 35700 14644 37996
rect 14700 36484 14756 40236
rect 15820 40180 15876 42140
rect 15820 40114 15876 40124
rect 15260 39508 15316 39518
rect 14924 39172 14980 39182
rect 14812 38834 14868 38846
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38276 14868 38782
rect 14812 37268 14868 38220
rect 14812 37202 14868 37212
rect 14924 38836 14980 39116
rect 14924 37266 14980 38780
rect 15260 38834 15316 39452
rect 15932 39358 15988 44268
rect 16044 44098 16100 44110
rect 16044 44046 16046 44098
rect 16098 44046 16100 44098
rect 16044 43652 16100 44046
rect 16044 43586 16100 43596
rect 16156 44100 16212 44110
rect 16380 44100 16436 47852
rect 16604 47460 16660 47470
rect 16492 47124 16548 47134
rect 16492 44548 16548 47068
rect 16604 46674 16660 47404
rect 16604 46622 16606 46674
rect 16658 46622 16660 46674
rect 16604 46610 16660 46622
rect 16716 46676 16772 47852
rect 16940 47852 17108 47908
rect 17276 48244 17332 48254
rect 16940 47796 16996 47852
rect 17276 47796 17332 48188
rect 16716 46610 16772 46620
rect 16828 47740 16996 47796
rect 17052 47740 17332 47796
rect 16716 46452 16772 46462
rect 16604 44548 16660 44558
rect 16492 44546 16660 44548
rect 16492 44494 16606 44546
rect 16658 44494 16660 44546
rect 16492 44492 16660 44494
rect 16604 44482 16660 44492
rect 16044 43428 16100 43438
rect 16044 43334 16100 43372
rect 16044 42644 16100 42654
rect 16044 42550 16100 42588
rect 16044 42420 16100 42430
rect 16044 41636 16100 42364
rect 16156 41970 16212 44044
rect 16268 44044 16436 44100
rect 16268 42308 16324 44044
rect 16380 43876 16436 43886
rect 16716 43876 16772 46396
rect 16828 44546 16884 47740
rect 16940 47124 16996 47134
rect 16940 46900 16996 47068
rect 16940 46834 16996 46844
rect 16940 46116 16996 46126
rect 16940 45780 16996 46060
rect 17052 45892 17108 47740
rect 17164 47572 17220 47582
rect 17164 47478 17220 47516
rect 17276 47460 17332 47470
rect 17276 47366 17332 47404
rect 17276 46900 17332 46910
rect 17276 46674 17332 46844
rect 17276 46622 17278 46674
rect 17330 46622 17332 46674
rect 17276 46610 17332 46622
rect 17388 46228 17444 49196
rect 17052 45826 17108 45836
rect 17164 46172 17444 46228
rect 16940 45686 16996 45724
rect 16828 44494 16830 44546
rect 16882 44494 16884 44546
rect 16828 44482 16884 44494
rect 16940 45444 16996 45454
rect 16940 44434 16996 45388
rect 17052 45106 17108 45118
rect 17052 45054 17054 45106
rect 17106 45054 17108 45106
rect 17052 44772 17108 45054
rect 17052 44706 17108 44716
rect 17164 44548 17220 46172
rect 17388 46002 17444 46014
rect 17388 45950 17390 46002
rect 17442 45950 17444 46002
rect 16940 44382 16942 44434
rect 16994 44382 16996 44434
rect 16940 44370 16996 44382
rect 17052 44492 17220 44548
rect 17276 44772 17332 44782
rect 16828 43876 16884 43886
rect 16716 43820 16828 43876
rect 16380 43650 16436 43820
rect 16380 43598 16382 43650
rect 16434 43598 16436 43650
rect 16380 43586 16436 43598
rect 16828 43650 16884 43820
rect 16828 43598 16830 43650
rect 16882 43598 16884 43650
rect 16828 43586 16884 43598
rect 16492 43428 16548 43438
rect 16492 43334 16548 43372
rect 16828 42308 16884 42318
rect 16324 42252 16436 42308
rect 16268 42242 16324 42252
rect 16156 41918 16158 41970
rect 16210 41918 16212 41970
rect 16156 41906 16212 41918
rect 16100 41580 16324 41636
rect 16044 41570 16100 41580
rect 16268 41412 16324 41580
rect 16380 41524 16436 42252
rect 16828 41970 16884 42252
rect 16828 41918 16830 41970
rect 16882 41918 16884 41970
rect 16828 41906 16884 41918
rect 16492 41858 16548 41870
rect 16492 41806 16494 41858
rect 16546 41806 16548 41858
rect 16492 41748 16548 41806
rect 16548 41692 16660 41748
rect 16492 41682 16548 41692
rect 16380 41468 16548 41524
rect 16268 41356 16436 41412
rect 16044 41300 16100 41310
rect 16044 41206 16100 41244
rect 16156 40180 16212 40190
rect 16156 39842 16212 40124
rect 16156 39790 16158 39842
rect 16210 39790 16212 39842
rect 16156 39778 16212 39790
rect 16268 39732 16324 39742
rect 16044 39508 16100 39518
rect 16044 39414 16100 39452
rect 15932 39302 16212 39358
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 15260 38388 15316 38782
rect 15820 39172 15876 39182
rect 15820 38834 15876 39116
rect 15820 38782 15822 38834
rect 15874 38782 15876 38834
rect 15820 38770 15876 38782
rect 15260 38322 15316 38332
rect 15372 38610 15428 38622
rect 15372 38558 15374 38610
rect 15426 38558 15428 38610
rect 15372 38276 15428 38558
rect 15372 38220 15764 38276
rect 15148 38162 15204 38174
rect 15148 38110 15150 38162
rect 15202 38110 15204 38162
rect 15036 38050 15092 38062
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37828 15092 37998
rect 15036 37762 15092 37772
rect 14924 37214 14926 37266
rect 14978 37214 14980 37266
rect 14924 37202 14980 37214
rect 15036 37156 15092 37166
rect 14924 36596 14980 36606
rect 14924 36502 14980 36540
rect 14700 36418 14756 36428
rect 14924 36260 14980 36270
rect 14924 35700 14980 36204
rect 14588 35644 14756 35700
rect 14476 34078 14478 34130
rect 14530 34078 14532 34130
rect 14476 34066 14532 34078
rect 14588 35476 14644 35486
rect 13916 33964 14420 34020
rect 13692 33628 13860 33684
rect 14028 33796 14084 33806
rect 13692 30212 13748 33628
rect 13916 33572 13972 33582
rect 13916 33478 13972 33516
rect 13804 33460 13860 33470
rect 13804 33346 13860 33404
rect 13804 33294 13806 33346
rect 13858 33294 13860 33346
rect 13804 33282 13860 33294
rect 13916 32340 13972 32350
rect 13916 32246 13972 32284
rect 13916 31780 13972 31790
rect 13916 30994 13972 31724
rect 13916 30942 13918 30994
rect 13970 30942 13972 30994
rect 13804 30436 13860 30446
rect 13804 30342 13860 30380
rect 13692 30156 13860 30212
rect 13580 29922 13636 29932
rect 13468 29586 13524 29596
rect 13692 29876 13748 29886
rect 13692 29652 13748 29820
rect 13692 29586 13748 29596
rect 13580 28756 13636 28766
rect 13356 28590 13358 28642
rect 13410 28590 13412 28642
rect 13356 28084 13412 28590
rect 13356 28018 13412 28028
rect 13468 28754 13636 28756
rect 13468 28702 13582 28754
rect 13634 28702 13636 28754
rect 13468 28700 13636 28702
rect 13020 27748 13076 27758
rect 13020 27654 13076 27692
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 27076 12964 27134
rect 12908 27010 12964 27020
rect 13020 27412 13076 27422
rect 12796 26238 12798 26290
rect 12850 26238 12852 26290
rect 12796 26226 12852 26238
rect 12908 26852 12964 26862
rect 12236 25730 12404 25732
rect 12236 25678 12238 25730
rect 12290 25678 12404 25730
rect 12236 25676 12404 25678
rect 12572 26180 12628 26190
rect 12236 25666 12292 25676
rect 12460 25396 12516 25406
rect 11900 21410 11956 21420
rect 12012 22540 12180 22596
rect 12236 24836 12292 24846
rect 12012 21700 12068 22540
rect 12124 22372 12180 22382
rect 12124 22278 12180 22316
rect 12124 21812 12180 21822
rect 12124 21718 12180 21756
rect 12012 20804 12068 21644
rect 12124 20804 12180 20814
rect 12012 20802 12180 20804
rect 12012 20750 12126 20802
rect 12178 20750 12180 20802
rect 12012 20748 12180 20750
rect 12124 20738 12180 20748
rect 11788 20626 11844 20636
rect 11564 20078 11566 20130
rect 11618 20078 11620 20130
rect 11564 20066 11620 20078
rect 11900 20468 11956 20478
rect 11788 19908 11844 19918
rect 11788 19814 11844 19852
rect 11452 18050 11508 18060
rect 11788 19234 11844 19246
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 11452 17892 11508 17902
rect 11452 17798 11508 17836
rect 11340 16046 11342 16098
rect 11394 16046 11396 16098
rect 11340 16034 11396 16046
rect 11340 14530 11396 14542
rect 11340 14478 11342 14530
rect 11394 14478 11396 14530
rect 11116 13458 11172 13468
rect 11228 13860 11284 13870
rect 11004 13300 11060 13310
rect 10892 12964 10948 12974
rect 10892 12870 10948 12908
rect 10892 10836 10948 10846
rect 10892 10742 10948 10780
rect 11004 10612 11060 13244
rect 11116 13074 11172 13086
rect 11116 13022 11118 13074
rect 11170 13022 11172 13074
rect 11116 11844 11172 13022
rect 11228 12178 11284 13804
rect 11340 13188 11396 14478
rect 11340 13122 11396 13132
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 11228 12114 11284 12126
rect 11676 12962 11732 12974
rect 11676 12910 11678 12962
rect 11730 12910 11732 12962
rect 11116 11778 11172 11788
rect 11564 11620 11620 11630
rect 11228 11506 11284 11518
rect 11228 11454 11230 11506
rect 11282 11454 11284 11506
rect 11116 11396 11172 11406
rect 11116 11302 11172 11340
rect 11004 10546 11060 10556
rect 11116 10836 11172 10846
rect 11004 10052 11060 10062
rect 11004 9958 11060 9996
rect 10780 9874 10836 9884
rect 11004 9380 11060 9390
rect 11004 9266 11060 9324
rect 11004 9214 11006 9266
rect 11058 9214 11060 9266
rect 11004 9202 11060 9214
rect 11004 8820 11060 8830
rect 10892 8260 10948 8270
rect 10892 8166 10948 8204
rect 10668 8082 10724 8092
rect 10556 7858 10612 7868
rect 10556 7476 10612 7486
rect 10556 6690 10612 7420
rect 10556 6638 10558 6690
rect 10610 6638 10612 6690
rect 10556 6626 10612 6638
rect 10668 7474 10724 7486
rect 10668 7422 10670 7474
rect 10722 7422 10724 7474
rect 10668 6468 10724 7422
rect 10668 6402 10724 6412
rect 10780 6916 10836 6926
rect 10780 6578 10836 6860
rect 10780 6526 10782 6578
rect 10834 6526 10836 6578
rect 10780 6244 10836 6526
rect 10780 6178 10836 6188
rect 10892 5908 10948 5918
rect 10892 5814 10948 5852
rect 10892 5348 10948 5358
rect 10444 5070 10446 5122
rect 10498 5070 10500 5122
rect 10444 5058 10500 5070
rect 10780 5124 10836 5134
rect 10556 5012 10612 5022
rect 10444 4564 10500 4574
rect 10444 4470 10500 4508
rect 10556 3388 10612 4956
rect 10668 4228 10724 4238
rect 10668 3554 10724 4172
rect 10668 3502 10670 3554
rect 10722 3502 10724 3554
rect 10668 3490 10724 3502
rect 10332 3332 10500 3388
rect 10556 3332 10724 3388
rect 10108 112 10164 3332
rect 10332 1202 10388 1214
rect 10332 1150 10334 1202
rect 10386 1150 10388 1202
rect 10332 196 10388 1150
rect 10444 1204 10500 3332
rect 10556 2996 10612 3006
rect 10668 2996 10724 3332
rect 10556 2994 10724 2996
rect 10556 2942 10558 2994
rect 10610 2942 10724 2994
rect 10556 2940 10724 2942
rect 10556 2930 10612 2940
rect 10780 2210 10836 5068
rect 10892 4226 10948 5292
rect 10892 4174 10894 4226
rect 10946 4174 10948 4226
rect 10892 4162 10948 4174
rect 11004 3388 11060 8764
rect 11116 7476 11172 10780
rect 11228 10612 11284 11454
rect 11452 10724 11508 10734
rect 11452 10630 11508 10668
rect 11340 10612 11396 10622
rect 11228 10610 11396 10612
rect 11228 10558 11342 10610
rect 11394 10558 11396 10610
rect 11228 10556 11396 10558
rect 11340 10546 11396 10556
rect 11564 10612 11620 11564
rect 11676 11508 11732 12910
rect 11788 12404 11844 19182
rect 11900 16212 11956 20412
rect 12124 19906 12180 19918
rect 12124 19854 12126 19906
rect 12178 19854 12180 19906
rect 12012 19796 12068 19806
rect 12012 19702 12068 19740
rect 12012 19460 12068 19470
rect 12124 19460 12180 19854
rect 12236 19908 12292 24780
rect 12348 22596 12404 22606
rect 12348 22148 12404 22540
rect 12348 22082 12404 22092
rect 12236 19842 12292 19852
rect 12068 19404 12180 19460
rect 12012 19394 12068 19404
rect 12460 19348 12516 25340
rect 12572 23716 12628 26124
rect 12796 25844 12852 25854
rect 12572 23492 12628 23660
rect 12572 23426 12628 23436
rect 12684 24276 12740 24286
rect 12124 19292 12516 19348
rect 12572 22370 12628 22382
rect 12572 22318 12574 22370
rect 12626 22318 12628 22370
rect 12012 19236 12068 19246
rect 12124 19236 12180 19292
rect 12012 19234 12180 19236
rect 12012 19182 12014 19234
rect 12066 19182 12180 19234
rect 12012 19180 12180 19182
rect 12012 19170 12068 19180
rect 12572 18788 12628 22318
rect 12684 21476 12740 24220
rect 12796 22708 12852 25788
rect 12908 25506 12964 26796
rect 13020 26290 13076 27356
rect 13132 27076 13188 27804
rect 13356 27860 13412 27870
rect 13468 27860 13524 28700
rect 13580 28690 13636 28700
rect 13692 28532 13748 28542
rect 13692 27970 13748 28476
rect 13692 27918 13694 27970
rect 13746 27918 13748 27970
rect 13692 27906 13748 27918
rect 13356 27858 13524 27860
rect 13356 27806 13358 27858
rect 13410 27806 13524 27858
rect 13356 27804 13524 27806
rect 13356 27794 13412 27804
rect 13244 27636 13300 27646
rect 13244 27634 13412 27636
rect 13244 27582 13246 27634
rect 13298 27582 13412 27634
rect 13244 27580 13412 27582
rect 13244 27570 13300 27580
rect 13244 27076 13300 27086
rect 13132 27074 13300 27076
rect 13132 27022 13246 27074
rect 13298 27022 13300 27074
rect 13132 27020 13300 27022
rect 13244 26852 13300 27020
rect 13244 26786 13300 26796
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 13020 26226 13076 26238
rect 13244 26292 13300 26302
rect 13356 26292 13412 27580
rect 13580 27076 13636 27086
rect 13692 27076 13748 27086
rect 13636 27074 13748 27076
rect 13636 27022 13694 27074
rect 13746 27022 13748 27074
rect 13636 27020 13748 27022
rect 13804 27076 13860 30156
rect 13916 29092 13972 30942
rect 13916 29026 13972 29036
rect 14028 28084 14084 33740
rect 14364 33458 14420 33964
rect 14364 33406 14366 33458
rect 14418 33406 14420 33458
rect 14364 33394 14420 33406
rect 14476 32452 14532 32462
rect 14476 31666 14532 32396
rect 14476 31614 14478 31666
rect 14530 31614 14532 31666
rect 14476 31108 14532 31614
rect 14588 31332 14644 35420
rect 14700 35252 14756 35644
rect 14924 35634 14980 35644
rect 14700 32564 14756 35196
rect 14812 35028 14868 35038
rect 14812 34934 14868 34972
rect 15036 34244 15092 37100
rect 15148 37044 15204 38110
rect 15148 36978 15204 36988
rect 15372 38052 15428 38062
rect 15372 37266 15428 37996
rect 15708 38050 15764 38220
rect 15708 37998 15710 38050
rect 15762 37998 15764 38050
rect 15708 37986 15764 37998
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 15260 36148 15316 36158
rect 14924 34188 15092 34244
rect 15148 36092 15260 36148
rect 14812 34132 14868 34142
rect 14812 34038 14868 34076
rect 14924 33572 14980 34188
rect 15036 34020 15092 34030
rect 15148 34020 15204 36092
rect 15260 36082 15316 36092
rect 15372 35140 15428 37214
rect 15820 37828 15876 37838
rect 15484 37044 15540 37054
rect 15484 36950 15540 36988
rect 15820 36708 15876 37772
rect 16044 37828 16100 37838
rect 16044 37734 16100 37772
rect 15932 37268 15988 37278
rect 15932 37174 15988 37212
rect 16044 36708 16100 36718
rect 15820 36706 16100 36708
rect 15820 36654 16046 36706
rect 16098 36654 16100 36706
rect 15820 36652 16100 36654
rect 16044 36642 16100 36652
rect 15596 36372 15652 36382
rect 15596 35588 15652 36316
rect 15820 36260 15876 36270
rect 15820 35700 15876 36204
rect 15820 35634 15876 35644
rect 15596 35522 15652 35532
rect 15036 34018 15204 34020
rect 15036 33966 15038 34018
rect 15090 33966 15204 34018
rect 15036 33964 15204 33966
rect 15260 35084 15428 35140
rect 15484 35474 15540 35486
rect 15484 35422 15486 35474
rect 15538 35422 15540 35474
rect 15036 33954 15092 33964
rect 14700 32498 14756 32508
rect 14812 33516 14980 33572
rect 14588 31266 14644 31276
rect 14812 31220 14868 33516
rect 15260 33460 15316 35084
rect 15372 34916 15428 34926
rect 15372 34692 15428 34860
rect 15372 34626 15428 34636
rect 15484 34130 15540 35422
rect 16156 35140 16212 39302
rect 16268 38388 16324 39676
rect 16268 38322 16324 38332
rect 15484 34078 15486 34130
rect 15538 34078 15540 34130
rect 15484 34066 15540 34078
rect 15708 34580 15764 34590
rect 15596 33908 15652 33918
rect 15372 33460 15428 33470
rect 15260 33404 15372 33460
rect 14924 33348 14980 33358
rect 14924 33254 14980 33292
rect 15148 33348 15204 33358
rect 15036 32564 15092 32574
rect 15036 32470 15092 32508
rect 14924 31892 14980 31902
rect 14924 31798 14980 31836
rect 14812 31164 14980 31220
rect 14476 31052 14868 31108
rect 14140 30996 14196 31006
rect 14140 30882 14196 30940
rect 14140 30830 14142 30882
rect 14194 30830 14196 30882
rect 14140 30818 14196 30830
rect 14588 30882 14644 30894
rect 14588 30830 14590 30882
rect 14642 30830 14644 30882
rect 14588 30436 14644 30830
rect 14588 30370 14644 30380
rect 14476 30212 14532 30222
rect 14364 29988 14420 29998
rect 13916 28028 14084 28084
rect 14140 29314 14196 29326
rect 14140 29262 14142 29314
rect 14194 29262 14196 29314
rect 13916 27524 13972 28028
rect 14028 27860 14084 27870
rect 14028 27766 14084 27804
rect 13916 27468 14084 27524
rect 13916 27300 13972 27310
rect 13916 27206 13972 27244
rect 13804 27020 13972 27076
rect 13580 26628 13636 27020
rect 13692 27010 13748 27020
rect 13580 26562 13636 26572
rect 13468 26292 13524 26302
rect 13356 26290 13524 26292
rect 13356 26238 13470 26290
rect 13522 26238 13524 26290
rect 13356 26236 13524 26238
rect 13244 26198 13300 26236
rect 13468 26226 13524 26236
rect 13580 26180 13636 26190
rect 12908 25454 12910 25506
rect 12962 25454 12964 25506
rect 12908 24162 12964 25454
rect 13132 26068 13188 26078
rect 13132 25284 13188 26012
rect 13468 25844 13524 25854
rect 13356 25620 13412 25630
rect 13244 25506 13300 25518
rect 13244 25454 13246 25506
rect 13298 25454 13300 25506
rect 13244 25396 13300 25454
rect 13244 25330 13300 25340
rect 13132 25218 13188 25228
rect 12908 24110 12910 24162
rect 12962 24110 12964 24162
rect 12908 24098 12964 24110
rect 12908 22932 12964 22942
rect 12908 22930 13300 22932
rect 12908 22878 12910 22930
rect 12962 22878 13300 22930
rect 12908 22876 13300 22878
rect 12908 22866 12964 22876
rect 12796 22652 12964 22708
rect 12796 22482 12852 22494
rect 12796 22430 12798 22482
rect 12850 22430 12852 22482
rect 12796 22148 12852 22430
rect 12796 22082 12852 22092
rect 12796 21476 12852 21486
rect 12684 21474 12852 21476
rect 12684 21422 12798 21474
rect 12850 21422 12852 21474
rect 12684 21420 12852 21422
rect 12796 21252 12852 21420
rect 12796 21186 12852 21196
rect 12908 21252 12964 22652
rect 13244 22482 13300 22876
rect 13244 22430 13246 22482
rect 13298 22430 13300 22482
rect 13244 22418 13300 22430
rect 13132 21812 13188 21822
rect 13132 21586 13188 21756
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 13132 21522 13188 21534
rect 13020 21252 13076 21262
rect 12908 21196 13020 21252
rect 12684 20914 12740 20926
rect 12684 20862 12686 20914
rect 12738 20862 12740 20914
rect 12684 20692 12740 20862
rect 12684 20244 12740 20636
rect 12684 20178 12740 20188
rect 12796 19236 12852 19246
rect 12796 19142 12852 19180
rect 12572 18732 12852 18788
rect 12684 18564 12740 18574
rect 12124 18452 12180 18462
rect 12124 18450 12628 18452
rect 12124 18398 12126 18450
rect 12178 18398 12628 18450
rect 12124 18396 12628 18398
rect 12124 18386 12180 18396
rect 12348 18228 12404 18238
rect 11900 16146 11956 16156
rect 12012 17780 12068 17790
rect 12012 16882 12068 17724
rect 12236 17668 12292 17678
rect 12236 17574 12292 17612
rect 12012 16830 12014 16882
rect 12066 16830 12068 16882
rect 11788 12338 11844 12348
rect 11900 14530 11956 14542
rect 11900 14478 11902 14530
rect 11954 14478 11956 14530
rect 11900 11788 11956 14478
rect 12012 12178 12068 16830
rect 12348 15428 12404 18172
rect 12348 15362 12404 15372
rect 12460 16098 12516 16110
rect 12460 16046 12462 16098
rect 12514 16046 12516 16098
rect 12124 15204 12180 15214
rect 12124 15110 12180 15148
rect 12348 14980 12404 14990
rect 12460 14980 12516 16046
rect 12404 14924 12516 14980
rect 12124 14532 12180 14542
rect 12124 14438 12180 14476
rect 12124 13972 12180 13982
rect 12124 13878 12180 13916
rect 12348 12962 12404 14924
rect 12572 14532 12628 18396
rect 12684 17890 12740 18508
rect 12684 17838 12686 17890
rect 12738 17838 12740 17890
rect 12684 17826 12740 17838
rect 12796 17444 12852 18732
rect 12908 18452 12964 21196
rect 13020 21186 13076 21196
rect 13132 20020 13188 20030
rect 12908 18386 12964 18396
rect 13020 20018 13188 20020
rect 13020 19966 13134 20018
rect 13186 19966 13188 20018
rect 13020 19964 13188 19966
rect 13020 19236 13076 19964
rect 13132 19954 13188 19964
rect 13356 19796 13412 25564
rect 13468 23828 13524 25788
rect 13468 23762 13524 23772
rect 13580 20580 13636 26124
rect 13692 23828 13748 23838
rect 13692 23380 13748 23772
rect 13692 23314 13748 23324
rect 13804 23492 13860 23502
rect 13804 23268 13860 23436
rect 13804 23202 13860 23212
rect 13804 22484 13860 22494
rect 13692 22372 13748 22382
rect 13692 21586 13748 22316
rect 13804 22370 13860 22428
rect 13804 22318 13806 22370
rect 13858 22318 13860 22370
rect 13804 22036 13860 22318
rect 13804 21970 13860 21980
rect 13916 21812 13972 27020
rect 14028 24724 14084 27468
rect 14140 26908 14196 29262
rect 14364 28980 14420 29932
rect 14476 29876 14532 30156
rect 14476 29810 14532 29820
rect 14588 30100 14644 30110
rect 14476 29426 14532 29438
rect 14476 29374 14478 29426
rect 14530 29374 14532 29426
rect 14476 29204 14532 29374
rect 14476 29138 14532 29148
rect 14364 28924 14532 28980
rect 14252 28642 14308 28654
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 14252 27748 14308 28590
rect 14252 27188 14308 27692
rect 14364 27188 14420 27198
rect 14252 27186 14420 27188
rect 14252 27134 14366 27186
rect 14418 27134 14420 27186
rect 14252 27132 14420 27134
rect 14140 26852 14308 26908
rect 14028 24722 14196 24724
rect 14028 24670 14030 24722
rect 14082 24670 14196 24722
rect 14028 24668 14196 24670
rect 14028 24658 14084 24668
rect 14140 23940 14196 24668
rect 14252 24388 14308 26852
rect 14364 25956 14420 27132
rect 14364 25890 14420 25900
rect 14364 25620 14420 25630
rect 14364 25506 14420 25564
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14252 24322 14308 24332
rect 14252 23940 14308 23950
rect 14140 23938 14308 23940
rect 14140 23886 14254 23938
rect 14306 23886 14308 23938
rect 14140 23884 14308 23886
rect 14140 23492 14196 23502
rect 14140 23042 14196 23436
rect 14140 22990 14142 23042
rect 14194 22990 14196 23042
rect 14140 22978 14196 22990
rect 13916 21746 13972 21756
rect 14252 21812 14308 23884
rect 14476 23492 14532 28924
rect 14588 28642 14644 30044
rect 14588 28590 14590 28642
rect 14642 28590 14644 28642
rect 14588 28578 14644 28590
rect 14700 29316 14756 29326
rect 14588 27860 14644 27870
rect 14588 27766 14644 27804
rect 14700 27746 14756 29260
rect 14700 27694 14702 27746
rect 14754 27694 14756 27746
rect 14700 27682 14756 27694
rect 14700 25620 14756 25630
rect 14700 24724 14756 25564
rect 14812 24948 14868 31052
rect 14924 30548 14980 31164
rect 14924 30434 14980 30492
rect 14924 30382 14926 30434
rect 14978 30382 14980 30434
rect 14924 30370 14980 30382
rect 15148 30994 15204 33292
rect 15260 33012 15316 33022
rect 15260 32788 15316 32956
rect 15260 32722 15316 32732
rect 15148 30942 15150 30994
rect 15202 30942 15204 30994
rect 15036 28308 15092 28318
rect 15036 27074 15092 28252
rect 15148 27972 15204 30942
rect 15260 30212 15316 30222
rect 15260 28644 15316 30156
rect 15260 28578 15316 28588
rect 15372 28532 15428 33404
rect 15484 32788 15540 32798
rect 15484 32674 15540 32732
rect 15484 32622 15486 32674
rect 15538 32622 15540 32674
rect 15484 32340 15540 32622
rect 15484 32274 15540 32284
rect 15372 28466 15428 28476
rect 15484 31892 15540 31902
rect 15148 27916 15316 27972
rect 15148 27748 15204 27758
rect 15148 27654 15204 27692
rect 15036 27022 15038 27074
rect 15090 27022 15092 27074
rect 15036 27010 15092 27022
rect 15260 26908 15316 27916
rect 15036 26852 15092 26862
rect 14812 24892 14924 24948
rect 14868 24836 14924 24892
rect 14868 24780 14980 24836
rect 14700 24668 14868 24724
rect 14588 24498 14644 24510
rect 14588 24446 14590 24498
rect 14642 24446 14644 24498
rect 14588 24388 14644 24446
rect 14588 24322 14644 24332
rect 14700 24050 14756 24062
rect 14700 23998 14702 24050
rect 14754 23998 14756 24050
rect 14700 23940 14756 23998
rect 14700 23874 14756 23884
rect 14476 23426 14532 23436
rect 14476 23268 14532 23278
rect 14476 23174 14532 23212
rect 14812 22372 14868 24668
rect 14812 22278 14868 22316
rect 14252 21746 14308 21756
rect 13692 21534 13694 21586
rect 13746 21534 13748 21586
rect 13692 21522 13748 21534
rect 13804 21700 13860 21710
rect 13804 21474 13860 21644
rect 14812 21586 14868 21598
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14252 21476 14308 21486
rect 13804 21422 13806 21474
rect 13858 21422 13860 21474
rect 13804 21410 13860 21422
rect 13916 21474 14308 21476
rect 13916 21422 14254 21474
rect 14306 21422 14308 21474
rect 13916 21420 14308 21422
rect 13804 21028 13860 21038
rect 13916 21028 13972 21420
rect 14252 21410 14308 21420
rect 14812 21252 14868 21534
rect 13804 21026 13972 21028
rect 13804 20974 13806 21026
rect 13858 20974 13972 21026
rect 13804 20972 13972 20974
rect 14252 21196 14868 21252
rect 13804 20962 13860 20972
rect 13580 20514 13636 20524
rect 14140 20244 14196 20254
rect 13580 19908 13636 19918
rect 13580 19814 13636 19852
rect 13020 18450 13076 19180
rect 13020 18398 13022 18450
rect 13074 18398 13076 18450
rect 13020 18228 13076 18398
rect 13244 19740 13412 19796
rect 13244 18452 13300 19740
rect 13356 19460 13412 19470
rect 13356 19366 13412 19404
rect 13468 19348 13524 19358
rect 13468 19254 13524 19292
rect 13244 18386 13300 18396
rect 13020 18162 13076 18172
rect 13356 18338 13412 18350
rect 13356 18286 13358 18338
rect 13410 18286 13412 18338
rect 13356 18116 13412 18286
rect 13244 18060 13412 18116
rect 12796 17378 12852 17388
rect 13020 17780 13076 17790
rect 13020 16322 13076 17724
rect 13244 17220 13300 18060
rect 13244 16772 13300 17164
rect 13356 17668 13412 17678
rect 13356 16994 13412 17612
rect 13804 17444 13860 17454
rect 13804 17442 13972 17444
rect 13804 17390 13806 17442
rect 13858 17390 13972 17442
rect 13804 17388 13972 17390
rect 13804 17378 13860 17388
rect 13356 16942 13358 16994
rect 13410 16942 13412 16994
rect 13356 16930 13412 16942
rect 13580 17220 13636 17230
rect 13468 16772 13524 16782
rect 13244 16716 13468 16772
rect 13468 16706 13524 16716
rect 13020 16270 13022 16322
rect 13074 16270 13076 16322
rect 13020 16258 13076 16270
rect 13580 16322 13636 17164
rect 13916 16996 13972 17388
rect 13804 16772 13860 16782
rect 13804 16678 13860 16716
rect 13580 16270 13582 16322
rect 13634 16270 13636 16322
rect 13580 16258 13636 16270
rect 13804 16436 13860 16446
rect 13356 16098 13412 16110
rect 13356 16046 13358 16098
rect 13410 16046 13412 16098
rect 12908 15986 12964 15998
rect 12908 15934 12910 15986
rect 12962 15934 12964 15986
rect 12908 15316 12964 15934
rect 13244 15764 13300 15774
rect 13132 15316 13188 15326
rect 12796 15202 12852 15214
rect 12796 15150 12798 15202
rect 12850 15150 12852 15202
rect 12796 14756 12852 15150
rect 12908 14980 12964 15260
rect 12908 14914 12964 14924
rect 13020 15314 13188 15316
rect 13020 15262 13134 15314
rect 13186 15262 13188 15314
rect 13020 15260 13188 15262
rect 12796 14690 12852 14700
rect 12572 14466 12628 14476
rect 12908 14532 12964 14542
rect 12908 14438 12964 14476
rect 12572 14308 12628 14318
rect 12348 12910 12350 12962
rect 12402 12910 12404 12962
rect 12348 12898 12404 12910
rect 12460 13188 12516 13198
rect 12012 12126 12014 12178
rect 12066 12126 12068 12178
rect 12012 12114 12068 12126
rect 12236 12404 12292 12414
rect 11676 11442 11732 11452
rect 11788 11732 11956 11788
rect 12012 11844 12068 11854
rect 11564 10518 11620 10556
rect 11676 11284 11732 11294
rect 11564 10164 11620 10174
rect 11452 10052 11508 10062
rect 11340 9940 11396 9950
rect 11340 9268 11396 9884
rect 11452 9716 11508 9996
rect 11452 9622 11508 9660
rect 11452 9268 11508 9278
rect 11340 9266 11508 9268
rect 11340 9214 11454 9266
rect 11506 9214 11508 9266
rect 11340 9212 11508 9214
rect 11452 9202 11508 9212
rect 11564 9042 11620 10108
rect 11564 8990 11566 9042
rect 11618 8990 11620 9042
rect 11564 8978 11620 8990
rect 11676 8820 11732 11228
rect 11788 11172 11844 11732
rect 11900 11508 11956 11518
rect 11900 11394 11956 11452
rect 11900 11342 11902 11394
rect 11954 11342 11956 11394
rect 11900 11330 11956 11342
rect 11788 11116 11956 11172
rect 11788 10388 11844 10398
rect 11788 10294 11844 10332
rect 11900 9604 11956 11116
rect 12012 9938 12068 11788
rect 12236 11394 12292 12348
rect 12236 11342 12238 11394
rect 12290 11342 12292 11394
rect 12236 11284 12292 11342
rect 12236 11218 12292 11228
rect 12348 11956 12404 11966
rect 12124 11172 12180 11182
rect 12124 10050 12180 11116
rect 12348 10948 12404 11900
rect 12348 10882 12404 10892
rect 12460 10724 12516 13132
rect 12460 10658 12516 10668
rect 12124 9998 12126 10050
rect 12178 9998 12180 10050
rect 12124 9986 12180 9998
rect 12348 10612 12404 10622
rect 12348 10052 12404 10556
rect 12572 10388 12628 14252
rect 13020 13972 13076 15260
rect 13132 15250 13188 15260
rect 13244 15148 13300 15708
rect 13020 13906 13076 13916
rect 13132 15092 13300 15148
rect 13132 13748 13188 15092
rect 13244 14868 13300 14878
rect 13244 14420 13300 14812
rect 13244 14354 13300 14364
rect 13244 13972 13300 13982
rect 13356 13972 13412 16046
rect 13468 15986 13524 15998
rect 13468 15934 13470 15986
rect 13522 15934 13524 15986
rect 13468 15652 13524 15934
rect 13468 15586 13524 15596
rect 13580 15764 13636 15774
rect 13580 15540 13636 15708
rect 13580 15474 13636 15484
rect 13580 15316 13636 15326
rect 13580 14196 13636 15260
rect 13804 15202 13860 16380
rect 13804 15150 13806 15202
rect 13858 15150 13860 15202
rect 13804 15138 13860 15150
rect 13804 14644 13860 14654
rect 13580 14130 13636 14140
rect 13692 14532 13748 14542
rect 13244 13970 13412 13972
rect 13244 13918 13246 13970
rect 13298 13918 13412 13970
rect 13244 13916 13412 13918
rect 13580 13972 13636 13982
rect 13244 13906 13300 13916
rect 13580 13878 13636 13916
rect 13356 13748 13412 13758
rect 13132 13692 13300 13748
rect 13132 12964 13188 12974
rect 13132 12870 13188 12908
rect 13020 12628 13076 12638
rect 13020 12180 13076 12572
rect 13244 12628 13300 13692
rect 13244 12562 13300 12572
rect 13020 12114 13076 12124
rect 13356 12290 13412 13692
rect 13356 12238 13358 12290
rect 13410 12238 13412 12290
rect 13132 11732 13188 11742
rect 12908 10610 12964 10622
rect 12908 10558 12910 10610
rect 12962 10558 12964 10610
rect 12908 10500 12964 10558
rect 12908 10434 12964 10444
rect 12572 10322 12628 10332
rect 12348 9996 12740 10052
rect 12012 9886 12014 9938
rect 12066 9886 12068 9938
rect 12012 9874 12068 9886
rect 12236 9940 12292 9950
rect 11900 9538 11956 9548
rect 11788 9380 11844 9390
rect 12236 9380 12292 9884
rect 12684 9938 12740 9996
rect 12684 9886 12686 9938
rect 12738 9886 12740 9938
rect 12684 9874 12740 9886
rect 12796 9940 12852 9950
rect 12796 9846 12852 9884
rect 13132 9716 13188 11676
rect 13132 9650 13188 9660
rect 13244 11394 13300 11406
rect 13244 11342 13246 11394
rect 13298 11342 13300 11394
rect 13244 10612 13300 11342
rect 11844 9324 12292 9380
rect 12572 9604 12628 9614
rect 12572 9380 12628 9548
rect 13244 9380 13300 10556
rect 12572 9324 12740 9380
rect 11788 9042 11844 9324
rect 11788 8990 11790 9042
rect 11842 8990 11844 9042
rect 11788 8978 11844 8990
rect 12236 8932 12292 8942
rect 12236 8930 12516 8932
rect 12236 8878 12238 8930
rect 12290 8878 12516 8930
rect 12236 8876 12516 8878
rect 12236 8866 12292 8876
rect 12124 8820 12180 8830
rect 11452 8764 11732 8820
rect 12012 8818 12180 8820
rect 12012 8766 12126 8818
rect 12178 8766 12180 8818
rect 12012 8764 12180 8766
rect 11340 7476 11396 7486
rect 11116 7474 11396 7476
rect 11116 7422 11342 7474
rect 11394 7422 11396 7474
rect 11116 7420 11396 7422
rect 11116 7140 11172 7420
rect 11340 7410 11396 7420
rect 11116 7074 11172 7084
rect 11228 7250 11284 7262
rect 11452 7252 11508 8764
rect 11564 8372 11620 8382
rect 11564 8370 11732 8372
rect 11564 8318 11566 8370
rect 11618 8318 11732 8370
rect 11564 8316 11732 8318
rect 11564 8306 11620 8316
rect 11228 7198 11230 7250
rect 11282 7198 11284 7250
rect 11228 6804 11284 7198
rect 11228 6738 11284 6748
rect 11340 7196 11508 7252
rect 11564 8148 11620 8158
rect 11116 6690 11172 6702
rect 11116 6638 11118 6690
rect 11170 6638 11172 6690
rect 11116 6468 11172 6638
rect 11116 6244 11172 6412
rect 11116 5124 11172 6188
rect 11116 5058 11172 5068
rect 11340 5122 11396 7196
rect 11564 6690 11620 8092
rect 11676 7476 11732 8316
rect 11788 8258 11844 8270
rect 11788 8206 11790 8258
rect 11842 8206 11844 8258
rect 11788 8036 11844 8206
rect 11788 7812 11844 7980
rect 11788 7746 11844 7756
rect 11900 8260 11956 8270
rect 11676 7410 11732 7420
rect 11900 7476 11956 8204
rect 12012 7588 12068 8764
rect 12124 8754 12180 8764
rect 12012 7522 12068 7532
rect 12124 8258 12180 8270
rect 12124 8206 12126 8258
rect 12178 8206 12180 8258
rect 11900 7382 11956 7420
rect 11564 6638 11566 6690
rect 11618 6638 11620 6690
rect 11564 6626 11620 6638
rect 11788 6802 11844 6814
rect 11788 6750 11790 6802
rect 11842 6750 11844 6802
rect 11788 6692 11844 6750
rect 11788 6626 11844 6636
rect 11452 6580 11508 6590
rect 11452 5906 11508 6524
rect 11900 6580 11956 6590
rect 11452 5854 11454 5906
rect 11506 5854 11508 5906
rect 11452 5842 11508 5854
rect 11676 6468 11732 6478
rect 11676 5906 11732 6412
rect 11676 5854 11678 5906
rect 11730 5854 11732 5906
rect 11676 5842 11732 5854
rect 11788 6020 11844 6030
rect 11340 5070 11342 5122
rect 11394 5070 11396 5122
rect 11340 5058 11396 5070
rect 11564 4452 11620 4462
rect 11564 4226 11620 4396
rect 11564 4174 11566 4226
rect 11618 4174 11620 4226
rect 11564 4162 11620 4174
rect 11228 4114 11284 4126
rect 11228 4062 11230 4114
rect 11282 4062 11284 4114
rect 11228 3892 11284 4062
rect 11228 3826 11284 3836
rect 11116 3780 11172 3790
rect 11116 3686 11172 3724
rect 11788 3388 11844 5964
rect 11900 5906 11956 6524
rect 12124 6244 12180 8206
rect 12236 7924 12292 7934
rect 12236 7586 12292 7868
rect 12236 7534 12238 7586
rect 12290 7534 12292 7586
rect 12236 6356 12292 7534
rect 12236 6290 12292 6300
rect 12348 7476 12404 7486
rect 12348 6690 12404 7420
rect 12460 7140 12516 8876
rect 12572 8372 12628 8382
rect 12572 8278 12628 8316
rect 12460 7074 12516 7084
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 12124 6178 12180 6188
rect 12012 6020 12068 6030
rect 12012 5926 12068 5964
rect 12236 6020 12292 6030
rect 11900 5854 11902 5906
rect 11954 5854 11956 5906
rect 11900 5842 11956 5854
rect 12124 5908 12180 5918
rect 12236 5908 12292 5964
rect 12124 5906 12292 5908
rect 12124 5854 12126 5906
rect 12178 5854 12292 5906
rect 12124 5852 12292 5854
rect 12124 5842 12180 5852
rect 12236 5236 12292 5246
rect 11900 5124 11956 5134
rect 11900 5030 11956 5068
rect 11900 4116 11956 4126
rect 11900 4022 11956 4060
rect 12236 3778 12292 5180
rect 12348 5124 12404 6638
rect 12684 6692 12740 9324
rect 13244 9314 13300 9324
rect 13356 11284 13412 12238
rect 13356 10164 13412 11228
rect 13580 13748 13636 13758
rect 13356 9714 13412 10108
rect 13356 9662 13358 9714
rect 13410 9662 13412 9714
rect 13132 9156 13188 9166
rect 13356 9156 13412 9662
rect 13132 9154 13412 9156
rect 13132 9102 13134 9154
rect 13186 9102 13412 9154
rect 13132 9100 13412 9102
rect 13468 10388 13524 10398
rect 13132 9090 13188 9100
rect 12796 8484 12852 8494
rect 12796 7362 12852 8428
rect 13244 8484 13300 8494
rect 13244 8263 13300 8428
rect 13244 8211 13246 8263
rect 13298 8211 13300 8263
rect 13132 7700 13188 7710
rect 13132 7474 13188 7644
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 13132 7410 13188 7422
rect 12796 7310 12798 7362
rect 12850 7310 12852 7362
rect 12796 7298 12852 7310
rect 13244 7364 13300 8211
rect 13244 7308 13412 7364
rect 13244 7140 13300 7150
rect 13244 6804 13300 7084
rect 13132 6748 13300 6804
rect 12796 6692 12852 6702
rect 12684 6690 12852 6692
rect 12684 6638 12798 6690
rect 12850 6638 12852 6690
rect 12684 6636 12852 6638
rect 12796 6626 12852 6636
rect 12908 6020 12964 6030
rect 12908 5926 12964 5964
rect 12684 5908 12740 5918
rect 12572 5906 12740 5908
rect 12572 5854 12686 5906
rect 12738 5854 12740 5906
rect 12572 5852 12740 5854
rect 12348 5058 12404 5068
rect 12460 5348 12516 5358
rect 12236 3726 12238 3778
rect 12290 3726 12292 3778
rect 11004 3332 11396 3388
rect 11788 3332 12068 3388
rect 11228 2772 11284 2782
rect 11228 2678 11284 2716
rect 10780 2158 10782 2210
rect 10834 2158 10836 2210
rect 10780 2146 10836 2158
rect 11340 2210 11396 3332
rect 12012 2770 12068 3332
rect 12012 2718 12014 2770
rect 12066 2718 12068 2770
rect 12012 2706 12068 2718
rect 12236 2772 12292 3726
rect 12236 2706 12292 2716
rect 12348 4900 12404 4910
rect 11564 2548 11620 2558
rect 11564 2546 11844 2548
rect 11564 2494 11566 2546
rect 11618 2494 11844 2546
rect 11564 2492 11844 2494
rect 11564 2482 11620 2492
rect 11340 2158 11342 2210
rect 11394 2158 11396 2210
rect 11340 2146 11396 2158
rect 10444 1138 10500 1148
rect 10556 1988 10612 1998
rect 10332 130 10388 140
rect 10556 112 10612 1932
rect 11564 1876 11620 1886
rect 11452 1652 11508 1662
rect 11564 1652 11620 1820
rect 11676 1652 11732 1662
rect 11564 1596 11676 1652
rect 11004 1540 11060 1550
rect 10892 978 10948 990
rect 10892 926 10894 978
rect 10946 926 10948 978
rect 10892 756 10948 926
rect 10892 690 10948 700
rect 11004 112 11060 1484
rect 11228 1092 11284 1102
rect 11228 998 11284 1036
rect 11452 112 11508 1596
rect 11676 1586 11732 1596
rect 11788 1202 11844 2492
rect 12236 2546 12292 2558
rect 12236 2494 12238 2546
rect 12290 2494 12292 2546
rect 12236 2212 12292 2494
rect 12236 2146 12292 2156
rect 12348 1988 12404 4844
rect 12460 2210 12516 5292
rect 12572 5346 12628 5852
rect 12684 5842 12740 5852
rect 13132 5794 13188 6748
rect 13356 6692 13412 7308
rect 13468 7362 13524 10332
rect 13580 9828 13636 13692
rect 13580 9762 13636 9772
rect 13692 12964 13748 14476
rect 13580 8818 13636 8830
rect 13580 8766 13582 8818
rect 13634 8766 13636 8818
rect 13580 8596 13636 8766
rect 13580 8530 13636 8540
rect 13692 8260 13748 12908
rect 13804 12180 13860 14588
rect 13916 13634 13972 16940
rect 14028 16100 14084 16110
rect 14028 16006 14084 16044
rect 13916 13582 13918 13634
rect 13970 13582 13972 13634
rect 13916 13570 13972 13582
rect 13916 13188 13972 13198
rect 13916 12962 13972 13132
rect 14140 13076 14196 20188
rect 14252 15764 14308 21196
rect 14924 21140 14980 24780
rect 14252 15698 14308 15708
rect 14364 21084 14980 21140
rect 15036 23268 15092 26796
rect 15148 26852 15316 26908
rect 15148 25060 15204 26852
rect 15372 26292 15428 26302
rect 15148 24994 15204 25004
rect 15260 26068 15316 26078
rect 15260 23604 15316 26012
rect 14364 16098 14420 21084
rect 14812 20916 14868 20926
rect 14812 20822 14868 20860
rect 14588 20804 14644 20814
rect 14476 20690 14532 20702
rect 14476 20638 14478 20690
rect 14530 20638 14532 20690
rect 14476 20132 14532 20638
rect 14476 20066 14532 20076
rect 14476 19236 14532 19246
rect 14476 19142 14532 19180
rect 14588 18450 14644 20748
rect 14812 20020 14868 20030
rect 14812 19926 14868 19964
rect 14924 19460 14980 19470
rect 15036 19460 15092 23212
rect 15148 23548 15316 23604
rect 15148 23044 15204 23548
rect 15372 23266 15428 26236
rect 15372 23214 15374 23266
rect 15426 23214 15428 23266
rect 15372 23202 15428 23214
rect 15484 23268 15540 31836
rect 15596 30212 15652 33852
rect 15596 30146 15652 30156
rect 15596 28644 15652 28654
rect 15596 25172 15652 28588
rect 15708 27858 15764 34524
rect 16156 34130 16212 35084
rect 16156 34078 16158 34130
rect 16210 34078 16212 34130
rect 16156 34066 16212 34078
rect 16268 37716 16324 37726
rect 16268 33908 16324 37660
rect 16156 33852 16324 33908
rect 16044 33572 16100 33582
rect 16044 33346 16100 33516
rect 16044 33294 16046 33346
rect 16098 33294 16100 33346
rect 16044 33236 16100 33294
rect 16044 33170 16100 33180
rect 15820 32564 15876 32574
rect 15820 32470 15876 32508
rect 16044 32452 16100 32462
rect 16044 31890 16100 32396
rect 16044 31838 16046 31890
rect 16098 31838 16100 31890
rect 16044 31826 16100 31838
rect 16156 31668 16212 33852
rect 16268 32564 16324 32574
rect 16268 32470 16324 32508
rect 15708 27806 15710 27858
rect 15762 27806 15764 27858
rect 15708 27794 15764 27806
rect 15820 31612 16212 31668
rect 15596 25106 15652 25116
rect 15708 24500 15764 24510
rect 15708 24406 15764 24444
rect 15820 23268 15876 31612
rect 16380 31332 16436 41356
rect 16492 37266 16548 41468
rect 16604 40292 16660 41692
rect 16940 41524 16996 41534
rect 16828 40964 16884 40974
rect 16828 40870 16884 40908
rect 16604 40226 16660 40236
rect 16716 40402 16772 40414
rect 16716 40350 16718 40402
rect 16770 40350 16772 40402
rect 16604 39172 16660 39182
rect 16604 38948 16660 39116
rect 16604 38834 16660 38892
rect 16604 38782 16606 38834
rect 16658 38782 16660 38834
rect 16604 38770 16660 38782
rect 16716 38668 16772 40350
rect 16940 39844 16996 41468
rect 16940 39778 16996 39788
rect 16492 37214 16494 37266
rect 16546 37214 16548 37266
rect 16492 34580 16548 37214
rect 16492 34514 16548 34524
rect 16604 38612 16772 38668
rect 16828 39508 16884 39518
rect 16604 32564 16660 38612
rect 16828 37044 16884 39452
rect 16828 36978 16884 36988
rect 17052 36596 17108 44492
rect 17276 43988 17332 44716
rect 17276 43922 17332 43932
rect 17164 43652 17220 43662
rect 17164 43538 17220 43596
rect 17164 43486 17166 43538
rect 17218 43486 17220 43538
rect 17164 41970 17220 43486
rect 17388 43316 17444 45950
rect 17388 43250 17444 43260
rect 17500 45444 17556 49756
rect 17724 48804 17780 50876
rect 17836 50708 17892 50718
rect 17836 50594 17892 50652
rect 17836 50542 17838 50594
rect 17890 50542 17892 50594
rect 17836 50484 17892 50542
rect 17836 50418 17892 50428
rect 17948 49476 18004 52110
rect 18284 52162 18340 52174
rect 18284 52110 18286 52162
rect 18338 52110 18340 52162
rect 18172 51716 18228 51726
rect 18172 50820 18228 51660
rect 18284 51492 18340 52110
rect 18284 51426 18340 51436
rect 18396 52052 18452 53116
rect 18396 51378 18452 51996
rect 18508 52276 18564 52286
rect 18508 51492 18564 52220
rect 18620 51828 18676 53788
rect 18844 53508 18900 54462
rect 18956 54404 19012 55246
rect 19404 55300 19460 56028
rect 19964 55972 20020 57344
rect 20412 56532 20468 57344
rect 20412 56466 20468 56476
rect 20636 56082 20692 56094
rect 20636 56030 20638 56082
rect 20690 56030 20692 56082
rect 19964 55906 20020 55916
rect 20412 55972 20468 55982
rect 20412 55878 20468 55916
rect 19516 55860 19572 55870
rect 19516 55766 19572 55804
rect 20188 55858 20244 55870
rect 20188 55806 20190 55858
rect 20242 55806 20244 55858
rect 20188 55522 20244 55806
rect 20188 55470 20190 55522
rect 20242 55470 20244 55522
rect 20188 55458 20244 55470
rect 20524 55524 20580 55534
rect 20636 55524 20692 56030
rect 20860 56084 20916 57344
rect 20860 56018 20916 56028
rect 20524 55522 20692 55524
rect 20524 55470 20526 55522
rect 20578 55470 20692 55522
rect 20524 55468 20692 55470
rect 20524 55458 20580 55468
rect 19516 55412 19572 55422
rect 19516 55318 19572 55356
rect 20860 55412 20916 55422
rect 20860 55318 20916 55356
rect 19740 55300 19796 55310
rect 19404 55234 19460 55244
rect 19628 55298 19796 55300
rect 19628 55246 19742 55298
rect 19794 55246 19796 55298
rect 19628 55244 19796 55246
rect 18956 54338 19012 54348
rect 19516 54292 19572 54302
rect 19628 54292 19684 55244
rect 19740 55234 19796 55244
rect 20300 55298 20356 55310
rect 20300 55246 20302 55298
rect 20354 55246 20356 55298
rect 20076 54964 20132 54974
rect 19740 54852 19796 54862
rect 19740 54402 19796 54796
rect 19740 54350 19742 54402
rect 19794 54350 19796 54402
rect 19740 54338 19796 54350
rect 19964 54514 20020 54526
rect 19964 54462 19966 54514
rect 20018 54462 20020 54514
rect 19516 54290 19684 54292
rect 19516 54238 19518 54290
rect 19570 54238 19684 54290
rect 19516 54236 19684 54238
rect 19292 54180 19348 54190
rect 19292 53954 19348 54124
rect 19516 54068 19572 54236
rect 19516 54002 19572 54012
rect 19964 54068 20020 54462
rect 20076 54068 20132 54908
rect 20300 54852 20356 55246
rect 21084 55298 21140 55310
rect 21084 55246 21086 55298
rect 21138 55246 21140 55298
rect 21084 55188 21140 55246
rect 20300 54786 20356 54796
rect 20860 55132 21140 55188
rect 20860 54290 20916 55132
rect 21308 54852 21364 57344
rect 21644 56420 21700 56430
rect 21644 56082 21700 56364
rect 21644 56030 21646 56082
rect 21698 56030 21700 56082
rect 21644 56018 21700 56030
rect 21532 55858 21588 55870
rect 21532 55806 21534 55858
rect 21586 55806 21588 55858
rect 21532 55636 21588 55806
rect 21756 55636 21812 57344
rect 22204 56756 22260 57344
rect 22204 56690 22260 56700
rect 22652 56532 22708 57344
rect 22540 56476 22708 56532
rect 21980 55972 22036 55982
rect 21980 55878 22036 55916
rect 21532 55580 21700 55636
rect 21532 55412 21588 55422
rect 20860 54238 20862 54290
rect 20914 54238 20916 54290
rect 20860 54180 20916 54238
rect 20860 54114 20916 54124
rect 20972 54796 21364 54852
rect 21420 55410 21588 55412
rect 21420 55358 21534 55410
rect 21586 55358 21588 55410
rect 21420 55356 21588 55358
rect 20076 54012 20468 54068
rect 19964 54002 20020 54012
rect 19292 53902 19294 53954
rect 19346 53902 19348 53954
rect 19292 53890 19348 53902
rect 20076 53844 20132 53854
rect 20076 53842 20244 53844
rect 20076 53790 20078 53842
rect 20130 53790 20244 53842
rect 20076 53788 20244 53790
rect 20076 53778 20132 53788
rect 18844 53442 18900 53452
rect 19516 53730 19572 53742
rect 19964 53732 20020 53742
rect 19516 53678 19518 53730
rect 19570 53678 19572 53730
rect 18732 52946 18788 52958
rect 18732 52894 18734 52946
rect 18786 52894 18788 52946
rect 18732 52612 18788 52894
rect 19292 52724 19348 52734
rect 19292 52630 19348 52668
rect 19516 52724 19572 53678
rect 19516 52658 19572 52668
rect 19628 53730 20020 53732
rect 19628 53678 19966 53730
rect 20018 53678 20020 53730
rect 19628 53676 20020 53678
rect 18732 52546 18788 52556
rect 19404 52612 19460 52622
rect 18956 52276 19012 52286
rect 18956 52182 19012 52220
rect 19180 52164 19236 52174
rect 19180 52070 19236 52108
rect 19404 52164 19460 52556
rect 19404 52098 19460 52108
rect 19516 52162 19572 52174
rect 19516 52110 19518 52162
rect 19570 52110 19572 52162
rect 19516 52052 19572 52110
rect 19516 51986 19572 51996
rect 18620 51762 18676 51772
rect 19516 51828 19572 51838
rect 18508 51426 18564 51436
rect 18396 51326 18398 51378
rect 18450 51326 18452 51378
rect 18172 50764 18340 50820
rect 17948 49252 18004 49420
rect 18060 50706 18116 50718
rect 18060 50654 18062 50706
rect 18114 50654 18116 50706
rect 18060 49364 18116 50654
rect 18172 50596 18228 50606
rect 18172 49810 18228 50540
rect 18172 49758 18174 49810
rect 18226 49758 18228 49810
rect 18172 49746 18228 49758
rect 18060 49308 18228 49364
rect 17948 49186 18004 49196
rect 18060 49138 18116 49150
rect 18060 49086 18062 49138
rect 18114 49086 18116 49138
rect 17612 48748 17780 48804
rect 17948 49026 18004 49038
rect 17948 48974 17950 49026
rect 18002 48974 18004 49026
rect 17612 48244 17668 48748
rect 17612 48178 17668 48188
rect 17724 48580 17780 48590
rect 17724 47458 17780 48524
rect 17724 47406 17726 47458
rect 17778 47406 17780 47458
rect 17724 47394 17780 47406
rect 17836 47460 17892 47470
rect 17164 41918 17166 41970
rect 17218 41918 17220 41970
rect 17164 41906 17220 41918
rect 17388 41300 17444 41310
rect 17388 41206 17444 41244
rect 17164 40964 17220 40974
rect 17164 40870 17220 40908
rect 17500 38834 17556 45388
rect 17724 45332 17780 45342
rect 17836 45332 17892 47404
rect 17948 46116 18004 48974
rect 18060 47682 18116 49086
rect 18172 48692 18228 49308
rect 18172 48626 18228 48636
rect 18060 47630 18062 47682
rect 18114 47630 18116 47682
rect 18060 47618 18116 47630
rect 18284 48242 18340 50764
rect 18396 50708 18452 51326
rect 18844 51378 18900 51390
rect 18844 51326 18846 51378
rect 18898 51326 18900 51378
rect 18620 51156 18676 51166
rect 18508 50708 18564 50718
rect 18396 50706 18564 50708
rect 18396 50654 18510 50706
rect 18562 50654 18564 50706
rect 18396 50652 18564 50654
rect 18508 50642 18564 50652
rect 18620 50428 18676 51100
rect 18844 50932 18900 51326
rect 18844 50866 18900 50876
rect 19292 50708 19348 50718
rect 18508 50372 18676 50428
rect 19068 50594 19124 50606
rect 19068 50542 19070 50594
rect 19122 50542 19124 50594
rect 18284 48190 18286 48242
rect 18338 48190 18340 48242
rect 18284 47348 18340 48190
rect 18396 49252 18452 49262
rect 18396 47684 18452 49196
rect 18396 47618 18452 47628
rect 18508 48468 18564 50372
rect 18284 47068 18340 47292
rect 17948 46050 18004 46060
rect 18060 47012 18340 47068
rect 17724 45330 17892 45332
rect 17724 45278 17726 45330
rect 17778 45278 17892 45330
rect 17724 45276 17892 45278
rect 17724 45266 17780 45276
rect 17836 44436 17892 44446
rect 17836 44324 17892 44380
rect 17612 44322 17892 44324
rect 17612 44270 17838 44322
rect 17890 44270 17892 44322
rect 17612 44268 17892 44270
rect 17612 42754 17668 44268
rect 17836 44258 17892 44268
rect 17724 43540 17780 43550
rect 18060 43540 18116 47012
rect 18172 46674 18228 46686
rect 18172 46622 18174 46674
rect 18226 46622 18228 46674
rect 18172 46452 18228 46622
rect 18172 46386 18228 46396
rect 18284 46340 18340 46350
rect 18508 46340 18564 48412
rect 18732 49924 18788 49934
rect 18732 49026 18788 49868
rect 19068 49700 19124 50542
rect 19180 49812 19236 49822
rect 19180 49718 19236 49756
rect 19068 49634 19124 49644
rect 18732 48974 18734 49026
rect 18786 48974 18788 49026
rect 18732 47460 18788 48974
rect 18844 49586 18900 49598
rect 18844 49534 18846 49586
rect 18898 49534 18900 49586
rect 18844 49028 18900 49534
rect 19180 49140 19236 49150
rect 18844 48962 18900 48972
rect 18956 49084 19180 49140
rect 17724 43538 18116 43540
rect 17724 43486 17726 43538
rect 17778 43486 18116 43538
rect 17724 43484 18116 43486
rect 18172 45780 18228 45790
rect 18284 45780 18340 46284
rect 18396 46284 18564 46340
rect 18620 47458 18788 47460
rect 18620 47406 18734 47458
rect 18786 47406 18788 47458
rect 18620 47404 18788 47406
rect 18396 45892 18452 46284
rect 18508 46116 18564 46126
rect 18508 46022 18564 46060
rect 18396 45836 18564 45892
rect 18228 45724 18340 45780
rect 18172 44324 18228 45724
rect 18284 44660 18340 44670
rect 18284 44546 18340 44604
rect 18284 44494 18286 44546
rect 18338 44494 18340 44546
rect 18284 44482 18340 44494
rect 18396 44548 18452 44558
rect 18396 44324 18452 44492
rect 18172 44268 18452 44324
rect 17724 43474 17780 43484
rect 17836 43316 17892 43326
rect 17836 43314 18004 43316
rect 17836 43262 17838 43314
rect 17890 43262 18004 43314
rect 17836 43260 18004 43262
rect 17836 43250 17892 43260
rect 17612 42702 17614 42754
rect 17666 42702 17668 42754
rect 17612 42690 17668 42702
rect 17724 42642 17780 42654
rect 17724 42590 17726 42642
rect 17778 42590 17780 42642
rect 17612 41972 17668 41982
rect 17612 41878 17668 41916
rect 17724 41300 17780 42590
rect 17724 41234 17780 41244
rect 17836 41746 17892 41758
rect 17836 41694 17838 41746
rect 17890 41694 17892 41746
rect 17836 40964 17892 41694
rect 17948 41298 18004 43260
rect 18060 42868 18116 42878
rect 18060 42774 18116 42812
rect 17948 41246 17950 41298
rect 18002 41246 18004 41298
rect 17948 41234 18004 41246
rect 17836 40898 17892 40908
rect 17500 38782 17502 38834
rect 17554 38782 17556 38834
rect 16828 36540 17108 36596
rect 17164 37716 17220 37726
rect 16828 36148 16884 36540
rect 16828 36082 16884 36092
rect 16940 36372 16996 36382
rect 17164 36372 17220 37660
rect 17388 37156 17444 37166
rect 17388 36706 17444 37100
rect 17500 36820 17556 38782
rect 18060 37604 18116 37614
rect 17612 37268 17668 37278
rect 17612 37174 17668 37212
rect 17500 36754 17556 36764
rect 17836 36820 17892 36830
rect 17388 36654 17390 36706
rect 17442 36654 17444 36706
rect 17388 36642 17444 36654
rect 16940 36370 17220 36372
rect 16940 36318 16942 36370
rect 16994 36318 17220 36370
rect 16940 36316 17220 36318
rect 16828 35140 16884 35150
rect 16604 32498 16660 32508
rect 16716 34692 16772 34702
rect 16492 32340 16548 32350
rect 16492 32246 16548 32284
rect 16716 31892 16772 34636
rect 16716 31826 16772 31836
rect 16380 31276 16660 31332
rect 16268 30994 16324 31006
rect 16268 30942 16270 30994
rect 16322 30942 16324 30994
rect 15932 30660 15988 30670
rect 15932 28980 15988 30604
rect 16044 30212 16100 30222
rect 16044 30118 16100 30156
rect 15932 28644 15988 28924
rect 15932 28578 15988 28588
rect 16268 28308 16324 30942
rect 16380 29314 16436 29326
rect 16380 29262 16382 29314
rect 16434 29262 16436 29314
rect 16380 28868 16436 29262
rect 16492 29202 16548 29214
rect 16492 29150 16494 29202
rect 16546 29150 16548 29202
rect 16492 29092 16548 29150
rect 16492 29026 16548 29036
rect 16380 28802 16436 28812
rect 16268 28242 16324 28252
rect 16492 28420 16548 28430
rect 16044 27748 16100 27758
rect 16044 27074 16100 27692
rect 16044 27022 16046 27074
rect 16098 27022 16100 27074
rect 16044 26516 16100 27022
rect 16044 26450 16100 26460
rect 16380 27188 16436 27198
rect 16044 25732 16100 25742
rect 15932 23716 15988 23726
rect 15932 23622 15988 23660
rect 15484 23212 15652 23268
rect 15820 23212 15988 23268
rect 15148 22978 15204 22988
rect 15484 23044 15540 23054
rect 15484 22950 15540 22988
rect 15260 22932 15316 22942
rect 15260 22838 15316 22876
rect 15372 22372 15428 22382
rect 15372 20018 15428 22316
rect 15372 19966 15374 20018
rect 15426 19966 15428 20018
rect 15372 19908 15428 19966
rect 15372 19842 15428 19852
rect 15484 20020 15540 20030
rect 14924 19458 15092 19460
rect 14924 19406 14926 19458
rect 14978 19406 15092 19458
rect 14924 19404 15092 19406
rect 14924 18564 14980 19404
rect 14924 18498 14980 18508
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14588 18386 14644 18398
rect 15036 18452 15092 18462
rect 15036 18358 15092 18396
rect 15484 18450 15540 19964
rect 15484 18398 15486 18450
rect 15538 18398 15540 18450
rect 15484 18386 15540 18398
rect 14924 18004 14980 18014
rect 14812 17892 14868 17902
rect 14364 16046 14366 16098
rect 14418 16046 14420 16098
rect 14364 15540 14420 16046
rect 14364 15474 14420 15484
rect 14476 17668 14532 17678
rect 14364 15314 14420 15326
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 14364 15204 14420 15262
rect 14364 15138 14420 15148
rect 14476 14530 14532 17612
rect 14700 16436 14756 16446
rect 14700 16212 14756 16380
rect 14700 16146 14756 16156
rect 14812 16210 14868 17836
rect 14924 17890 14980 17948
rect 14924 17838 14926 17890
rect 14978 17838 14980 17890
rect 14924 17826 14980 17838
rect 15260 17444 15316 17454
rect 14924 17220 14980 17230
rect 14924 17106 14980 17164
rect 14924 17054 14926 17106
rect 14978 17054 14980 17106
rect 14924 17042 14980 17054
rect 15260 16660 15316 17388
rect 15484 17108 15540 17118
rect 15484 17014 15540 17052
rect 15372 16884 15428 16922
rect 15372 16818 15428 16828
rect 15596 16772 15652 23212
rect 15820 23044 15876 23054
rect 15708 23042 15876 23044
rect 15708 22990 15822 23042
rect 15874 22990 15876 23042
rect 15708 22988 15876 22990
rect 15708 22372 15764 22988
rect 15820 22978 15876 22988
rect 15708 22306 15764 22316
rect 15820 22370 15876 22382
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15820 21812 15876 22318
rect 15820 21746 15876 21756
rect 15820 21588 15876 21598
rect 15708 21252 15764 21262
rect 15708 18452 15764 21196
rect 15820 20468 15876 21532
rect 15820 20402 15876 20412
rect 15820 18452 15876 18462
rect 15708 18450 15876 18452
rect 15708 18398 15822 18450
rect 15874 18398 15876 18450
rect 15708 18396 15876 18398
rect 15820 18386 15876 18396
rect 15932 17892 15988 23212
rect 16044 22594 16100 25676
rect 16044 22542 16046 22594
rect 16098 22542 16100 22594
rect 16044 22530 16100 22542
rect 16156 25620 16212 25630
rect 16156 22482 16212 25564
rect 16380 25060 16436 27132
rect 16492 25508 16548 28364
rect 16604 27860 16660 31276
rect 16828 31106 16884 35084
rect 16940 34802 16996 36316
rect 17276 35700 17332 35710
rect 16940 34750 16942 34802
rect 16994 34750 16996 34802
rect 16940 33236 16996 34750
rect 17164 35252 17220 35262
rect 17052 34132 17108 34142
rect 17052 34038 17108 34076
rect 17164 33796 17220 35196
rect 17164 33730 17220 33740
rect 17276 35026 17332 35644
rect 17276 34974 17278 35026
rect 17330 34974 17332 35026
rect 16940 33234 17108 33236
rect 16940 33182 16942 33234
rect 16994 33182 17108 33234
rect 16940 33180 17108 33182
rect 16940 33170 16996 33180
rect 16940 32452 16996 32462
rect 16940 32358 16996 32396
rect 16828 31054 16830 31106
rect 16882 31054 16884 31106
rect 16828 30884 16884 31054
rect 16828 30548 16884 30828
rect 16716 30492 16884 30548
rect 16940 31332 16996 31342
rect 16716 30436 16772 30492
rect 16716 30370 16772 30380
rect 16828 30322 16884 30334
rect 16828 30270 16830 30322
rect 16882 30270 16884 30322
rect 16828 30212 16884 30270
rect 16940 30322 16996 31276
rect 16940 30270 16942 30322
rect 16994 30270 16996 30322
rect 16940 30258 16996 30270
rect 16716 30156 16884 30212
rect 16716 29092 16772 30156
rect 16828 29986 16884 29998
rect 16828 29934 16830 29986
rect 16882 29934 16884 29986
rect 16828 29204 16884 29934
rect 16828 29138 16884 29148
rect 16940 29876 16996 29886
rect 16716 29026 16772 29036
rect 16940 28642 16996 29820
rect 16940 28590 16942 28642
rect 16994 28590 16996 28642
rect 16940 27972 16996 28590
rect 16940 27906 16996 27916
rect 16716 27860 16772 27870
rect 16604 27858 16772 27860
rect 16604 27806 16718 27858
rect 16770 27806 16772 27858
rect 16604 27804 16772 27806
rect 16604 27636 16660 27804
rect 16716 27794 16772 27804
rect 16604 27570 16660 27580
rect 16604 27188 16660 27198
rect 16604 26068 16660 27132
rect 17052 26628 17108 33180
rect 17164 30994 17220 31006
rect 17164 30942 17166 30994
rect 17218 30942 17220 30994
rect 17164 30212 17220 30942
rect 17276 30660 17332 34974
rect 17388 35588 17444 35598
rect 17388 33458 17444 35532
rect 17388 33406 17390 33458
rect 17442 33406 17444 33458
rect 17388 32452 17444 33406
rect 17612 33796 17668 33806
rect 17388 32386 17444 32396
rect 17500 32562 17556 32574
rect 17500 32510 17502 32562
rect 17554 32510 17556 32562
rect 17500 32116 17556 32510
rect 17500 32050 17556 32060
rect 17612 30994 17668 33740
rect 17836 31780 17892 36764
rect 17836 31714 17892 31724
rect 17948 36148 18004 36158
rect 17948 31444 18004 36092
rect 18060 35588 18116 37548
rect 18060 35522 18116 35532
rect 18060 35028 18116 35038
rect 18060 34244 18116 34972
rect 18060 34178 18116 34188
rect 17948 31388 18116 31444
rect 17836 31332 17892 31342
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17612 30930 17668 30942
rect 17724 30996 17780 31006
rect 17276 30604 17444 30660
rect 17164 30146 17220 30156
rect 17276 30436 17332 30446
rect 17388 30436 17444 30604
rect 17388 30380 17556 30436
rect 17164 29421 17220 29433
rect 17164 29369 17166 29421
rect 17218 29369 17220 29421
rect 17164 28532 17220 29369
rect 17164 27188 17220 28476
rect 17164 27122 17220 27132
rect 17276 26908 17332 30380
rect 17388 30210 17444 30222
rect 17388 30158 17390 30210
rect 17442 30158 17444 30210
rect 17388 29876 17444 30158
rect 17388 29810 17444 29820
rect 17388 28756 17444 28766
rect 17500 28756 17556 30380
rect 17388 28754 17556 28756
rect 17388 28702 17390 28754
rect 17442 28702 17556 28754
rect 17388 28700 17556 28702
rect 17388 28196 17444 28700
rect 17388 28130 17444 28140
rect 17500 27972 17556 27982
rect 17500 27878 17556 27916
rect 17612 27076 17668 27086
rect 17276 26852 17444 26908
rect 17388 26786 17444 26796
rect 17612 26628 17668 27020
rect 17052 26572 17444 26628
rect 16940 26460 17332 26516
rect 16828 26292 16884 26302
rect 16828 26198 16884 26236
rect 16604 26002 16660 26012
rect 16492 25442 16548 25452
rect 16828 25956 16884 25966
rect 16716 25394 16772 25406
rect 16716 25342 16718 25394
rect 16770 25342 16772 25394
rect 16716 25284 16772 25342
rect 16380 24994 16436 25004
rect 16492 25228 16772 25284
rect 16492 25172 16548 25228
rect 16268 24500 16324 24510
rect 16268 23154 16324 24444
rect 16492 24052 16548 25116
rect 16828 24724 16884 25900
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 16268 23090 16324 23102
rect 16380 23996 16548 24052
rect 16604 24610 16660 24622
rect 16604 24558 16606 24610
rect 16658 24558 16660 24610
rect 16156 22430 16158 22482
rect 16210 22430 16212 22482
rect 16156 22418 16212 22430
rect 16268 22260 16324 22270
rect 16156 21812 16212 21822
rect 16044 20916 16100 20926
rect 16156 20916 16212 21756
rect 16268 21700 16324 22204
rect 16268 21634 16324 21644
rect 16380 21476 16436 23996
rect 16604 23548 16660 24558
rect 16716 24052 16772 24062
rect 16828 24052 16884 24668
rect 16716 24050 16884 24052
rect 16716 23998 16718 24050
rect 16770 23998 16884 24050
rect 16716 23996 16884 23998
rect 16716 23986 16772 23996
rect 16940 23548 16996 26460
rect 17276 26402 17332 26460
rect 17276 26350 17278 26402
rect 17330 26350 17332 26402
rect 17276 26338 17332 26350
rect 17052 26290 17108 26302
rect 17052 26238 17054 26290
rect 17106 26238 17108 26290
rect 17052 25732 17108 26238
rect 17052 25666 17108 25676
rect 17052 25506 17108 25518
rect 17052 25454 17054 25506
rect 17106 25454 17108 25506
rect 17052 24722 17108 25454
rect 17052 24670 17054 24722
rect 17106 24670 17108 24722
rect 17052 24500 17108 24670
rect 17052 23938 17108 24444
rect 17052 23886 17054 23938
rect 17106 23886 17108 23938
rect 17052 23874 17108 23886
rect 17164 25508 17220 25518
rect 16604 23492 16772 23548
rect 16940 23492 17108 23548
rect 16492 23212 16660 23268
rect 16492 23156 16548 23212
rect 16492 23090 16548 23100
rect 16604 23154 16660 23212
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16604 23090 16660 23102
rect 16044 20914 16212 20916
rect 16044 20862 16046 20914
rect 16098 20862 16212 20914
rect 16044 20860 16212 20862
rect 16268 21420 16436 21476
rect 16492 21474 16548 21486
rect 16492 21422 16494 21474
rect 16546 21422 16548 21474
rect 16044 20850 16100 20860
rect 16156 20468 16212 20478
rect 16044 19460 16100 19470
rect 16044 19366 16100 19404
rect 16044 18340 16100 18350
rect 16156 18340 16212 20412
rect 16268 19572 16324 21420
rect 16268 19506 16324 19516
rect 16380 21140 16436 21150
rect 16268 18788 16324 18798
rect 16268 18564 16324 18732
rect 16268 18498 16324 18508
rect 16044 18338 16212 18340
rect 16044 18286 16046 18338
rect 16098 18286 16212 18338
rect 16044 18284 16212 18286
rect 16044 18274 16100 18284
rect 15932 17826 15988 17836
rect 16268 18228 16324 18238
rect 16044 17668 16100 17678
rect 16044 17574 16100 17612
rect 16156 17556 16212 17566
rect 16156 16994 16212 17500
rect 16156 16942 16158 16994
rect 16210 16942 16212 16994
rect 16156 16930 16212 16942
rect 15596 16706 15652 16716
rect 15260 16594 15316 16604
rect 15484 16658 15540 16670
rect 15484 16606 15486 16658
rect 15538 16606 15540 16658
rect 14812 16158 14814 16210
rect 14866 16158 14868 16210
rect 14812 16146 14868 16158
rect 15484 15876 15540 16606
rect 16044 16212 16100 16222
rect 16044 16118 16100 16156
rect 15596 15876 15652 15886
rect 15484 15820 15596 15876
rect 14812 15316 14868 15326
rect 14476 14478 14478 14530
rect 14530 14478 14532 14530
rect 14364 14420 14420 14430
rect 14364 13634 14420 14364
rect 14364 13582 14366 13634
rect 14418 13582 14420 13634
rect 14364 13570 14420 13582
rect 14476 13188 14532 14478
rect 14476 13122 14532 13132
rect 14588 15314 14868 15316
rect 14588 15262 14814 15314
rect 14866 15262 14868 15314
rect 14588 15260 14868 15262
rect 14252 13076 14308 13086
rect 14140 13074 14308 13076
rect 14140 13022 14254 13074
rect 14306 13022 14308 13074
rect 14140 13020 14308 13022
rect 14252 13010 14308 13020
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12898 13972 12910
rect 14140 12292 14196 12302
rect 13804 12124 13972 12180
rect 13804 11954 13860 11966
rect 13804 11902 13806 11954
rect 13858 11902 13860 11954
rect 13804 11458 13860 11902
rect 13916 11844 13972 12124
rect 13916 11778 13972 11788
rect 13804 11402 14084 11458
rect 13804 11282 13860 11294
rect 13804 11230 13806 11282
rect 13858 11230 13860 11282
rect 13804 10836 13860 11230
rect 13916 11172 13972 11182
rect 13916 11078 13972 11116
rect 14028 10836 14084 11402
rect 13804 10770 13860 10780
rect 13916 10780 14084 10836
rect 13804 9938 13860 9950
rect 13804 9886 13806 9938
rect 13858 9886 13860 9938
rect 13804 9828 13860 9886
rect 13804 9762 13860 9772
rect 13916 8484 13972 10780
rect 14028 10610 14084 10622
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 14028 10164 14084 10558
rect 14028 10098 14084 10108
rect 14140 9268 14196 12236
rect 14588 11458 14644 15260
rect 14812 15250 14868 15260
rect 14924 15204 14980 15214
rect 14812 15092 14980 15148
rect 14812 14642 14868 15092
rect 14812 14590 14814 14642
rect 14866 14590 14868 14642
rect 14812 14578 14868 14590
rect 14924 14980 14980 14990
rect 14812 13860 14868 13870
rect 14924 13860 14980 14924
rect 14812 13858 14980 13860
rect 14812 13806 14814 13858
rect 14866 13806 14980 13858
rect 14812 13804 14980 13806
rect 15036 14196 15092 14206
rect 14812 13794 14868 13804
rect 14700 12180 14756 12190
rect 14700 11620 14756 12124
rect 14924 11954 14980 11966
rect 14924 11902 14926 11954
rect 14978 11902 14980 11954
rect 14700 11564 14868 11620
rect 14812 11506 14868 11564
rect 14364 11394 14420 11406
rect 14588 11402 14756 11458
rect 14812 11454 14814 11506
rect 14866 11454 14868 11506
rect 14812 11442 14868 11454
rect 14364 11342 14366 11394
rect 14418 11342 14420 11394
rect 14364 11284 14420 11342
rect 14364 10948 14420 11228
rect 14588 11284 14644 11294
rect 14588 10948 14644 11228
rect 14364 10882 14420 10892
rect 14476 10892 14644 10948
rect 14476 10500 14532 10892
rect 14700 10724 14756 11402
rect 14924 10836 14980 11902
rect 15036 11620 15092 14140
rect 15596 13972 15652 15820
rect 15820 15316 15876 15326
rect 15708 15314 15876 15316
rect 15708 15262 15822 15314
rect 15874 15262 15876 15314
rect 15708 15260 15876 15262
rect 15708 14420 15764 15260
rect 15820 15250 15876 15260
rect 16156 15204 16212 15214
rect 15708 14354 15764 14364
rect 15820 14756 15876 14766
rect 15260 13746 15316 13758
rect 15260 13694 15262 13746
rect 15314 13694 15316 13746
rect 15036 11554 15092 11564
rect 15148 13524 15204 13534
rect 15036 11396 15092 11406
rect 15148 11396 15204 13468
rect 15260 13188 15316 13694
rect 15596 13746 15652 13916
rect 15596 13694 15598 13746
rect 15650 13694 15652 13746
rect 15596 13682 15652 13694
rect 15820 13634 15876 14700
rect 16156 14532 16212 15148
rect 15820 13582 15822 13634
rect 15874 13582 15876 13634
rect 15820 13570 15876 13582
rect 15932 14476 16212 14532
rect 15260 13122 15316 13132
rect 15372 13300 15428 13310
rect 15372 12964 15428 13244
rect 15484 13188 15540 13198
rect 15484 13094 15540 13132
rect 15372 12908 15540 12964
rect 15372 12068 15428 12078
rect 15260 12066 15428 12068
rect 15260 12014 15374 12066
rect 15426 12014 15428 12066
rect 15260 12012 15428 12014
rect 15260 11732 15316 12012
rect 15372 12002 15428 12012
rect 15484 11788 15540 12908
rect 15820 12962 15876 12974
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15708 12178 15764 12190
rect 15708 12126 15710 12178
rect 15762 12126 15764 12178
rect 15260 11666 15316 11676
rect 15372 11732 15540 11788
rect 15596 11844 15652 11854
rect 15372 11620 15428 11732
rect 15372 11554 15428 11564
rect 15596 11620 15652 11788
rect 15708 11732 15764 12126
rect 15708 11666 15764 11676
rect 15596 11554 15652 11564
rect 15148 11340 15652 11396
rect 15036 11284 15092 11340
rect 15036 11228 15428 11284
rect 15372 10836 15428 11228
rect 15484 10836 15540 10846
rect 15372 10780 15484 10836
rect 14924 10770 14980 10780
rect 15484 10770 15540 10780
rect 14700 10658 14756 10668
rect 15596 10624 15652 11340
rect 14588 10612 14644 10622
rect 14588 10518 14644 10556
rect 14924 10612 14980 10622
rect 14140 9212 14308 9268
rect 14140 9044 14196 9054
rect 13916 8428 14084 8484
rect 13916 8260 13972 8270
rect 13692 8258 13972 8260
rect 13692 8206 13918 8258
rect 13970 8206 13972 8258
rect 13692 8204 13972 8206
rect 13916 8194 13972 8204
rect 13468 7310 13470 7362
rect 13522 7310 13524 7362
rect 13468 7298 13524 7310
rect 13580 7476 13636 7486
rect 14028 7476 14084 8428
rect 13580 6916 13636 7420
rect 13916 7420 14084 7476
rect 13580 6850 13636 6860
rect 13804 7250 13860 7262
rect 13804 7198 13806 7250
rect 13858 7198 13860 7250
rect 13804 6916 13860 7198
rect 13804 6850 13860 6860
rect 13804 6692 13860 6702
rect 13356 6690 13860 6692
rect 13356 6638 13806 6690
rect 13858 6638 13860 6690
rect 13356 6636 13860 6638
rect 13804 6626 13860 6636
rect 13132 5742 13134 5794
rect 13186 5742 13188 5794
rect 13132 5684 13188 5742
rect 12572 5294 12574 5346
rect 12626 5294 12628 5346
rect 12572 5282 12628 5294
rect 13020 5628 13188 5684
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 12908 5236 12964 5246
rect 12684 5124 12740 5134
rect 12684 5030 12740 5068
rect 12908 4452 12964 5180
rect 13020 4564 13076 5628
rect 13132 5124 13188 5134
rect 13132 5030 13188 5068
rect 13244 5012 13300 5854
rect 13916 5124 13972 7420
rect 14028 7252 14084 7262
rect 14028 7158 14084 7196
rect 14140 6132 14196 8988
rect 14252 8484 14308 9212
rect 14252 8418 14308 8428
rect 14252 7364 14308 7374
rect 14252 7270 14308 7308
rect 14364 7362 14420 7374
rect 14364 7310 14366 7362
rect 14418 7310 14420 7362
rect 14364 7028 14420 7310
rect 14476 7364 14532 10444
rect 14924 10050 14980 10556
rect 15260 10612 15316 10622
rect 15372 10612 15652 10624
rect 15260 10610 15652 10612
rect 15260 10558 15262 10610
rect 15314 10568 15652 10610
rect 15708 10612 15764 10622
rect 15314 10558 15428 10568
rect 15260 10556 15428 10558
rect 15260 10546 15316 10556
rect 15708 10518 15764 10556
rect 15484 10500 15540 10510
rect 14924 9998 14926 10050
rect 14978 9998 14980 10050
rect 14924 9986 14980 9998
rect 15036 10386 15092 10398
rect 15036 10334 15038 10386
rect 15090 10334 15092 10386
rect 14588 9828 14644 9838
rect 14588 8148 14644 9772
rect 14700 9044 14756 9054
rect 14700 8950 14756 8988
rect 15036 8708 15092 10334
rect 15372 10388 15428 10398
rect 14924 8652 15092 8708
rect 15260 10052 15316 10062
rect 15260 9154 15316 9996
rect 15260 9102 15262 9154
rect 15314 9102 15316 9154
rect 14924 8372 14980 8652
rect 15148 8372 15204 8382
rect 14924 8306 14980 8316
rect 15036 8370 15204 8372
rect 15036 8318 15150 8370
rect 15202 8318 15204 8370
rect 15036 8316 15204 8318
rect 14700 8260 14756 8270
rect 14700 8166 14756 8204
rect 14588 8082 14644 8092
rect 14924 7812 14980 7822
rect 14476 7298 14532 7308
rect 14812 7588 14868 7598
rect 14812 7362 14868 7532
rect 14924 7474 14980 7756
rect 14924 7422 14926 7474
rect 14978 7422 14980 7474
rect 14924 7410 14980 7422
rect 14812 7310 14814 7362
rect 14866 7310 14868 7362
rect 14812 7298 14868 7310
rect 14588 7252 14644 7262
rect 14588 7250 14756 7252
rect 14588 7198 14590 7250
rect 14642 7198 14756 7250
rect 14588 7196 14756 7198
rect 14588 7186 14644 7196
rect 14364 6962 14420 6972
rect 14476 7140 14532 7150
rect 14476 6914 14532 7084
rect 14476 6862 14478 6914
rect 14530 6862 14532 6914
rect 14476 6850 14532 6862
rect 14588 6804 14644 6814
rect 14588 6710 14644 6748
rect 14252 6690 14308 6702
rect 14252 6638 14254 6690
rect 14306 6638 14308 6690
rect 14252 6468 14308 6638
rect 14700 6580 14756 7196
rect 15036 7028 15092 8316
rect 15148 8306 15204 8316
rect 15260 7028 15316 9102
rect 15372 8258 15428 10332
rect 15484 9828 15540 10444
rect 15596 10052 15652 10062
rect 15596 9958 15652 9996
rect 15708 10052 15764 10062
rect 15820 10052 15876 12910
rect 15932 12180 15988 14476
rect 16268 14420 16324 18172
rect 16380 15148 16436 21084
rect 16492 20468 16548 21422
rect 16492 20402 16548 20412
rect 16492 20018 16548 20030
rect 16492 19966 16494 20018
rect 16546 19966 16548 20018
rect 16492 19908 16548 19966
rect 16492 19842 16548 19852
rect 16716 19908 16772 23492
rect 17052 23426 17108 23436
rect 16828 22930 16884 22942
rect 16828 22878 16830 22930
rect 16882 22878 16884 22930
rect 16828 22708 16884 22878
rect 16828 22642 16884 22652
rect 17052 22932 17108 22942
rect 16940 22482 16996 22494
rect 16940 22430 16942 22482
rect 16994 22430 16996 22482
rect 16940 22372 16996 22430
rect 16828 21586 16884 21598
rect 16828 21534 16830 21586
rect 16882 21534 16884 21586
rect 16828 20804 16884 21534
rect 16828 20738 16884 20748
rect 16716 19842 16772 19852
rect 16828 20018 16884 20030
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16604 19572 16660 19582
rect 16492 16772 16548 16782
rect 16492 16678 16548 16716
rect 16492 16212 16548 16222
rect 16492 15316 16548 16156
rect 16492 15250 16548 15260
rect 16604 15204 16660 19516
rect 16828 19460 16884 19966
rect 16716 19404 16828 19460
rect 16716 18450 16772 19404
rect 16828 19394 16884 19404
rect 16828 19236 16884 19246
rect 16940 19236 16996 22316
rect 17052 20692 17108 22876
rect 17164 22596 17220 25452
rect 17388 25284 17444 26572
rect 17612 26562 17668 26572
rect 17724 26292 17780 30940
rect 17836 30882 17892 31276
rect 17836 30830 17838 30882
rect 17890 30830 17892 30882
rect 17836 30818 17892 30830
rect 17948 31220 18004 31230
rect 17948 30434 18004 31164
rect 17948 30382 17950 30434
rect 18002 30382 18004 30434
rect 17836 29428 17892 29438
rect 17836 29334 17892 29372
rect 17948 27972 18004 30382
rect 17948 27906 18004 27916
rect 17948 27636 18004 27646
rect 17948 27542 18004 27580
rect 18060 27076 18116 31388
rect 18060 27010 18116 27020
rect 18172 28980 18228 44268
rect 18284 43426 18340 43438
rect 18284 43374 18286 43426
rect 18338 43374 18340 43426
rect 18284 42644 18340 43374
rect 18284 41970 18340 42588
rect 18284 41918 18286 41970
rect 18338 41918 18340 41970
rect 18284 41906 18340 41918
rect 18508 41636 18564 45836
rect 18620 44436 18676 47404
rect 18732 47394 18788 47404
rect 18844 48018 18900 48030
rect 18844 47966 18846 48018
rect 18898 47966 18900 48018
rect 18844 46676 18900 47966
rect 18956 47012 19012 49084
rect 19180 49046 19236 49084
rect 19180 48020 19236 48030
rect 19180 47926 19236 47964
rect 19068 47908 19124 47918
rect 19068 47570 19124 47852
rect 19068 47518 19070 47570
rect 19122 47518 19124 47570
rect 19068 47124 19124 47518
rect 19068 47058 19124 47068
rect 18956 46946 19012 46956
rect 19180 46900 19236 46910
rect 19292 46900 19348 50652
rect 19516 50596 19572 51772
rect 19628 51268 19684 53676
rect 19964 53666 20020 53676
rect 20076 53508 20132 53518
rect 19852 53506 20132 53508
rect 19852 53454 20078 53506
rect 20130 53454 20132 53506
rect 19852 53452 20132 53454
rect 19740 52722 19796 52734
rect 19740 52670 19742 52722
rect 19794 52670 19796 52722
rect 19740 52612 19796 52670
rect 19740 52546 19796 52556
rect 19740 51716 19796 51726
rect 19740 51380 19796 51660
rect 19852 51604 19908 53452
rect 20076 53442 20132 53452
rect 19964 53284 20020 53294
rect 19964 53058 20020 53228
rect 20076 53172 20132 53182
rect 20076 53078 20132 53116
rect 19964 53006 19966 53058
rect 20018 53006 20020 53058
rect 19964 52994 20020 53006
rect 20188 52948 20244 53788
rect 19964 52162 20020 52174
rect 19964 52110 19966 52162
rect 20018 52110 20020 52162
rect 19964 51828 20020 52110
rect 19964 51762 20020 51772
rect 19852 51548 20020 51604
rect 19852 51380 19908 51390
rect 19740 51378 19908 51380
rect 19740 51326 19854 51378
rect 19906 51326 19908 51378
rect 19740 51324 19908 51326
rect 19852 51314 19908 51324
rect 19628 51202 19684 51212
rect 19964 51044 20020 51548
rect 19964 50978 20020 50988
rect 19516 50530 19572 50540
rect 20076 50594 20132 50606
rect 20076 50542 20078 50594
rect 20130 50542 20132 50594
rect 20076 50372 20132 50542
rect 19964 50148 20020 50158
rect 19964 50036 20020 50092
rect 19852 49980 20020 50036
rect 19404 49698 19460 49710
rect 19404 49646 19406 49698
rect 19458 49646 19460 49698
rect 19404 47460 19460 49646
rect 19740 49700 19796 49710
rect 19852 49700 19908 49980
rect 20076 49812 20132 50316
rect 20188 50260 20244 52892
rect 20412 52162 20468 54012
rect 20524 53956 20580 53966
rect 20524 52948 20580 53900
rect 20860 53956 20916 53966
rect 20972 53956 21028 54796
rect 21196 54516 21252 54526
rect 21196 54402 21252 54460
rect 21196 54350 21198 54402
rect 21250 54350 21252 54402
rect 21196 54338 21252 54350
rect 21420 53956 21476 55356
rect 21532 55346 21588 55356
rect 21644 55300 21700 55580
rect 21756 55570 21812 55580
rect 21868 55858 21924 55870
rect 21868 55806 21870 55858
rect 21922 55806 21924 55858
rect 21868 55524 21924 55806
rect 22316 55858 22372 55870
rect 22316 55806 22318 55858
rect 22370 55806 22372 55858
rect 22204 55524 22260 55534
rect 22316 55524 22372 55806
rect 22540 55860 22596 56476
rect 22652 55972 22708 55982
rect 22652 55878 22708 55916
rect 23100 55972 23156 57344
rect 23548 56756 23604 57344
rect 23100 55906 23156 55916
rect 23324 56700 23604 56756
rect 23324 55970 23380 56700
rect 23996 56644 24052 57344
rect 23996 56588 24276 56644
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 23324 55918 23326 55970
rect 23378 55918 23380 55970
rect 23324 55906 23380 55918
rect 24220 55970 24276 56588
rect 24220 55918 24222 55970
rect 24274 55918 24276 55970
rect 24220 55906 24276 55918
rect 24444 56532 24500 57344
rect 24892 57092 24948 57344
rect 24892 57036 25060 57092
rect 22540 55794 22596 55804
rect 22988 55860 23044 55870
rect 24444 55860 24500 56476
rect 24892 56868 24948 56878
rect 24556 56308 24612 56318
rect 24556 56082 24612 56252
rect 24556 56030 24558 56082
rect 24610 56030 24612 56082
rect 24556 56018 24612 56030
rect 24892 55970 24948 56812
rect 24892 55918 24894 55970
rect 24946 55918 24948 55970
rect 24892 55906 24948 55918
rect 22988 55766 23044 55804
rect 24332 55804 24500 55860
rect 25004 55860 25060 57036
rect 25340 56980 25396 57344
rect 25340 56914 25396 56924
rect 25116 56420 25172 56430
rect 25116 56082 25172 56364
rect 25788 56196 25844 57344
rect 25788 56140 26068 56196
rect 25116 56030 25118 56082
rect 25170 56030 25172 56082
rect 25116 56018 25172 56030
rect 25788 55972 25844 55982
rect 25788 55878 25844 55916
rect 25340 55860 25396 55870
rect 25004 55804 25172 55860
rect 24332 55748 24388 55804
rect 24220 55692 24388 55748
rect 24464 55692 24728 55702
rect 21868 55468 22036 55524
rect 21756 55300 21812 55310
rect 21644 55244 21756 55300
rect 21756 55206 21812 55244
rect 21756 54740 21812 54750
rect 21756 54514 21812 54684
rect 21980 54516 22036 55468
rect 22204 55522 22372 55524
rect 22204 55470 22206 55522
rect 22258 55470 22372 55522
rect 22204 55468 22372 55470
rect 23212 55524 23268 55534
rect 22204 55458 22260 55468
rect 22876 55410 22932 55422
rect 22876 55358 22878 55410
rect 22930 55358 22932 55410
rect 22540 55300 22596 55310
rect 22540 55206 22596 55244
rect 22876 55076 22932 55358
rect 23100 55300 23156 55310
rect 22876 55010 22932 55020
rect 22988 55298 23156 55300
rect 22988 55246 23102 55298
rect 23154 55246 23156 55298
rect 22988 55244 23156 55246
rect 21756 54462 21758 54514
rect 21810 54462 21812 54514
rect 21756 54450 21812 54462
rect 21868 54460 22036 54516
rect 20860 53954 21028 53956
rect 20860 53902 20862 53954
rect 20914 53902 21028 53954
rect 20860 53900 21028 53902
rect 21084 53900 21476 53956
rect 21532 54290 21588 54302
rect 21532 54238 21534 54290
rect 21586 54238 21588 54290
rect 20860 53890 20916 53900
rect 20636 53732 20692 53742
rect 21084 53732 21140 53900
rect 20636 53730 21140 53732
rect 20636 53678 20638 53730
rect 20690 53678 21140 53730
rect 20636 53676 21140 53678
rect 20636 53666 20692 53676
rect 21196 53620 21252 53630
rect 21196 53526 21252 53564
rect 21532 53620 21588 54238
rect 21532 53554 21588 53564
rect 21756 53842 21812 53854
rect 21756 53790 21758 53842
rect 21810 53790 21812 53842
rect 20860 52948 20916 52958
rect 20524 52946 20916 52948
rect 20524 52894 20862 52946
rect 20914 52894 20916 52946
rect 20524 52892 20916 52894
rect 20860 52882 20916 52892
rect 21644 52948 21700 52958
rect 21644 52854 21700 52892
rect 20636 52722 20692 52734
rect 20636 52670 20638 52722
rect 20690 52670 20692 52722
rect 20636 52388 20692 52670
rect 21308 52724 21364 52734
rect 21308 52722 21700 52724
rect 21308 52670 21310 52722
rect 21362 52670 21700 52722
rect 21308 52668 21700 52670
rect 21308 52658 21364 52668
rect 20636 52322 20692 52332
rect 20860 52276 20916 52286
rect 20860 52182 20916 52220
rect 21196 52274 21252 52286
rect 21196 52222 21198 52274
rect 21250 52222 21252 52274
rect 20412 52110 20414 52162
rect 20466 52110 20468 52162
rect 20412 52098 20468 52110
rect 20524 52162 20580 52174
rect 20524 52110 20526 52162
rect 20578 52110 20580 52162
rect 20524 51940 20580 52110
rect 20524 51874 20580 51884
rect 20636 52052 20692 52062
rect 20636 51716 20692 51996
rect 20748 52052 20804 52062
rect 20748 52050 21140 52052
rect 20748 51998 20750 52050
rect 20802 51998 21140 52050
rect 20748 51996 21140 51998
rect 20748 51986 20804 51996
rect 20636 51660 20804 51716
rect 20748 51492 20804 51660
rect 20972 51492 21028 51502
rect 20748 51490 21028 51492
rect 20748 51438 20974 51490
rect 21026 51438 21028 51490
rect 20748 51436 21028 51438
rect 20972 51426 21028 51436
rect 20636 51380 20692 51390
rect 21084 51380 21140 51996
rect 21196 51492 21252 52222
rect 21532 52164 21588 52174
rect 21532 52070 21588 52108
rect 21420 52052 21476 52062
rect 21196 51436 21364 51492
rect 21084 51324 21252 51380
rect 20636 51286 20692 51324
rect 20748 51268 20804 51278
rect 20748 50706 20804 51212
rect 20748 50654 20750 50706
rect 20802 50654 20804 50706
rect 20748 50428 20804 50654
rect 20188 50194 20244 50204
rect 20412 50372 20804 50428
rect 20860 51154 20916 51166
rect 20860 51102 20862 51154
rect 20914 51102 20916 51154
rect 19796 49644 19908 49700
rect 19964 49700 20020 49710
rect 19740 49634 19796 49644
rect 19964 49606 20020 49644
rect 19628 49252 19684 49262
rect 19404 47394 19460 47404
rect 19516 48018 19572 48030
rect 19516 47966 19518 48018
rect 19570 47966 19572 48018
rect 19180 46898 19348 46900
rect 19180 46846 19182 46898
rect 19234 46846 19348 46898
rect 19180 46844 19348 46846
rect 19404 47124 19460 47134
rect 19180 46834 19236 46844
rect 18620 44370 18676 44380
rect 18732 46620 18900 46676
rect 18732 41860 18788 46620
rect 18844 46452 18900 46462
rect 18844 46450 19348 46452
rect 18844 46398 18846 46450
rect 18898 46398 19348 46450
rect 18844 46396 19348 46398
rect 18844 46386 18900 46396
rect 18956 46116 19012 46126
rect 18844 44882 18900 44894
rect 18844 44830 18846 44882
rect 18898 44830 18900 44882
rect 18844 42196 18900 44830
rect 18956 43316 19012 46060
rect 19292 46002 19348 46396
rect 19404 46228 19460 47068
rect 19404 46162 19460 46172
rect 19292 45950 19294 46002
rect 19346 45950 19348 46002
rect 19292 45938 19348 45950
rect 19404 45890 19460 45902
rect 19404 45838 19406 45890
rect 19458 45838 19460 45890
rect 19068 45668 19124 45678
rect 19068 44324 19124 45612
rect 19292 45106 19348 45118
rect 19292 45054 19294 45106
rect 19346 45054 19348 45106
rect 19292 44548 19348 45054
rect 19292 44482 19348 44492
rect 19404 44546 19460 45838
rect 19404 44494 19406 44546
rect 19458 44494 19460 44546
rect 19404 44482 19460 44494
rect 19068 44268 19460 44324
rect 19068 44100 19124 44110
rect 19068 43538 19124 44044
rect 19068 43486 19070 43538
rect 19122 43486 19124 43538
rect 19068 43474 19124 43486
rect 18956 43260 19124 43316
rect 18844 42140 19012 42196
rect 18732 41794 18788 41804
rect 18956 41748 19012 42140
rect 19068 41972 19124 43260
rect 19068 41878 19124 41916
rect 19292 42530 19348 42542
rect 19292 42478 19294 42530
rect 19346 42478 19348 42530
rect 18844 41692 19012 41748
rect 18508 41580 18788 41636
rect 18508 41300 18564 41310
rect 18508 41186 18564 41244
rect 18508 41134 18510 41186
rect 18562 41134 18564 41186
rect 18396 40516 18452 40526
rect 18508 40516 18564 41134
rect 18396 40514 18564 40516
rect 18396 40462 18398 40514
rect 18450 40462 18564 40514
rect 18396 40460 18564 40462
rect 18396 40450 18452 40460
rect 18508 39618 18564 40460
rect 18508 39566 18510 39618
rect 18562 39566 18564 39618
rect 18508 39554 18564 39566
rect 18620 40964 18676 40974
rect 18284 38834 18340 38846
rect 18284 38782 18286 38834
rect 18338 38782 18340 38834
rect 18284 37716 18340 38782
rect 18284 37650 18340 37660
rect 18508 38612 18564 38622
rect 18396 37604 18452 37614
rect 18284 37266 18340 37278
rect 18284 37214 18286 37266
rect 18338 37214 18340 37266
rect 18284 37044 18340 37214
rect 18284 36978 18340 36988
rect 18284 31780 18340 31790
rect 18284 31686 18340 31724
rect 18396 30996 18452 37548
rect 18508 37156 18564 38556
rect 18508 37090 18564 37100
rect 18508 36258 18564 36270
rect 18508 36206 18510 36258
rect 18562 36206 18564 36258
rect 18508 36148 18564 36206
rect 18508 36082 18564 36092
rect 18620 35364 18676 40908
rect 18732 38164 18788 41580
rect 18844 41076 18900 41692
rect 18844 40740 18900 41020
rect 18956 41298 19012 41310
rect 18956 41246 18958 41298
rect 19010 41246 19012 41298
rect 18956 40852 19012 41246
rect 19292 41300 19348 42478
rect 19292 41234 19348 41244
rect 19012 40796 19348 40852
rect 18956 40786 19012 40796
rect 18844 40674 18900 40684
rect 19180 40404 19236 40414
rect 18844 40292 18900 40302
rect 18844 40198 18900 40236
rect 19068 40068 19124 40078
rect 18844 39732 18900 39742
rect 18900 39676 19012 39732
rect 18844 39638 18900 39676
rect 18844 38724 18900 38762
rect 18844 38658 18900 38668
rect 18844 38164 18900 38174
rect 18732 38162 18900 38164
rect 18732 38110 18846 38162
rect 18898 38110 18900 38162
rect 18732 38108 18900 38110
rect 18732 36708 18788 38108
rect 18844 38098 18900 38108
rect 18844 37156 18900 37166
rect 18956 37156 19012 39676
rect 18844 37154 19012 37156
rect 18844 37102 18846 37154
rect 18898 37102 19012 37154
rect 18844 37100 19012 37102
rect 18844 36932 18900 37100
rect 18844 36866 18900 36876
rect 18732 36652 18900 36708
rect 18620 35298 18676 35308
rect 18508 35252 18564 35262
rect 18508 34690 18564 35196
rect 18620 35140 18676 35150
rect 18844 35140 18900 36652
rect 18956 36596 19012 36606
rect 19068 36596 19124 40012
rect 19180 37380 19236 40348
rect 19292 38612 19348 40796
rect 19292 38546 19348 38556
rect 19180 37314 19236 37324
rect 19292 38050 19348 38062
rect 19292 37998 19294 38050
rect 19346 37998 19348 38050
rect 18956 36594 19124 36596
rect 18956 36542 18958 36594
rect 19010 36542 19124 36594
rect 18956 36540 19124 36542
rect 18956 36530 19012 36540
rect 19068 36036 19124 36540
rect 19292 36484 19348 37998
rect 19404 37156 19460 44268
rect 19516 41524 19572 47966
rect 19628 44100 19684 49196
rect 20076 49028 20132 49756
rect 19964 48972 20132 49028
rect 20188 49252 20244 49262
rect 19740 48804 19796 48814
rect 19740 47236 19796 48748
rect 19964 48468 20020 48972
rect 19964 48402 20020 48412
rect 19852 48020 19908 48030
rect 20076 48020 20132 48030
rect 19852 47926 19908 47964
rect 19964 48018 20132 48020
rect 19964 47966 20078 48018
rect 20130 47966 20132 48018
rect 19964 47964 20132 47966
rect 19740 47170 19796 47180
rect 19852 47572 19908 47582
rect 19852 46674 19908 47516
rect 19964 47460 20020 47964
rect 20076 47954 20132 47964
rect 19964 47394 20020 47404
rect 20076 47236 20132 47246
rect 20076 46900 20132 47180
rect 20076 46834 20132 46844
rect 19852 46622 19854 46674
rect 19906 46622 19908 46674
rect 19852 46610 19908 46622
rect 19964 46562 20020 46574
rect 19964 46510 19966 46562
rect 20018 46510 20020 46562
rect 19964 46116 20020 46510
rect 19964 46050 20020 46060
rect 20076 46452 20132 46462
rect 19628 44034 19684 44044
rect 19740 45892 19796 45902
rect 19516 41458 19572 41468
rect 19628 43540 19684 43550
rect 19628 42644 19684 43484
rect 19740 43092 19796 45836
rect 19964 45892 20020 45902
rect 20076 45892 20132 46396
rect 19964 45890 20132 45892
rect 19964 45838 19966 45890
rect 20018 45838 20132 45890
rect 19964 45836 20132 45838
rect 19964 45826 20020 45836
rect 19964 44772 20020 44782
rect 19852 43540 19908 43550
rect 19852 43446 19908 43484
rect 19964 43428 20020 44716
rect 20188 44548 20244 49196
rect 20300 48804 20356 48814
rect 20300 48710 20356 48748
rect 20300 47572 20356 47582
rect 20300 47478 20356 47516
rect 20300 46788 20356 46798
rect 20300 46114 20356 46732
rect 20300 46062 20302 46114
rect 20354 46062 20356 46114
rect 20300 46050 20356 46062
rect 20188 44492 20356 44548
rect 20076 44212 20132 44222
rect 20076 44118 20132 44156
rect 19964 43204 20020 43372
rect 19740 43026 19796 43036
rect 19852 43148 20020 43204
rect 19740 42868 19796 42878
rect 19852 42868 19908 43148
rect 20188 43092 20244 43102
rect 19740 42866 19908 42868
rect 19740 42814 19742 42866
rect 19794 42814 19908 42866
rect 19740 42812 19908 42814
rect 19964 43036 20188 43092
rect 19740 42802 19796 42812
rect 19516 41076 19572 41086
rect 19516 40404 19572 41020
rect 19516 40338 19572 40348
rect 19628 38668 19684 42588
rect 19740 42308 19796 42318
rect 19740 40292 19796 42252
rect 19964 41972 20020 43036
rect 20188 43026 20244 43036
rect 20076 42756 20132 42766
rect 20076 42754 20244 42756
rect 20076 42702 20078 42754
rect 20130 42702 20244 42754
rect 20076 42700 20244 42702
rect 20076 42690 20132 42700
rect 19740 40226 19796 40236
rect 19852 41970 20020 41972
rect 19852 41918 19966 41970
rect 20018 41918 20020 41970
rect 19852 41916 20020 41918
rect 19852 40068 19908 41916
rect 19964 41906 20020 41916
rect 20188 41972 20244 42700
rect 20188 41410 20244 41916
rect 20188 41358 20190 41410
rect 20242 41358 20244 41410
rect 20188 41346 20244 41358
rect 19964 40404 20020 40414
rect 19964 40310 20020 40348
rect 19852 40002 19908 40012
rect 20076 40068 20132 40078
rect 20076 39842 20132 40012
rect 20076 39790 20078 39842
rect 20130 39790 20132 39842
rect 20076 39778 20132 39790
rect 20300 38668 20356 44492
rect 20412 43428 20468 50372
rect 20524 50260 20580 50270
rect 20524 48020 20580 50204
rect 20748 48916 20804 48926
rect 20748 48822 20804 48860
rect 20636 48692 20692 48702
rect 20636 48242 20692 48636
rect 20748 48468 20804 48478
rect 20860 48468 20916 51102
rect 21084 51154 21140 51166
rect 21084 51102 21086 51154
rect 21138 51102 21140 51154
rect 21084 51044 21140 51102
rect 21196 51154 21252 51324
rect 21196 51102 21198 51154
rect 21250 51102 21252 51154
rect 21196 51090 21252 51102
rect 21084 50978 21140 50988
rect 21084 50596 21140 50606
rect 21084 49924 21140 50540
rect 21084 49830 21140 49868
rect 21196 50594 21252 50606
rect 21196 50542 21198 50594
rect 21250 50542 21252 50594
rect 21084 49028 21140 49038
rect 21196 49028 21252 50542
rect 21084 49026 21252 49028
rect 21084 48974 21086 49026
rect 21138 48974 21252 49026
rect 21084 48972 21252 48974
rect 20748 48466 20916 48468
rect 20748 48414 20750 48466
rect 20802 48414 20916 48466
rect 20748 48412 20916 48414
rect 20972 48916 21028 48926
rect 20748 48402 20804 48412
rect 20636 48190 20638 48242
rect 20690 48190 20692 48242
rect 20636 48178 20692 48190
rect 20748 48020 20804 48030
rect 20524 48018 20804 48020
rect 20524 47966 20750 48018
rect 20802 47966 20804 48018
rect 20524 47964 20804 47966
rect 20748 47954 20804 47964
rect 20524 47348 20580 47358
rect 20524 47068 20580 47292
rect 20748 47346 20804 47358
rect 20748 47294 20750 47346
rect 20802 47294 20804 47346
rect 20748 47236 20804 47294
rect 20748 47170 20804 47180
rect 20524 47012 20692 47068
rect 20636 46004 20692 47012
rect 20748 46900 20804 46910
rect 20748 46806 20804 46844
rect 20860 46676 20916 46686
rect 20860 46582 20916 46620
rect 20748 46564 20804 46574
rect 20748 46470 20804 46508
rect 20748 46004 20804 46014
rect 20636 46002 20804 46004
rect 20636 45950 20750 46002
rect 20802 45950 20804 46002
rect 20636 45948 20804 45950
rect 20524 45780 20580 45790
rect 20524 44434 20580 45724
rect 20524 44382 20526 44434
rect 20578 44382 20580 44434
rect 20524 44324 20580 44382
rect 20524 44258 20580 44268
rect 20636 44884 20692 44894
rect 20412 43362 20468 43372
rect 20636 43764 20692 44828
rect 20524 42754 20580 42766
rect 20524 42702 20526 42754
rect 20578 42702 20580 42754
rect 20524 42644 20580 42702
rect 20524 42578 20580 42588
rect 20636 42420 20692 43708
rect 20748 43540 20804 45948
rect 20748 43474 20804 43484
rect 20972 43092 21028 48860
rect 21084 48804 21140 48972
rect 21084 47458 21140 48748
rect 21084 47406 21086 47458
rect 21138 47406 21140 47458
rect 21084 45890 21140 47406
rect 21308 46788 21364 51436
rect 21420 49476 21476 51996
rect 21532 51828 21588 51838
rect 21532 51044 21588 51772
rect 21532 50594 21588 50988
rect 21532 50542 21534 50594
rect 21586 50542 21588 50594
rect 21532 50530 21588 50542
rect 21532 49812 21588 49822
rect 21532 49698 21588 49756
rect 21532 49646 21534 49698
rect 21586 49646 21588 49698
rect 21532 49634 21588 49646
rect 21420 49410 21476 49420
rect 21644 49364 21700 52668
rect 21756 51604 21812 53790
rect 21868 52500 21924 54460
rect 22092 54402 22148 54414
rect 22092 54350 22094 54402
rect 22146 54350 22148 54402
rect 21980 54290 22036 54302
rect 21980 54238 21982 54290
rect 22034 54238 22036 54290
rect 21980 53844 22036 54238
rect 22092 54068 22148 54350
rect 22428 54404 22484 54414
rect 22428 54310 22484 54348
rect 22092 54002 22148 54012
rect 22764 54290 22820 54302
rect 22764 54238 22766 54290
rect 22818 54238 22820 54290
rect 21980 53778 22036 53788
rect 22652 53842 22708 53854
rect 22652 53790 22654 53842
rect 22706 53790 22708 53842
rect 22092 53732 22148 53742
rect 22092 53638 22148 53676
rect 22428 53618 22484 53630
rect 22428 53566 22430 53618
rect 22482 53566 22484 53618
rect 22092 53508 22148 53518
rect 21980 52836 22036 52846
rect 21980 52742 22036 52780
rect 21868 52444 22036 52500
rect 21756 51538 21812 51548
rect 21868 51492 21924 51502
rect 21868 51398 21924 51436
rect 21756 51380 21812 51390
rect 21756 50932 21812 51324
rect 21756 50866 21812 50876
rect 21756 50708 21812 50718
rect 21756 50614 21812 50652
rect 21644 49298 21700 49308
rect 21756 49138 21812 49150
rect 21756 49086 21758 49138
rect 21810 49086 21812 49138
rect 21532 49028 21588 49038
rect 21420 49026 21588 49028
rect 21420 48974 21534 49026
rect 21586 48974 21588 49026
rect 21420 48972 21588 48974
rect 21756 49028 21812 49086
rect 21868 49028 21924 49038
rect 21756 48972 21868 49028
rect 21420 47124 21476 48972
rect 21532 48962 21588 48972
rect 21868 48962 21924 48972
rect 21980 48916 22036 52444
rect 22092 52388 22148 53452
rect 22428 53508 22484 53566
rect 22428 53442 22484 53452
rect 22652 52948 22708 53790
rect 22764 53508 22820 54238
rect 22988 53956 23044 55244
rect 23100 55234 23156 55244
rect 23100 54292 23156 54302
rect 23100 54198 23156 54236
rect 22764 53442 22820 53452
rect 22876 53900 23044 53956
rect 23100 53956 23156 53966
rect 22652 52882 22708 52892
rect 22428 52836 22484 52846
rect 22316 52724 22372 52734
rect 22316 52630 22372 52668
rect 22092 52322 22148 52332
rect 22316 52164 22372 52174
rect 22428 52164 22484 52780
rect 22764 52388 22820 52398
rect 22764 52294 22820 52332
rect 22316 52162 22484 52164
rect 22316 52110 22318 52162
rect 22370 52110 22484 52162
rect 22316 52108 22484 52110
rect 22316 51492 22372 52108
rect 22316 51426 22372 51436
rect 22316 51154 22372 51166
rect 22316 51102 22318 51154
rect 22370 51102 22372 51154
rect 22316 50820 22372 51102
rect 22316 50754 22372 50764
rect 22764 51156 22820 51166
rect 22764 50932 22820 51100
rect 22428 50596 22484 50606
rect 22428 50594 22708 50596
rect 22428 50542 22430 50594
rect 22482 50542 22708 50594
rect 22428 50540 22708 50542
rect 22428 50530 22484 50540
rect 22652 50036 22708 50540
rect 22764 50594 22820 50876
rect 22764 50542 22766 50594
rect 22818 50542 22820 50594
rect 22764 50530 22820 50542
rect 21980 48850 22036 48860
rect 22428 50034 22708 50036
rect 22428 49982 22654 50034
rect 22706 49982 22708 50034
rect 22428 49980 22708 49982
rect 22428 49026 22484 49980
rect 22652 49970 22708 49980
rect 22428 48974 22430 49026
rect 22482 48974 22484 49026
rect 21980 48468 22036 48478
rect 21644 48244 21700 48254
rect 21420 47058 21476 47068
rect 21532 48242 21700 48244
rect 21532 48190 21646 48242
rect 21698 48190 21700 48242
rect 21532 48188 21700 48190
rect 21532 47068 21588 48188
rect 21644 48178 21700 48188
rect 21756 47572 21812 47582
rect 21756 47570 21924 47572
rect 21756 47518 21758 47570
rect 21810 47518 21924 47570
rect 21756 47516 21924 47518
rect 21756 47506 21812 47516
rect 21644 47458 21700 47470
rect 21644 47406 21646 47458
rect 21698 47406 21700 47458
rect 21644 47348 21700 47406
rect 21868 47460 21924 47516
rect 21868 47394 21924 47404
rect 21644 47282 21700 47292
rect 21980 47124 22036 48412
rect 22092 48132 22148 48142
rect 22092 48038 22148 48076
rect 22428 47458 22484 48974
rect 22764 49140 22820 49150
rect 22764 49026 22820 49084
rect 22764 48974 22766 49026
rect 22818 48974 22820 49026
rect 22652 48804 22708 48814
rect 22428 47406 22430 47458
rect 22482 47406 22484 47458
rect 21756 47068 22036 47124
rect 22316 47236 22372 47246
rect 21532 47012 21700 47068
rect 21084 45838 21086 45890
rect 21138 45838 21140 45890
rect 21084 45826 21140 45838
rect 21196 46732 21364 46788
rect 20860 43036 21028 43092
rect 20636 42354 20692 42364
rect 20748 42866 20804 42878
rect 20748 42814 20750 42866
rect 20802 42814 20804 42866
rect 20636 41300 20692 41310
rect 20748 41300 20804 42814
rect 20860 42756 20916 43036
rect 21196 42980 21252 46732
rect 21644 46676 21700 47012
rect 20860 42690 20916 42700
rect 20972 42924 21252 42980
rect 21308 46674 21700 46676
rect 21308 46622 21646 46674
rect 21698 46622 21700 46674
rect 21308 46620 21700 46622
rect 20636 41298 20804 41300
rect 20636 41246 20638 41298
rect 20690 41246 20804 41298
rect 20636 41244 20804 41246
rect 20860 41972 20916 41982
rect 20636 41234 20692 41244
rect 20860 39618 20916 41916
rect 20972 41636 21028 42924
rect 20972 41570 21028 41580
rect 20972 41186 21028 41198
rect 20972 41134 20974 41186
rect 21026 41134 21028 41186
rect 20972 40068 21028 41134
rect 20972 40002 21028 40012
rect 21084 40292 21140 40302
rect 20860 39566 20862 39618
rect 20914 39566 20916 39618
rect 20860 39554 20916 39566
rect 20524 39506 20580 39518
rect 20524 39454 20526 39506
rect 20578 39454 20580 39506
rect 20524 38668 20580 39454
rect 19628 38612 19796 38668
rect 19628 38050 19684 38062
rect 19628 37998 19630 38050
rect 19682 37998 19684 38050
rect 19628 37940 19684 37998
rect 19628 37874 19684 37884
rect 19404 37090 19460 37100
rect 19404 36484 19460 36494
rect 19292 36482 19460 36484
rect 19292 36430 19406 36482
rect 19458 36430 19460 36482
rect 19292 36428 19460 36430
rect 19404 36148 19460 36428
rect 19740 36484 19796 38612
rect 19964 38612 20020 38622
rect 20300 38612 20468 38668
rect 20524 38612 20692 38668
rect 19964 38610 20244 38612
rect 19964 38558 19966 38610
rect 20018 38558 20244 38610
rect 19964 38556 20244 38558
rect 19964 38546 20020 38556
rect 19740 36390 19796 36428
rect 19852 38162 19908 38174
rect 19852 38110 19854 38162
rect 19906 38110 19908 38162
rect 19404 36082 19460 36092
rect 19068 35980 19348 36036
rect 18676 35084 18900 35140
rect 19180 35140 19236 35150
rect 18620 35074 18676 35084
rect 19068 35028 19124 35038
rect 18508 34638 18510 34690
rect 18562 34638 18564 34690
rect 18508 34020 18564 34638
rect 18844 35026 19124 35028
rect 18844 34974 19070 35026
rect 19122 34974 19124 35026
rect 18844 34972 19124 34974
rect 18620 34132 18676 34142
rect 18620 34038 18676 34076
rect 18844 34132 18900 34972
rect 19068 34962 19124 34972
rect 19180 35026 19236 35084
rect 19180 34974 19182 35026
rect 19234 34974 19236 35026
rect 19180 34962 19236 34974
rect 19068 34692 19124 34702
rect 19068 34598 19124 34636
rect 19068 34468 19124 34478
rect 19068 34354 19124 34412
rect 19068 34302 19070 34354
rect 19122 34302 19124 34354
rect 19068 34290 19124 34302
rect 19292 34244 19348 35980
rect 19852 35924 19908 38110
rect 20188 38164 20244 38556
rect 20300 38164 20356 38174
rect 20188 38162 20356 38164
rect 20188 38110 20302 38162
rect 20354 38110 20356 38162
rect 20188 38108 20356 38110
rect 19964 38052 20020 38062
rect 19964 37490 20020 37996
rect 19964 37438 19966 37490
rect 20018 37438 20020 37490
rect 19964 37426 20020 37438
rect 19404 35868 19908 35924
rect 19964 36594 20020 36606
rect 19964 36542 19966 36594
rect 20018 36542 20020 36594
rect 19404 35140 19460 35868
rect 19964 35700 20020 36542
rect 20300 36596 20356 38108
rect 20412 36820 20468 38612
rect 20412 36764 20580 36820
rect 20412 36596 20468 36606
rect 20300 36594 20468 36596
rect 20300 36542 20414 36594
rect 20466 36542 20468 36594
rect 20300 36540 20468 36542
rect 20076 35700 20132 35710
rect 19964 35698 20132 35700
rect 19964 35646 20078 35698
rect 20130 35646 20132 35698
rect 19964 35644 20132 35646
rect 20076 35634 20132 35644
rect 19404 35074 19460 35084
rect 19516 35586 19572 35598
rect 19516 35534 19518 35586
rect 19570 35534 19572 35586
rect 19516 34468 19572 35534
rect 19740 35586 19796 35598
rect 19740 35534 19742 35586
rect 19794 35534 19796 35586
rect 19740 35364 19796 35534
rect 19740 35298 19796 35308
rect 19852 35474 19908 35486
rect 19852 35422 19854 35474
rect 19906 35422 19908 35474
rect 19628 35140 19684 35150
rect 19852 35140 19908 35422
rect 19628 35138 19908 35140
rect 19628 35086 19630 35138
rect 19682 35086 19908 35138
rect 19628 35084 19908 35086
rect 19628 35074 19684 35084
rect 20412 35028 20468 36540
rect 20412 34962 20468 34972
rect 19740 34916 19796 34926
rect 19628 34914 19796 34916
rect 19628 34862 19742 34914
rect 19794 34862 19796 34914
rect 19628 34860 19796 34862
rect 19628 34692 19684 34860
rect 19740 34850 19796 34860
rect 19964 34914 20020 34926
rect 19964 34862 19966 34914
rect 20018 34862 20020 34914
rect 19628 34626 19684 34636
rect 19852 34804 19908 34814
rect 19852 34580 19908 34748
rect 19516 34402 19572 34412
rect 19740 34524 19908 34580
rect 19292 34188 19572 34244
rect 18844 34066 18900 34076
rect 18508 33926 18564 33964
rect 18956 34020 19012 34030
rect 19404 34020 19460 34030
rect 18956 34018 19460 34020
rect 18956 33966 18958 34018
rect 19010 33966 19406 34018
rect 19458 33966 19460 34018
rect 18956 33964 19460 33966
rect 18508 33572 18564 33582
rect 18956 33572 19012 33964
rect 19404 33954 19460 33964
rect 19516 33684 19572 34188
rect 19628 34132 19684 34142
rect 19628 34038 19684 34076
rect 19516 33628 19684 33684
rect 18508 33570 19012 33572
rect 18508 33518 18510 33570
rect 18562 33518 19012 33570
rect 18508 33516 19012 33518
rect 18508 33506 18564 33516
rect 19516 33460 19572 33470
rect 18620 32788 18676 32798
rect 18508 32564 18564 32574
rect 18508 32470 18564 32508
rect 18396 30930 18452 30940
rect 18508 30994 18564 31006
rect 18508 30942 18510 30994
rect 18562 30942 18564 30994
rect 18508 30436 18564 30942
rect 18508 29426 18564 30380
rect 18508 29374 18510 29426
rect 18562 29374 18564 29426
rect 18508 29362 18564 29374
rect 18172 26292 18228 28924
rect 18620 28980 18676 32732
rect 18844 32676 18900 32686
rect 18620 28914 18676 28924
rect 18732 31668 18788 31678
rect 18508 28868 18564 28878
rect 18508 28644 18564 28812
rect 18732 28756 18788 31612
rect 18844 31220 18900 32620
rect 19516 32564 19572 33404
rect 19404 31780 19460 31790
rect 19516 31780 19572 32508
rect 19404 31778 19572 31780
rect 19404 31726 19406 31778
rect 19458 31726 19572 31778
rect 19404 31724 19572 31726
rect 19404 31714 19460 31724
rect 18844 31154 18900 31164
rect 19180 31556 19236 31566
rect 18844 30996 18900 31006
rect 18844 30902 18900 30940
rect 18508 28578 18564 28588
rect 18620 28700 18788 28756
rect 18844 30548 18900 30558
rect 18508 27860 18564 27870
rect 18396 27412 18452 27422
rect 18284 27076 18340 27086
rect 18284 26404 18340 27020
rect 18396 26964 18452 27356
rect 18396 26898 18452 26908
rect 18396 26404 18452 26414
rect 18284 26402 18452 26404
rect 18284 26350 18398 26402
rect 18450 26350 18452 26402
rect 18284 26348 18452 26350
rect 17724 26236 17892 26292
rect 18172 26236 18340 26292
rect 17612 26180 17668 26190
rect 17612 26086 17668 26124
rect 17500 26068 17556 26078
rect 17500 25974 17556 26012
rect 17724 26066 17780 26078
rect 17724 26014 17726 26066
rect 17778 26014 17780 26066
rect 17724 25844 17780 26014
rect 17500 25788 17780 25844
rect 17500 25508 17556 25788
rect 17724 25620 17780 25630
rect 17724 25526 17780 25564
rect 17500 25442 17556 25452
rect 17612 25506 17668 25518
rect 17612 25454 17614 25506
rect 17666 25454 17668 25506
rect 17612 25396 17668 25454
rect 17836 25396 17892 26236
rect 18172 25506 18228 25518
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 17612 25340 18116 25396
rect 17388 25228 18004 25284
rect 17388 24722 17444 24734
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17276 23716 17332 23726
rect 17276 23154 17332 23660
rect 17276 23102 17278 23154
rect 17330 23102 17332 23154
rect 17276 23090 17332 23102
rect 17388 22932 17444 24670
rect 17612 24500 17668 24510
rect 17612 24498 17892 24500
rect 17612 24446 17614 24498
rect 17666 24446 17892 24498
rect 17612 24444 17892 24446
rect 17612 24434 17668 24444
rect 17724 24052 17780 24062
rect 17612 24050 17780 24052
rect 17612 23998 17726 24050
rect 17778 23998 17780 24050
rect 17612 23996 17780 23998
rect 17500 23940 17556 23950
rect 17500 23846 17556 23884
rect 17388 22876 17556 22932
rect 17388 22708 17444 22718
rect 17276 22596 17332 22606
rect 17164 22594 17332 22596
rect 17164 22542 17278 22594
rect 17330 22542 17332 22594
rect 17164 22540 17332 22542
rect 17276 22530 17332 22540
rect 17388 22594 17444 22652
rect 17388 22542 17390 22594
rect 17442 22542 17444 22594
rect 17388 22530 17444 22542
rect 17164 22370 17220 22382
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 17164 21812 17220 22318
rect 17164 20914 17220 21756
rect 17500 21812 17556 22876
rect 17612 22708 17668 23996
rect 17724 23986 17780 23996
rect 17836 23380 17892 24444
rect 17836 23314 17892 23324
rect 17948 23044 18004 25228
rect 18060 23492 18116 25340
rect 18172 24722 18228 25454
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 18172 23938 18228 24670
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18172 23716 18228 23886
rect 18172 23650 18228 23660
rect 18060 23426 18116 23436
rect 18060 23156 18116 23166
rect 18060 23062 18116 23100
rect 17612 22642 17668 22652
rect 17836 22988 18004 23044
rect 17500 21746 17556 21756
rect 17276 21588 17332 21598
rect 17276 21586 17556 21588
rect 17276 21534 17278 21586
rect 17330 21534 17556 21586
rect 17276 21532 17556 21534
rect 17276 21522 17332 21532
rect 17164 20862 17166 20914
rect 17218 20862 17220 20914
rect 17164 20850 17220 20862
rect 17388 21364 17444 21374
rect 17276 20692 17332 20702
rect 17052 20690 17332 20692
rect 17052 20638 17278 20690
rect 17330 20638 17332 20690
rect 17052 20636 17332 20638
rect 17276 20626 17332 20636
rect 17276 20468 17332 20478
rect 17164 20132 17220 20142
rect 17164 19460 17220 20076
rect 17164 19394 17220 19404
rect 16828 19234 16996 19236
rect 16828 19182 16830 19234
rect 16882 19182 16996 19234
rect 16828 19180 16996 19182
rect 16828 19170 16884 19180
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18386 16772 18398
rect 17164 18452 17220 18462
rect 17164 18358 17220 18396
rect 16828 17948 17108 18004
rect 16716 17666 16772 17678
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 16884 16772 17614
rect 16828 17220 16884 17948
rect 16940 17780 16996 17790
rect 16940 17686 16996 17724
rect 17052 17778 17108 17948
rect 17052 17726 17054 17778
rect 17106 17726 17108 17778
rect 17052 17714 17108 17726
rect 17164 17778 17220 17790
rect 17164 17726 17166 17778
rect 17218 17726 17220 17778
rect 16828 17154 16884 17164
rect 16940 17554 16996 17566
rect 16940 17502 16942 17554
rect 16994 17502 16996 17554
rect 16716 16818 16772 16828
rect 16940 16100 16996 17502
rect 17164 17108 17220 17726
rect 17164 17042 17220 17052
rect 16940 16034 16996 16044
rect 17052 16772 17108 16782
rect 16380 15092 16548 15148
rect 16604 15138 16660 15148
rect 16716 15988 16772 15998
rect 16268 14364 16436 14420
rect 16044 14308 16100 14318
rect 16380 14308 16436 14364
rect 16044 14306 16324 14308
rect 16044 14254 16046 14306
rect 16098 14254 16324 14306
rect 16044 14252 16324 14254
rect 16044 14242 16100 14252
rect 16268 13746 16324 14252
rect 16380 14242 16436 14252
rect 16268 13694 16270 13746
rect 16322 13694 16324 13746
rect 16268 13682 16324 13694
rect 15932 12114 15988 12124
rect 16044 13074 16100 13086
rect 16044 13022 16046 13074
rect 16098 13022 16100 13074
rect 16044 11396 16100 13022
rect 16156 12964 16212 12974
rect 16156 12962 16436 12964
rect 16156 12910 16158 12962
rect 16210 12910 16436 12962
rect 16156 12908 16436 12910
rect 16156 12898 16212 12908
rect 16156 12178 16212 12190
rect 16156 12126 16158 12178
rect 16210 12126 16212 12178
rect 16156 11844 16212 12126
rect 16380 12066 16436 12908
rect 16492 12740 16548 15092
rect 16716 13748 16772 15932
rect 17052 15540 17108 16716
rect 16828 15202 16884 15214
rect 16828 15150 16830 15202
rect 16882 15150 16884 15202
rect 16828 13972 16884 15150
rect 17052 14530 17108 15484
rect 17164 15316 17220 15326
rect 17164 15222 17220 15260
rect 17052 14478 17054 14530
rect 17106 14478 17108 14530
rect 17052 14466 17108 14478
rect 16828 13906 16884 13916
rect 16828 13748 16884 13758
rect 16716 13746 16884 13748
rect 16716 13694 16830 13746
rect 16882 13694 16884 13746
rect 16716 13692 16884 13694
rect 16828 13682 16884 13692
rect 17276 12964 17332 20412
rect 17388 16324 17444 21308
rect 17500 19906 17556 21532
rect 17612 21364 17668 21374
rect 17612 21270 17668 21308
rect 17836 20998 17892 22988
rect 18060 22708 18116 22718
rect 17948 22260 18004 22270
rect 17948 22166 18004 22204
rect 18060 21476 18116 22652
rect 18060 21410 18116 21420
rect 17724 20942 17892 20998
rect 17948 21364 18004 21374
rect 17612 20132 17668 20142
rect 17612 20018 17668 20076
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17612 19954 17668 19966
rect 17500 19854 17502 19906
rect 17554 19854 17556 19906
rect 17500 19842 17556 19854
rect 17724 17668 17780 20942
rect 17836 20804 17892 20814
rect 17836 20710 17892 20748
rect 17948 20580 18004 21308
rect 18172 20916 18228 20926
rect 18172 20822 18228 20860
rect 17948 20514 18004 20524
rect 18060 20020 18116 20030
rect 18060 19926 18116 19964
rect 18060 19572 18116 19582
rect 18060 19348 18116 19516
rect 17948 19346 18116 19348
rect 17948 19294 18062 19346
rect 18114 19294 18116 19346
rect 17948 19292 18116 19294
rect 17948 18228 18004 19292
rect 18060 19282 18116 19292
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 17948 18162 18004 18172
rect 17388 16258 17444 16268
rect 17612 17612 17780 17668
rect 18060 17666 18116 17678
rect 18060 17614 18062 17666
rect 18114 17614 18116 17666
rect 17500 14980 17556 14990
rect 17500 14754 17556 14924
rect 17500 14702 17502 14754
rect 17554 14702 17556 14754
rect 17500 14690 17556 14702
rect 17500 14196 17556 14206
rect 17164 12962 17332 12964
rect 17164 12910 17278 12962
rect 17330 12910 17332 12962
rect 17164 12908 17332 12910
rect 16492 12674 16548 12684
rect 16716 12850 16772 12862
rect 16716 12798 16718 12850
rect 16770 12798 16772 12850
rect 16380 12014 16382 12066
rect 16434 12014 16436 12066
rect 16380 12002 16436 12014
rect 16716 11788 16772 12798
rect 16828 12738 16884 12750
rect 16828 12686 16830 12738
rect 16882 12686 16884 12738
rect 16828 12292 16884 12686
rect 16828 12236 17108 12292
rect 16156 11778 16212 11788
rect 16492 11732 16772 11788
rect 16828 12066 16884 12078
rect 16828 12014 16830 12066
rect 16882 12014 16884 12066
rect 16380 11396 16436 11406
rect 16044 11340 16212 11396
rect 16044 11170 16100 11182
rect 16044 11118 16046 11170
rect 16098 11118 16100 11170
rect 16044 10948 16100 11118
rect 16156 11172 16212 11340
rect 16156 11106 16212 11116
rect 15708 10050 15876 10052
rect 15708 9998 15710 10050
rect 15762 9998 15876 10050
rect 15708 9996 15876 9998
rect 15932 10892 16100 10948
rect 16268 11060 16324 11070
rect 15932 10052 15988 10892
rect 16044 10498 16100 10510
rect 16044 10446 16046 10498
rect 16098 10446 16100 10498
rect 16044 10276 16100 10446
rect 16268 10276 16324 11004
rect 16380 10722 16436 11340
rect 16380 10670 16382 10722
rect 16434 10670 16436 10722
rect 16380 10658 16436 10670
rect 16044 10220 16324 10276
rect 16044 10052 16100 10062
rect 15932 9996 16044 10052
rect 15708 9986 15764 9996
rect 16044 9986 16100 9996
rect 16492 10052 16548 11732
rect 16604 11172 16660 11182
rect 16604 10276 16660 11116
rect 16716 10836 16772 10846
rect 16716 10610 16772 10780
rect 16716 10558 16718 10610
rect 16770 10558 16772 10610
rect 16716 10500 16772 10558
rect 16828 10612 16884 12014
rect 16828 10546 16884 10556
rect 16940 11172 16996 11182
rect 16716 10434 16772 10444
rect 16940 10276 16996 11116
rect 17052 10388 17108 12236
rect 17164 11282 17220 12908
rect 17276 12898 17332 12908
rect 17388 13972 17444 13982
rect 17388 11396 17444 13916
rect 17500 12964 17556 14140
rect 17500 12178 17556 12908
rect 17500 12126 17502 12178
rect 17554 12126 17556 12178
rect 17500 12114 17556 12126
rect 17612 11732 17668 17612
rect 17724 17108 17780 17118
rect 17724 17014 17780 17052
rect 17836 16660 17892 16670
rect 17836 16100 17892 16604
rect 17724 15314 17780 15326
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 14532 17780 15262
rect 17836 15202 17892 16044
rect 18060 15540 18116 17614
rect 18172 15988 18228 15998
rect 18172 15894 18228 15932
rect 18060 15484 18228 15540
rect 18172 15316 18228 15484
rect 18172 15250 18228 15260
rect 17836 15150 17838 15202
rect 17890 15150 17892 15202
rect 17836 15138 17892 15150
rect 17948 15204 18004 15214
rect 17724 14466 17780 14476
rect 17836 13748 17892 13758
rect 17388 11330 17444 11340
rect 17500 11676 17668 11732
rect 17724 13746 17892 13748
rect 17724 13694 17838 13746
rect 17890 13694 17892 13746
rect 17724 13692 17892 13694
rect 17164 11230 17166 11282
rect 17218 11230 17220 11282
rect 17164 10500 17220 11230
rect 17500 10948 17556 11676
rect 17500 10882 17556 10892
rect 17612 11506 17668 11518
rect 17612 11454 17614 11506
rect 17666 11454 17668 11506
rect 17276 10836 17332 10846
rect 17276 10622 17332 10780
rect 17276 10570 17278 10622
rect 17330 10570 17332 10622
rect 17276 10558 17332 10570
rect 17164 10444 17332 10500
rect 17052 10332 17220 10388
rect 16604 10220 16772 10276
rect 16940 10220 17108 10276
rect 16492 9986 16548 9996
rect 16156 9940 16212 9950
rect 16156 9846 16212 9884
rect 15484 9772 15596 9828
rect 15540 9716 15596 9772
rect 15932 9826 15988 9838
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15540 9660 15652 9716
rect 15596 9042 15652 9660
rect 15708 9714 15764 9726
rect 15708 9662 15710 9714
rect 15762 9662 15764 9714
rect 15708 9492 15764 9662
rect 15820 9492 15876 9502
rect 15708 9436 15820 9492
rect 15820 9426 15876 9436
rect 15596 8990 15598 9042
rect 15650 8990 15652 9042
rect 15596 8978 15652 8990
rect 15708 8820 15764 8830
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 15372 8194 15428 8206
rect 15596 8260 15652 8270
rect 14924 6972 15092 7028
rect 15148 6972 15316 7028
rect 14924 6802 14980 6972
rect 14924 6750 14926 6802
rect 14978 6750 14980 6802
rect 14924 6738 14980 6750
rect 15036 6802 15092 6814
rect 15036 6750 15038 6802
rect 15090 6750 15092 6802
rect 14700 6514 14756 6524
rect 14252 6402 14308 6412
rect 15036 6244 15092 6750
rect 13580 5012 13636 5022
rect 13244 4956 13524 5012
rect 13468 4788 13524 4956
rect 13580 4918 13636 4956
rect 13020 4498 13076 4508
rect 13244 4732 13524 4788
rect 12908 4338 12964 4396
rect 12908 4286 12910 4338
rect 12962 4286 12964 4338
rect 12908 4274 12964 4286
rect 13020 3780 13076 3790
rect 13020 3686 13076 3724
rect 12684 3668 12740 3678
rect 12684 3574 12740 3612
rect 13244 3388 13300 4732
rect 13468 4340 13524 4350
rect 13356 4228 13412 4238
rect 13356 4134 13412 4172
rect 13468 3554 13524 4284
rect 13468 3502 13470 3554
rect 13522 3502 13524 3554
rect 13468 3490 13524 3502
rect 13580 4228 13636 4238
rect 13580 3388 13636 4172
rect 13916 4228 13972 5068
rect 13916 4162 13972 4172
rect 14028 6076 14196 6132
rect 14364 6188 15092 6244
rect 14028 4004 14084 6076
rect 14140 5908 14196 5918
rect 14140 5906 14308 5908
rect 14140 5854 14142 5906
rect 14194 5854 14308 5906
rect 14140 5852 14308 5854
rect 14140 5842 14196 5852
rect 14140 5236 14196 5246
rect 14140 5122 14196 5180
rect 14140 5070 14142 5122
rect 14194 5070 14196 5122
rect 14140 5058 14196 5070
rect 14028 3938 14084 3948
rect 14252 3780 14308 5852
rect 14252 3714 14308 3724
rect 14364 5906 14420 6188
rect 14476 6020 14532 6030
rect 14476 5926 14532 5964
rect 14364 5854 14366 5906
rect 14418 5854 14420 5906
rect 13692 3668 13748 3678
rect 13692 3666 14196 3668
rect 13692 3614 13694 3666
rect 13746 3614 14196 3666
rect 13692 3612 14196 3614
rect 13692 3602 13748 3612
rect 13244 3332 13524 3388
rect 13580 3332 13748 3388
rect 13020 3108 13076 3118
rect 13020 2770 13076 3052
rect 13020 2718 13022 2770
rect 13074 2718 13076 2770
rect 13020 2706 13076 2718
rect 12796 2548 12852 2558
rect 12796 2454 12852 2492
rect 12460 2158 12462 2210
rect 12514 2158 12516 2210
rect 12460 2146 12516 2158
rect 13468 2210 13524 3332
rect 13468 2158 13470 2210
rect 13522 2158 13524 2210
rect 13468 2146 13524 2158
rect 13580 2772 13636 2782
rect 13580 2098 13636 2716
rect 13580 2046 13582 2098
rect 13634 2046 13636 2098
rect 13580 2034 13636 2046
rect 12348 1922 12404 1932
rect 12908 1988 12964 1998
rect 12908 1894 12964 1932
rect 13468 1764 13524 1774
rect 11788 1150 11790 1202
rect 11842 1150 11844 1202
rect 11788 1138 11844 1150
rect 12348 1652 12404 1662
rect 11564 978 11620 990
rect 11564 926 11566 978
rect 11618 926 11620 978
rect 11564 868 11620 926
rect 11564 802 11620 812
rect 11900 756 11956 766
rect 11900 112 11956 700
rect 12348 112 12404 1596
rect 13244 1652 13300 1662
rect 12796 1316 12852 1326
rect 12572 1204 12628 1214
rect 12572 1110 12628 1148
rect 12796 112 12852 1260
rect 13244 112 13300 1596
rect 7644 18 7700 28
rect 7840 0 7952 112
rect 8288 0 8400 112
rect 8736 0 8848 112
rect 9184 0 9296 112
rect 9632 0 9744 112
rect 10080 0 10192 112
rect 10528 0 10640 112
rect 10976 0 11088 112
rect 11424 0 11536 112
rect 11872 0 11984 112
rect 12320 0 12432 112
rect 12768 0 12880 112
rect 13216 0 13328 112
rect 13468 84 13524 1708
rect 13692 1090 13748 3332
rect 13804 2884 13860 2894
rect 13804 2790 13860 2828
rect 13916 2436 13972 2446
rect 13916 2210 13972 2380
rect 13916 2158 13918 2210
rect 13970 2158 13972 2210
rect 13916 2146 13972 2158
rect 14140 1986 14196 3612
rect 14252 3332 14308 3342
rect 14252 2658 14308 3276
rect 14252 2606 14254 2658
rect 14306 2606 14308 2658
rect 14252 2436 14308 2606
rect 14252 2370 14308 2380
rect 14140 1934 14142 1986
rect 14194 1934 14196 1986
rect 14140 1922 14196 1934
rect 14252 1988 14308 1998
rect 14252 1202 14308 1932
rect 14364 1764 14420 5854
rect 14588 5796 14644 5806
rect 14588 5702 14644 5740
rect 14924 5794 14980 5806
rect 14924 5742 14926 5794
rect 14978 5742 14980 5794
rect 14588 5572 14644 5582
rect 14588 5346 14644 5516
rect 14588 5294 14590 5346
rect 14642 5294 14644 5346
rect 14588 5282 14644 5294
rect 14924 5572 14980 5742
rect 14476 5236 14532 5246
rect 14476 3554 14532 5180
rect 14700 4900 14756 4910
rect 14588 4564 14644 4574
rect 14588 4470 14644 4508
rect 14476 3502 14478 3554
rect 14530 3502 14532 3554
rect 14476 2884 14532 3502
rect 14476 2818 14532 2828
rect 14700 3220 14756 4844
rect 14924 4116 14980 5516
rect 15148 5012 15204 6972
rect 15260 6804 15316 6814
rect 15260 6710 15316 6748
rect 15484 6690 15540 6702
rect 15484 6638 15486 6690
rect 15538 6638 15540 6690
rect 15036 4452 15092 4462
rect 15148 4452 15204 4956
rect 15036 4450 15204 4452
rect 15036 4398 15038 4450
rect 15090 4398 15204 4450
rect 15036 4396 15204 4398
rect 15260 6356 15316 6366
rect 15260 5906 15316 6300
rect 15484 6020 15540 6638
rect 15596 6356 15652 8204
rect 15708 6916 15764 8764
rect 15932 8708 15988 9774
rect 16604 9826 16660 9838
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16044 9716 16100 9726
rect 16044 9380 16100 9660
rect 16268 9604 16324 9614
rect 16044 9314 16100 9324
rect 16156 9548 16268 9604
rect 16156 9042 16212 9548
rect 16268 9538 16324 9548
rect 16156 8990 16158 9042
rect 16210 8990 16212 9042
rect 16156 8978 16212 8990
rect 16268 9380 16324 9390
rect 16268 8930 16324 9324
rect 16604 9380 16660 9774
rect 16716 9658 16772 10220
rect 16828 9828 16884 9866
rect 16828 9762 16884 9772
rect 16940 9826 16996 9838
rect 16940 9774 16942 9826
rect 16994 9774 16996 9826
rect 16940 9716 16996 9774
rect 16716 9602 16884 9658
rect 16940 9650 16996 9660
rect 16604 9314 16660 9324
rect 16716 9044 16772 9054
rect 16716 8950 16772 8988
rect 16268 8878 16270 8930
rect 16322 8878 16324 8930
rect 16268 8866 16324 8878
rect 15932 8652 16660 8708
rect 16604 8482 16660 8652
rect 16604 8430 16606 8482
rect 16658 8430 16660 8482
rect 16604 8418 16660 8430
rect 16828 8482 16884 9602
rect 16828 8430 16830 8482
rect 16882 8430 16884 8482
rect 16828 8418 16884 8430
rect 16940 8372 16996 8382
rect 16940 8278 16996 8316
rect 15820 8258 15876 8270
rect 15820 8206 15822 8258
rect 15874 8206 15876 8258
rect 15820 7364 15876 8206
rect 16268 8260 16324 8270
rect 16156 8146 16212 8158
rect 16156 8094 16158 8146
rect 16210 8094 16212 8146
rect 16156 7476 16212 8094
rect 16156 7410 16212 7420
rect 16268 7474 16324 8204
rect 17052 7812 17108 10220
rect 17164 9826 17220 10332
rect 17164 9774 17166 9826
rect 17218 9774 17220 9826
rect 17164 9762 17220 9774
rect 17276 9828 17332 10444
rect 17388 10386 17444 10398
rect 17388 10334 17390 10386
rect 17442 10334 17444 10386
rect 17388 9828 17444 10334
rect 17500 9828 17556 9838
rect 17388 9826 17556 9828
rect 17388 9774 17502 9826
rect 17554 9774 17556 9826
rect 17388 9772 17556 9774
rect 17276 9762 17332 9772
rect 17500 9762 17556 9772
rect 17052 7746 17108 7756
rect 17276 9042 17332 9054
rect 17276 8990 17278 9042
rect 17330 8990 17332 9042
rect 16268 7422 16270 7474
rect 16322 7422 16324 7474
rect 16268 7410 16324 7422
rect 16716 7588 16772 7598
rect 16716 7474 16772 7532
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16716 7410 16772 7422
rect 15820 7298 15876 7308
rect 15932 7362 15988 7374
rect 15932 7310 15934 7362
rect 15986 7310 15988 7362
rect 15932 7028 15988 7310
rect 16492 7364 16548 7374
rect 15932 6962 15988 6972
rect 16268 7252 16324 7262
rect 15820 6916 15876 6926
rect 15708 6914 15876 6916
rect 15708 6862 15822 6914
rect 15874 6862 15876 6914
rect 15708 6860 15876 6862
rect 15820 6850 15876 6860
rect 15932 6804 15988 6814
rect 15932 6710 15988 6748
rect 15708 6692 15764 6702
rect 15708 6598 15764 6636
rect 16156 6690 16212 6702
rect 16156 6638 16158 6690
rect 16210 6638 16212 6690
rect 15596 6290 15652 6300
rect 15932 6578 15988 6590
rect 15932 6526 15934 6578
rect 15986 6526 15988 6578
rect 15932 6356 15988 6526
rect 15932 6290 15988 6300
rect 15484 5954 15540 5964
rect 15820 6020 15876 6030
rect 15260 5854 15262 5906
rect 15314 5854 15316 5906
rect 15260 4788 15316 5854
rect 15820 5906 15876 5964
rect 15820 5854 15822 5906
rect 15874 5854 15876 5906
rect 15820 5842 15876 5854
rect 15932 5796 15988 5806
rect 15932 5702 15988 5740
rect 16156 5124 16212 6638
rect 16268 6020 16324 7196
rect 16268 5954 16324 5964
rect 16156 5058 16212 5068
rect 16492 5906 16548 7308
rect 16940 7250 16996 7262
rect 16940 7198 16942 7250
rect 16994 7198 16996 7250
rect 16716 6802 16772 6814
rect 16716 6750 16718 6802
rect 16770 6750 16772 6802
rect 16492 5854 16494 5906
rect 16546 5854 16548 5906
rect 15708 4900 15764 4910
rect 16492 4900 16548 5854
rect 16604 6692 16660 6702
rect 16604 5346 16660 6636
rect 16716 6132 16772 6750
rect 16940 6132 16996 7198
rect 17052 6692 17108 6702
rect 17052 6598 17108 6636
rect 17164 6580 17220 6590
rect 16940 6076 17108 6132
rect 16716 6066 16772 6076
rect 16604 5294 16606 5346
rect 16658 5294 16660 5346
rect 16604 5282 16660 5294
rect 15036 4386 15092 4396
rect 14924 4050 14980 4060
rect 14924 3668 14980 3678
rect 14924 3574 14980 3612
rect 15260 3388 15316 4732
rect 15484 4898 16548 4900
rect 15484 4846 15710 4898
rect 15762 4846 16548 4898
rect 15484 4844 16548 4846
rect 16828 5234 16884 5246
rect 16828 5182 16830 5234
rect 16882 5182 16884 5234
rect 15484 4338 15540 4844
rect 15708 4834 15764 4844
rect 16604 4788 16660 4798
rect 16268 4564 16324 4574
rect 15484 4286 15486 4338
rect 15538 4286 15540 4338
rect 15484 4274 15540 4286
rect 15932 4340 15988 4350
rect 15932 4246 15988 4284
rect 16044 4116 16100 4126
rect 16268 4116 16324 4508
rect 16604 4338 16660 4732
rect 16828 4564 16884 5182
rect 16940 5236 16996 5246
rect 17052 5236 17108 6076
rect 17164 5906 17220 6524
rect 17164 5854 17166 5906
rect 17218 5854 17220 5906
rect 17164 5842 17220 5854
rect 16940 5234 17108 5236
rect 16940 5182 16942 5234
rect 16994 5182 17108 5234
rect 16940 5180 17108 5182
rect 16940 5170 16996 5180
rect 16828 4498 16884 4508
rect 16940 5012 16996 5022
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 16044 4114 16212 4116
rect 16044 4062 16046 4114
rect 16098 4062 16212 4114
rect 16044 4060 16212 4062
rect 16044 4050 16100 4060
rect 15932 3780 15988 3790
rect 15932 3444 15988 3724
rect 16156 3556 16212 4060
rect 16156 3490 16212 3500
rect 16044 3444 16100 3454
rect 15932 3442 16100 3444
rect 15932 3390 16046 3442
rect 16098 3390 16100 3442
rect 15932 3388 16100 3390
rect 15260 3332 15428 3388
rect 16044 3378 16100 3388
rect 14700 2660 14756 3164
rect 15372 2994 15428 3332
rect 15372 2942 15374 2994
rect 15426 2942 15428 2994
rect 15372 2930 15428 2942
rect 15820 3332 15876 3342
rect 14700 2594 14756 2604
rect 15596 2772 15652 2782
rect 15260 2324 15316 2334
rect 14924 2212 14980 2222
rect 14924 2118 14980 2156
rect 15260 2210 15316 2268
rect 15260 2158 15262 2210
rect 15314 2158 15316 2210
rect 15260 2146 15316 2158
rect 15596 2210 15652 2716
rect 15820 2658 15876 3276
rect 16156 2996 16212 3006
rect 16156 2770 16212 2940
rect 16156 2718 16158 2770
rect 16210 2718 16212 2770
rect 16156 2706 16212 2718
rect 15820 2606 15822 2658
rect 15874 2606 15876 2658
rect 15820 2594 15876 2606
rect 15596 2158 15598 2210
rect 15650 2158 15652 2210
rect 15596 2146 15652 2158
rect 14588 2100 14644 2110
rect 14588 2006 14644 2044
rect 16156 2100 16212 2110
rect 16268 2100 16324 4060
rect 16828 4004 16884 4014
rect 16716 3780 16772 3790
rect 16604 3556 16660 3566
rect 16604 3462 16660 3500
rect 16156 2098 16324 2100
rect 16156 2046 16158 2098
rect 16210 2046 16324 2098
rect 16156 2044 16324 2046
rect 16492 3444 16548 3454
rect 16156 2034 16212 2044
rect 14364 1698 14420 1708
rect 16044 1764 16100 1774
rect 16044 1670 16100 1708
rect 14252 1150 14254 1202
rect 14306 1150 14308 1202
rect 14252 1138 14308 1150
rect 14588 1652 14644 1662
rect 13692 1038 13694 1090
rect 13746 1038 13748 1090
rect 13692 1026 13748 1038
rect 14140 980 14196 990
rect 13692 868 13748 878
rect 13692 112 13748 812
rect 14140 112 14196 924
rect 14588 112 14644 1596
rect 15036 1652 15092 1662
rect 15036 112 15092 1596
rect 15932 1652 15988 1662
rect 15484 1204 15540 1214
rect 15484 1110 15540 1148
rect 15148 978 15204 990
rect 15148 926 15150 978
rect 15202 926 15204 978
rect 15148 756 15204 926
rect 15148 690 15204 700
rect 15484 756 15540 766
rect 15484 112 15540 700
rect 15932 112 15988 1596
rect 16380 1652 16436 1662
rect 16268 978 16324 990
rect 16268 926 16270 978
rect 16322 926 16324 978
rect 16268 532 16324 926
rect 16268 466 16324 476
rect 16380 112 16436 1596
rect 16492 1202 16548 3388
rect 16604 2884 16660 2894
rect 16716 2884 16772 3724
rect 16828 3388 16884 3948
rect 16940 3778 16996 4956
rect 17276 4338 17332 8990
rect 17500 9044 17556 9054
rect 17500 8950 17556 8988
rect 17388 8260 17444 8270
rect 17388 8166 17444 8204
rect 17500 8146 17556 8158
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 17388 7364 17444 7374
rect 17388 7270 17444 7308
rect 17500 6690 17556 8094
rect 17612 8148 17668 11454
rect 17724 11172 17780 13692
rect 17836 13682 17892 13692
rect 17836 13300 17892 13310
rect 17836 13186 17892 13244
rect 17836 13134 17838 13186
rect 17890 13134 17892 13186
rect 17836 13122 17892 13134
rect 17948 11284 18004 15148
rect 17948 11218 18004 11228
rect 18172 14532 18228 14542
rect 17724 11106 17780 11116
rect 17836 10612 17892 10622
rect 17836 10518 17892 10556
rect 18060 10052 18116 10062
rect 17724 9940 17780 9950
rect 17724 9846 17780 9884
rect 17836 9826 17892 9838
rect 17836 9774 17838 9826
rect 17890 9774 17892 9826
rect 17836 9716 17892 9774
rect 18060 9826 18116 9996
rect 18060 9774 18062 9826
rect 18114 9774 18116 9826
rect 18060 9762 18116 9774
rect 17836 9650 17892 9660
rect 18172 9380 18228 14476
rect 18060 9324 18228 9380
rect 18060 8484 18116 9324
rect 18284 9268 18340 26236
rect 18396 23548 18452 26348
rect 18508 25732 18564 27804
rect 18508 25666 18564 25676
rect 18620 25508 18676 28700
rect 18732 27076 18788 27086
rect 18732 26982 18788 27020
rect 18844 26178 18900 30492
rect 19068 30436 19124 30446
rect 19068 30342 19124 30380
rect 18956 30324 19012 30334
rect 18956 27188 19012 30268
rect 19180 29988 19236 31500
rect 19628 30884 19684 33628
rect 19628 30818 19684 30828
rect 19740 30324 19796 34524
rect 19964 34132 20020 34862
rect 20188 34914 20244 34926
rect 20188 34862 20190 34914
rect 20242 34862 20244 34914
rect 19964 34066 20020 34076
rect 20076 34130 20132 34142
rect 20076 34078 20078 34130
rect 20130 34078 20132 34130
rect 19852 33906 19908 33918
rect 19852 33854 19854 33906
rect 19906 33854 19908 33906
rect 19852 33796 19908 33854
rect 19852 33730 19908 33740
rect 20076 33572 20132 34078
rect 20188 33796 20244 34862
rect 20524 34916 20580 36764
rect 20636 35140 20692 38612
rect 21084 38050 21140 40236
rect 21084 37998 21086 38050
rect 21138 37998 21140 38050
rect 21084 37604 21140 37998
rect 21084 37538 21140 37548
rect 21308 38948 21364 46620
rect 21644 46610 21700 46620
rect 21756 46340 21812 47068
rect 22092 46564 22148 46574
rect 22092 46470 22148 46508
rect 21532 46284 21812 46340
rect 21532 43876 21588 46284
rect 21756 46116 21812 46126
rect 21756 46022 21812 46060
rect 21980 46116 22036 46126
rect 21644 45892 21700 45902
rect 21980 45892 22036 46060
rect 21644 45890 22036 45892
rect 21644 45838 21646 45890
rect 21698 45838 22036 45890
rect 21644 45836 22036 45838
rect 21644 45668 21700 45836
rect 21644 45602 21700 45612
rect 21980 45668 22036 45678
rect 21644 45108 21700 45118
rect 21644 44546 21700 45052
rect 21644 44494 21646 44546
rect 21698 44494 21700 44546
rect 21644 44482 21700 44494
rect 21532 43820 21812 43876
rect 21644 43428 21700 43438
rect 21420 42754 21476 42766
rect 21420 42702 21422 42754
rect 21474 42702 21476 42754
rect 21420 40404 21476 42702
rect 21644 41972 21700 43372
rect 21756 43316 21812 43820
rect 21756 43250 21812 43260
rect 21868 43540 21924 43550
rect 21756 43092 21812 43102
rect 21756 42754 21812 43036
rect 21756 42702 21758 42754
rect 21810 42702 21812 42754
rect 21756 42690 21812 42702
rect 21644 41970 21812 41972
rect 21644 41918 21646 41970
rect 21698 41918 21812 41970
rect 21644 41916 21812 41918
rect 21644 41906 21700 41916
rect 21644 41298 21700 41310
rect 21644 41246 21646 41298
rect 21698 41246 21700 41298
rect 21420 40338 21476 40348
rect 21532 41186 21588 41198
rect 21532 41134 21534 41186
rect 21586 41134 21588 41186
rect 21532 39842 21588 41134
rect 21644 40628 21700 41246
rect 21644 40562 21700 40572
rect 21532 39790 21534 39842
rect 21586 39790 21588 39842
rect 21532 39778 21588 39790
rect 21308 37044 21364 38892
rect 21420 39618 21476 39630
rect 21420 39566 21422 39618
rect 21474 39566 21476 39618
rect 21420 38668 21476 39566
rect 21644 38724 21700 38762
rect 21420 38612 21588 38668
rect 20972 36820 21028 36830
rect 20972 36482 21028 36764
rect 20972 36430 20974 36482
rect 21026 36430 21028 36482
rect 20972 36418 21028 36430
rect 20636 35074 20692 35084
rect 21084 36148 21140 36158
rect 20524 34850 20580 34860
rect 20972 35028 21028 35038
rect 20748 34804 20804 34814
rect 20748 34710 20804 34748
rect 20524 34132 20580 34142
rect 20524 34038 20580 34076
rect 20860 34132 20916 34142
rect 20860 34038 20916 34076
rect 20748 34020 20804 34030
rect 20748 33926 20804 33964
rect 20188 33730 20244 33740
rect 20636 33796 20692 33806
rect 20524 33572 20580 33582
rect 20076 33570 20580 33572
rect 20076 33518 20526 33570
rect 20578 33518 20580 33570
rect 20076 33516 20580 33518
rect 20524 33506 20580 33516
rect 19964 33348 20020 33358
rect 20636 33348 20692 33740
rect 20972 33458 21028 34972
rect 20972 33406 20974 33458
rect 21026 33406 21028 33458
rect 20972 33394 21028 33406
rect 21084 34914 21140 36092
rect 21308 35308 21364 36988
rect 21084 34862 21086 34914
rect 21138 34862 21140 34914
rect 19964 33254 20020 33292
rect 20412 33334 20692 33348
rect 20412 33282 20414 33334
rect 20466 33292 20692 33334
rect 21084 33348 21140 34862
rect 20466 33282 20468 33292
rect 21084 33282 21140 33292
rect 21196 35252 21364 35308
rect 20412 32116 20468 33282
rect 20748 33124 20804 33134
rect 20412 32060 20580 32116
rect 20412 31892 20468 31902
rect 20188 31890 20468 31892
rect 20188 31838 20414 31890
rect 20466 31838 20468 31890
rect 20188 31836 20468 31838
rect 19964 31778 20020 31790
rect 19964 31726 19966 31778
rect 20018 31726 20020 31778
rect 19852 30996 19908 31006
rect 19852 30660 19908 30940
rect 19852 30594 19908 30604
rect 19740 30258 19796 30268
rect 19964 30436 20020 31726
rect 19628 30212 19684 30222
rect 19180 29922 19236 29932
rect 19516 30098 19572 30110
rect 19516 30046 19518 30098
rect 19570 30046 19572 30098
rect 19516 29988 19572 30046
rect 19516 29922 19572 29932
rect 19180 29428 19236 29466
rect 19180 29362 19236 29372
rect 19628 29426 19684 30156
rect 19964 30210 20020 30380
rect 19964 30158 19966 30210
rect 20018 30158 20020 30210
rect 19964 30146 20020 30158
rect 20076 30884 20132 30894
rect 19628 29374 19630 29426
rect 19682 29374 19684 29426
rect 19628 29362 19684 29374
rect 19852 30100 19908 30110
rect 19068 29316 19124 29326
rect 19068 29222 19124 29260
rect 19180 29204 19236 29214
rect 19068 28868 19124 28878
rect 19068 28774 19124 28812
rect 19180 28866 19236 29148
rect 19852 29204 19908 30044
rect 20076 29540 20132 30828
rect 19852 29138 19908 29148
rect 19964 29538 20132 29540
rect 19964 29486 20078 29538
rect 20130 29486 20132 29538
rect 19964 29484 20132 29486
rect 19180 28814 19182 28866
rect 19234 28814 19236 28866
rect 19180 28802 19236 28814
rect 19404 28868 19460 28878
rect 19852 28868 19908 28878
rect 19404 28866 19908 28868
rect 19404 28814 19406 28866
rect 19458 28814 19854 28866
rect 19906 28814 19908 28866
rect 19404 28812 19908 28814
rect 19404 28802 19460 28812
rect 19852 28802 19908 28812
rect 19516 28644 19572 28654
rect 19292 28532 19348 28542
rect 19292 28438 19348 28476
rect 19516 28420 19572 28588
rect 19628 28644 19684 28654
rect 19628 28642 19908 28644
rect 19628 28590 19630 28642
rect 19682 28590 19908 28642
rect 19628 28588 19908 28590
rect 19628 28578 19684 28588
rect 19516 28364 19796 28420
rect 19180 27972 19236 27982
rect 19068 27860 19124 27870
rect 19068 27766 19124 27804
rect 19180 27298 19236 27916
rect 19404 27972 19460 27982
rect 19404 27636 19460 27916
rect 19628 27860 19684 27870
rect 19628 27766 19684 27804
rect 19740 27858 19796 28364
rect 19740 27806 19742 27858
rect 19794 27806 19796 27858
rect 19740 27794 19796 27806
rect 19404 27570 19460 27580
rect 19852 27634 19908 28588
rect 19852 27582 19854 27634
rect 19906 27582 19908 27634
rect 19852 27570 19908 27582
rect 19964 27412 20020 29484
rect 20076 29474 20132 29484
rect 20076 29092 20132 29102
rect 20076 28866 20132 29036
rect 20076 28814 20078 28866
rect 20130 28814 20132 28866
rect 20076 28802 20132 28814
rect 20188 28754 20244 31836
rect 20412 31826 20468 31836
rect 20524 31220 20580 32060
rect 20636 31778 20692 31790
rect 20636 31726 20638 31778
rect 20690 31726 20692 31778
rect 20636 31332 20692 31726
rect 20748 31556 20804 33068
rect 20748 31490 20804 31500
rect 20860 32676 20916 32686
rect 21196 32676 21252 35252
rect 20860 32674 21252 32676
rect 20860 32622 20862 32674
rect 20914 32622 21252 32674
rect 20860 32620 21252 32622
rect 21420 35140 21476 35150
rect 21420 32676 21476 35084
rect 20636 31266 20692 31276
rect 20524 31154 20580 31164
rect 20860 31108 20916 32620
rect 21420 32610 21476 32620
rect 21308 32452 21364 32462
rect 21308 32358 21364 32396
rect 21196 32004 21252 32014
rect 20860 31014 20916 31052
rect 20972 31778 21028 31790
rect 20972 31726 20974 31778
rect 21026 31726 21028 31778
rect 20188 28702 20190 28754
rect 20242 28702 20244 28754
rect 20188 28690 20244 28702
rect 20300 30884 20356 30894
rect 20076 28532 20132 28542
rect 20300 28532 20356 30828
rect 20524 30322 20580 30334
rect 20524 30270 20526 30322
rect 20578 30270 20580 30322
rect 20412 30210 20468 30222
rect 20412 30158 20414 30210
rect 20466 30158 20468 30210
rect 20412 29988 20468 30158
rect 20412 29922 20468 29932
rect 20076 27858 20132 28476
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 20076 27794 20132 27806
rect 20188 28476 20356 28532
rect 20524 28532 20580 30270
rect 20972 30212 21028 31726
rect 21196 30882 21252 31948
rect 21196 30830 21198 30882
rect 21250 30830 21252 30882
rect 21196 30818 21252 30830
rect 21420 31666 21476 31678
rect 21420 31614 21422 31666
rect 21474 31614 21476 31666
rect 21420 31220 21476 31614
rect 21308 30770 21364 30782
rect 21308 30718 21310 30770
rect 21362 30718 21364 30770
rect 20972 30118 21028 30156
rect 21196 30212 21252 30222
rect 21196 29988 21252 30156
rect 21196 29922 21252 29932
rect 20860 29426 20916 29438
rect 20860 29374 20862 29426
rect 20914 29374 20916 29426
rect 20636 29316 20692 29326
rect 20636 29222 20692 29260
rect 20748 29202 20804 29214
rect 20748 29150 20750 29202
rect 20802 29150 20804 29202
rect 20748 28868 20804 29150
rect 20748 28802 20804 28812
rect 20636 28756 20692 28766
rect 20636 28662 20692 28700
rect 20860 28644 20916 29374
rect 21084 29426 21140 29438
rect 21084 29374 21086 29426
rect 21138 29374 21140 29426
rect 20860 28578 20916 28588
rect 20972 28756 21028 28766
rect 20972 28642 21028 28700
rect 20972 28590 20974 28642
rect 21026 28590 21028 28642
rect 19180 27246 19182 27298
rect 19234 27246 19236 27298
rect 19180 27234 19236 27246
rect 19404 27356 20020 27412
rect 20076 27524 20132 27534
rect 18956 27122 19012 27132
rect 18844 26126 18846 26178
rect 18898 26126 18900 26178
rect 18844 26114 18900 26126
rect 19180 27076 19236 27086
rect 18732 25508 18788 25518
rect 18620 25506 18788 25508
rect 18620 25454 18734 25506
rect 18786 25454 18788 25506
rect 18620 25452 18788 25454
rect 18732 25442 18788 25452
rect 18956 25396 19012 25406
rect 18844 24948 18900 24958
rect 18844 24722 18900 24892
rect 18844 24670 18846 24722
rect 18898 24670 18900 24722
rect 18844 24658 18900 24670
rect 18844 23940 18900 23950
rect 18956 23940 19012 25340
rect 18844 23938 19012 23940
rect 18844 23886 18846 23938
rect 18898 23886 19012 23938
rect 18844 23884 19012 23886
rect 19180 23940 19236 27020
rect 19404 25396 19460 27356
rect 19852 27188 19908 27198
rect 19740 26404 19796 26414
rect 19404 25330 19460 25340
rect 19516 26068 19572 26078
rect 18396 23492 18676 23548
rect 18396 22708 18452 22718
rect 18396 22594 18452 22652
rect 18396 22542 18398 22594
rect 18450 22542 18452 22594
rect 18396 22530 18452 22542
rect 18396 22260 18452 22270
rect 18396 21586 18452 22204
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18396 19684 18452 21534
rect 18508 21812 18564 21822
rect 18508 20244 18564 21756
rect 18620 20468 18676 23492
rect 18844 23156 18900 23884
rect 18844 23090 18900 23100
rect 18956 23156 19012 23166
rect 18956 23154 19124 23156
rect 18956 23102 18958 23154
rect 19010 23102 19124 23154
rect 18956 23100 19124 23102
rect 18956 23090 19012 23100
rect 18620 20402 18676 20412
rect 18732 23044 18788 23054
rect 18508 20130 18564 20188
rect 18508 20078 18510 20130
rect 18562 20078 18564 20130
rect 18508 20066 18564 20078
rect 18732 20132 18788 22988
rect 18844 21364 18900 21374
rect 18844 20692 18900 21308
rect 18844 20626 18900 20636
rect 18732 20076 18900 20132
rect 18508 19684 18564 19694
rect 18396 19628 18508 19684
rect 18396 19460 18452 19470
rect 18396 19234 18452 19404
rect 18396 19182 18398 19234
rect 18450 19182 18452 19234
rect 18396 19170 18452 19182
rect 18396 17220 18452 17230
rect 18396 16994 18452 17164
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 18396 16930 18452 16942
rect 18508 16772 18564 19628
rect 18396 16716 18564 16772
rect 18732 17332 18788 17342
rect 18396 14532 18452 16716
rect 18508 16212 18564 16222
rect 18508 16118 18564 16156
rect 18508 15314 18564 15326
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 14756 18564 15262
rect 18732 15316 18788 17276
rect 18844 16770 18900 20076
rect 18956 19908 19012 19918
rect 18956 19348 19012 19852
rect 18956 19282 19012 19292
rect 18956 17892 19012 17902
rect 18956 17666 19012 17836
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18956 16884 19012 17614
rect 18956 16818 19012 16828
rect 18844 16718 18846 16770
rect 18898 16718 18900 16770
rect 18844 16706 18900 16718
rect 18956 15428 19012 15438
rect 18844 15316 18900 15326
rect 18732 15314 18900 15316
rect 18732 15262 18846 15314
rect 18898 15262 18900 15314
rect 18732 15260 18900 15262
rect 18844 15250 18900 15260
rect 18956 14868 19012 15372
rect 19068 15148 19124 23100
rect 19180 17892 19236 23884
rect 19292 24388 19348 24398
rect 19292 19460 19348 24332
rect 19404 23380 19460 23390
rect 19404 23286 19460 23324
rect 19404 23156 19460 23166
rect 19404 22148 19460 23100
rect 19516 22930 19572 26012
rect 19740 26068 19796 26348
rect 19740 26002 19796 26012
rect 19740 25508 19796 25518
rect 19740 25414 19796 25452
rect 19628 24724 19684 24734
rect 19628 24630 19684 24668
rect 19740 24500 19796 24510
rect 19740 23940 19796 24444
rect 19740 23156 19796 23884
rect 19740 23090 19796 23100
rect 19516 22878 19518 22930
rect 19570 22878 19572 22930
rect 19516 22866 19572 22878
rect 19628 22930 19684 22942
rect 19628 22878 19630 22930
rect 19682 22878 19684 22930
rect 19628 22484 19684 22878
rect 19628 22418 19684 22428
rect 19740 22932 19796 22942
rect 19516 22372 19572 22382
rect 19516 22278 19572 22316
rect 19404 22092 19572 22148
rect 19292 19394 19348 19404
rect 19404 20578 19460 20590
rect 19404 20526 19406 20578
rect 19458 20526 19460 20578
rect 19404 19348 19460 20526
rect 19404 19282 19460 19292
rect 19180 17826 19236 17836
rect 19292 19122 19348 19134
rect 19292 19070 19294 19122
rect 19346 19070 19348 19122
rect 19292 17220 19348 19070
rect 19292 17154 19348 17164
rect 19404 18116 19460 18126
rect 19516 18116 19572 22092
rect 19460 18060 19572 18116
rect 19628 20132 19684 20142
rect 19068 15092 19236 15148
rect 18620 14756 18676 14766
rect 18508 14754 18676 14756
rect 18508 14702 18622 14754
rect 18674 14702 18676 14754
rect 18508 14700 18676 14702
rect 18620 14690 18676 14700
rect 18956 14644 19012 14812
rect 19068 14644 19124 14654
rect 18956 14642 19124 14644
rect 18956 14590 19070 14642
rect 19122 14590 19124 14642
rect 18956 14588 19124 14590
rect 19068 14578 19124 14588
rect 18396 14466 18452 14476
rect 19068 13970 19124 13982
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 18620 13860 18676 13870
rect 19068 13860 19124 13918
rect 18620 13858 19124 13860
rect 18620 13806 18622 13858
rect 18674 13806 19124 13858
rect 18620 13804 19124 13806
rect 18620 13794 18676 13804
rect 18732 13634 18788 13646
rect 18732 13582 18734 13634
rect 18786 13582 18788 13634
rect 18508 13524 18564 13534
rect 18508 13430 18564 13468
rect 18620 13076 18676 13086
rect 18508 12404 18564 12414
rect 18396 12180 18452 12190
rect 18396 12086 18452 12124
rect 18508 11172 18564 12348
rect 18508 11106 18564 11116
rect 18508 10612 18564 10622
rect 18508 10518 18564 10556
rect 18060 8418 18116 8428
rect 18172 9212 18340 9268
rect 18396 9268 18452 9278
rect 17948 8370 18004 8382
rect 17948 8318 17950 8370
rect 18002 8318 18004 8370
rect 17948 8260 18004 8318
rect 17948 8194 18004 8204
rect 17612 8082 17668 8092
rect 18060 8148 18116 8158
rect 17500 6638 17502 6690
rect 17554 6638 17556 6690
rect 17500 5124 17556 6638
rect 17612 7812 17668 7822
rect 17612 5796 17668 7756
rect 17948 7474 18004 7486
rect 17948 7422 17950 7474
rect 18002 7422 18004 7474
rect 17948 7140 18004 7422
rect 17948 7074 18004 7084
rect 18060 6804 18116 8092
rect 18060 6710 18116 6748
rect 17948 6132 18004 6142
rect 17948 5906 18004 6076
rect 17948 5854 17950 5906
rect 18002 5854 18004 5906
rect 17948 5842 18004 5854
rect 17612 5740 17780 5796
rect 17612 5124 17668 5134
rect 17500 5122 17668 5124
rect 17500 5070 17614 5122
rect 17666 5070 17668 5122
rect 17500 5068 17668 5070
rect 17276 4286 17278 4338
rect 17330 4286 17332 4338
rect 17276 4274 17332 4286
rect 17500 4788 17556 4798
rect 16940 3726 16942 3778
rect 16994 3726 16996 3778
rect 16940 3714 16996 3726
rect 17052 4116 17108 4126
rect 17052 3666 17108 4060
rect 17052 3614 17054 3666
rect 17106 3614 17108 3666
rect 17052 3602 17108 3614
rect 17164 3554 17220 3566
rect 17164 3502 17166 3554
rect 17218 3502 17220 3554
rect 16828 3332 17108 3388
rect 16604 2882 16772 2884
rect 16604 2830 16606 2882
rect 16658 2830 16772 2882
rect 16604 2828 16772 2830
rect 16604 2818 16660 2828
rect 16716 2660 16772 2670
rect 16716 2566 16772 2604
rect 17052 2210 17108 3332
rect 17164 2660 17220 3502
rect 17500 3388 17556 4732
rect 17612 3556 17668 5068
rect 17724 4228 17780 5740
rect 18172 5684 18228 9212
rect 17948 5628 18228 5684
rect 18284 9044 18340 9054
rect 18396 9044 18452 9212
rect 18284 9042 18452 9044
rect 18284 8990 18286 9042
rect 18338 8990 18452 9042
rect 18284 8988 18452 8990
rect 18620 9044 18676 13020
rect 18732 11620 18788 13582
rect 19068 13524 19124 13534
rect 18956 12852 19012 12862
rect 18956 12758 19012 12796
rect 19068 12402 19124 13468
rect 19180 12852 19236 15092
rect 19292 13746 19348 13758
rect 19292 13694 19294 13746
rect 19346 13694 19348 13746
rect 19292 13636 19348 13694
rect 19292 13570 19348 13580
rect 19404 13076 19460 18060
rect 19516 17666 19572 17678
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19516 17108 19572 17614
rect 19516 17042 19572 17052
rect 19628 16324 19684 20076
rect 19740 19572 19796 22876
rect 19852 20804 19908 27132
rect 19964 26066 20020 26078
rect 19964 26014 19966 26066
rect 20018 26014 20020 26066
rect 19964 25620 20020 26014
rect 19964 25554 20020 25564
rect 19964 24724 20020 24734
rect 19964 22932 20020 24668
rect 19964 22866 20020 22876
rect 19964 22484 20020 22494
rect 20076 22484 20132 27468
rect 20188 27076 20244 28476
rect 20524 28466 20580 28476
rect 20972 28308 21028 28590
rect 20300 28252 21028 28308
rect 20300 27298 20356 28252
rect 20748 28084 20804 28094
rect 21084 28084 21140 29374
rect 20748 28082 21140 28084
rect 20748 28030 20750 28082
rect 20802 28030 21140 28082
rect 20748 28028 21140 28030
rect 21196 28644 21252 28654
rect 20748 28018 20804 28028
rect 20636 27860 20692 27870
rect 21196 27860 21252 28588
rect 21308 28532 21364 30718
rect 21420 29876 21476 31164
rect 21532 30884 21588 38612
rect 21644 35140 21700 38668
rect 21756 37940 21812 41916
rect 21868 40516 21924 43484
rect 21980 42308 22036 45612
rect 21980 42242 22036 42252
rect 22204 45106 22260 45118
rect 22204 45054 22206 45106
rect 22258 45054 22260 45106
rect 22204 44322 22260 45054
rect 22204 44270 22206 44322
rect 22258 44270 22260 44322
rect 22204 44212 22260 44270
rect 22204 43538 22260 44156
rect 22204 43486 22206 43538
rect 22258 43486 22260 43538
rect 21980 41972 22036 41982
rect 21980 41878 22036 41916
rect 21980 41748 22036 41758
rect 21980 40740 22036 41692
rect 22092 41300 22148 41310
rect 22092 41206 22148 41244
rect 21980 40674 22036 40684
rect 21980 40516 22036 40526
rect 21868 40514 22036 40516
rect 21868 40462 21982 40514
rect 22034 40462 22036 40514
rect 21868 40460 22036 40462
rect 21868 38052 21924 40460
rect 21980 40450 22036 40460
rect 22092 40404 22148 40414
rect 22092 39618 22148 40348
rect 22204 40180 22260 43486
rect 22316 42308 22372 47180
rect 22428 45890 22484 47406
rect 22540 48356 22596 48366
rect 22540 46564 22596 48300
rect 22540 46498 22596 46508
rect 22428 45838 22430 45890
rect 22482 45838 22484 45890
rect 22428 45826 22484 45838
rect 22652 45444 22708 48748
rect 22764 47684 22820 48974
rect 22764 47618 22820 47628
rect 22764 47458 22820 47470
rect 22764 47406 22766 47458
rect 22818 47406 22820 47458
rect 22764 46900 22820 47406
rect 22764 46834 22820 46844
rect 22764 45892 22820 45902
rect 22764 45798 22820 45836
rect 22540 44996 22596 45006
rect 22540 44902 22596 44940
rect 22428 44660 22484 44670
rect 22428 44212 22484 44604
rect 22428 44146 22484 44156
rect 22540 44436 22596 44446
rect 22316 42242 22372 42252
rect 22428 43764 22484 43774
rect 22316 41972 22372 41982
rect 22316 40402 22372 41916
rect 22428 40516 22484 43708
rect 22540 42532 22596 44380
rect 22652 43540 22708 45388
rect 22764 44434 22820 44446
rect 22764 44382 22766 44434
rect 22818 44382 22820 44434
rect 22764 44324 22820 44382
rect 22764 44258 22820 44268
rect 22652 43484 22820 43540
rect 22652 43316 22708 43326
rect 22652 43222 22708 43260
rect 22764 42754 22820 43484
rect 22764 42702 22766 42754
rect 22818 42702 22820 42754
rect 22764 42690 22820 42702
rect 22540 42476 22820 42532
rect 22540 41972 22596 41982
rect 22540 41878 22596 41916
rect 22652 41746 22708 41758
rect 22652 41694 22654 41746
rect 22706 41694 22708 41746
rect 22652 41186 22708 41694
rect 22764 41300 22820 42476
rect 22764 41234 22820 41244
rect 22652 41134 22654 41186
rect 22706 41134 22708 41186
rect 22652 41122 22708 41134
rect 22428 40450 22484 40460
rect 22764 40516 22820 40526
rect 22764 40404 22820 40460
rect 22316 40350 22318 40402
rect 22370 40350 22372 40402
rect 22316 40338 22372 40350
rect 22652 40402 22820 40404
rect 22652 40350 22766 40402
rect 22818 40350 22820 40402
rect 22652 40348 22820 40350
rect 22652 40292 22708 40348
rect 22764 40338 22820 40348
rect 22652 40226 22708 40236
rect 22876 40180 22932 53900
rect 22988 53732 23044 53742
rect 22988 53638 23044 53676
rect 23100 53508 23156 53900
rect 22988 53452 23156 53508
rect 22988 43988 23044 53452
rect 23100 53284 23156 53294
rect 23100 53170 23156 53228
rect 23100 53118 23102 53170
rect 23154 53118 23156 53170
rect 23100 53106 23156 53118
rect 23100 51380 23156 51390
rect 23100 51044 23156 51324
rect 23100 44660 23156 50988
rect 23212 49252 23268 55468
rect 23548 55412 23604 55422
rect 23548 55318 23604 55356
rect 23772 55300 23828 55310
rect 23660 55298 23828 55300
rect 23660 55246 23774 55298
rect 23826 55246 23828 55298
rect 23660 55244 23828 55246
rect 23436 54292 23492 54302
rect 23436 54198 23492 54236
rect 23660 53956 23716 55244
rect 23772 55234 23828 55244
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 23772 54740 23828 54750
rect 23772 54514 23828 54684
rect 23772 54462 23774 54514
rect 23826 54462 23828 54514
rect 23772 54450 23828 54462
rect 23884 54292 23940 54302
rect 23884 54198 23940 54236
rect 24108 54290 24164 54302
rect 24108 54238 24110 54290
rect 24162 54238 24164 54290
rect 23436 53900 23716 53956
rect 23324 53842 23380 53854
rect 23324 53790 23326 53842
rect 23378 53790 23380 53842
rect 23324 53620 23380 53790
rect 23324 53554 23380 53564
rect 23436 52836 23492 53900
rect 24108 53844 24164 54238
rect 24108 53778 24164 53788
rect 23212 49186 23268 49196
rect 23324 52780 23492 52836
rect 23548 53730 23604 53742
rect 23548 53678 23550 53730
rect 23602 53678 23604 53730
rect 23324 48468 23380 52780
rect 23548 52500 23604 53678
rect 24220 53620 24276 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 24556 55410 24612 55422
rect 24556 55358 24558 55410
rect 24610 55358 24612 55410
rect 24556 54628 24612 55358
rect 24780 55298 24836 55310
rect 24780 55246 24782 55298
rect 24834 55246 24836 55298
rect 24780 55188 24836 55246
rect 24780 55122 24836 55132
rect 24556 54562 24612 54572
rect 24444 54292 24500 54302
rect 24444 54290 25060 54292
rect 24444 54238 24446 54290
rect 24498 54238 25060 54290
rect 24444 54236 25060 54238
rect 24444 54226 24500 54236
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 24444 53732 24500 53742
rect 24220 53554 24276 53564
rect 24332 53730 24500 53732
rect 24332 53678 24446 53730
rect 24498 53678 24500 53730
rect 24332 53676 24500 53678
rect 24220 53396 24276 53406
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24108 53172 24164 53182
rect 23548 52434 23604 52444
rect 23660 52948 23716 52958
rect 23660 52276 23716 52892
rect 23660 52210 23716 52220
rect 23884 52276 23940 52286
rect 23884 52182 23940 52220
rect 24108 51940 24164 53116
rect 24220 52948 24276 53340
rect 24220 52882 24276 52892
rect 24220 52722 24276 52734
rect 24220 52670 24222 52722
rect 24274 52670 24276 52722
rect 24220 52164 24276 52670
rect 24220 52098 24276 52108
rect 24332 52052 24388 53676
rect 24444 53666 24500 53676
rect 24668 53732 24724 53742
rect 24668 53638 24724 53676
rect 24780 53730 24836 53742
rect 24780 53678 24782 53730
rect 24834 53678 24836 53730
rect 24780 53172 24836 53678
rect 25004 53730 25060 54236
rect 25004 53678 25006 53730
rect 25058 53678 25060 53730
rect 25004 53172 25060 53678
rect 25116 53396 25172 55804
rect 25340 55410 25396 55804
rect 25340 55358 25342 55410
rect 25394 55358 25396 55410
rect 25340 55346 25396 55358
rect 25452 55858 25508 55870
rect 25452 55806 25454 55858
rect 25506 55806 25508 55858
rect 25116 53330 25172 53340
rect 25340 54180 25396 54190
rect 25004 53116 25284 53172
rect 24780 53106 24836 53116
rect 24892 53060 24948 53070
rect 24668 52946 24724 52958
rect 24668 52894 24670 52946
rect 24722 52894 24724 52946
rect 24668 52836 24724 52894
rect 24668 52770 24724 52780
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 24892 52274 24948 53004
rect 25228 53058 25284 53116
rect 25228 53006 25230 53058
rect 25282 53006 25284 53058
rect 25228 52994 25284 53006
rect 24892 52222 24894 52274
rect 24946 52222 24948 52274
rect 24892 52210 24948 52222
rect 25004 52948 25060 52958
rect 25340 52948 25396 54124
rect 25452 53956 25508 55806
rect 25676 55858 25732 55870
rect 25676 55806 25678 55858
rect 25730 55806 25732 55858
rect 25676 55524 25732 55806
rect 25676 55468 25844 55524
rect 25676 55298 25732 55310
rect 25676 55246 25678 55298
rect 25730 55246 25732 55298
rect 25676 54516 25732 55246
rect 25676 54450 25732 54460
rect 25564 54290 25620 54302
rect 25564 54238 25566 54290
rect 25618 54238 25620 54290
rect 25564 54180 25620 54238
rect 25564 54114 25620 54124
rect 25676 53956 25732 53966
rect 25452 53954 25732 53956
rect 25452 53902 25678 53954
rect 25730 53902 25732 53954
rect 25452 53900 25732 53902
rect 25676 53890 25732 53900
rect 25788 53844 25844 55468
rect 26012 54740 26068 56140
rect 26124 55858 26180 55870
rect 26124 55806 26126 55858
rect 26178 55806 26180 55858
rect 26124 55636 26180 55806
rect 26124 55570 26180 55580
rect 26236 55524 26292 57344
rect 26684 56868 26740 57344
rect 26684 56802 26740 56812
rect 26908 56082 26964 56094
rect 26908 56030 26910 56082
rect 26962 56030 26964 56082
rect 26908 55972 26964 56030
rect 27132 56084 27188 57344
rect 27132 56018 27188 56028
rect 26908 55906 26964 55916
rect 26460 55860 26516 55870
rect 26460 55766 26516 55804
rect 27132 55858 27188 55870
rect 27132 55806 27134 55858
rect 27186 55806 27188 55858
rect 26236 55458 26292 55468
rect 26572 55412 26628 55422
rect 26572 55410 26740 55412
rect 26572 55358 26574 55410
rect 26626 55358 26740 55410
rect 26572 55356 26740 55358
rect 26572 55346 26628 55356
rect 26348 55298 26404 55310
rect 26348 55246 26350 55298
rect 26402 55246 26404 55298
rect 26012 54684 26292 54740
rect 26124 54514 26180 54526
rect 26124 54462 26126 54514
rect 26178 54462 26180 54514
rect 26124 54404 26180 54462
rect 26124 54338 26180 54348
rect 25788 53778 25844 53788
rect 25452 53732 25508 53742
rect 25676 53732 25732 53742
rect 25452 53638 25508 53676
rect 25564 53676 25676 53732
rect 25340 52892 25508 52948
rect 24332 51996 24612 52052
rect 24108 51884 24276 51940
rect 23804 51772 24068 51782
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 23804 51706 24068 51716
rect 23772 51604 23828 51614
rect 23436 51154 23492 51166
rect 23436 51102 23438 51154
rect 23490 51102 23492 51154
rect 23436 51044 23492 51102
rect 23436 50978 23492 50988
rect 23772 50596 23828 51548
rect 23996 51604 24052 51614
rect 23996 51378 24052 51548
rect 23996 51326 23998 51378
rect 24050 51326 24052 51378
rect 23996 51314 24052 51326
rect 24220 51266 24276 51884
rect 24220 51214 24222 51266
rect 24274 51214 24276 51266
rect 24220 51202 24276 51214
rect 24332 51268 24388 51278
rect 24332 51174 24388 51212
rect 24556 51156 24612 51996
rect 25004 51604 25060 52892
rect 25340 52724 25396 52734
rect 25340 52630 25396 52668
rect 25228 52276 25284 52286
rect 25228 52164 25284 52220
rect 25004 51538 25060 51548
rect 25116 52162 25284 52164
rect 25116 52110 25230 52162
rect 25282 52110 25284 52162
rect 25116 52108 25284 52110
rect 24668 51380 24724 51390
rect 24668 51286 24724 51324
rect 25004 51380 25060 51390
rect 24556 51100 24948 51156
rect 24108 51044 24164 51054
rect 24108 50820 24164 50988
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 24108 50754 24164 50764
rect 24892 50708 24948 51100
rect 24444 50652 24948 50708
rect 25004 50708 25060 51324
rect 23772 50594 24388 50596
rect 23772 50542 23774 50594
rect 23826 50542 24388 50594
rect 23772 50540 24388 50542
rect 23772 50530 23828 50540
rect 24332 50484 24388 50540
rect 24332 50418 24388 50428
rect 23436 50260 23492 50270
rect 23660 50260 23716 50270
rect 23492 50204 23604 50260
rect 23436 50194 23492 50204
rect 23436 50036 23492 50046
rect 23436 49698 23492 49980
rect 23436 49646 23438 49698
rect 23490 49646 23492 49698
rect 23436 49588 23492 49646
rect 23436 49522 23492 49532
rect 23548 49476 23604 50204
rect 23660 49812 23716 50204
rect 23804 50204 24068 50214
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 24220 50148 24276 50158
rect 23996 50036 24052 50046
rect 24220 50036 24276 50092
rect 24052 49980 24276 50036
rect 23996 49970 24052 49980
rect 23772 49812 23828 49822
rect 23660 49810 23828 49812
rect 23660 49758 23774 49810
rect 23826 49758 23828 49810
rect 23660 49756 23828 49758
rect 23772 49746 23828 49756
rect 24220 49810 24276 49822
rect 24220 49758 24222 49810
rect 24274 49758 24276 49810
rect 23548 49410 23604 49420
rect 24220 49476 24276 49758
rect 24444 49698 24500 50652
rect 25004 50594 25060 50652
rect 25004 50542 25006 50594
rect 25058 50542 25060 50594
rect 25004 50530 25060 50542
rect 25116 51378 25172 52108
rect 25228 52098 25284 52108
rect 25452 51940 25508 52892
rect 25116 51326 25118 51378
rect 25170 51326 25172 51378
rect 24556 50484 24612 50522
rect 24556 50372 24948 50428
rect 24444 49646 24446 49698
rect 24498 49646 24500 49698
rect 24444 49634 24500 49646
rect 24220 49410 24276 49420
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 23324 48402 23380 48412
rect 23436 49140 23492 49150
rect 23324 48018 23380 48030
rect 23324 47966 23326 48018
rect 23378 47966 23380 48018
rect 23324 47684 23380 47966
rect 23324 47618 23380 47628
rect 23324 46900 23380 46910
rect 23324 46806 23380 46844
rect 23100 44604 23380 44660
rect 22988 43932 23268 43988
rect 23100 41858 23156 41870
rect 23100 41806 23102 41858
rect 23154 41806 23156 41858
rect 22988 41188 23044 41198
rect 22988 40290 23044 41132
rect 23100 40404 23156 41806
rect 23100 40338 23156 40348
rect 22988 40238 22990 40290
rect 23042 40238 23044 40290
rect 22988 40226 23044 40238
rect 22204 40124 22484 40180
rect 22092 39566 22094 39618
rect 22146 39566 22148 39618
rect 22092 39554 22148 39566
rect 21868 38050 22036 38052
rect 21868 37998 21870 38050
rect 21922 37998 22036 38050
rect 21868 37996 22036 37998
rect 21868 37986 21924 37996
rect 21756 37874 21812 37884
rect 21868 36820 21924 36830
rect 21756 36372 21812 36382
rect 21756 35810 21812 36316
rect 21756 35758 21758 35810
rect 21810 35758 21812 35810
rect 21756 35746 21812 35758
rect 21868 35588 21924 36764
rect 21868 35522 21924 35532
rect 21644 35074 21700 35084
rect 21756 35026 21812 35038
rect 21756 34974 21758 35026
rect 21810 34974 21812 35026
rect 21644 34914 21700 34926
rect 21644 34862 21646 34914
rect 21698 34862 21700 34914
rect 21644 34020 21700 34862
rect 21756 34132 21812 34974
rect 21756 34066 21812 34076
rect 21644 33954 21700 33964
rect 21868 33684 21924 33694
rect 21756 33348 21812 33358
rect 21756 33254 21812 33292
rect 21532 30818 21588 30828
rect 21644 32676 21700 32686
rect 21644 30660 21700 32620
rect 21868 32676 21924 33628
rect 21980 33460 22036 37996
rect 22316 37940 22372 37950
rect 22204 37266 22260 37278
rect 22204 37214 22206 37266
rect 22258 37214 22260 37266
rect 22092 36484 22148 36494
rect 22092 36390 22148 36428
rect 22204 36372 22260 37214
rect 22204 36306 22260 36316
rect 22092 35588 22148 35598
rect 22092 35494 22148 35532
rect 22204 35028 22260 35038
rect 22204 34934 22260 34972
rect 21980 33404 22148 33460
rect 21868 32610 21924 32620
rect 21980 33236 22036 33246
rect 21980 31892 22036 33180
rect 21980 31826 22036 31836
rect 21644 30594 21700 30604
rect 21756 31108 21812 31118
rect 21644 30436 21700 30446
rect 21420 28642 21476 29820
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21420 28578 21476 28590
rect 21532 30380 21644 30436
rect 21532 30210 21588 30380
rect 21644 30370 21700 30380
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 21308 28466 21364 28476
rect 20636 27766 20692 27804
rect 21084 27804 21252 27860
rect 20972 27636 21028 27646
rect 20860 27634 21028 27636
rect 20860 27582 20974 27634
rect 21026 27582 21028 27634
rect 20860 27580 21028 27582
rect 20300 27246 20302 27298
rect 20354 27246 20356 27298
rect 20300 27234 20356 27246
rect 20524 27412 20580 27422
rect 20524 27188 20580 27356
rect 20860 27300 20916 27580
rect 20972 27570 21028 27580
rect 20524 27122 20580 27132
rect 20636 27244 20916 27300
rect 20972 27412 21028 27422
rect 20188 27020 20356 27076
rect 20300 22540 20356 27020
rect 20524 26964 20580 26974
rect 20524 26740 20580 26908
rect 20524 26674 20580 26684
rect 20636 26292 20692 27244
rect 20748 27076 20804 27086
rect 20972 27076 21028 27356
rect 20748 27074 21028 27076
rect 20748 27022 20750 27074
rect 20802 27022 21028 27074
rect 20748 27020 21028 27022
rect 21084 27074 21140 27804
rect 21308 27748 21364 27758
rect 21308 27746 21476 27748
rect 21308 27694 21310 27746
rect 21362 27694 21476 27746
rect 21308 27692 21476 27694
rect 21308 27682 21364 27692
rect 21084 27022 21086 27074
rect 21138 27022 21140 27074
rect 20748 27010 20804 27020
rect 20972 26740 21028 26750
rect 20524 26236 20692 26292
rect 20860 26516 20916 26526
rect 20412 25732 20468 25742
rect 20412 22798 20468 25676
rect 20524 25396 20580 26236
rect 20860 26180 20916 26460
rect 20972 26290 21028 26684
rect 20972 26238 20974 26290
rect 21026 26238 21028 26290
rect 20972 26226 21028 26238
rect 21084 26292 21140 27022
rect 21196 27634 21252 27646
rect 21196 27582 21198 27634
rect 21250 27582 21252 27634
rect 21196 26516 21252 27582
rect 21308 27524 21364 27534
rect 21308 27188 21364 27468
rect 21308 27122 21364 27132
rect 21196 26450 21252 26460
rect 21308 26852 21364 26862
rect 21308 26402 21364 26796
rect 21308 26350 21310 26402
rect 21362 26350 21364 26402
rect 21308 26338 21364 26350
rect 21196 26292 21252 26302
rect 21084 26236 21196 26292
rect 20748 26178 20916 26180
rect 20748 26126 20862 26178
rect 20914 26126 20916 26178
rect 20748 26124 20916 26126
rect 20636 26066 20692 26078
rect 20636 26014 20638 26066
rect 20690 26014 20692 26066
rect 20636 25732 20692 26014
rect 20636 25666 20692 25676
rect 20636 25508 20692 25518
rect 20636 25414 20692 25452
rect 20524 25330 20580 25340
rect 20524 24948 20580 24958
rect 20524 23156 20580 24892
rect 20524 23090 20580 23100
rect 20636 24610 20692 24622
rect 20636 24558 20638 24610
rect 20690 24558 20692 24610
rect 20412 22742 20580 22798
rect 20300 22484 20468 22540
rect 19964 22482 20132 22484
rect 19964 22430 19966 22482
rect 20018 22430 20132 22482
rect 19964 22428 20132 22430
rect 19964 22418 20020 22428
rect 20300 22372 20356 22382
rect 20076 22370 20356 22372
rect 20076 22318 20302 22370
rect 20354 22318 20356 22370
rect 20076 22316 20356 22318
rect 19964 21812 20020 21822
rect 20076 21812 20132 22316
rect 20300 22306 20356 22316
rect 19964 21810 20132 21812
rect 19964 21758 19966 21810
rect 20018 21758 20132 21810
rect 19964 21756 20132 21758
rect 19964 21746 20020 21756
rect 19852 20738 19908 20748
rect 19964 20802 20020 20814
rect 19964 20750 19966 20802
rect 20018 20750 20020 20802
rect 19964 20468 20020 20750
rect 19964 20402 20020 20412
rect 19740 19506 19796 19516
rect 20300 19460 20356 19470
rect 20300 19366 20356 19404
rect 19740 19236 19796 19246
rect 20076 19236 20132 19246
rect 19740 19234 20020 19236
rect 19740 19182 19742 19234
rect 19794 19182 20020 19234
rect 19740 19180 20020 19182
rect 19740 19170 19796 19180
rect 19964 17106 20020 19180
rect 20076 19142 20132 19180
rect 20412 18788 20468 22484
rect 20524 22484 20580 22742
rect 20524 22418 20580 22428
rect 20636 22036 20692 24558
rect 20748 24050 20804 26124
rect 20860 26114 20916 26124
rect 21084 26068 21140 26236
rect 21196 26226 21252 26236
rect 20972 26012 21140 26068
rect 20972 25620 21028 26012
rect 21308 25956 21364 25966
rect 20972 25506 21028 25564
rect 21196 25620 21252 25630
rect 20972 25454 20974 25506
rect 21026 25454 21028 25506
rect 20972 25442 21028 25454
rect 21084 25508 21140 25518
rect 21084 24834 21140 25452
rect 21084 24782 21086 24834
rect 21138 24782 21140 24834
rect 21084 24770 21140 24782
rect 20748 23998 20750 24050
rect 20802 23998 20804 24050
rect 20748 23156 20804 23998
rect 20860 24610 20916 24622
rect 20860 24558 20862 24610
rect 20914 24558 20916 24610
rect 20860 24162 20916 24558
rect 21196 24388 21252 25564
rect 21308 25508 21364 25900
rect 21420 25620 21476 27692
rect 21532 27412 21588 30158
rect 21644 30212 21700 30222
rect 21644 28980 21700 30156
rect 21756 29538 21812 31052
rect 22092 30996 22148 33404
rect 22316 32788 22372 37884
rect 22428 35700 22484 40124
rect 22764 40124 22932 40180
rect 22540 39956 22596 39966
rect 22540 39844 22596 39900
rect 22540 39788 22708 39844
rect 22540 39620 22596 39630
rect 22540 39526 22596 39564
rect 22652 37268 22708 39788
rect 22764 38274 22820 40124
rect 22764 38222 22766 38274
rect 22818 38222 22820 38274
rect 22764 38210 22820 38222
rect 22876 38610 22932 38622
rect 22876 38558 22878 38610
rect 22930 38558 22932 38610
rect 22876 37940 22932 38558
rect 22876 37874 22932 37884
rect 23100 37826 23156 37838
rect 23100 37774 23102 37826
rect 23154 37774 23156 37826
rect 22652 37212 22932 37268
rect 22540 37156 22596 37166
rect 22540 37062 22596 37100
rect 22428 34130 22484 35644
rect 22428 34078 22430 34130
rect 22482 34078 22484 34130
rect 22428 34066 22484 34078
rect 22764 37044 22820 37054
rect 22764 34914 22820 36988
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22652 33572 22708 33582
rect 22316 32722 22372 32732
rect 22540 33348 22596 33358
rect 22428 32338 22484 32350
rect 22428 32286 22430 32338
rect 22482 32286 22484 32338
rect 22428 31892 22484 32286
rect 22428 31826 22484 31836
rect 22092 30930 22148 30940
rect 22316 31666 22372 31678
rect 22316 31614 22318 31666
rect 22370 31614 22372 31666
rect 22316 30100 22372 31614
rect 22428 31220 22484 31230
rect 22428 31126 22484 31164
rect 22316 30034 22372 30044
rect 21756 29486 21758 29538
rect 21810 29486 21812 29538
rect 21756 29474 21812 29486
rect 21868 29540 21924 29550
rect 21644 28924 21812 28980
rect 21532 27346 21588 27356
rect 21644 28754 21700 28766
rect 21644 28702 21646 28754
rect 21698 28702 21700 28754
rect 21532 27188 21588 27198
rect 21532 27074 21588 27132
rect 21532 27022 21534 27074
rect 21586 27022 21588 27074
rect 21532 27010 21588 27022
rect 21644 26516 21700 28702
rect 21756 27524 21812 28924
rect 21868 27972 21924 29484
rect 22092 29316 22148 29326
rect 22092 29222 22148 29260
rect 22204 28756 22260 28766
rect 22092 28644 22148 28654
rect 22092 28550 22148 28588
rect 22092 27972 22148 27982
rect 21868 27970 22036 27972
rect 21868 27918 21870 27970
rect 21922 27918 22036 27970
rect 21868 27916 22036 27918
rect 21868 27906 21924 27916
rect 21756 27458 21812 27468
rect 21756 27186 21812 27198
rect 21756 27134 21758 27186
rect 21810 27134 21812 27186
rect 21756 26740 21812 27134
rect 21756 26674 21812 26684
rect 21868 27188 21924 27198
rect 21644 26460 21812 26516
rect 21644 26292 21700 26302
rect 21644 26198 21700 26236
rect 21644 25674 21700 25686
rect 21644 25622 21646 25674
rect 21698 25622 21700 25674
rect 21644 25620 21700 25622
rect 21420 25564 21700 25620
rect 21308 25494 21476 25508
rect 21308 25452 21422 25494
rect 21420 25442 21422 25452
rect 21474 25442 21476 25494
rect 21420 25430 21476 25442
rect 21196 24322 21252 24332
rect 21308 24722 21364 24734
rect 21308 24670 21310 24722
rect 21362 24670 21364 24722
rect 21308 24276 21364 24670
rect 21644 24722 21700 24734
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21644 24612 21700 24670
rect 21644 24546 21700 24556
rect 21308 24210 21364 24220
rect 21644 24388 21700 24398
rect 20860 24110 20862 24162
rect 20914 24110 20916 24162
rect 20860 24052 20916 24110
rect 21644 24162 21700 24332
rect 21644 24110 21646 24162
rect 21698 24110 21700 24162
rect 21644 24098 21700 24110
rect 20860 23986 20916 23996
rect 21420 24052 21476 24090
rect 21420 23986 21476 23996
rect 21756 24050 21812 26460
rect 21868 26404 21924 27132
rect 21868 26338 21924 26348
rect 21756 23998 21758 24050
rect 21810 23998 21812 24050
rect 21756 23986 21812 23998
rect 21308 23938 21364 23950
rect 21308 23886 21310 23938
rect 21362 23886 21364 23938
rect 21980 23946 22036 27916
rect 22092 26292 22148 27916
rect 22204 27186 22260 28700
rect 22540 28644 22596 33292
rect 22652 33346 22708 33516
rect 22652 33294 22654 33346
rect 22706 33294 22708 33346
rect 22652 33282 22708 33294
rect 22652 31890 22708 31902
rect 22652 31838 22654 31890
rect 22706 31838 22708 31890
rect 22652 31108 22708 31838
rect 22652 30548 22708 31052
rect 22652 30482 22708 30492
rect 22652 30212 22708 30222
rect 22764 30212 22820 34862
rect 22652 30210 22820 30212
rect 22652 30158 22654 30210
rect 22706 30158 22820 30210
rect 22652 30156 22820 30158
rect 22652 30146 22708 30156
rect 22652 28644 22708 28654
rect 22540 28642 22708 28644
rect 22540 28590 22654 28642
rect 22706 28590 22708 28642
rect 22540 28588 22708 28590
rect 22652 28578 22708 28588
rect 22316 28196 22372 28206
rect 22316 27634 22372 28140
rect 22316 27582 22318 27634
rect 22370 27582 22372 27634
rect 22316 27412 22372 27582
rect 22316 27346 22372 27356
rect 22204 27134 22206 27186
rect 22258 27134 22260 27186
rect 22204 27122 22260 27134
rect 22428 27074 22484 27086
rect 22428 27022 22430 27074
rect 22482 27022 22484 27074
rect 22428 26908 22484 27022
rect 22764 27074 22820 30156
rect 22764 27022 22766 27074
rect 22818 27022 22820 27074
rect 22764 27010 22820 27022
rect 22428 26852 22708 26908
rect 22204 26292 22260 26302
rect 22092 26290 22260 26292
rect 22092 26238 22206 26290
rect 22258 26238 22260 26290
rect 22092 26236 22260 26238
rect 22204 25956 22260 26236
rect 22204 25890 22260 25900
rect 22316 26066 22372 26078
rect 22652 26068 22708 26852
rect 22764 26178 22820 26190
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 22764 26068 22820 26126
rect 22316 26014 22318 26066
rect 22370 26014 22372 26066
rect 22316 25844 22372 26014
rect 22316 25778 22372 25788
rect 22428 26012 22820 26068
rect 22316 25508 22372 25518
rect 22428 25508 22484 26012
rect 22652 25508 22708 25518
rect 22316 25506 22484 25508
rect 22316 25454 22318 25506
rect 22370 25454 22484 25506
rect 22316 25452 22484 25454
rect 22540 25506 22708 25508
rect 22540 25454 22654 25506
rect 22706 25454 22708 25506
rect 22540 25452 22708 25454
rect 22316 25442 22372 25452
rect 22540 24948 22596 25452
rect 22652 25442 22708 25452
rect 22540 24882 22596 24892
rect 22652 25172 22708 25182
rect 22204 24500 22260 24510
rect 22204 24498 22484 24500
rect 22204 24446 22206 24498
rect 22258 24446 22484 24498
rect 22204 24444 22484 24446
rect 22204 24434 22260 24444
rect 22428 24052 22484 24444
rect 22428 23996 22596 24052
rect 22204 23946 22260 23950
rect 21980 23938 22260 23946
rect 21980 23890 22206 23938
rect 20748 23090 20804 23100
rect 21084 23828 21140 23838
rect 20748 22932 20804 22942
rect 20748 22370 20804 22876
rect 20972 22596 21028 22606
rect 20972 22502 21028 22540
rect 20748 22318 20750 22370
rect 20802 22318 20804 22370
rect 20748 22260 20804 22318
rect 20748 22194 20804 22204
rect 20636 21980 20916 22036
rect 20748 21586 20804 21598
rect 20748 21534 20750 21586
rect 20802 21534 20804 21586
rect 20524 21252 20580 21262
rect 20524 21026 20580 21196
rect 20524 20974 20526 21026
rect 20578 20974 20580 21026
rect 20524 20962 20580 20974
rect 20748 20468 20804 21534
rect 20860 21588 20916 21980
rect 20972 21588 21028 21598
rect 20860 21532 20972 21588
rect 20972 21522 21028 21532
rect 21084 20818 21140 23772
rect 21308 23828 21364 23886
rect 22204 23886 22206 23890
rect 22258 23886 22260 23938
rect 22204 23874 22260 23886
rect 21308 23762 21364 23772
rect 21868 23828 21924 23838
rect 21196 23716 21252 23726
rect 21196 21474 21252 23660
rect 21532 23716 21588 23726
rect 21588 23660 21812 23716
rect 21308 23492 21364 23502
rect 21308 22708 21364 23436
rect 21532 23266 21588 23660
rect 21532 23214 21534 23266
rect 21586 23214 21588 23266
rect 21532 23202 21588 23214
rect 21756 23156 21812 23660
rect 21868 23380 21924 23772
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 21868 23314 21924 23324
rect 22092 23492 22148 23502
rect 21644 23100 21812 23156
rect 21532 22708 21588 22718
rect 21308 22652 21532 22708
rect 21644 22708 21700 23100
rect 21868 23042 21924 23054
rect 21868 22990 21870 23042
rect 21922 22990 21924 23042
rect 21644 22652 21812 22708
rect 21532 22642 21588 22652
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21196 21422 21198 21474
rect 21250 21422 21252 21474
rect 21196 21410 21252 21422
rect 21420 21252 21476 21262
rect 21476 21196 21700 21252
rect 21420 21186 21476 21196
rect 21644 21026 21700 21196
rect 21644 20974 21646 21026
rect 21698 20974 21700 21026
rect 21644 20962 21700 20974
rect 21084 20762 21252 20818
rect 20748 20402 20804 20412
rect 20860 20692 20916 20702
rect 20748 19348 20804 19358
rect 20748 19254 20804 19292
rect 20412 18722 20468 18732
rect 20412 18564 20468 18574
rect 20300 18452 20356 18462
rect 20188 17892 20244 17902
rect 20188 17798 20244 17836
rect 19964 17054 19966 17106
rect 20018 17054 20020 17106
rect 19964 17042 20020 17054
rect 20076 17220 20132 17230
rect 19628 16258 19684 16268
rect 19964 16884 20020 16894
rect 19740 16100 19796 16110
rect 19740 16006 19796 16044
rect 19852 15764 19908 15774
rect 19852 15314 19908 15708
rect 19852 15262 19854 15314
rect 19906 15262 19908 15314
rect 19852 15250 19908 15262
rect 19740 14868 19796 14878
rect 19404 13010 19460 13020
rect 19516 14530 19572 14542
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19516 14084 19572 14478
rect 19404 12852 19460 12862
rect 19180 12850 19460 12852
rect 19180 12798 19406 12850
rect 19458 12798 19460 12850
rect 19180 12796 19460 12798
rect 19068 12350 19070 12402
rect 19122 12350 19124 12402
rect 19068 12180 19124 12350
rect 19068 12114 19124 12124
rect 19180 12068 19236 12078
rect 19180 11974 19236 12012
rect 18732 11554 18788 11564
rect 18844 11732 18900 11742
rect 18732 11396 18788 11406
rect 18844 11396 18900 11676
rect 18732 11394 18900 11396
rect 18732 11342 18734 11394
rect 18786 11342 18900 11394
rect 18732 11340 18900 11342
rect 19180 11396 19236 11406
rect 18732 11330 18788 11340
rect 19180 11282 19236 11340
rect 19180 11230 19182 11282
rect 19234 11230 19236 11282
rect 19180 11172 19236 11230
rect 19180 11106 19236 11116
rect 18956 10612 19012 10622
rect 18732 9716 18788 9726
rect 18788 9660 18900 9716
rect 18732 9622 18788 9660
rect 17724 4172 17892 4228
rect 17612 3490 17668 3500
rect 17500 3332 17780 3388
rect 17276 2884 17332 2894
rect 17276 2790 17332 2828
rect 17500 2884 17556 2894
rect 17164 2594 17220 2604
rect 17052 2158 17054 2210
rect 17106 2158 17108 2210
rect 17052 2146 17108 2158
rect 16492 1150 16494 1202
rect 16546 1150 16548 1202
rect 16492 1138 16548 1150
rect 16716 2098 16772 2110
rect 16716 2046 16718 2098
rect 16770 2046 16772 2098
rect 16716 1204 16772 2046
rect 16716 1138 16772 1148
rect 16828 1652 16884 1662
rect 16828 112 16884 1596
rect 17276 1652 17332 1662
rect 17276 112 17332 1596
rect 17500 1202 17556 2828
rect 17724 2548 17780 3332
rect 17724 2454 17780 2492
rect 17612 2324 17668 2334
rect 17612 1874 17668 2268
rect 17724 2100 17780 2110
rect 17724 2006 17780 2044
rect 17612 1822 17614 1874
rect 17666 1822 17668 1874
rect 17612 1810 17668 1822
rect 17836 1764 17892 4172
rect 17948 2884 18004 5628
rect 18284 5572 18340 8988
rect 18620 8978 18676 8988
rect 18844 9044 18900 9660
rect 18844 8978 18900 8988
rect 18396 8484 18452 8494
rect 18396 6804 18452 8428
rect 18620 8372 18676 8382
rect 18396 6748 18564 6804
rect 18508 6580 18564 6748
rect 18620 6692 18676 8316
rect 18620 6626 18676 6636
rect 18956 7474 19012 10556
rect 19068 10164 19124 10174
rect 19068 9380 19124 10108
rect 19068 9314 19124 9324
rect 19180 9938 19236 9950
rect 19180 9886 19182 9938
rect 19234 9886 19236 9938
rect 19180 9716 19236 9886
rect 19180 8484 19236 9660
rect 19180 8418 19236 8428
rect 19068 8260 19124 8270
rect 19068 8166 19124 8204
rect 18956 7422 18958 7474
rect 19010 7422 19012 7474
rect 18060 5516 18340 5572
rect 18396 6524 18564 6580
rect 18396 5908 18452 6524
rect 18060 4338 18116 5516
rect 18172 5348 18228 5358
rect 18396 5348 18452 5852
rect 18172 5346 18452 5348
rect 18172 5294 18174 5346
rect 18226 5294 18452 5346
rect 18172 5292 18452 5294
rect 18508 6356 18564 6366
rect 18956 6356 19012 7422
rect 19292 7812 19348 12796
rect 19404 12786 19460 12796
rect 19516 11732 19572 14028
rect 19516 11394 19572 11676
rect 19628 13746 19684 13758
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 19628 11954 19684 13694
rect 19740 13748 19796 14812
rect 19964 14530 20020 16828
rect 20076 14868 20132 17164
rect 20188 16548 20244 16558
rect 20188 16210 20244 16492
rect 20188 16158 20190 16210
rect 20242 16158 20244 16210
rect 20188 16146 20244 16158
rect 20300 15988 20356 18396
rect 20412 17892 20468 18508
rect 20412 17826 20468 17836
rect 20860 18562 20916 20636
rect 21084 20692 21140 20702
rect 21084 20130 21140 20636
rect 21084 20078 21086 20130
rect 21138 20078 21140 20130
rect 21084 20066 21140 20078
rect 20860 18510 20862 18562
rect 20914 18510 20916 18562
rect 20412 17668 20468 17678
rect 20748 17668 20804 17678
rect 20412 17666 20692 17668
rect 20412 17614 20414 17666
rect 20466 17614 20692 17666
rect 20412 17612 20692 17614
rect 20412 17602 20468 17612
rect 20524 16100 20580 16110
rect 20636 16100 20692 17612
rect 20748 17574 20804 17612
rect 20860 17220 20916 18510
rect 21196 18228 21252 20762
rect 21532 20020 21588 20030
rect 21420 19906 21476 19918
rect 21420 19854 21422 19906
rect 21474 19854 21476 19906
rect 21308 19572 21364 19582
rect 21308 19234 21364 19516
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 21308 19170 21364 19182
rect 21420 19236 21476 19854
rect 21532 19572 21588 19964
rect 21532 19506 21588 19516
rect 21420 19170 21476 19180
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21308 18228 21364 18238
rect 21196 18226 21364 18228
rect 21196 18174 21310 18226
rect 21362 18174 21364 18226
rect 21196 18172 21364 18174
rect 21308 17668 21364 18172
rect 21532 18228 21588 19182
rect 21756 19236 21812 22652
rect 21868 20580 21924 22990
rect 21980 22484 22036 22494
rect 21980 22370 22036 22428
rect 21980 22318 21982 22370
rect 22034 22318 22036 22370
rect 21980 22306 22036 22318
rect 21868 20514 21924 20524
rect 21756 19170 21812 19180
rect 21532 18162 21588 18172
rect 21308 17602 21364 17612
rect 21196 17556 21252 17566
rect 21196 17462 21252 17500
rect 20860 17154 20916 17164
rect 21756 17220 21812 17230
rect 21756 16996 21812 17164
rect 21756 16994 22036 16996
rect 21756 16942 21758 16994
rect 21810 16942 22036 16994
rect 21756 16940 22036 16942
rect 21756 16930 21812 16940
rect 21308 16884 21364 16894
rect 21196 16324 21252 16334
rect 21196 16230 21252 16268
rect 20972 16100 21028 16110
rect 20636 16098 21028 16100
rect 20636 16046 20974 16098
rect 21026 16046 21028 16098
rect 20636 16044 21028 16046
rect 20524 16006 20580 16044
rect 20412 15988 20468 15998
rect 20300 15932 20412 15988
rect 20412 15876 20468 15932
rect 20412 15820 20804 15876
rect 20748 15314 20804 15820
rect 20748 15262 20750 15314
rect 20802 15262 20804 15314
rect 20748 15250 20804 15262
rect 20076 14802 20132 14812
rect 20972 14868 21028 16044
rect 21308 15988 21364 16828
rect 21196 15932 21364 15988
rect 21532 16548 21588 16558
rect 20972 14802 21028 14812
rect 21084 15204 21140 15214
rect 20076 14644 20132 14654
rect 20076 14642 20244 14644
rect 20076 14590 20078 14642
rect 20130 14590 20244 14642
rect 20076 14588 20244 14590
rect 20076 14578 20132 14588
rect 19964 14478 19966 14530
rect 20018 14478 20020 14530
rect 19852 14308 19908 14318
rect 19852 13858 19908 14252
rect 19852 13806 19854 13858
rect 19906 13806 19908 13858
rect 19852 13794 19908 13806
rect 19964 13748 20020 14478
rect 19964 13692 20132 13748
rect 19740 13682 19796 13692
rect 19740 13524 19796 13534
rect 19740 13430 19796 13468
rect 19964 13522 20020 13534
rect 19964 13470 19966 13522
rect 20018 13470 20020 13522
rect 19628 11902 19630 11954
rect 19682 11902 19684 11954
rect 19628 11508 19684 11902
rect 19740 12962 19796 12974
rect 19740 12910 19742 12962
rect 19794 12910 19796 12962
rect 19740 11732 19796 12910
rect 19964 12290 20020 13470
rect 20076 12404 20132 13692
rect 20188 13188 20244 14588
rect 20636 14532 20692 14542
rect 20636 13860 20692 14476
rect 20748 14532 20804 14542
rect 20748 14530 20916 14532
rect 20748 14478 20750 14530
rect 20802 14478 20916 14530
rect 20748 14476 20916 14478
rect 20748 14466 20804 14476
rect 20188 13122 20244 13132
rect 20300 13858 20692 13860
rect 20300 13806 20638 13858
rect 20690 13806 20692 13858
rect 20300 13804 20692 13806
rect 20188 12964 20244 12974
rect 20188 12870 20244 12908
rect 20300 12898 20356 13804
rect 20636 13794 20692 13804
rect 20748 13524 20804 13534
rect 20860 13524 20916 14476
rect 21084 14530 21140 15148
rect 21084 14478 21086 14530
rect 21138 14478 21140 14530
rect 21084 14466 21140 14478
rect 20972 14084 21028 14094
rect 20972 13746 21028 14028
rect 20972 13694 20974 13746
rect 21026 13694 21028 13746
rect 20972 13682 21028 13694
rect 21084 13524 21140 13534
rect 20860 13468 21084 13524
rect 20412 13076 20468 13086
rect 20412 13074 20692 13076
rect 20412 13022 20414 13074
rect 20466 13022 20692 13074
rect 20412 13020 20692 13022
rect 20412 13010 20468 13020
rect 20300 12842 20468 12898
rect 20076 12348 20244 12404
rect 19964 12238 19966 12290
rect 20018 12238 20020 12290
rect 19964 12226 20020 12238
rect 19852 12180 19908 12190
rect 19852 12086 19908 12124
rect 20076 12180 20132 12190
rect 20076 12086 20132 12124
rect 20188 11788 20244 12348
rect 19740 11666 19796 11676
rect 19852 11732 20244 11788
rect 20300 12068 20356 12078
rect 19852 11508 19908 11732
rect 20188 11620 20244 11630
rect 20188 11526 20244 11564
rect 19628 11442 19684 11452
rect 19740 11452 19908 11508
rect 19516 11342 19518 11394
rect 19570 11342 19572 11394
rect 19516 11330 19572 11342
rect 19404 10610 19460 10622
rect 19404 10558 19406 10610
rect 19458 10558 19460 10610
rect 19404 10052 19460 10558
rect 19404 9986 19460 9996
rect 19292 7476 19348 7756
rect 19292 7410 19348 7420
rect 19516 8148 19572 8158
rect 19740 8148 19796 11452
rect 19964 11394 20020 11406
rect 19964 11342 19966 11394
rect 20018 11342 20020 11394
rect 19964 10836 20020 11342
rect 19964 10770 20020 10780
rect 20076 10948 20132 10958
rect 19964 8372 20020 8382
rect 19516 8146 19796 8148
rect 19516 8094 19518 8146
rect 19570 8094 19796 8146
rect 19516 8092 19796 8094
rect 19852 8258 19908 8270
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19180 6692 19236 6702
rect 19180 6598 19236 6636
rect 19516 6580 19572 8092
rect 19852 7476 19908 8206
rect 19516 6514 19572 6524
rect 19740 6690 19796 6702
rect 19740 6638 19742 6690
rect 19794 6638 19796 6690
rect 19740 6356 19796 6638
rect 19852 6692 19908 7420
rect 19852 6626 19908 6636
rect 18956 6300 19796 6356
rect 18172 5282 18228 5292
rect 18396 5012 18452 5022
rect 18060 4286 18062 4338
rect 18114 4286 18116 4338
rect 18060 4274 18116 4286
rect 18284 4452 18340 4462
rect 18172 3556 18228 3566
rect 18172 3462 18228 3500
rect 17948 2818 18004 2828
rect 18060 2660 18116 2670
rect 18060 2100 18116 2604
rect 18284 2324 18340 4396
rect 18396 4340 18452 4956
rect 18396 4274 18452 4284
rect 18508 3556 18564 6300
rect 18956 6132 19012 6142
rect 18508 3490 18564 3500
rect 18620 5236 18676 5246
rect 18620 4450 18676 5180
rect 18956 4788 19012 6076
rect 19740 5908 19796 5918
rect 19292 5906 19796 5908
rect 19292 5854 19742 5906
rect 19794 5854 19796 5906
rect 19292 5852 19796 5854
rect 19964 5908 20020 8316
rect 20076 8148 20132 10892
rect 20076 8082 20132 8092
rect 20188 10052 20244 10062
rect 20188 8260 20244 9996
rect 20300 10050 20356 12012
rect 20300 9998 20302 10050
rect 20354 9998 20356 10050
rect 20300 9986 20356 9998
rect 20300 8260 20356 8270
rect 20188 8258 20356 8260
rect 20188 8206 20302 8258
rect 20354 8206 20356 8258
rect 20188 8204 20356 8206
rect 20188 7364 20244 8204
rect 20300 8194 20356 8204
rect 20188 7298 20244 7308
rect 20076 7252 20132 7262
rect 20076 6130 20132 7196
rect 20076 6078 20078 6130
rect 20130 6078 20132 6130
rect 20076 6066 20132 6078
rect 20188 6692 20244 6702
rect 19964 5852 20132 5908
rect 19292 5348 19348 5852
rect 19740 5842 19796 5852
rect 19852 5682 19908 5694
rect 19852 5630 19854 5682
rect 19906 5630 19908 5682
rect 18956 4722 19012 4732
rect 19068 5346 19348 5348
rect 19068 5294 19294 5346
rect 19346 5294 19348 5346
rect 19068 5292 19348 5294
rect 18620 4398 18622 4450
rect 18674 4398 18676 4450
rect 18508 3332 18564 3342
rect 18284 2268 18452 2324
rect 18060 2034 18116 2044
rect 18284 2100 18340 2110
rect 18284 2006 18340 2044
rect 17948 1988 18004 1998
rect 17948 1894 18004 1932
rect 17500 1150 17502 1202
rect 17554 1150 17556 1202
rect 17500 1138 17556 1150
rect 17724 1708 17892 1764
rect 18060 1764 18116 1774
rect 17724 112 17780 1708
rect 18060 1090 18116 1708
rect 18060 1038 18062 1090
rect 18114 1038 18116 1090
rect 18060 1026 18116 1038
rect 18172 1652 18228 1662
rect 18172 112 18228 1596
rect 18396 756 18452 2268
rect 18508 980 18564 3276
rect 18620 2884 18676 4398
rect 19068 4450 19124 5292
rect 19292 5282 19348 5292
rect 19628 5572 19684 5582
rect 19180 5124 19236 5134
rect 19180 4562 19236 5068
rect 19628 4788 19684 5516
rect 19740 5124 19796 5134
rect 19740 5030 19796 5068
rect 19628 4732 19796 4788
rect 19180 4510 19182 4562
rect 19234 4510 19236 4562
rect 19180 4498 19236 4510
rect 19068 4398 19070 4450
rect 19122 4398 19124 4450
rect 19068 4386 19124 4398
rect 18956 4228 19012 4238
rect 18732 4116 18788 4126
rect 18732 4114 18900 4116
rect 18732 4062 18734 4114
rect 18786 4062 18900 4114
rect 18732 4060 18900 4062
rect 18732 4050 18788 4060
rect 18732 3668 18788 3678
rect 18732 3574 18788 3612
rect 18844 3444 18900 4060
rect 18844 3378 18900 3388
rect 18956 3108 19012 4172
rect 19628 4114 19684 4126
rect 19628 4062 19630 4114
rect 19682 4062 19684 4114
rect 19628 3780 19684 4062
rect 19628 3714 19684 3724
rect 18956 3042 19012 3052
rect 18620 2818 18676 2828
rect 19068 2772 19124 2782
rect 18844 2546 18900 2558
rect 18844 2494 18846 2546
rect 18898 2494 18900 2546
rect 18620 2436 18676 2446
rect 18620 1764 18676 2380
rect 18844 2436 18900 2494
rect 18732 1988 18788 1998
rect 18844 1988 18900 2380
rect 18788 1932 18900 1988
rect 19068 1986 19124 2716
rect 19516 2772 19572 2782
rect 19292 2212 19348 2222
rect 19292 2118 19348 2156
rect 19068 1934 19070 1986
rect 19122 1934 19124 1986
rect 18732 1894 18788 1932
rect 19068 1922 19124 1934
rect 19180 1988 19236 1998
rect 18620 1708 18788 1764
rect 18732 1204 18788 1708
rect 19180 1426 19236 1932
rect 19516 1988 19572 2716
rect 19516 1922 19572 1932
rect 19740 1764 19796 4732
rect 19852 4338 19908 5630
rect 19964 5682 20020 5694
rect 19964 5630 19966 5682
rect 20018 5630 20020 5682
rect 19964 5572 20020 5630
rect 19964 5506 20020 5516
rect 20076 5348 20132 5852
rect 19964 5292 20132 5348
rect 19964 4900 20020 5292
rect 20188 5122 20244 6636
rect 20412 6020 20468 12842
rect 20636 12402 20692 13020
rect 20636 12350 20638 12402
rect 20690 12350 20692 12402
rect 20636 12338 20692 12350
rect 20748 12290 20804 13468
rect 20972 13076 21028 13086
rect 20748 12238 20750 12290
rect 20802 12238 20804 12290
rect 20748 12226 20804 12238
rect 20860 12962 20916 12974
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20860 12852 20916 12910
rect 20748 11508 20804 11518
rect 20748 9266 20804 11452
rect 20860 11394 20916 12796
rect 20972 12178 21028 13020
rect 21084 12962 21140 13468
rect 21084 12910 21086 12962
rect 21138 12910 21140 12962
rect 21084 12898 21140 12910
rect 20972 12126 20974 12178
rect 21026 12126 21028 12178
rect 20972 12068 21028 12126
rect 20972 12002 21028 12012
rect 20860 11342 20862 11394
rect 20914 11342 20916 11394
rect 20860 11330 20916 11342
rect 21196 11394 21252 15932
rect 21532 15652 21588 16492
rect 21756 16324 21812 16334
rect 21532 15586 21588 15596
rect 21644 16100 21700 16110
rect 21308 15540 21364 15550
rect 21308 15202 21364 15484
rect 21644 15316 21700 16044
rect 21756 15652 21812 16268
rect 21756 15586 21812 15596
rect 21868 16098 21924 16110
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 15540 21924 16046
rect 21868 15474 21924 15484
rect 21644 15260 21924 15316
rect 21308 15150 21310 15202
rect 21362 15150 21364 15202
rect 21308 15138 21364 15150
rect 21756 14868 21812 14878
rect 21308 14532 21364 14542
rect 21308 14438 21364 14476
rect 21420 13748 21476 13758
rect 21420 13654 21476 13692
rect 21644 13522 21700 13534
rect 21644 13470 21646 13522
rect 21698 13470 21700 13522
rect 21196 11342 21198 11394
rect 21250 11342 21252 11394
rect 20748 9214 20750 9266
rect 20802 9214 20804 9266
rect 20748 9202 20804 9214
rect 20860 11172 20916 11182
rect 20524 8372 20580 8382
rect 20524 8278 20580 8316
rect 20636 7812 20692 7822
rect 20636 7586 20692 7756
rect 20636 7534 20638 7586
rect 20690 7534 20692 7586
rect 20636 6692 20692 7534
rect 20636 6626 20692 6636
rect 20860 7140 20916 11116
rect 20972 10724 21028 10734
rect 20972 10630 21028 10668
rect 21196 10612 21252 11342
rect 21196 10546 21252 10556
rect 21308 12964 21364 12974
rect 21308 11732 21364 12908
rect 21532 12964 21588 12974
rect 21532 12870 21588 12908
rect 21308 11284 21364 11676
rect 20972 8260 21028 8270
rect 20972 8166 21028 8204
rect 20972 7476 21028 7486
rect 21308 7476 21364 11228
rect 21420 12852 21476 12862
rect 21420 12178 21476 12796
rect 21420 12126 21422 12178
rect 21474 12126 21476 12178
rect 21420 10724 21476 12126
rect 21420 10658 21476 10668
rect 21532 12516 21588 12526
rect 21420 10388 21476 10398
rect 21532 10388 21588 12460
rect 21644 12180 21700 13470
rect 21644 12114 21700 12124
rect 21756 11172 21812 14812
rect 21868 13748 21924 15260
rect 21868 13682 21924 13692
rect 21980 12292 22036 16940
rect 22092 16436 22148 23436
rect 22316 23380 22372 23774
rect 22316 23314 22372 23324
rect 22540 23156 22596 23996
rect 22540 23090 22596 23100
rect 22652 22036 22708 25116
rect 22764 24948 22820 24958
rect 22764 24724 22820 24892
rect 22764 24162 22820 24668
rect 22764 24110 22766 24162
rect 22818 24110 22820 24162
rect 22764 24098 22820 24110
rect 22204 21980 22708 22036
rect 22764 23604 22820 23614
rect 22764 22708 22820 23548
rect 22204 21812 22260 21980
rect 22204 21746 22260 21756
rect 22428 21812 22484 21822
rect 22764 21812 22820 22652
rect 22428 21810 22820 21812
rect 22428 21758 22430 21810
rect 22482 21758 22820 21810
rect 22428 21756 22820 21758
rect 22428 21746 22484 21756
rect 22764 21028 22820 21038
rect 22876 21028 22932 37212
rect 23100 37044 23156 37774
rect 23100 36978 23156 36988
rect 22988 36372 23044 36382
rect 22988 35588 23044 36316
rect 22988 35522 23044 35532
rect 23100 35476 23156 35486
rect 22988 33906 23044 33918
rect 22988 33854 22990 33906
rect 23042 33854 23044 33906
rect 22988 27412 23044 33854
rect 23100 32562 23156 35420
rect 23100 32510 23102 32562
rect 23154 32510 23156 32562
rect 23100 32498 23156 32510
rect 23100 30996 23156 31006
rect 23100 30902 23156 30940
rect 22988 27188 23044 27356
rect 22988 27122 23044 27132
rect 23100 29316 23156 29326
rect 22988 26180 23044 26190
rect 22988 23716 23044 26124
rect 23100 24388 23156 29260
rect 23100 24322 23156 24332
rect 22988 23650 23044 23660
rect 23100 23156 23156 23166
rect 23100 23062 23156 23100
rect 22988 22372 23044 22382
rect 22988 22278 23044 22316
rect 23212 21812 23268 43932
rect 23324 41972 23380 44604
rect 23436 43092 23492 49084
rect 23660 49140 23716 49150
rect 23548 48468 23604 48478
rect 23548 46564 23604 48412
rect 23548 46498 23604 46508
rect 23660 47460 23716 49084
rect 23772 49026 23828 49038
rect 23772 48974 23774 49026
rect 23826 48974 23828 49026
rect 23772 48804 23828 48974
rect 23772 48738 23828 48748
rect 24220 48692 24276 48702
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 23804 48570 24068 48580
rect 23996 48242 24052 48254
rect 23996 48190 23998 48242
rect 24050 48190 24052 48242
rect 23772 47460 23828 47470
rect 23660 47458 23828 47460
rect 23660 47406 23774 47458
rect 23826 47406 23828 47458
rect 23660 47404 23828 47406
rect 23660 46228 23716 47404
rect 23772 47394 23828 47404
rect 23996 47236 24052 48190
rect 24220 47796 24276 48636
rect 24220 47730 24276 47740
rect 24332 48132 24388 48142
rect 24332 47236 24388 48076
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 24444 47236 24500 47246
rect 23996 47180 24276 47236
rect 24332 47180 24444 47236
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 24220 47012 24276 47180
rect 24444 47170 24500 47180
rect 24668 47234 24724 47246
rect 24668 47182 24670 47234
rect 24722 47182 24724 47234
rect 23884 46676 23940 46686
rect 24220 46676 24276 46956
rect 23884 46674 24276 46676
rect 23884 46622 23886 46674
rect 23938 46622 24276 46674
rect 23884 46620 24276 46622
rect 24444 46676 24500 46686
rect 23884 46340 23940 46620
rect 24444 46562 24500 46620
rect 24444 46510 24446 46562
rect 24498 46510 24500 46562
rect 24444 46498 24500 46510
rect 24668 46452 24724 47182
rect 24892 47068 24948 50372
rect 25004 50148 25060 50158
rect 25004 49140 25060 50092
rect 25116 49810 25172 51326
rect 25116 49758 25118 49810
rect 25170 49758 25172 49810
rect 25116 49746 25172 49758
rect 25228 51884 25508 51940
rect 25564 51940 25620 53676
rect 25676 53666 25732 53676
rect 25900 53730 25956 53742
rect 25900 53678 25902 53730
rect 25954 53678 25956 53730
rect 25788 53620 25844 53630
rect 25788 53526 25844 53564
rect 25900 52948 25956 53678
rect 26124 53730 26180 53742
rect 26124 53678 26126 53730
rect 26178 53678 26180 53730
rect 26124 53172 26180 53678
rect 26236 53284 26292 54684
rect 26348 53956 26404 55246
rect 26572 54516 26628 54526
rect 26348 53890 26404 53900
rect 26460 54404 26516 54414
rect 26348 53732 26404 53742
rect 26348 53638 26404 53676
rect 26236 53218 26292 53228
rect 26124 53106 26180 53116
rect 25900 52882 25956 52892
rect 26348 52836 26404 52846
rect 26460 52836 26516 54348
rect 26572 53844 26628 54460
rect 26684 53956 26740 55356
rect 26908 55300 26964 55310
rect 26908 55206 26964 55244
rect 27132 54852 27188 55806
rect 27468 55860 27524 55870
rect 27244 55412 27300 55422
rect 27244 55410 27412 55412
rect 27244 55358 27246 55410
rect 27298 55358 27412 55410
rect 27244 55356 27412 55358
rect 27244 55346 27300 55356
rect 27132 54786 27188 54796
rect 27020 54514 27076 54526
rect 27020 54462 27022 54514
rect 27074 54462 27076 54514
rect 27020 54068 27076 54462
rect 27244 54292 27300 54302
rect 27244 54198 27300 54236
rect 27020 54012 27300 54068
rect 26684 53900 26964 53956
rect 26572 53788 26740 53844
rect 26572 53618 26628 53630
rect 26572 53566 26574 53618
rect 26626 53566 26628 53618
rect 26572 53172 26628 53566
rect 26572 53106 26628 53116
rect 26404 52780 26516 52836
rect 25788 52722 25844 52734
rect 25788 52670 25790 52722
rect 25842 52670 25844 52722
rect 25676 52500 25732 52510
rect 25676 52162 25732 52444
rect 25676 52110 25678 52162
rect 25730 52110 25732 52162
rect 25676 52098 25732 52110
rect 25564 51884 25732 51940
rect 25116 49252 25172 49262
rect 25116 49158 25172 49196
rect 25004 49074 25060 49084
rect 25004 47460 25060 47470
rect 25004 47366 25060 47404
rect 24892 47012 25172 47068
rect 24668 46386 24724 46396
rect 25004 46340 25060 46350
rect 23884 46274 23940 46284
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 23660 46162 23716 46172
rect 25004 46116 25060 46284
rect 23772 46060 25060 46116
rect 23772 45780 23828 46060
rect 23884 45892 23940 45902
rect 23884 45798 23940 45836
rect 23548 45724 23828 45780
rect 24892 45778 24948 45790
rect 24892 45726 24894 45778
rect 24946 45726 24948 45778
rect 23548 44436 23604 45724
rect 23660 45612 24500 45668
rect 23660 45556 23716 45612
rect 23660 45490 23716 45500
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 24332 45444 24388 45454
rect 23772 45220 23828 45230
rect 23660 45164 23772 45220
rect 23660 44772 23716 45164
rect 23772 45154 23828 45164
rect 24220 45220 24276 45230
rect 24332 45220 24388 45388
rect 24220 45218 24388 45220
rect 24220 45166 24222 45218
rect 24274 45166 24388 45218
rect 24220 45164 24388 45166
rect 24220 45154 24276 45164
rect 24444 44996 24500 45612
rect 24668 45108 24724 45118
rect 24668 45014 24724 45052
rect 24444 44930 24500 44940
rect 23660 44706 23716 44716
rect 23772 44882 23828 44894
rect 23772 44830 23774 44882
rect 23826 44830 23828 44882
rect 23772 44660 23828 44830
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 23772 44604 24164 44660
rect 24464 44650 24728 44660
rect 24108 44578 24164 44604
rect 24108 44522 24276 44578
rect 23884 44436 23940 44446
rect 23548 44434 23940 44436
rect 23548 44382 23886 44434
rect 23938 44382 23940 44434
rect 23548 44380 23940 44382
rect 24220 44436 24276 44522
rect 24220 44380 24612 44436
rect 23884 44370 23940 44380
rect 23996 44100 24052 44110
rect 24220 44100 24276 44110
rect 24052 44044 24220 44100
rect 23996 44034 24052 44044
rect 24220 44034 24276 44044
rect 23436 43026 23492 43036
rect 23548 43988 23604 43998
rect 23324 40964 23380 41916
rect 23548 41636 23604 43932
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 24220 43876 24276 43886
rect 24220 43764 24276 43820
rect 23660 43708 24276 43764
rect 23660 41970 23716 43708
rect 24556 43538 24612 44380
rect 24780 44324 24836 44334
rect 24780 44100 24836 44268
rect 24780 44034 24836 44044
rect 24892 44210 24948 45726
rect 24892 44158 24894 44210
rect 24946 44158 24948 44210
rect 24892 43988 24948 44158
rect 24892 43922 24948 43932
rect 25004 45106 25060 45118
rect 25004 45054 25006 45106
rect 25058 45054 25060 45106
rect 24556 43486 24558 43538
rect 24610 43486 24612 43538
rect 24556 43474 24612 43486
rect 25004 43540 25060 45054
rect 25004 43446 25060 43484
rect 24220 43426 24276 43438
rect 24220 43374 24222 43426
rect 24274 43374 24276 43426
rect 23772 43314 23828 43326
rect 23772 43262 23774 43314
rect 23826 43262 23828 43314
rect 23772 43092 23828 43262
rect 23772 43026 23828 43036
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 24220 42084 24276 43374
rect 24332 43428 24388 43438
rect 24332 43092 24388 43372
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 24332 43026 24388 43036
rect 25116 42980 25172 47012
rect 25228 45108 25284 51884
rect 25452 51378 25508 51390
rect 25452 51326 25454 51378
rect 25506 51326 25508 51378
rect 25340 50708 25396 50718
rect 25340 50594 25396 50652
rect 25340 50542 25342 50594
rect 25394 50542 25396 50594
rect 25340 50530 25396 50542
rect 25452 50428 25508 51326
rect 25564 51268 25620 51278
rect 25564 50818 25620 51212
rect 25676 51266 25732 51884
rect 25676 51214 25678 51266
rect 25730 51214 25732 51266
rect 25676 51202 25732 51214
rect 25564 50766 25566 50818
rect 25618 50766 25620 50818
rect 25564 50754 25620 50766
rect 25340 50372 25508 50428
rect 25340 47796 25396 50372
rect 25564 50260 25620 50270
rect 25564 49810 25620 50204
rect 25564 49758 25566 49810
rect 25618 49758 25620 49810
rect 25452 48804 25508 48814
rect 25452 48710 25508 48748
rect 25564 48468 25620 49758
rect 25788 49138 25844 52670
rect 25900 52388 25956 52398
rect 26348 52388 26404 52780
rect 25900 52294 25956 52332
rect 26124 52332 26404 52388
rect 26124 52052 26180 52332
rect 26012 51996 26180 52052
rect 26236 52164 26292 52174
rect 25900 50932 25956 50942
rect 25900 50484 25956 50876
rect 25900 50418 25956 50428
rect 25788 49086 25790 49138
rect 25842 49086 25844 49138
rect 25788 49074 25844 49086
rect 25564 48402 25620 48412
rect 25676 49028 25732 49038
rect 25564 48020 25620 48030
rect 25564 47926 25620 47964
rect 25340 47740 25508 47796
rect 25340 47572 25396 47582
rect 25340 47478 25396 47516
rect 25340 46228 25396 46238
rect 25340 46114 25396 46172
rect 25340 46062 25342 46114
rect 25394 46062 25396 46114
rect 25340 45780 25396 46062
rect 25340 45714 25396 45724
rect 25452 45220 25508 47740
rect 25676 47570 25732 48972
rect 25676 47518 25678 47570
rect 25730 47518 25732 47570
rect 25676 47506 25732 47518
rect 25900 49028 25956 49038
rect 25452 45154 25508 45164
rect 25564 46450 25620 46462
rect 25564 46398 25566 46450
rect 25618 46398 25620 46450
rect 25228 45052 25396 45108
rect 25228 44884 25284 44894
rect 25228 44790 25284 44828
rect 25228 44660 25284 44670
rect 25228 44434 25284 44604
rect 25228 44382 25230 44434
rect 25282 44382 25284 44434
rect 25228 44370 25284 44382
rect 24220 42018 24276 42028
rect 24780 42924 25172 42980
rect 25228 43314 25284 43326
rect 25228 43262 25230 43314
rect 25282 43262 25284 43314
rect 23660 41918 23662 41970
rect 23714 41918 23716 41970
rect 23660 41906 23716 41918
rect 24780 41970 24836 42924
rect 25228 42420 25284 43262
rect 25228 42354 25284 42364
rect 24780 41918 24782 41970
rect 24834 41918 24836 41970
rect 24780 41748 24836 41918
rect 24780 41682 24836 41692
rect 25004 41972 25060 41982
rect 23548 41570 23604 41580
rect 24220 41636 24276 41646
rect 23884 41524 23940 41534
rect 23660 41188 23716 41198
rect 23660 41094 23716 41132
rect 23884 40964 23940 41468
rect 23324 40908 23716 40964
rect 23436 40404 23492 40414
rect 23436 40310 23492 40348
rect 23548 40292 23604 40302
rect 23436 40068 23492 40078
rect 23324 38724 23380 38734
rect 23324 38164 23380 38668
rect 23324 38098 23380 38108
rect 23324 36036 23380 36046
rect 23324 35922 23380 35980
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 23324 35588 23380 35598
rect 23324 33628 23380 35532
rect 23436 34020 23492 40012
rect 23548 39618 23604 40236
rect 23548 39566 23550 39618
rect 23602 39566 23604 39618
rect 23548 39172 23604 39566
rect 23548 39106 23604 39116
rect 23548 38948 23604 38958
rect 23548 38854 23604 38892
rect 23548 38052 23604 38062
rect 23548 37958 23604 37996
rect 23436 33954 23492 33964
rect 23548 36484 23604 36494
rect 23660 36484 23716 40908
rect 23884 40898 23940 40908
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 23772 40516 23828 40526
rect 23772 39508 23828 40460
rect 23772 39442 23828 39452
rect 24108 40404 24164 40414
rect 24220 40404 24276 41580
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 24108 40402 24276 40404
rect 24108 40350 24110 40402
rect 24162 40350 24276 40402
rect 24108 40348 24276 40350
rect 24444 40852 24500 40862
rect 24108 39508 24164 40348
rect 24220 40180 24276 40190
rect 24444 40180 24500 40796
rect 25004 40402 25060 41916
rect 25228 41188 25284 41198
rect 25340 41188 25396 45052
rect 25564 44324 25620 46398
rect 25676 46340 25732 46350
rect 25676 45106 25732 46284
rect 25676 45054 25678 45106
rect 25730 45054 25732 45106
rect 25676 45042 25732 45054
rect 25564 44258 25620 44268
rect 25900 44212 25956 48972
rect 25900 44146 25956 44156
rect 25676 43428 25732 43438
rect 25676 43334 25732 43372
rect 25452 41970 25508 41982
rect 25452 41918 25454 41970
rect 25506 41918 25508 41970
rect 25452 41300 25508 41918
rect 25900 41748 25956 41758
rect 25900 41654 25956 41692
rect 25452 41244 25844 41300
rect 25340 41132 25508 41188
rect 25004 40350 25006 40402
rect 25058 40350 25060 40402
rect 25004 40338 25060 40350
rect 25116 40404 25172 40414
rect 24276 40124 24500 40180
rect 24892 40292 24948 40302
rect 24220 40114 24276 40124
rect 24464 40012 24728 40022
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 24108 39442 24164 39452
rect 24332 39620 24388 39630
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 23804 39162 24068 39172
rect 23772 38836 23828 38846
rect 23772 38500 23828 38780
rect 23996 38836 24052 38846
rect 23996 38722 24052 38780
rect 23996 38670 23998 38722
rect 24050 38670 24052 38722
rect 23996 38612 24052 38670
rect 23996 38546 24052 38556
rect 23772 38434 23828 38444
rect 23884 38164 23940 38174
rect 23884 38070 23940 38108
rect 24332 37716 24388 39564
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 24220 37604 24276 37614
rect 24220 37156 24276 37548
rect 24220 37062 24276 37100
rect 23772 37042 23828 37054
rect 23772 36990 23774 37042
rect 23826 36990 23828 37042
rect 23772 36820 23828 36990
rect 23772 36754 23828 36764
rect 24332 36596 24388 37660
rect 24556 37940 24612 37950
rect 24556 37266 24612 37884
rect 24892 37604 24948 40236
rect 25116 38948 25172 40348
rect 25228 39732 25284 41132
rect 25228 39666 25284 39676
rect 25340 40964 25396 40974
rect 25116 38882 25172 38892
rect 24892 37538 24948 37548
rect 25116 38610 25172 38622
rect 25116 38558 25118 38610
rect 25170 38558 25172 38610
rect 25004 37268 25060 37278
rect 24556 37214 24558 37266
rect 24610 37214 24612 37266
rect 24556 37156 24612 37214
rect 24556 37090 24612 37100
rect 24892 37266 25060 37268
rect 24892 37214 25006 37266
rect 25058 37214 25060 37266
rect 24892 37212 25060 37214
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24556 36596 24612 36606
rect 24332 36594 24612 36596
rect 24332 36542 24558 36594
rect 24610 36542 24612 36594
rect 24332 36540 24612 36542
rect 24556 36530 24612 36540
rect 23604 36428 23716 36484
rect 24892 36484 24948 37212
rect 25004 37202 25060 37212
rect 25116 37268 25172 38558
rect 23324 33572 23492 33628
rect 23324 30212 23380 30222
rect 23324 29650 23380 30156
rect 23324 29598 23326 29650
rect 23378 29598 23380 29650
rect 23324 29586 23380 29598
rect 23436 29540 23492 33572
rect 23436 29474 23492 29484
rect 23436 27860 23492 27870
rect 23436 27766 23492 27804
rect 23324 26290 23380 26302
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 25172 23380 26238
rect 23324 25106 23380 25116
rect 23436 26180 23492 26190
rect 23324 24498 23380 24510
rect 23324 24446 23326 24498
rect 23378 24446 23380 24498
rect 23324 23268 23380 24446
rect 23324 23202 23380 23212
rect 23436 23044 23492 26124
rect 23548 25508 23604 36428
rect 24892 36418 24948 36428
rect 25004 36484 25060 36494
rect 25116 36484 25172 37212
rect 25228 38164 25284 38174
rect 25228 37154 25284 38108
rect 25228 37102 25230 37154
rect 25282 37102 25284 37154
rect 25228 37090 25284 37102
rect 25004 36482 25172 36484
rect 25004 36430 25006 36482
rect 25058 36430 25172 36482
rect 25004 36428 25172 36430
rect 25004 36418 25060 36428
rect 23660 36316 24500 36372
rect 23660 36260 23716 36316
rect 23660 36194 23716 36204
rect 24444 36148 24500 36316
rect 24892 36260 24948 36270
rect 24668 36204 24892 36260
rect 24668 36148 24724 36204
rect 24892 36194 24948 36204
rect 23804 36092 24068 36102
rect 24444 36092 24724 36148
rect 25228 36148 25284 36158
rect 23660 36036 23716 36046
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 24892 36036 24948 36046
rect 23660 35700 23716 35980
rect 23996 35700 24052 35710
rect 23660 35644 23828 35700
rect 23772 35588 23828 35644
rect 23996 35698 24612 35700
rect 23996 35646 23998 35698
rect 24050 35646 24612 35698
rect 23996 35644 24612 35646
rect 23996 35634 24052 35644
rect 23772 35522 23828 35532
rect 23772 35252 23828 35262
rect 23772 34916 23828 35196
rect 23772 34850 23828 34860
rect 23884 34914 23940 34926
rect 23884 34862 23886 34914
rect 23938 34862 23940 34914
rect 23884 34692 23940 34862
rect 24332 34804 24388 35644
rect 24444 35476 24500 35514
rect 24556 35476 24612 35644
rect 24668 35476 24724 35486
rect 24556 35420 24668 35476
rect 24444 35410 24500 35420
rect 24668 35410 24724 35420
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24332 34748 24836 34804
rect 23660 34636 23884 34692
rect 23660 31332 23716 34636
rect 23884 34626 23940 34636
rect 24556 34580 24612 34590
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 24556 34020 24612 34524
rect 24332 34018 24612 34020
rect 24332 33966 24558 34018
rect 24610 33966 24612 34018
rect 24332 33964 24612 33966
rect 23884 33908 23940 33918
rect 23884 33460 23940 33852
rect 24108 33908 24164 33918
rect 24108 33814 24164 33852
rect 24332 33796 24388 33964
rect 24556 33954 24612 33964
rect 24780 33908 24836 34748
rect 24892 34130 24948 35980
rect 24892 34078 24894 34130
rect 24946 34078 24948 34130
rect 24892 34066 24948 34078
rect 25116 35364 25172 35374
rect 25116 34804 25172 35308
rect 25228 34914 25284 36092
rect 25228 34862 25230 34914
rect 25282 34862 25284 34914
rect 25228 34850 25284 34862
rect 25116 34132 25172 34748
rect 25340 34804 25396 40908
rect 25452 38500 25508 41132
rect 25788 41186 25844 41244
rect 26012 41188 26068 51996
rect 26124 50596 26180 50606
rect 26124 44548 26180 50540
rect 26236 50594 26292 52108
rect 26348 52162 26404 52174
rect 26348 52110 26350 52162
rect 26402 52110 26404 52162
rect 26348 51380 26404 52110
rect 26348 51286 26404 51324
rect 26460 51716 26516 51726
rect 26460 51044 26516 51660
rect 26684 51492 26740 53788
rect 26796 53730 26852 53742
rect 26796 53678 26798 53730
rect 26850 53678 26852 53730
rect 26796 53508 26852 53678
rect 26796 53442 26852 53452
rect 26908 52948 26964 53900
rect 27132 53844 27188 53854
rect 26908 52882 26964 52892
rect 27020 53730 27076 53742
rect 27020 53678 27022 53730
rect 27074 53678 27076 53730
rect 26908 52722 26964 52734
rect 26908 52670 26910 52722
rect 26962 52670 26964 52722
rect 26908 52612 26964 52670
rect 27020 52724 27076 53678
rect 27020 52658 27076 52668
rect 26908 52546 26964 52556
rect 26908 52388 26964 52398
rect 26908 52162 26964 52332
rect 26908 52110 26910 52162
rect 26962 52110 26964 52162
rect 26908 52098 26964 52110
rect 26572 51436 26740 51492
rect 26796 51716 26852 51726
rect 26572 51156 26628 51436
rect 26796 51378 26852 51660
rect 26796 51326 26798 51378
rect 26850 51326 26852 51378
rect 26796 51314 26852 51326
rect 26572 51100 26852 51156
rect 26460 50988 26740 51044
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 26236 50530 26292 50542
rect 26572 50594 26628 50606
rect 26572 50542 26574 50594
rect 26626 50542 26628 50594
rect 26572 50428 26628 50542
rect 26348 50372 26628 50428
rect 26236 49140 26292 49150
rect 26236 49046 26292 49084
rect 26236 48242 26292 48254
rect 26236 48190 26238 48242
rect 26290 48190 26292 48242
rect 26236 47012 26292 48190
rect 26236 46786 26292 46956
rect 26236 46734 26238 46786
rect 26290 46734 26292 46786
rect 26236 46340 26292 46734
rect 26236 46274 26292 46284
rect 26348 46116 26404 50372
rect 26460 49924 26516 49934
rect 26460 49810 26516 49868
rect 26460 49758 26462 49810
rect 26514 49758 26516 49810
rect 26460 49588 26516 49758
rect 26460 49522 26516 49532
rect 26684 49364 26740 50988
rect 26684 49298 26740 49308
rect 26796 49252 26852 51100
rect 26796 49186 26852 49196
rect 27020 49026 27076 49038
rect 27020 48974 27022 49026
rect 27074 48974 27076 49026
rect 26684 48914 26740 48926
rect 26684 48862 26686 48914
rect 26738 48862 26740 48914
rect 26684 48692 26740 48862
rect 26684 48626 26740 48636
rect 26348 46050 26404 46060
rect 26460 48356 26516 48366
rect 26460 45892 26516 48300
rect 26572 48132 26628 48142
rect 26572 48038 26628 48076
rect 27020 47460 27076 48974
rect 26796 47458 27076 47460
rect 26796 47406 27022 47458
rect 27074 47406 27076 47458
rect 26796 47404 27076 47406
rect 26684 47348 26740 47358
rect 26684 47124 26740 47292
rect 26684 47058 26740 47068
rect 26796 46900 26852 47404
rect 27020 47394 27076 47404
rect 26796 46834 26852 46844
rect 26684 46450 26740 46462
rect 26684 46398 26686 46450
rect 26738 46398 26740 46450
rect 26684 46004 26740 46398
rect 26684 45948 27076 46004
rect 26124 44482 26180 44492
rect 26236 45836 26516 45892
rect 25788 41134 25790 41186
rect 25842 41134 25844 41186
rect 25676 39396 25732 39406
rect 25676 39060 25732 39340
rect 25676 38994 25732 39004
rect 25452 37380 25508 38444
rect 25452 37314 25508 37324
rect 25676 37268 25732 37278
rect 25676 37174 25732 37212
rect 25564 37044 25620 37054
rect 25340 34738 25396 34748
rect 25452 36932 25508 36942
rect 25452 36482 25508 36876
rect 25564 36706 25620 36988
rect 25564 36654 25566 36706
rect 25618 36654 25620 36706
rect 25564 36642 25620 36654
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 25340 34132 25396 34142
rect 25116 34130 25396 34132
rect 25116 34078 25342 34130
rect 25394 34078 25396 34130
rect 25116 34076 25396 34078
rect 25340 34066 25396 34076
rect 25452 34020 25508 36430
rect 25564 35476 25620 35486
rect 25564 35382 25620 35420
rect 25676 35026 25732 35038
rect 25676 34974 25678 35026
rect 25730 34974 25732 35026
rect 25676 34916 25732 34974
rect 25676 34850 25732 34860
rect 25564 34020 25620 34030
rect 25452 34018 25620 34020
rect 25452 33966 25566 34018
rect 25618 33966 25620 34018
rect 25452 33964 25620 33966
rect 25564 33954 25620 33964
rect 24780 33852 24948 33908
rect 24332 33730 24388 33740
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 23884 33394 23940 33404
rect 24220 33012 24276 33022
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 24220 32788 24276 32956
rect 24108 32732 24276 32788
rect 23884 32562 23940 32574
rect 23884 32510 23886 32562
rect 23938 32510 23940 32562
rect 23884 32116 23940 32510
rect 24108 32562 24164 32732
rect 24444 32564 24500 32574
rect 24108 32510 24110 32562
rect 24162 32510 24164 32562
rect 24108 32498 24164 32510
rect 24332 32562 24500 32564
rect 24332 32510 24446 32562
rect 24498 32510 24500 32562
rect 24332 32508 24500 32510
rect 23884 32050 23940 32060
rect 23884 31780 23940 31790
rect 23884 31686 23940 31724
rect 23804 31388 24068 31398
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23660 29652 23716 31276
rect 23884 30996 23940 31006
rect 23884 30902 23940 30940
rect 24108 30996 24164 31006
rect 24108 30994 24276 30996
rect 24108 30942 24110 30994
rect 24162 30942 24276 30994
rect 24108 30940 24276 30942
rect 24108 30930 24164 30940
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 23660 29596 23828 29652
rect 23660 29092 23716 29102
rect 23660 28756 23716 29036
rect 23660 28642 23716 28700
rect 23660 28590 23662 28642
rect 23714 28590 23716 28642
rect 23660 28578 23716 28590
rect 23772 28420 23828 29596
rect 23996 29540 24052 29550
rect 23996 29446 24052 29484
rect 23660 28364 23828 28420
rect 23660 27076 23716 28364
rect 24220 28308 24276 30940
rect 24332 30212 24388 32508
rect 24444 32498 24500 32508
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24556 32004 24612 32014
rect 24556 31220 24612 31948
rect 24668 31668 24724 31678
rect 24668 31574 24724 31612
rect 24556 30994 24612 31164
rect 24556 30942 24558 30994
rect 24610 30942 24612 30994
rect 24556 30930 24612 30942
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 24332 30146 24388 30156
rect 24444 29316 24500 29326
rect 24332 29260 24444 29316
rect 24332 28532 24388 29260
rect 24444 29222 24500 29260
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 24332 28466 24388 28476
rect 24892 28532 24948 33852
rect 25116 33572 25172 33582
rect 25116 33348 25172 33516
rect 25116 33282 25172 33292
rect 25452 33124 25508 33134
rect 25004 33012 25060 33022
rect 25004 32228 25060 32956
rect 25340 33012 25396 33022
rect 25340 32562 25396 32956
rect 25340 32510 25342 32562
rect 25394 32510 25396 32562
rect 25004 32162 25060 32172
rect 25116 32338 25172 32350
rect 25116 32286 25118 32338
rect 25170 32286 25172 32338
rect 25004 31780 25060 31790
rect 25116 31780 25172 32286
rect 25228 31892 25284 31902
rect 25228 31798 25284 31836
rect 25004 31778 25172 31780
rect 25004 31726 25006 31778
rect 25058 31726 25172 31778
rect 25004 31724 25172 31726
rect 25004 31714 25060 31724
rect 25228 30996 25284 31006
rect 25228 30902 25284 30940
rect 25116 30884 25172 30894
rect 25116 30790 25172 30828
rect 25116 29092 25172 29102
rect 25116 28756 25172 29036
rect 25116 28690 25172 28700
rect 24892 28466 24948 28476
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24220 28242 24276 28252
rect 25340 28198 25396 32510
rect 25452 30212 25508 33068
rect 25676 32562 25732 32574
rect 25676 32510 25678 32562
rect 25730 32510 25732 32562
rect 25676 32004 25732 32510
rect 25676 31938 25732 31948
rect 25564 31890 25620 31902
rect 25564 31838 25566 31890
rect 25618 31838 25620 31890
rect 25564 30884 25620 31838
rect 25564 30818 25620 30828
rect 25676 30994 25732 31006
rect 25676 30942 25678 30994
rect 25730 30942 25732 30994
rect 25676 30324 25732 30942
rect 25676 30258 25732 30268
rect 25452 30146 25508 30156
rect 25676 30100 25732 30110
rect 25676 30006 25732 30044
rect 23804 28186 24068 28196
rect 24892 28142 25396 28198
rect 25564 29202 25620 29214
rect 25564 29150 25566 29202
rect 25618 29150 25620 29202
rect 24780 28084 24836 28094
rect 24220 27860 24276 27870
rect 24220 27766 24276 27804
rect 24780 27858 24836 28028
rect 24780 27806 24782 27858
rect 24834 27806 24836 27858
rect 23884 27746 23940 27758
rect 23884 27694 23886 27746
rect 23938 27694 23940 27746
rect 23884 27412 23940 27694
rect 24780 27748 24836 27806
rect 24780 27682 24836 27692
rect 24892 27746 24948 28142
rect 25564 27858 25620 29150
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25564 27794 25620 27806
rect 25676 28868 25732 28878
rect 24892 27694 24894 27746
rect 24946 27694 24948 27746
rect 24892 27682 24948 27694
rect 23884 27346 23940 27356
rect 24220 27524 24276 27534
rect 24892 27524 24948 27534
rect 23772 27076 23828 27086
rect 23660 27074 23828 27076
rect 23660 27022 23774 27074
rect 23826 27022 23828 27074
rect 23660 27020 23828 27022
rect 23660 26964 23716 27020
rect 23772 27010 23828 27020
rect 23660 26898 23716 26908
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 24220 26628 24276 27468
rect 24464 27468 24728 27478
rect 24332 27412 24388 27422
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24332 27300 24388 27356
rect 24892 27300 24948 27468
rect 24332 27244 24948 27300
rect 25116 27300 25172 27310
rect 25004 27188 25060 27198
rect 25004 26628 25060 27132
rect 25116 26852 25172 27244
rect 25116 26786 25172 26796
rect 25564 27076 25620 27086
rect 25004 26572 25396 26628
rect 24220 26562 24276 26572
rect 24332 26290 24388 26302
rect 24332 26238 24334 26290
rect 24386 26238 24388 26290
rect 24220 26180 24276 26190
rect 24332 26180 24388 26238
rect 24276 26124 24388 26180
rect 24444 26180 24500 26190
rect 24220 26114 24276 26124
rect 24444 26068 24500 26124
rect 25004 26180 25060 26190
rect 25004 26086 25060 26124
rect 24332 26012 24500 26068
rect 24892 26066 24948 26078
rect 24892 26014 24894 26066
rect 24946 26014 24948 26066
rect 24332 25844 24388 26012
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24332 25778 24388 25788
rect 24780 25732 24836 25742
rect 24892 25732 24948 26014
rect 24892 25676 25172 25732
rect 24780 25638 24836 25676
rect 23660 25508 23716 25518
rect 23548 25506 23716 25508
rect 23548 25454 23662 25506
rect 23714 25454 23716 25506
rect 23548 25452 23716 25454
rect 23548 25060 23604 25070
rect 23548 24276 23604 25004
rect 23548 24210 23604 24220
rect 22764 21026 22932 21028
rect 22764 20974 22766 21026
rect 22818 20974 22932 21026
rect 22764 20972 22932 20974
rect 22988 21756 23268 21812
rect 23324 22988 23492 23044
rect 23548 23044 23604 23054
rect 22764 20962 22820 20972
rect 22316 20692 22372 20702
rect 22316 20598 22372 20636
rect 22204 20580 22260 20590
rect 22204 16770 22260 20524
rect 22652 20580 22708 20590
rect 22652 20130 22708 20524
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22652 20066 22708 20078
rect 22428 20020 22484 20030
rect 22204 16718 22206 16770
rect 22258 16718 22260 16770
rect 22204 16660 22260 16718
rect 22204 16594 22260 16604
rect 22316 19908 22372 19918
rect 22316 19234 22372 19852
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 22092 16380 22260 16436
rect 22092 14530 22148 14542
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 14420 22148 14478
rect 22092 14354 22148 14364
rect 22092 13634 22148 13646
rect 22092 13582 22094 13634
rect 22146 13582 22148 13634
rect 22092 13524 22148 13582
rect 22092 13458 22148 13468
rect 21980 12236 22148 12292
rect 21980 12068 22036 12078
rect 21980 11974 22036 12012
rect 21756 11106 21812 11116
rect 21980 11844 22036 11854
rect 21420 10386 21588 10388
rect 21420 10334 21422 10386
rect 21474 10334 21588 10386
rect 21420 10332 21588 10334
rect 21868 10948 21924 10958
rect 21420 8036 21476 10332
rect 21868 10052 21924 10892
rect 21868 9986 21924 9996
rect 21532 9940 21588 9950
rect 21532 8258 21588 9884
rect 21532 8206 21534 8258
rect 21586 8206 21588 8258
rect 21532 8194 21588 8206
rect 21756 9940 21812 9950
rect 21756 8820 21812 9884
rect 21868 8820 21924 8830
rect 21756 8818 21924 8820
rect 21756 8766 21870 8818
rect 21922 8766 21924 8818
rect 21756 8764 21924 8766
rect 21420 7980 21588 8036
rect 21420 7476 21476 7486
rect 21028 7420 21252 7476
rect 21308 7474 21476 7476
rect 21308 7422 21422 7474
rect 21474 7422 21476 7474
rect 21308 7420 21476 7422
rect 20972 7382 21028 7420
rect 20860 6690 20916 7084
rect 20860 6638 20862 6690
rect 20914 6638 20916 6690
rect 20860 6626 20916 6638
rect 21196 6690 21252 7420
rect 21420 7410 21476 7420
rect 21532 7252 21588 7980
rect 21196 6638 21198 6690
rect 21250 6638 21252 6690
rect 21196 6626 21252 6638
rect 21420 7196 21588 7252
rect 21644 7252 21700 7262
rect 20412 5292 20468 5964
rect 20748 5908 20804 5918
rect 20748 5906 21364 5908
rect 20748 5854 20750 5906
rect 20802 5854 21364 5906
rect 20748 5852 21364 5854
rect 20748 5842 20804 5852
rect 20636 5684 20692 5694
rect 20188 5070 20190 5122
rect 20242 5070 20244 5122
rect 20188 5058 20244 5070
rect 20300 5236 20468 5292
rect 20524 5682 20692 5684
rect 20524 5630 20638 5682
rect 20690 5630 20692 5682
rect 20524 5628 20692 5630
rect 20524 5292 20580 5628
rect 20636 5618 20692 5628
rect 20860 5684 20916 5694
rect 20860 5682 21028 5684
rect 20860 5630 20862 5682
rect 20914 5630 21028 5682
rect 20860 5628 21028 5630
rect 20860 5618 20916 5628
rect 20972 5572 21028 5628
rect 20860 5460 20916 5470
rect 20524 5236 20692 5292
rect 20300 5124 20356 5236
rect 20300 5058 20356 5068
rect 20524 5124 20580 5162
rect 20636 5124 20692 5236
rect 20748 5234 20804 5246
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 5124 20804 5182
rect 20636 5068 20804 5124
rect 20524 5058 20580 5068
rect 19964 4844 20132 4900
rect 19852 4286 19854 4338
rect 19906 4286 19908 4338
rect 19852 4274 19908 4286
rect 19964 4340 20020 4350
rect 19964 4246 20020 4284
rect 20076 4338 20132 4844
rect 20748 4676 20804 4686
rect 20748 4562 20804 4620
rect 20748 4510 20750 4562
rect 20802 4510 20804 4562
rect 20076 4286 20078 4338
rect 20130 4286 20132 4338
rect 20076 4274 20132 4286
rect 20636 4340 20692 4350
rect 20188 4116 20244 4126
rect 19852 3668 19908 3678
rect 19852 3574 19908 3612
rect 19964 2660 20020 2670
rect 19964 2566 20020 2604
rect 19852 2546 19908 2558
rect 19852 2494 19854 2546
rect 19906 2494 19908 2546
rect 19852 2436 19908 2494
rect 20076 2548 20132 2558
rect 20076 2454 20132 2492
rect 19852 2370 19908 2380
rect 19852 1988 19908 1998
rect 19852 1894 19908 1932
rect 19740 1708 20020 1764
rect 19180 1374 19182 1426
rect 19234 1374 19236 1426
rect 19180 1362 19236 1374
rect 19516 1428 19572 1438
rect 18732 1138 18788 1148
rect 18508 914 18564 924
rect 18396 700 18676 756
rect 18620 112 18676 700
rect 19068 420 19124 430
rect 19068 112 19124 364
rect 19516 112 19572 1372
rect 19964 112 20020 1708
rect 20188 1204 20244 4060
rect 20524 3556 20580 3566
rect 20636 3556 20692 4284
rect 20524 3554 20692 3556
rect 20524 3502 20526 3554
rect 20578 3502 20692 3554
rect 20524 3500 20692 3502
rect 20748 3554 20804 4510
rect 20860 3668 20916 5404
rect 20972 5236 21028 5516
rect 20972 5170 21028 5180
rect 21084 5682 21140 5694
rect 21084 5630 21086 5682
rect 21138 5630 21140 5682
rect 21084 4788 21140 5630
rect 21084 4722 21140 4732
rect 21308 4340 21364 5852
rect 21420 5796 21476 7196
rect 21644 7158 21700 7196
rect 21756 6580 21812 8764
rect 21868 8754 21924 8764
rect 21980 7476 22036 11788
rect 22092 7588 22148 12236
rect 22204 11732 22260 16380
rect 22316 16100 22372 19182
rect 22428 18450 22484 19964
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22428 18386 22484 18398
rect 22764 18116 22820 18126
rect 22316 16034 22372 16044
rect 22428 16884 22484 16894
rect 22428 16098 22484 16828
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22428 16034 22484 16046
rect 22764 15988 22820 18060
rect 22988 16884 23044 21756
rect 23100 21586 23156 21598
rect 23100 21534 23102 21586
rect 23154 21534 23156 21586
rect 23100 21364 23156 21534
rect 23100 20916 23156 21308
rect 23100 20850 23156 20860
rect 23212 20692 23268 20702
rect 23100 19908 23156 19918
rect 23100 19814 23156 19852
rect 23100 18564 23156 18574
rect 23212 18564 23268 20636
rect 23324 19796 23380 22988
rect 23548 22950 23604 22988
rect 23436 22036 23492 22046
rect 23436 20356 23492 21980
rect 23548 21476 23604 21486
rect 23548 21382 23604 21420
rect 23660 21028 23716 25452
rect 24556 25506 24612 25518
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 24444 25172 24500 25182
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 24444 24948 24500 25116
rect 23996 24892 24500 24948
rect 23996 24834 24052 24892
rect 23996 24782 23998 24834
rect 24050 24782 24052 24834
rect 23996 24770 24052 24782
rect 24444 24724 24500 24734
rect 24444 24610 24500 24668
rect 24444 24558 24446 24610
rect 24498 24558 24500 24610
rect 24444 24546 24500 24558
rect 24556 24612 24612 25454
rect 25004 25506 25060 25518
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 24556 24546 24612 24556
rect 24892 25394 24948 25406
rect 24892 25342 24894 25394
rect 24946 25342 24948 25394
rect 24464 24332 24728 24342
rect 24220 24276 24276 24286
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 23884 23940 23940 23950
rect 23884 23846 23940 23884
rect 23804 23548 24068 23558
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 24220 23492 24276 24220
rect 24556 24052 24612 24062
rect 24556 23828 24612 23996
rect 24556 23762 24612 23772
rect 24220 23426 24276 23436
rect 23884 23156 23940 23166
rect 23884 23062 23940 23100
rect 24220 23156 24276 23166
rect 24444 23156 24500 23166
rect 24220 22932 24276 23100
rect 24220 22866 24276 22876
rect 24332 23154 24500 23156
rect 24332 23102 24446 23154
rect 24498 23102 24500 23154
rect 24332 23100 24500 23102
rect 24332 22596 24388 23100
rect 24444 23090 24500 23100
rect 24892 23044 24948 25342
rect 25004 25396 25060 25454
rect 25004 25330 25060 25340
rect 25116 23380 25172 25676
rect 25228 25508 25284 25518
rect 25228 25414 25284 25452
rect 25116 23314 25172 23324
rect 25228 25172 25284 25182
rect 25004 23268 25060 23278
rect 25004 23154 25060 23212
rect 25228 23156 25284 25116
rect 25340 24724 25396 26572
rect 25564 24946 25620 27020
rect 25564 24894 25566 24946
rect 25618 24894 25620 24946
rect 25564 24882 25620 24894
rect 25340 24658 25396 24668
rect 25676 24164 25732 28812
rect 25452 24108 25732 24164
rect 25452 23548 25508 24108
rect 25004 23102 25006 23154
rect 25058 23102 25060 23154
rect 25004 23090 25060 23102
rect 25116 23100 25284 23156
rect 25340 23492 25508 23548
rect 25564 23826 25620 23838
rect 25564 23774 25566 23826
rect 25618 23774 25620 23826
rect 25564 23604 25620 23774
rect 25564 23538 25620 23548
rect 25676 23716 25732 23726
rect 24892 22978 24948 22988
rect 24556 22932 24612 22942
rect 24780 22932 24836 22942
rect 24556 22930 24780 22932
rect 24556 22878 24558 22930
rect 24610 22878 24780 22930
rect 24556 22876 24780 22878
rect 24556 22866 24612 22876
rect 24780 22866 24836 22876
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24332 22530 24388 22540
rect 24556 22036 24612 22046
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 24556 21588 24612 21980
rect 25116 21868 25172 23100
rect 25004 21812 25172 21868
rect 25228 22932 25284 22942
rect 24556 21522 24612 21532
rect 24780 21588 24836 21598
rect 24780 21494 24836 21532
rect 24892 21476 24948 21486
rect 23548 20972 23716 21028
rect 24332 21252 24388 21262
rect 24332 21028 24388 21196
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 24892 21028 24948 21420
rect 24332 20972 24948 21028
rect 23548 20468 23604 20972
rect 23660 20804 23716 20814
rect 23660 20580 23716 20748
rect 23884 20804 23940 20814
rect 23884 20710 23940 20748
rect 24556 20692 24612 20702
rect 23660 20524 24276 20580
rect 23548 20412 23716 20468
rect 23436 20290 23492 20300
rect 23436 20020 23492 20030
rect 23436 19926 23492 19964
rect 23324 19740 23492 19796
rect 23100 18562 23268 18564
rect 23100 18510 23102 18562
rect 23154 18510 23268 18562
rect 23100 18508 23268 18510
rect 23100 18340 23156 18508
rect 23100 18274 23156 18284
rect 22988 16818 23044 16828
rect 23324 16884 23380 16894
rect 23324 16790 23380 16828
rect 23324 16548 23380 16558
rect 23436 16548 23492 19740
rect 23380 16492 23492 16548
rect 23548 18226 23604 18238
rect 23548 18174 23550 18226
rect 23602 18174 23604 18226
rect 23548 18004 23604 18174
rect 23100 16212 23156 16222
rect 22764 15932 23044 15988
rect 22428 15540 22484 15550
rect 22428 15446 22484 15484
rect 22204 11666 22260 11676
rect 22316 14532 22372 14542
rect 22204 11508 22260 11518
rect 22204 11394 22260 11452
rect 22204 11342 22206 11394
rect 22258 11342 22260 11394
rect 22204 10948 22260 11342
rect 22204 10882 22260 10892
rect 22204 10724 22260 10734
rect 22204 9826 22260 10668
rect 22316 10500 22372 14476
rect 22764 13746 22820 15932
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22316 10434 22372 10444
rect 22428 12964 22484 12974
rect 22204 9774 22206 9826
rect 22258 9774 22260 9826
rect 22204 9762 22260 9774
rect 22316 9044 22372 9054
rect 22316 8950 22372 8988
rect 22316 8260 22372 8270
rect 22092 7532 22260 7588
rect 21980 7420 22148 7476
rect 21756 6514 21812 6524
rect 21868 6802 21924 6814
rect 21868 6750 21870 6802
rect 21922 6750 21924 6802
rect 21868 6130 21924 6750
rect 21980 6804 22036 6814
rect 21980 6690 22036 6748
rect 21980 6638 21982 6690
rect 22034 6638 22036 6690
rect 21980 6626 22036 6638
rect 21868 6078 21870 6130
rect 21922 6078 21924 6130
rect 21868 6066 21924 6078
rect 21420 5730 21476 5740
rect 21532 6018 21588 6030
rect 21532 5966 21534 6018
rect 21586 5966 21588 6018
rect 21420 5124 21476 5134
rect 21420 5030 21476 5068
rect 21532 4676 21588 5966
rect 21868 5908 21924 5918
rect 21644 5684 21700 5694
rect 21644 5682 21812 5684
rect 21644 5630 21646 5682
rect 21698 5630 21812 5682
rect 21644 5628 21812 5630
rect 21644 5618 21700 5628
rect 21756 5572 21812 5628
rect 21756 5506 21812 5516
rect 21532 4610 21588 4620
rect 21644 5460 21700 5470
rect 20972 4338 21364 4340
rect 20972 4286 21310 4338
rect 21362 4286 21364 4338
rect 20972 4284 21364 4286
rect 20972 3892 21028 4284
rect 21308 4274 21364 4284
rect 21532 4452 21588 4462
rect 21084 4116 21140 4126
rect 21084 4114 21252 4116
rect 21084 4062 21086 4114
rect 21138 4062 21252 4114
rect 21084 4060 21252 4062
rect 21084 4050 21140 4060
rect 20972 3836 21140 3892
rect 20972 3668 21028 3678
rect 20860 3666 21028 3668
rect 20860 3614 20974 3666
rect 21026 3614 21028 3666
rect 20860 3612 21028 3614
rect 21084 3668 21140 3836
rect 21196 3780 21252 4060
rect 21420 4114 21476 4126
rect 21420 4062 21422 4114
rect 21474 4062 21476 4114
rect 21196 3724 21364 3780
rect 21084 3612 21252 3668
rect 20972 3602 21028 3612
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20524 3490 20580 3500
rect 20748 3490 20804 3502
rect 21196 3554 21252 3612
rect 21196 3502 21198 3554
rect 21250 3502 21252 3554
rect 21196 3490 21252 3502
rect 20860 3444 20916 3454
rect 20300 2884 20356 2894
rect 20300 1986 20356 2828
rect 20860 2772 20916 3388
rect 21084 3444 21140 3454
rect 21308 3388 21364 3724
rect 21084 3350 21140 3388
rect 21196 3332 21364 3388
rect 21196 2996 21252 3332
rect 21084 2940 21252 2996
rect 20972 2772 21028 2782
rect 20860 2770 21028 2772
rect 20860 2718 20974 2770
rect 21026 2718 21028 2770
rect 20860 2716 21028 2718
rect 20972 2706 21028 2716
rect 20748 2658 20804 2670
rect 20748 2606 20750 2658
rect 20802 2606 20804 2658
rect 20748 2548 20804 2606
rect 21084 2548 21140 2940
rect 21196 2772 21252 2782
rect 21196 2678 21252 2716
rect 21308 2770 21364 2782
rect 21308 2718 21310 2770
rect 21362 2718 21364 2770
rect 20748 2492 21140 2548
rect 21196 2548 21252 2558
rect 20748 2436 20804 2492
rect 20748 2370 20804 2380
rect 20300 1934 20302 1986
rect 20354 1934 20356 1986
rect 20300 1922 20356 1934
rect 20412 1652 20468 1662
rect 20300 1204 20356 1214
rect 20188 1202 20356 1204
rect 20188 1150 20302 1202
rect 20354 1150 20356 1202
rect 20188 1148 20356 1150
rect 20300 1138 20356 1148
rect 20412 112 20468 1596
rect 20860 1540 20916 1550
rect 20636 978 20692 990
rect 20636 926 20638 978
rect 20690 926 20692 978
rect 20636 532 20692 926
rect 20636 466 20692 476
rect 20860 112 20916 1484
rect 21084 1204 21140 1214
rect 21196 1204 21252 2492
rect 21308 2324 21364 2718
rect 21420 2772 21476 4062
rect 21532 3332 21588 4396
rect 21644 4338 21700 5404
rect 21644 4286 21646 4338
rect 21698 4286 21700 4338
rect 21644 4274 21700 4286
rect 21756 4788 21812 4798
rect 21644 3780 21700 3790
rect 21644 3686 21700 3724
rect 21756 3668 21812 4732
rect 21756 3574 21812 3612
rect 21868 3388 21924 5852
rect 21980 5124 22036 5134
rect 22092 5124 22148 7420
rect 21980 5122 22148 5124
rect 21980 5070 21982 5122
rect 22034 5070 22148 5122
rect 21980 5068 22148 5070
rect 21980 5058 22036 5068
rect 22092 4340 22148 4350
rect 22092 4246 22148 4284
rect 22204 3892 22260 7532
rect 22316 7474 22372 8204
rect 22316 7422 22318 7474
rect 22370 7422 22372 7474
rect 22316 6692 22372 7422
rect 22428 7476 22484 12908
rect 22540 12962 22596 12974
rect 22540 12910 22542 12962
rect 22594 12910 22596 12962
rect 22540 12068 22596 12910
rect 22652 12964 22708 12974
rect 22652 12516 22708 12908
rect 22652 12450 22708 12460
rect 22540 12002 22596 12012
rect 22764 11844 22820 13694
rect 22764 11778 22820 11788
rect 22876 15764 22932 15774
rect 22876 11620 22932 15708
rect 22988 15652 23044 15932
rect 23100 15764 23156 16156
rect 23100 15698 23156 15708
rect 23212 16098 23268 16110
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 22988 15586 23044 15596
rect 23212 15204 23268 16046
rect 23212 15138 23268 15148
rect 23100 13636 23156 13646
rect 22988 13188 23044 13198
rect 22988 13074 23044 13132
rect 23100 13186 23156 13580
rect 23100 13134 23102 13186
rect 23154 13134 23156 13186
rect 23100 13122 23156 13134
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 22988 13010 23044 13022
rect 23212 13076 23268 13086
rect 23212 12982 23268 13020
rect 23100 12180 23156 12190
rect 23100 12086 23156 12124
rect 23324 12068 23380 16492
rect 23548 16212 23604 17948
rect 23548 16146 23604 16156
rect 23436 15876 23492 15886
rect 23436 13076 23492 15820
rect 23436 13010 23492 13020
rect 23548 15764 23604 15774
rect 23548 12292 23604 15708
rect 23660 13748 23716 20412
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 24220 20356 24276 20524
rect 24556 20468 24612 20636
rect 24780 20692 24836 20972
rect 24780 20626 24836 20636
rect 24892 20802 24948 20814
rect 24892 20750 24894 20802
rect 24946 20750 24948 20802
rect 24892 20580 24948 20750
rect 24892 20514 24948 20524
rect 24556 20402 24612 20412
rect 24220 20132 24276 20300
rect 23996 20076 24276 20132
rect 23996 20018 24052 20076
rect 23996 19966 23998 20018
rect 24050 19966 24052 20018
rect 23996 19954 24052 19966
rect 24780 20020 24836 20030
rect 24780 20018 24948 20020
rect 24780 19966 24782 20018
rect 24834 19966 24948 20018
rect 24780 19964 24948 19966
rect 24780 19954 24836 19964
rect 24220 19908 24276 19918
rect 24108 19852 24220 19908
rect 24108 19794 24164 19852
rect 24220 19842 24276 19852
rect 24108 19742 24110 19794
rect 24162 19742 24164 19794
rect 24108 19572 24164 19742
rect 24108 19506 24164 19516
rect 24220 19684 24276 19694
rect 24220 18900 24276 19628
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 24892 19348 24948 19964
rect 24668 19292 24948 19348
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24220 18834 24276 18844
rect 24332 19236 24388 19246
rect 23804 18778 24068 18788
rect 24220 17444 24276 17454
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 23772 17108 23828 17118
rect 23772 16994 23828 17052
rect 23772 16942 23774 16994
rect 23826 16942 23828 16994
rect 23772 16930 23828 16942
rect 24108 16884 24164 16894
rect 24108 16790 24164 16828
rect 24108 16436 24164 16446
rect 24108 15988 24164 16380
rect 24108 15922 24164 15932
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 23660 13746 23828 13748
rect 23660 13694 23662 13746
rect 23714 13694 23828 13746
rect 23660 13692 23828 13694
rect 23660 13682 23716 13692
rect 23660 13300 23716 13310
rect 23660 12404 23716 13244
rect 23772 13188 23828 13692
rect 23772 13122 23828 13132
rect 24220 12628 24276 17388
rect 24332 15316 24388 19180
rect 24668 18674 24724 19292
rect 24668 18622 24670 18674
rect 24722 18622 24724 18674
rect 24668 18610 24724 18622
rect 24892 19124 24948 19134
rect 25004 19124 25060 21812
rect 25116 20580 25172 20590
rect 25116 19908 25172 20524
rect 25116 19842 25172 19852
rect 24892 19122 25060 19124
rect 24892 19070 24894 19122
rect 24946 19070 25060 19122
rect 24892 19068 25060 19070
rect 24892 18452 24948 19068
rect 24892 18386 24948 18396
rect 25004 18788 25060 18798
rect 24892 18116 24948 18126
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 24892 17892 24948 18060
rect 24556 17836 24948 17892
rect 24556 16882 24612 17836
rect 24556 16830 24558 16882
rect 24610 16830 24612 16882
rect 24556 16818 24612 16830
rect 24668 17442 24724 17454
rect 24668 17390 24670 17442
rect 24722 17390 24724 17442
rect 24668 16884 24724 17390
rect 24668 16818 24724 16828
rect 24780 17332 24836 17342
rect 24780 16770 24836 17276
rect 24780 16718 24782 16770
rect 24834 16718 24836 16770
rect 24780 16706 24836 16718
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 24892 16212 24948 16222
rect 24444 15316 24500 15326
rect 24332 15314 24500 15316
rect 24332 15262 24446 15314
rect 24498 15262 24500 15314
rect 24332 15260 24500 15262
rect 24444 15148 24500 15260
rect 24332 15092 24500 15148
rect 24892 15202 24948 16156
rect 24892 15150 24894 15202
rect 24946 15150 24948 15202
rect 24892 15138 24948 15150
rect 24332 14420 24388 15092
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 25004 14756 25060 18732
rect 25116 17668 25172 17678
rect 25116 15876 25172 17612
rect 25228 17332 25284 22876
rect 25340 21476 25396 23492
rect 25676 23154 25732 23660
rect 25676 23102 25678 23154
rect 25730 23102 25732 23154
rect 25676 23090 25732 23102
rect 25788 22708 25844 41134
rect 25900 41132 26068 41188
rect 26124 43988 26180 43998
rect 25900 28378 25956 41132
rect 26124 41076 26180 43932
rect 26236 41636 26292 45836
rect 26908 45778 26964 45790
rect 26908 45726 26910 45778
rect 26962 45726 26964 45778
rect 26460 45668 26516 45678
rect 26460 45666 26852 45668
rect 26460 45614 26462 45666
rect 26514 45614 26852 45666
rect 26460 45612 26852 45614
rect 26460 45602 26516 45612
rect 26348 45106 26404 45118
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26348 43540 26404 45054
rect 26348 43446 26404 43484
rect 26460 44098 26516 44110
rect 26460 44046 26462 44098
rect 26514 44046 26516 44098
rect 26460 43092 26516 44046
rect 26460 43026 26516 43036
rect 26348 42756 26404 42766
rect 26348 42084 26404 42700
rect 26796 42754 26852 45612
rect 26908 44210 26964 45726
rect 27020 45108 27076 45948
rect 27020 45042 27076 45052
rect 26908 44158 26910 44210
rect 26962 44158 26964 44210
rect 26908 43764 26964 44158
rect 26908 43698 26964 43708
rect 26796 42702 26798 42754
rect 26850 42702 26852 42754
rect 26796 42690 26852 42702
rect 26460 42642 26516 42654
rect 26460 42590 26462 42642
rect 26514 42590 26516 42642
rect 26460 42308 26516 42590
rect 26460 42242 26516 42252
rect 26348 42028 26516 42084
rect 26236 41570 26292 41580
rect 26348 41860 26404 41870
rect 26348 41410 26404 41804
rect 26348 41358 26350 41410
rect 26402 41358 26404 41410
rect 26348 41346 26404 41358
rect 26236 41298 26292 41310
rect 26236 41246 26238 41298
rect 26290 41246 26292 41298
rect 26236 41188 26292 41246
rect 26236 41122 26292 41132
rect 26012 41020 26180 41076
rect 26012 38050 26068 41020
rect 26236 40964 26292 40974
rect 26236 40404 26292 40908
rect 26236 40310 26292 40348
rect 26460 39844 26516 42028
rect 27020 41746 27076 41758
rect 27020 41694 27022 41746
rect 27074 41694 27076 41746
rect 26348 39788 26516 39844
rect 26572 41300 26628 41310
rect 26236 39732 26292 39742
rect 26236 39172 26292 39676
rect 26236 39106 26292 39116
rect 26236 38836 26292 38846
rect 26236 38742 26292 38780
rect 26012 37998 26014 38050
rect 26066 37998 26068 38050
rect 26012 37604 26068 37998
rect 26012 37538 26068 37548
rect 26236 38388 26292 38398
rect 26012 37156 26068 37166
rect 26012 36594 26068 37100
rect 26012 36542 26014 36594
rect 26066 36542 26068 36594
rect 26012 36530 26068 36542
rect 26124 35700 26180 35710
rect 26124 35606 26180 35644
rect 26012 35588 26068 35598
rect 26012 34130 26068 35532
rect 26012 34078 26014 34130
rect 26066 34078 26068 34130
rect 26012 34066 26068 34078
rect 26124 33348 26180 33358
rect 26124 32674 26180 33292
rect 26124 32622 26126 32674
rect 26178 32622 26180 32674
rect 26012 31668 26068 31678
rect 26012 30322 26068 31612
rect 26124 31444 26180 32622
rect 26236 32116 26292 38332
rect 26348 37268 26404 39788
rect 26460 39508 26516 39518
rect 26572 39508 26628 41244
rect 26684 40180 26740 40190
rect 26684 40086 26740 40124
rect 26796 39956 26852 39966
rect 26684 39508 26740 39518
rect 26572 39452 26684 39508
rect 26460 39414 26516 39452
rect 26684 39442 26740 39452
rect 26460 39172 26516 39182
rect 26460 38274 26516 39116
rect 26684 39172 26740 39182
rect 26684 38722 26740 39116
rect 26684 38670 26686 38722
rect 26738 38670 26740 38722
rect 26684 38658 26740 38670
rect 26460 38222 26462 38274
rect 26514 38222 26516 38274
rect 26460 38210 26516 38222
rect 26460 37268 26516 37278
rect 26348 37266 26516 37268
rect 26348 37214 26462 37266
rect 26514 37214 26516 37266
rect 26348 37212 26516 37214
rect 26460 37156 26516 37212
rect 26460 37090 26516 37100
rect 26796 36484 26852 39900
rect 26908 39620 26964 39630
rect 27020 39620 27076 41694
rect 26908 39618 27076 39620
rect 26908 39566 26910 39618
rect 26962 39566 27076 39618
rect 26908 39564 27076 39566
rect 26908 39554 26964 39564
rect 26796 36390 26852 36428
rect 26908 37716 26964 37726
rect 26684 36148 26740 36158
rect 26684 35586 26740 36092
rect 26684 35534 26686 35586
rect 26738 35534 26740 35586
rect 26684 35522 26740 35534
rect 26796 34690 26852 34702
rect 26796 34638 26798 34690
rect 26850 34638 26852 34690
rect 26684 34244 26740 34254
rect 26684 34130 26740 34188
rect 26684 34078 26686 34130
rect 26738 34078 26740 34130
rect 26684 34066 26740 34078
rect 26796 34132 26852 34638
rect 26796 34066 26852 34076
rect 26572 33236 26628 33246
rect 26236 32050 26292 32060
rect 26460 33234 26628 33236
rect 26460 33182 26574 33234
rect 26626 33182 26628 33234
rect 26460 33180 26628 33182
rect 26460 31668 26516 33180
rect 26572 33170 26628 33180
rect 26124 31378 26180 31388
rect 26348 31666 26516 31668
rect 26348 31614 26462 31666
rect 26514 31614 26516 31666
rect 26348 31612 26516 31614
rect 26124 31220 26180 31230
rect 26124 31106 26180 31164
rect 26124 31054 26126 31106
rect 26178 31054 26180 31106
rect 26124 31042 26180 31054
rect 26348 30884 26404 31612
rect 26460 31602 26516 31612
rect 26572 32116 26628 32126
rect 26012 30270 26014 30322
rect 26066 30270 26068 30322
rect 26012 28868 26068 30270
rect 26012 28802 26068 28812
rect 26124 30828 26404 30884
rect 26012 28532 26068 28570
rect 26012 28466 26068 28476
rect 25900 28322 26068 28378
rect 25900 27858 25956 27870
rect 25900 27806 25902 27858
rect 25954 27806 25956 27858
rect 25900 25732 25956 27806
rect 25900 25666 25956 25676
rect 25900 23944 25956 23956
rect 25900 23940 25902 23944
rect 25954 23940 25956 23944
rect 25900 23852 25956 23884
rect 25788 22642 25844 22652
rect 26012 22372 26068 28322
rect 26124 27188 26180 30828
rect 26236 29540 26292 29550
rect 26236 29446 26292 29484
rect 26572 29314 26628 32060
rect 26908 31948 26964 37660
rect 27132 37380 27188 53788
rect 27244 51940 27300 54012
rect 27356 53508 27412 55356
rect 27468 54292 27524 55804
rect 27580 55524 27636 57344
rect 27804 56308 27860 56318
rect 27580 55458 27636 55468
rect 27692 55636 27748 55646
rect 27580 55298 27636 55310
rect 27580 55246 27582 55298
rect 27634 55246 27636 55298
rect 27580 54516 27636 55246
rect 27580 54450 27636 54460
rect 27468 53844 27524 54236
rect 27468 53778 27524 53788
rect 27580 54290 27636 54302
rect 27580 54238 27582 54290
rect 27634 54238 27636 54290
rect 27356 53442 27412 53452
rect 27356 53060 27412 53070
rect 27356 52966 27412 53004
rect 27580 52836 27636 54238
rect 27692 53620 27748 55580
rect 27804 54068 27860 56252
rect 27916 55860 27972 55870
rect 27916 55766 27972 55804
rect 28028 55524 28084 57344
rect 28252 56644 28308 56654
rect 28028 55458 28084 55468
rect 28140 56196 28196 56206
rect 27916 55410 27972 55422
rect 27916 55358 27918 55410
rect 27970 55358 27972 55410
rect 27916 54516 27972 55358
rect 28140 55412 28196 56140
rect 28252 55970 28308 56588
rect 28252 55918 28254 55970
rect 28306 55918 28308 55970
rect 28252 55906 28308 55918
rect 28252 55412 28308 55422
rect 28140 55410 28308 55412
rect 28140 55358 28254 55410
rect 28306 55358 28308 55410
rect 28140 55356 28308 55358
rect 28252 55346 28308 55356
rect 28476 54628 28532 57344
rect 28700 56082 28756 56094
rect 28924 56084 28980 57344
rect 28700 56030 28702 56082
rect 28754 56030 28756 56082
rect 28588 55298 28644 55310
rect 28588 55246 28590 55298
rect 28642 55246 28644 55298
rect 28588 54740 28644 55246
rect 28588 54674 28644 54684
rect 28364 54572 28532 54628
rect 28700 54628 28756 56030
rect 28812 56028 28980 56084
rect 28812 55188 28868 56028
rect 28924 55860 28980 55870
rect 29260 55860 29316 55870
rect 28924 55858 29316 55860
rect 28924 55806 28926 55858
rect 28978 55806 29262 55858
rect 29314 55806 29316 55858
rect 28924 55804 29316 55806
rect 28924 55794 28980 55804
rect 29260 55794 29316 55804
rect 29260 55636 29316 55646
rect 29036 55412 29092 55422
rect 29036 55410 29204 55412
rect 29036 55358 29038 55410
rect 29090 55358 29204 55410
rect 29036 55356 29204 55358
rect 29036 55346 29092 55356
rect 28812 55122 28868 55132
rect 28924 55298 28980 55310
rect 28924 55246 28926 55298
rect 28978 55246 28980 55298
rect 27916 54460 28196 54516
rect 27916 54292 27972 54302
rect 27916 54198 27972 54236
rect 27804 54002 27860 54012
rect 28028 53842 28084 53854
rect 28028 53790 28030 53842
rect 28082 53790 28084 53842
rect 27804 53732 27860 53742
rect 27804 53638 27860 53676
rect 27692 53554 27748 53564
rect 27580 52770 27636 52780
rect 27916 53284 27972 53294
rect 27244 51874 27300 51884
rect 27356 52612 27412 52622
rect 27356 49028 27412 52556
rect 27804 52500 27860 52510
rect 27692 51492 27748 51502
rect 27692 51378 27748 51436
rect 27692 51326 27694 51378
rect 27746 51326 27748 51378
rect 27692 51156 27748 51326
rect 27692 51090 27748 51100
rect 27804 51044 27860 52444
rect 27804 50978 27860 50988
rect 27916 52162 27972 53228
rect 27916 52110 27918 52162
rect 27970 52110 27972 52162
rect 27580 50932 27636 50942
rect 27468 50708 27524 50718
rect 27468 49028 27524 50652
rect 27580 50594 27636 50876
rect 27580 50542 27582 50594
rect 27634 50542 27636 50594
rect 27580 50530 27636 50542
rect 27692 49140 27748 49150
rect 27692 49046 27748 49084
rect 27580 49028 27636 49038
rect 27468 49026 27636 49028
rect 27468 48974 27582 49026
rect 27634 48974 27636 49026
rect 27468 48972 27636 48974
rect 27356 48962 27412 48972
rect 27580 48916 27636 48972
rect 27580 48850 27636 48860
rect 27692 48804 27748 48814
rect 27244 48020 27300 48030
rect 27244 45890 27300 47964
rect 27692 47682 27748 48748
rect 27692 47630 27694 47682
rect 27746 47630 27748 47682
rect 27692 47618 27748 47630
rect 27804 48018 27860 48030
rect 27804 47966 27806 48018
rect 27858 47966 27860 48018
rect 27804 47572 27860 47966
rect 27804 47506 27860 47516
rect 27244 45838 27246 45890
rect 27298 45838 27300 45890
rect 27244 45826 27300 45838
rect 27356 47460 27412 47470
rect 27356 45106 27412 47404
rect 27580 47460 27636 47470
rect 27580 47366 27636 47404
rect 27916 47068 27972 52110
rect 28028 49588 28084 53790
rect 28028 49522 28084 49532
rect 28140 48132 28196 54460
rect 28252 52948 28308 52958
rect 28252 49476 28308 52892
rect 28252 49410 28308 49420
rect 28364 49252 28420 54572
rect 28700 54562 28756 54572
rect 28924 54516 28980 55246
rect 28924 54450 28980 54460
rect 29036 55074 29092 55086
rect 29036 55022 29038 55074
rect 29090 55022 29092 55074
rect 28476 54402 28532 54414
rect 28476 54350 28478 54402
rect 28530 54350 28532 54402
rect 28476 54180 28532 54350
rect 28588 54292 28644 54302
rect 28588 54290 28756 54292
rect 28588 54238 28590 54290
rect 28642 54238 28756 54290
rect 28588 54236 28756 54238
rect 28588 54226 28644 54236
rect 28476 54114 28532 54124
rect 28476 53956 28532 53966
rect 28476 53284 28532 53900
rect 28476 53218 28532 53228
rect 28588 53618 28644 53630
rect 28588 53566 28590 53618
rect 28642 53566 28644 53618
rect 28588 53060 28644 53566
rect 28700 53396 28756 54236
rect 28700 53330 28756 53340
rect 28812 54290 28868 54302
rect 28812 54238 28814 54290
rect 28866 54238 28868 54290
rect 28588 52948 28644 53004
rect 28588 52892 28756 52948
rect 28588 52722 28644 52734
rect 28588 52670 28590 52722
rect 28642 52670 28644 52722
rect 28588 52164 28644 52670
rect 28700 52388 28756 52892
rect 28812 52388 28868 54238
rect 29036 54068 29092 55022
rect 29148 54964 29204 55356
rect 29148 54898 29204 54908
rect 29148 54740 29204 54750
rect 29148 54646 29204 54684
rect 29036 54012 29204 54068
rect 29036 53842 29092 53854
rect 29036 53790 29038 53842
rect 29090 53790 29092 53842
rect 29036 52724 29092 53790
rect 29036 52658 29092 52668
rect 28812 52332 29092 52388
rect 28700 52164 28756 52332
rect 28924 52164 28980 52174
rect 28700 52162 28980 52164
rect 28700 52110 28926 52162
rect 28978 52110 28980 52162
rect 28700 52108 28980 52110
rect 28588 51940 28644 52108
rect 28924 52098 28980 52108
rect 28588 51884 28980 51940
rect 28700 51604 28756 51614
rect 28700 51510 28756 51548
rect 28588 51492 28644 51502
rect 28588 51378 28644 51436
rect 28588 51326 28590 51378
rect 28642 51326 28644 51378
rect 28588 51314 28644 51326
rect 28700 51154 28756 51166
rect 28700 51102 28702 51154
rect 28754 51102 28756 51154
rect 28588 51044 28644 51054
rect 28588 50706 28644 50988
rect 28588 50654 28590 50706
rect 28642 50654 28644 50706
rect 28588 50642 28644 50654
rect 28700 50260 28756 51102
rect 28924 50594 28980 51884
rect 29036 51716 29092 52332
rect 29148 51716 29204 54012
rect 29260 53732 29316 55580
rect 29372 55524 29428 57344
rect 29372 55458 29428 55468
rect 29484 56196 29540 56206
rect 29484 55412 29540 56140
rect 29596 55860 29652 55870
rect 29596 55766 29652 55804
rect 29820 55748 29876 57344
rect 30268 56084 30324 57344
rect 30604 57092 30660 57102
rect 30268 56018 30324 56028
rect 30380 56532 30436 56542
rect 29932 55972 29988 55982
rect 29932 55878 29988 55916
rect 30268 55860 30324 55870
rect 30268 55766 30324 55804
rect 29820 55682 29876 55692
rect 29484 55346 29540 55356
rect 29820 55412 29876 55422
rect 29820 55318 29876 55356
rect 29596 55300 29652 55310
rect 29596 55206 29652 55244
rect 30268 55298 30324 55310
rect 30268 55246 30270 55298
rect 30322 55246 30324 55298
rect 30268 54740 30324 55246
rect 30268 54674 30324 54684
rect 29260 53666 29316 53676
rect 29372 54628 29428 54638
rect 29372 52948 29428 54572
rect 29372 52882 29428 52892
rect 29484 54514 29540 54526
rect 29484 54462 29486 54514
rect 29538 54462 29540 54514
rect 29484 52500 29540 54462
rect 30156 54514 30212 54526
rect 30156 54462 30158 54514
rect 30210 54462 30212 54514
rect 30044 54404 30100 54414
rect 29484 52434 29540 52444
rect 29596 54402 30100 54404
rect 29596 54350 30046 54402
rect 30098 54350 30100 54402
rect 29596 54348 30100 54350
rect 29484 52274 29540 52286
rect 29484 52222 29486 52274
rect 29538 52222 29540 52274
rect 29372 52164 29428 52174
rect 29148 51660 29316 51716
rect 29036 51650 29092 51660
rect 29148 51268 29204 51278
rect 29148 51174 29204 51212
rect 29260 51044 29316 51660
rect 29372 51380 29428 52108
rect 29484 52052 29540 52222
rect 29484 51986 29540 51996
rect 29484 51380 29540 51390
rect 29372 51378 29540 51380
rect 29372 51326 29486 51378
rect 29538 51326 29540 51378
rect 29372 51324 29540 51326
rect 29484 51314 29540 51324
rect 29260 50978 29316 50988
rect 29484 51156 29540 51166
rect 28924 50542 28926 50594
rect 28978 50542 28980 50594
rect 28924 50530 28980 50542
rect 29372 50932 29428 50942
rect 29372 50594 29428 50876
rect 29372 50542 29374 50594
rect 29426 50542 29428 50594
rect 28700 50194 28756 50204
rect 28140 48066 28196 48076
rect 28252 49196 28420 49252
rect 28924 50036 28980 50046
rect 28252 47908 28308 49196
rect 27468 47012 27524 47022
rect 27468 45892 27524 46956
rect 27468 45826 27524 45836
rect 27580 47012 27972 47068
rect 28028 47852 28308 47908
rect 28364 49026 28420 49038
rect 28364 48974 28366 49026
rect 28418 48974 28420 49026
rect 27356 45054 27358 45106
rect 27410 45054 27412 45106
rect 27244 44324 27300 44334
rect 27244 44230 27300 44268
rect 27244 43540 27300 43550
rect 27356 43540 27412 45054
rect 27580 44772 27636 47012
rect 28028 46788 28084 47852
rect 28140 47684 28196 47694
rect 28140 47570 28196 47628
rect 28140 47518 28142 47570
rect 28194 47518 28196 47570
rect 28140 47506 28196 47518
rect 28252 47572 28308 47582
rect 28252 47012 28308 47516
rect 28364 47458 28420 48974
rect 28364 47406 28366 47458
rect 28418 47406 28420 47458
rect 28364 47394 28420 47406
rect 28476 49028 28532 49038
rect 28700 49028 28756 49038
rect 28476 47068 28532 48972
rect 28140 46956 28308 47012
rect 28420 47012 28532 47068
rect 28588 49026 28756 49028
rect 28588 48974 28702 49026
rect 28754 48974 28756 49026
rect 28588 48972 28756 48974
rect 28140 46900 28196 46956
rect 28140 46834 28196 46844
rect 28420 46900 28476 47012
rect 28420 46834 28476 46844
rect 27692 46732 28084 46788
rect 27692 46116 27748 46732
rect 28588 46564 28644 48972
rect 28700 48962 28756 48972
rect 28700 47458 28756 47470
rect 28700 47406 28702 47458
rect 28754 47406 28756 47458
rect 28700 47348 28756 47406
rect 28700 47282 28756 47292
rect 28924 46900 28980 49980
rect 29036 48916 29092 48926
rect 29036 47012 29092 48860
rect 29372 48804 29428 50542
rect 29372 48738 29428 48748
rect 29484 47460 29540 51100
rect 29596 50818 29652 54348
rect 30044 54338 30100 54348
rect 30156 53954 30212 54462
rect 30156 53902 30158 53954
rect 30210 53902 30212 53954
rect 30156 53890 30212 53902
rect 29820 52948 29876 52958
rect 29596 50766 29598 50818
rect 29650 50766 29652 50818
rect 29596 50754 29652 50766
rect 29708 52722 29764 52734
rect 29708 52670 29710 52722
rect 29762 52670 29764 52722
rect 29708 49924 29764 52670
rect 29820 50708 29876 52892
rect 30268 52946 30324 52958
rect 30268 52894 30270 52946
rect 30322 52894 30324 52946
rect 30156 52500 30212 52510
rect 29820 50642 29876 50652
rect 29932 52388 29988 52398
rect 29708 49858 29764 49868
rect 29820 50372 29876 50382
rect 29820 49810 29876 50316
rect 29820 49758 29822 49810
rect 29874 49758 29876 49810
rect 29820 49746 29876 49758
rect 29596 49700 29652 49710
rect 29596 49606 29652 49644
rect 29708 49586 29764 49598
rect 29708 49534 29710 49586
rect 29762 49534 29764 49586
rect 29708 49252 29764 49534
rect 29708 49196 29876 49252
rect 29708 49026 29764 49038
rect 29708 48974 29710 49026
rect 29762 48974 29764 49026
rect 29708 48692 29764 48974
rect 29708 48626 29764 48636
rect 29820 47572 29876 49196
rect 29820 47506 29876 47516
rect 29708 47460 29764 47470
rect 29484 47404 29708 47460
rect 29708 47366 29764 47404
rect 29932 47236 29988 52332
rect 30044 51378 30100 51390
rect 30044 51326 30046 51378
rect 30098 51326 30100 51378
rect 30044 50596 30100 51326
rect 30156 51266 30212 52444
rect 30268 52164 30324 52894
rect 30268 52098 30324 52108
rect 30156 51214 30158 51266
rect 30210 51214 30212 51266
rect 30156 51202 30212 51214
rect 30380 50932 30436 56476
rect 30492 56196 30548 56206
rect 30492 55636 30548 56140
rect 30604 56082 30660 57036
rect 30604 56030 30606 56082
rect 30658 56030 30660 56082
rect 30604 56018 30660 56030
rect 30492 55580 30660 55636
rect 30492 55412 30548 55422
rect 30492 55318 30548 55356
rect 30604 52500 30660 55580
rect 30716 55524 30772 57344
rect 30940 55858 30996 55870
rect 30940 55806 30942 55858
rect 30994 55806 30996 55858
rect 30940 55748 30996 55806
rect 30940 55682 30996 55692
rect 31164 55524 31220 57344
rect 30716 55458 30772 55468
rect 31052 55468 31220 55524
rect 31388 56868 31444 56878
rect 30828 55410 30884 55422
rect 30828 55358 30830 55410
rect 30882 55358 30884 55410
rect 30828 55300 30884 55358
rect 30828 55234 30884 55244
rect 31052 55076 31108 55468
rect 31164 55300 31220 55310
rect 31164 55206 31220 55244
rect 30604 52434 30660 52444
rect 30716 55020 31108 55076
rect 30380 50866 30436 50876
rect 30604 51938 30660 51950
rect 30604 51886 30606 51938
rect 30658 51886 30660 51938
rect 30604 51378 30660 51886
rect 30604 51326 30606 51378
rect 30658 51326 30660 51378
rect 30492 50820 30548 50830
rect 30044 50530 30100 50540
rect 30268 50596 30324 50606
rect 30268 50502 30324 50540
rect 30380 49924 30436 49934
rect 30044 49810 30100 49822
rect 30044 49758 30046 49810
rect 30098 49758 30100 49810
rect 30044 48356 30100 49758
rect 30268 49812 30324 49822
rect 30268 49718 30324 49756
rect 30380 48804 30436 49868
rect 30492 49252 30548 50764
rect 30604 50596 30660 51326
rect 30604 50530 30660 50540
rect 30716 50428 30772 55020
rect 31276 54628 31332 54638
rect 30940 54572 31276 54628
rect 30940 54514 30996 54572
rect 31276 54562 31332 54572
rect 30940 54462 30942 54514
rect 30994 54462 30996 54514
rect 30940 54450 30996 54462
rect 31164 54402 31220 54414
rect 31164 54350 31166 54402
rect 31218 54350 31220 54402
rect 31164 54292 31220 54350
rect 31388 54292 31444 56812
rect 31612 56308 31668 57344
rect 32060 57204 32116 57344
rect 32060 57138 32116 57148
rect 31612 56242 31668 56252
rect 31724 56756 31780 56766
rect 31500 56196 31556 56206
rect 31500 55410 31556 56140
rect 31724 56084 31780 56700
rect 31500 55358 31502 55410
rect 31554 55358 31556 55410
rect 31500 55346 31556 55358
rect 31612 56028 31780 56084
rect 31836 56532 31892 56542
rect 31612 54404 31668 56028
rect 31724 55860 31780 55870
rect 31724 55766 31780 55804
rect 31836 55410 31892 56476
rect 32508 56084 32564 57344
rect 32508 56018 32564 56028
rect 32732 55972 32788 55982
rect 32732 55878 32788 55916
rect 32060 55860 32116 55870
rect 32060 55858 32340 55860
rect 32060 55806 32062 55858
rect 32114 55806 32340 55858
rect 32060 55804 32340 55806
rect 32060 55794 32116 55804
rect 31836 55358 31838 55410
rect 31890 55358 31892 55410
rect 31836 55346 31892 55358
rect 31836 54404 31892 54414
rect 31612 54402 31892 54404
rect 31612 54350 31838 54402
rect 31890 54350 31892 54402
rect 31612 54348 31892 54350
rect 31836 54338 31892 54348
rect 31164 54236 31444 54292
rect 31500 54290 31556 54302
rect 31500 54238 31502 54290
rect 31554 54238 31556 54290
rect 31500 53956 31556 54238
rect 31388 53900 31556 53956
rect 31948 53956 32004 53966
rect 30828 53842 30884 53854
rect 30828 53790 30830 53842
rect 30882 53790 30884 53842
rect 30828 53620 30884 53790
rect 31276 53844 31332 53854
rect 30828 53554 30884 53564
rect 31164 53730 31220 53742
rect 31164 53678 31166 53730
rect 31218 53678 31220 53730
rect 31164 53508 31220 53678
rect 31164 53442 31220 53452
rect 31276 53172 31332 53788
rect 31164 53116 31332 53172
rect 30940 52836 30996 52846
rect 30940 52742 30996 52780
rect 31164 52386 31220 53116
rect 31164 52334 31166 52386
rect 31218 52334 31220 52386
rect 31164 52322 31220 52334
rect 31276 52722 31332 52734
rect 31276 52670 31278 52722
rect 31330 52670 31332 52722
rect 30828 52164 30884 52174
rect 31052 52164 31108 52174
rect 30884 52108 30996 52164
rect 30828 52098 30884 52108
rect 30828 50596 30884 50606
rect 30828 50502 30884 50540
rect 30604 50372 30772 50428
rect 30604 49476 30660 50372
rect 30940 49924 30996 52108
rect 31052 52070 31108 52108
rect 31164 51380 31220 51390
rect 31164 51286 31220 51324
rect 31276 50148 31332 52670
rect 31276 50082 31332 50092
rect 31388 50036 31444 53900
rect 31836 53842 31892 53854
rect 31836 53790 31838 53842
rect 31890 53790 31892 53842
rect 31500 53732 31556 53742
rect 31500 53638 31556 53676
rect 31724 53732 31780 53742
rect 31500 53508 31556 53518
rect 31500 52724 31556 53452
rect 31724 53170 31780 53676
rect 31724 53118 31726 53170
rect 31778 53118 31780 53170
rect 31724 53106 31780 53118
rect 31836 53172 31892 53790
rect 31836 53106 31892 53116
rect 31500 52658 31556 52668
rect 31612 52946 31668 52958
rect 31612 52894 31614 52946
rect 31666 52894 31668 52946
rect 31500 52276 31556 52286
rect 31500 52182 31556 52220
rect 31612 50708 31668 52894
rect 31836 52948 31892 52958
rect 31948 52948 32004 53900
rect 32172 53620 32228 53630
rect 32060 53172 32116 53182
rect 32060 53078 32116 53116
rect 32172 53170 32228 53564
rect 32172 53118 32174 53170
rect 32226 53118 32228 53170
rect 32172 53106 32228 53118
rect 31836 52946 32004 52948
rect 31836 52894 31838 52946
rect 31890 52894 32004 52946
rect 31836 52892 32004 52894
rect 31836 52882 31892 52892
rect 31612 50428 31668 50652
rect 31836 52274 31892 52286
rect 31836 52222 31838 52274
rect 31890 52222 31892 52274
rect 31388 49970 31444 49980
rect 31500 50372 31668 50428
rect 31724 50594 31780 50606
rect 31724 50542 31726 50594
rect 31778 50542 31780 50594
rect 30940 49858 30996 49868
rect 30716 49700 30772 49710
rect 30716 49698 31444 49700
rect 30716 49646 30718 49698
rect 30770 49646 31444 49698
rect 30716 49644 31444 49646
rect 30716 49634 30772 49644
rect 30604 49420 30996 49476
rect 30604 49252 30660 49262
rect 30492 49250 30660 49252
rect 30492 49198 30606 49250
rect 30658 49198 30660 49250
rect 30492 49196 30660 49198
rect 30604 49186 30660 49196
rect 30828 49252 30884 49262
rect 30828 49158 30884 49196
rect 30492 49028 30548 49038
rect 30492 48934 30548 48972
rect 30380 48748 30548 48804
rect 30156 48356 30212 48366
rect 30044 48300 30156 48356
rect 29036 46946 29092 46956
rect 29596 47180 29988 47236
rect 28812 46844 28980 46900
rect 29260 46900 29316 46910
rect 29596 46900 29652 47180
rect 29260 46898 29652 46900
rect 29260 46846 29262 46898
rect 29314 46846 29652 46898
rect 29260 46844 29652 46846
rect 28812 46738 28868 46844
rect 29260 46834 29316 46844
rect 29148 46788 29204 46798
rect 28588 46498 28644 46508
rect 28700 46682 28868 46738
rect 28980 46786 29204 46788
rect 28980 46734 29150 46786
rect 29202 46734 29204 46786
rect 28980 46732 29204 46734
rect 27692 46050 27748 46060
rect 27804 46450 27860 46462
rect 27804 46398 27806 46450
rect 27858 46398 27860 46450
rect 27580 44706 27636 44716
rect 27692 45890 27748 45902
rect 27692 45838 27694 45890
rect 27746 45838 27748 45890
rect 27692 44322 27748 45838
rect 27692 44270 27694 44322
rect 27746 44270 27748 44322
rect 27244 43538 27412 43540
rect 27244 43486 27246 43538
rect 27298 43486 27412 43538
rect 27244 43484 27412 43486
rect 27468 43540 27524 43550
rect 27244 43428 27300 43484
rect 27244 43362 27300 43372
rect 27468 42978 27524 43484
rect 27468 42926 27470 42978
rect 27522 42926 27524 42978
rect 27468 42914 27524 42926
rect 27244 42754 27300 42766
rect 27692 42756 27748 44270
rect 27804 44324 27860 46398
rect 28028 46228 28084 46238
rect 27916 46116 27972 46154
rect 28028 46116 28084 46172
rect 28028 46060 28644 46116
rect 27916 46050 27972 46060
rect 28588 46004 28644 46060
rect 28588 45938 28644 45948
rect 28364 45892 28420 45902
rect 28364 45798 28420 45836
rect 28700 45332 28756 46682
rect 28700 45266 28756 45276
rect 28812 46564 28868 46574
rect 28700 45108 28756 45118
rect 28588 44884 28644 44894
rect 28364 44882 28644 44884
rect 28364 44830 28590 44882
rect 28642 44830 28644 44882
rect 28364 44828 28644 44830
rect 27916 44660 27972 44670
rect 27916 44546 27972 44604
rect 27916 44494 27918 44546
rect 27970 44494 27972 44546
rect 27916 44482 27972 44494
rect 27804 44258 27860 44268
rect 28252 43540 28308 43550
rect 27916 43092 27972 43102
rect 27916 42866 27972 43036
rect 27916 42814 27918 42866
rect 27970 42814 27972 42866
rect 27916 42802 27972 42814
rect 27244 42702 27246 42754
rect 27298 42702 27300 42754
rect 27244 42084 27300 42702
rect 27244 42018 27300 42028
rect 27356 42700 27748 42756
rect 27356 39844 27412 42700
rect 27692 42308 27748 42318
rect 27692 41076 27748 42252
rect 28140 41636 28196 41646
rect 27916 41076 27972 41086
rect 27692 41074 27972 41076
rect 27692 41022 27918 41074
rect 27970 41022 27972 41074
rect 27692 41020 27972 41022
rect 27468 40962 27524 40974
rect 27468 40910 27470 40962
rect 27522 40910 27524 40962
rect 27468 40180 27524 40910
rect 27468 40114 27524 40124
rect 27468 39844 27524 39854
rect 27356 39842 27524 39844
rect 27356 39790 27470 39842
rect 27522 39790 27524 39842
rect 27356 39788 27524 39790
rect 27468 39778 27524 39788
rect 27244 39620 27300 39630
rect 27692 39620 27748 41020
rect 27916 41010 27972 41020
rect 27804 40180 27860 40190
rect 28028 40180 28084 40190
rect 27804 40178 27972 40180
rect 27804 40126 27806 40178
rect 27858 40126 27972 40178
rect 27804 40124 27972 40126
rect 27804 40114 27860 40124
rect 27244 39526 27300 39564
rect 27356 39564 27748 39620
rect 27132 37314 27188 37324
rect 27244 37268 27300 37278
rect 27244 37174 27300 37212
rect 27020 37156 27076 37166
rect 27020 33908 27076 37100
rect 27356 35308 27412 39564
rect 27804 38612 27860 38622
rect 27804 38518 27860 38556
rect 27916 38052 27972 40124
rect 28028 39618 28084 40124
rect 28028 39566 28030 39618
rect 28082 39566 28084 39618
rect 28028 39554 28084 39566
rect 28140 38500 28196 41580
rect 28140 38434 28196 38444
rect 27916 37986 27972 37996
rect 28252 37940 28308 43484
rect 28364 41186 28420 44828
rect 28588 44818 28644 44828
rect 28476 44324 28532 44334
rect 28476 44230 28532 44268
rect 28700 43988 28756 45052
rect 28700 43650 28756 43932
rect 28700 43598 28702 43650
rect 28754 43598 28756 43650
rect 28700 43586 28756 43598
rect 28588 43428 28644 43438
rect 28476 42644 28532 42654
rect 28476 41636 28532 42588
rect 28476 41570 28532 41580
rect 28364 41134 28366 41186
rect 28418 41134 28420 41186
rect 28364 41122 28420 41134
rect 28588 40180 28644 43372
rect 28700 42756 28756 42766
rect 28700 42662 28756 42700
rect 28700 42084 28756 42094
rect 28700 41188 28756 42028
rect 28812 41524 28868 46508
rect 28980 46452 29036 46732
rect 29148 46722 29204 46732
rect 29596 46674 29652 46844
rect 29596 46622 29598 46674
rect 29650 46622 29652 46674
rect 29596 46610 29652 46622
rect 30044 47124 30100 47134
rect 29148 46564 29204 46574
rect 28980 46396 29092 46452
rect 28812 41458 28868 41468
rect 28924 45890 28980 45902
rect 28924 45838 28926 45890
rect 28978 45838 28980 45890
rect 28924 44322 28980 45838
rect 29036 45892 29092 46396
rect 29036 45826 29092 45836
rect 28924 44270 28926 44322
rect 28978 44270 28980 44322
rect 28924 41410 28980 44270
rect 28924 41358 28926 41410
rect 28978 41358 28980 41410
rect 28924 41346 28980 41358
rect 29036 45332 29092 45342
rect 28700 41186 28868 41188
rect 28700 41134 28702 41186
rect 28754 41134 28868 41186
rect 28700 41132 28868 41134
rect 28700 41122 28756 41132
rect 28588 40114 28644 40124
rect 28700 40740 28756 40750
rect 28700 40516 28756 40684
rect 28700 39618 28756 40460
rect 28700 39566 28702 39618
rect 28754 39566 28756 39618
rect 28700 39554 28756 39566
rect 28700 39172 28756 39182
rect 28140 37938 28308 37940
rect 28140 37886 28254 37938
rect 28306 37886 28308 37938
rect 28140 37884 28308 37886
rect 27580 37828 27636 37838
rect 27580 37826 27748 37828
rect 27580 37774 27582 37826
rect 27634 37774 27748 37826
rect 27580 37772 27748 37774
rect 27580 37762 27636 37772
rect 27244 35252 27412 35308
rect 27468 36484 27524 36494
rect 27244 34802 27300 35252
rect 27244 34750 27246 34802
rect 27298 34750 27300 34802
rect 27244 34692 27300 34750
rect 27244 34626 27300 34636
rect 27020 33842 27076 33852
rect 27132 33796 27188 33806
rect 27020 33348 27076 33358
rect 27132 33348 27188 33740
rect 27020 33346 27188 33348
rect 27020 33294 27022 33346
rect 27074 33294 27188 33346
rect 27020 33292 27188 33294
rect 27356 33346 27412 33358
rect 27356 33294 27358 33346
rect 27410 33294 27412 33346
rect 27020 33282 27076 33292
rect 27356 32340 27412 33294
rect 27468 32452 27524 36428
rect 27580 36482 27636 36494
rect 27580 36430 27582 36482
rect 27634 36430 27636 36482
rect 27580 35252 27636 36430
rect 27580 35186 27636 35196
rect 27692 34914 27748 37772
rect 27804 35476 27860 35486
rect 27804 35474 27972 35476
rect 27804 35422 27806 35474
rect 27858 35422 27972 35474
rect 27804 35420 27972 35422
rect 27804 35410 27860 35420
rect 27692 34862 27694 34914
rect 27746 34862 27748 34914
rect 27692 34850 27748 34862
rect 27580 34130 27636 34142
rect 27580 34078 27582 34130
rect 27634 34078 27636 34130
rect 27580 33908 27636 34078
rect 27580 33684 27636 33852
rect 27580 33618 27636 33628
rect 27580 33458 27636 33470
rect 27580 33406 27582 33458
rect 27634 33406 27636 33458
rect 27580 32900 27636 33406
rect 27916 33460 27972 35420
rect 28028 34916 28084 34926
rect 28028 34822 28084 34860
rect 28028 33460 28084 33470
rect 27916 33458 28084 33460
rect 27916 33406 28030 33458
rect 28082 33406 28084 33458
rect 27916 33404 28084 33406
rect 28028 33394 28084 33404
rect 27580 32834 27636 32844
rect 28140 32676 28196 37884
rect 28252 37874 28308 37884
rect 28588 38836 28644 38846
rect 28700 38836 28756 39116
rect 28812 39060 28868 41132
rect 28924 41076 28980 41086
rect 28924 40514 28980 41020
rect 28924 40462 28926 40514
rect 28978 40462 28980 40514
rect 28924 40450 28980 40462
rect 29036 39172 29092 45276
rect 29148 44212 29204 46508
rect 29708 46452 29764 46462
rect 29708 46358 29764 46396
rect 29932 46450 29988 46462
rect 29932 46398 29934 46450
rect 29986 46398 29988 46450
rect 29932 46340 29988 46398
rect 29932 46274 29988 46284
rect 29932 45892 29988 45902
rect 30044 45892 30100 47068
rect 29932 45890 30100 45892
rect 29932 45838 29934 45890
rect 29986 45838 30100 45890
rect 29932 45836 30100 45838
rect 29820 44994 29876 45006
rect 29820 44942 29822 44994
rect 29874 44942 29876 44994
rect 29596 44884 29652 44894
rect 29596 44660 29652 44828
rect 29596 44604 29764 44660
rect 29148 44146 29204 44156
rect 29148 43314 29204 43326
rect 29148 43262 29150 43314
rect 29202 43262 29204 43314
rect 29148 42532 29204 43262
rect 29148 42466 29204 42476
rect 29372 43316 29428 43326
rect 29372 42084 29428 43260
rect 29596 43316 29652 43326
rect 29484 43092 29540 43102
rect 29484 42754 29540 43036
rect 29484 42702 29486 42754
rect 29538 42702 29540 42754
rect 29484 42690 29540 42702
rect 29372 40290 29428 42028
rect 29596 41186 29652 43260
rect 29596 41134 29598 41186
rect 29650 41134 29652 41186
rect 29596 41122 29652 41134
rect 29372 40238 29374 40290
rect 29426 40238 29428 40290
rect 29372 39284 29428 40238
rect 29036 39106 29092 39116
rect 29148 39228 29428 39284
rect 29484 39618 29540 39630
rect 29484 39566 29486 39618
rect 29538 39566 29540 39618
rect 28812 39004 28980 39060
rect 28644 38834 28756 38836
rect 28644 38782 28702 38834
rect 28754 38782 28756 38834
rect 28644 38780 28756 38782
rect 28476 37380 28532 37390
rect 28476 37286 28532 37324
rect 28364 37268 28420 37278
rect 28252 35026 28308 35038
rect 28252 34974 28254 35026
rect 28306 34974 28308 35026
rect 28252 33684 28308 34974
rect 28252 33618 28308 33628
rect 28140 32620 28308 32676
rect 27468 32386 27524 32396
rect 28140 32452 28196 32462
rect 26908 31892 27076 31948
rect 26908 31780 26964 31790
rect 26908 31686 26964 31724
rect 26908 31220 26964 31230
rect 26796 31108 26852 31118
rect 26796 30994 26852 31052
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30930 26852 30942
rect 26684 30882 26740 30894
rect 26684 30830 26686 30882
rect 26738 30830 26740 30882
rect 26684 30436 26740 30830
rect 26684 30370 26740 30380
rect 26572 29262 26574 29314
rect 26626 29262 26628 29314
rect 26572 29250 26628 29262
rect 26684 29316 26740 29326
rect 26460 28868 26516 28878
rect 26460 28774 26516 28812
rect 26124 27122 26180 27132
rect 26236 28532 26292 28542
rect 26236 28196 26292 28476
rect 26236 26402 26292 28140
rect 26460 27972 26516 27982
rect 26348 27300 26404 27310
rect 26348 26964 26404 27244
rect 26348 26898 26404 26908
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 26236 26338 26292 26350
rect 26124 26290 26180 26302
rect 26124 26238 26126 26290
rect 26178 26238 26180 26290
rect 26124 25506 26180 26238
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 25172 26180 25454
rect 26124 25106 26180 25116
rect 26236 25396 26292 25406
rect 26236 24834 26292 25340
rect 26236 24782 26238 24834
rect 26290 24782 26292 24834
rect 26124 24724 26180 24734
rect 26124 23268 26180 24668
rect 26124 23202 26180 23212
rect 26012 22306 26068 22316
rect 26124 22372 26180 22382
rect 26236 22372 26292 24782
rect 26460 24276 26516 27916
rect 26572 27188 26628 27198
rect 26572 27094 26628 27132
rect 26572 26180 26628 26190
rect 26572 26086 26628 26124
rect 26572 25732 26628 25742
rect 26684 25732 26740 29260
rect 26908 27524 26964 31164
rect 27020 30324 27076 31892
rect 27356 31778 27412 32284
rect 27356 31726 27358 31778
rect 27410 31726 27412 31778
rect 27356 31714 27412 31726
rect 27468 31890 27524 31902
rect 27468 31838 27470 31890
rect 27522 31838 27524 31890
rect 27468 31556 27524 31838
rect 27916 31778 27972 31790
rect 27916 31726 27918 31778
rect 27970 31726 27972 31778
rect 27468 31500 27748 31556
rect 27468 30996 27524 31006
rect 27468 30902 27524 30940
rect 27692 30660 27748 31500
rect 27804 30772 27860 30782
rect 27804 30678 27860 30716
rect 27692 30594 27748 30604
rect 27244 30436 27300 30446
rect 27916 30436 27972 31726
rect 27244 30434 27972 30436
rect 27244 30382 27246 30434
rect 27298 30382 27972 30434
rect 27244 30380 27972 30382
rect 28028 30996 28084 31006
rect 27244 30370 27300 30380
rect 27020 28084 27076 30268
rect 27804 30212 27860 30222
rect 27020 28018 27076 28028
rect 27244 30100 27300 30110
rect 26908 27458 26964 27468
rect 27020 27858 27076 27870
rect 27020 27806 27022 27858
rect 27074 27806 27076 27858
rect 26908 27076 26964 27114
rect 26908 27010 26964 27020
rect 27020 26908 27076 27806
rect 26908 26852 27076 26908
rect 27132 27524 27188 27534
rect 26572 25730 26740 25732
rect 26572 25678 26574 25730
rect 26626 25678 26740 25730
rect 26572 25676 26740 25678
rect 26572 25666 26628 25676
rect 26684 25508 26740 25676
rect 26684 25442 26740 25452
rect 26796 25732 26852 25742
rect 26796 25284 26852 25676
rect 26572 25228 26852 25284
rect 26572 24276 26628 25228
rect 26684 24500 26740 24510
rect 26684 24406 26740 24444
rect 26572 24220 26740 24276
rect 26460 24210 26516 24220
rect 26572 24052 26628 24062
rect 26460 24050 26628 24052
rect 26460 23998 26574 24050
rect 26626 23998 26628 24050
rect 26460 23996 26628 23998
rect 26348 23940 26404 23950
rect 26348 23846 26404 23884
rect 26124 22370 26292 22372
rect 26124 22318 26126 22370
rect 26178 22318 26292 22370
rect 26124 22316 26292 22318
rect 26124 22306 26180 22316
rect 25452 21812 25508 21822
rect 25452 21588 25508 21756
rect 25452 21586 25844 21588
rect 25452 21534 25454 21586
rect 25506 21534 25844 21586
rect 25452 21532 25844 21534
rect 25452 21522 25508 21532
rect 25340 21410 25396 21420
rect 25676 21364 25732 21374
rect 25564 21252 25620 21262
rect 25340 20916 25396 20926
rect 25564 20916 25620 21196
rect 25340 20802 25396 20860
rect 25340 20750 25342 20802
rect 25394 20750 25396 20802
rect 25340 20738 25396 20750
rect 25452 20914 25620 20916
rect 25452 20862 25566 20914
rect 25618 20862 25620 20914
rect 25452 20860 25620 20862
rect 25340 20018 25396 20030
rect 25340 19966 25342 20018
rect 25394 19966 25396 20018
rect 25340 19908 25396 19966
rect 25452 20020 25508 20860
rect 25564 20850 25620 20860
rect 25452 19954 25508 19964
rect 25564 20132 25620 20142
rect 25340 19842 25396 19852
rect 25340 19684 25396 19694
rect 25340 19460 25396 19628
rect 25340 19458 25508 19460
rect 25340 19406 25342 19458
rect 25394 19406 25508 19458
rect 25340 19404 25508 19406
rect 25340 19394 25396 19404
rect 25452 18564 25508 19404
rect 25564 19124 25620 20076
rect 25564 19058 25620 19068
rect 25452 18498 25508 18508
rect 25676 18340 25732 21308
rect 25788 20356 25844 21532
rect 26124 21476 26180 21486
rect 25900 21364 25956 21374
rect 26124 21364 26180 21420
rect 25900 21362 26180 21364
rect 25900 21310 25902 21362
rect 25954 21310 26180 21362
rect 25900 21308 26180 21310
rect 25900 21298 25956 21308
rect 26124 20804 26180 20814
rect 26124 20710 26180 20748
rect 25788 20290 25844 20300
rect 26236 20244 26292 22316
rect 26460 21812 26516 23996
rect 26572 23986 26628 23996
rect 26684 23492 26740 24220
rect 26908 23716 26964 26852
rect 26684 23426 26740 23436
rect 26796 23660 26964 23716
rect 27020 23938 27076 23950
rect 27020 23886 27022 23938
rect 27074 23886 27076 23938
rect 26684 23154 26740 23166
rect 26684 23102 26686 23154
rect 26738 23102 26740 23154
rect 26684 23044 26740 23102
rect 26684 22978 26740 22988
rect 26460 21746 26516 21756
rect 26572 22482 26628 22494
rect 26572 22430 26574 22482
rect 26626 22430 26628 22482
rect 26572 21028 26628 22430
rect 26796 22036 26852 23660
rect 25452 18284 25732 18340
rect 26124 20188 26292 20244
rect 26348 20972 26628 21028
rect 26684 21140 26740 21150
rect 26124 18340 26180 20188
rect 26236 20020 26292 20030
rect 26236 19926 26292 19964
rect 26236 19796 26292 19806
rect 26236 19236 26292 19740
rect 26348 19348 26404 20972
rect 26348 19282 26404 19292
rect 26572 20802 26628 20814
rect 26572 20750 26574 20802
rect 26626 20750 26628 20802
rect 26572 19908 26628 20750
rect 26684 20692 26740 21084
rect 26684 20626 26740 20636
rect 26236 19170 26292 19180
rect 26460 19236 26516 19246
rect 26460 19142 26516 19180
rect 26348 18788 26404 18798
rect 26236 18452 26292 18462
rect 26236 18358 26292 18396
rect 25228 17276 25396 17332
rect 25228 16884 25284 16894
rect 25228 16790 25284 16828
rect 25116 15810 25172 15820
rect 24668 14700 25060 14756
rect 24668 14642 24724 14700
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14578 24724 14590
rect 25004 14532 25060 14542
rect 24332 14354 24388 14364
rect 24780 14530 25060 14532
rect 24780 14478 25006 14530
rect 25058 14478 25060 14530
rect 24780 14476 25060 14478
rect 24780 14084 24836 14476
rect 25004 14466 25060 14476
rect 25116 14532 25172 14542
rect 24332 14028 24836 14084
rect 24892 14084 24948 14094
rect 24332 13970 24388 14028
rect 24332 13918 24334 13970
rect 24386 13918 24388 13970
rect 24332 13906 24388 13918
rect 24892 13748 24948 14028
rect 24892 13682 24948 13692
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24668 12740 24724 12750
rect 24668 12738 25060 12740
rect 24668 12686 24670 12738
rect 24722 12686 25060 12738
rect 24668 12684 25060 12686
rect 24668 12674 24724 12684
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24220 12562 24276 12572
rect 24444 12628 24500 12638
rect 23804 12506 24068 12516
rect 23660 12348 24052 12404
rect 23548 12236 23716 12292
rect 22876 11554 22932 11564
rect 23100 11956 23156 11966
rect 22540 10948 22596 10958
rect 22540 10834 22596 10892
rect 22540 10782 22542 10834
rect 22594 10782 22596 10834
rect 22540 10770 22596 10782
rect 22540 10500 22596 10510
rect 22540 8258 22596 10444
rect 22988 10500 23044 10538
rect 22988 10434 23044 10444
rect 22988 10276 23044 10286
rect 22764 10052 22820 10062
rect 22764 9958 22820 9996
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22540 8194 22596 8206
rect 22764 8148 22820 8158
rect 22652 7476 22708 7486
rect 22428 7474 22708 7476
rect 22428 7422 22654 7474
rect 22706 7422 22708 7474
rect 22428 7420 22708 7422
rect 22652 7410 22708 7420
rect 22764 7252 22820 8092
rect 22652 7196 22820 7252
rect 22428 6692 22484 6702
rect 22316 6690 22484 6692
rect 22316 6638 22430 6690
rect 22482 6638 22484 6690
rect 22316 6636 22484 6638
rect 22316 5124 22372 6636
rect 22428 6626 22484 6636
rect 22652 6018 22708 7196
rect 22876 7028 22932 7038
rect 22876 6692 22932 6972
rect 22652 5966 22654 6018
rect 22706 5966 22708 6018
rect 22652 5954 22708 5966
rect 22764 6690 22932 6692
rect 22764 6638 22878 6690
rect 22930 6638 22932 6690
rect 22764 6636 22932 6638
rect 22764 5348 22820 6636
rect 22876 6626 22932 6636
rect 22316 5058 22372 5068
rect 22652 5292 22820 5348
rect 22876 5796 22932 5806
rect 22652 4452 22708 5292
rect 22764 5124 22820 5134
rect 22764 5030 22820 5068
rect 22652 4396 22820 4452
rect 22316 4116 22372 4126
rect 22652 4116 22708 4126
rect 22316 4114 22596 4116
rect 22316 4062 22318 4114
rect 22370 4062 22596 4114
rect 22316 4060 22596 4062
rect 22316 4050 22372 4060
rect 22204 3836 22372 3892
rect 22316 3554 22372 3836
rect 22316 3502 22318 3554
rect 22370 3502 22372 3554
rect 21868 3332 22148 3388
rect 21532 3266 21588 3276
rect 21868 2772 21924 2782
rect 21420 2706 21476 2716
rect 21532 2770 21924 2772
rect 21532 2718 21870 2770
rect 21922 2718 21924 2770
rect 21532 2716 21924 2718
rect 21532 2546 21588 2716
rect 21868 2706 21924 2716
rect 21532 2494 21534 2546
rect 21586 2494 21588 2546
rect 21532 2482 21588 2494
rect 21308 2258 21364 2268
rect 21420 2436 21476 2446
rect 21420 1986 21476 2380
rect 21420 1934 21422 1986
rect 21474 1934 21476 1986
rect 21420 1764 21476 1934
rect 21420 1698 21476 1708
rect 21980 1764 22036 1774
rect 22092 1764 22148 3332
rect 22204 3332 22260 3342
rect 22204 2994 22260 3276
rect 22204 2942 22206 2994
rect 22258 2942 22260 2994
rect 22204 2930 22260 2942
rect 22316 1986 22372 3502
rect 22540 3388 22596 4060
rect 22652 4022 22708 4060
rect 22764 4004 22820 4396
rect 22764 3938 22820 3948
rect 22652 3892 22708 3902
rect 22652 3666 22708 3836
rect 22652 3614 22654 3666
rect 22706 3614 22708 3666
rect 22652 3602 22708 3614
rect 22540 3332 22820 3388
rect 22764 2884 22820 3332
rect 22876 3220 22932 5740
rect 22988 4338 23044 10220
rect 23100 9268 23156 11900
rect 23324 11844 23380 12012
rect 23548 12068 23604 12078
rect 23548 11974 23604 12012
rect 23324 11788 23604 11844
rect 23436 11508 23492 11518
rect 23324 10948 23380 10958
rect 23324 10610 23380 10892
rect 23324 10558 23326 10610
rect 23378 10558 23380 10610
rect 23324 10546 23380 10558
rect 23436 10500 23492 11452
rect 23436 10434 23492 10444
rect 23100 9202 23156 9212
rect 23436 9044 23492 9054
rect 23324 7588 23380 7598
rect 23324 6356 23380 7532
rect 23436 6804 23492 8988
rect 23548 7476 23604 11788
rect 23660 10612 23716 12236
rect 23884 12180 23940 12190
rect 23884 12086 23940 12124
rect 23996 12068 24052 12348
rect 24444 12178 24500 12572
rect 24444 12126 24446 12178
rect 24498 12126 24500 12178
rect 24444 12114 24500 12126
rect 25004 12178 25060 12684
rect 25004 12126 25006 12178
rect 25058 12126 25060 12178
rect 25004 12114 25060 12126
rect 23996 12002 24052 12012
rect 24556 11956 24612 11966
rect 24332 11954 24612 11956
rect 24332 11902 24558 11954
rect 24610 11902 24612 11954
rect 24332 11900 24612 11902
rect 23772 11844 23828 11854
rect 24332 11844 24388 11900
rect 24556 11890 24612 11900
rect 23772 11172 23828 11788
rect 23772 11106 23828 11116
rect 24220 11788 24388 11844
rect 24464 11788 24728 11798
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23772 10612 23828 10622
rect 23660 10610 23828 10612
rect 23660 10558 23774 10610
rect 23826 10558 23828 10610
rect 23660 10556 23828 10558
rect 23772 10546 23828 10556
rect 23884 10612 23940 10622
rect 23884 10050 23940 10556
rect 23996 10388 24052 10398
rect 23996 10294 24052 10332
rect 23884 9998 23886 10050
rect 23938 9998 23940 10050
rect 23884 9986 23940 9998
rect 23804 9436 24068 9446
rect 23660 9380 23716 9390
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 23660 9044 23716 9324
rect 23660 8978 23716 8988
rect 23884 9042 23940 9054
rect 23884 8990 23886 9042
rect 23938 8990 23940 9042
rect 23884 8260 23940 8990
rect 23884 8194 23940 8204
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 23660 7476 23716 7486
rect 23548 7474 23716 7476
rect 23548 7422 23662 7474
rect 23714 7422 23716 7474
rect 23548 7420 23716 7422
rect 23660 7410 23716 7420
rect 23548 6804 23604 6814
rect 23436 6748 23548 6804
rect 23436 6580 23492 6590
rect 23436 6486 23492 6524
rect 23324 6300 23492 6356
rect 23100 6132 23156 6142
rect 23100 5794 23156 6076
rect 23100 5742 23102 5794
rect 23154 5742 23156 5794
rect 23100 5730 23156 5742
rect 22988 4286 22990 4338
rect 23042 4286 23044 4338
rect 22988 4274 23044 4286
rect 22876 3154 22932 3164
rect 23436 3220 23492 6300
rect 23548 4338 23604 6748
rect 23660 6802 23716 6814
rect 23660 6750 23662 6802
rect 23714 6750 23716 6802
rect 23660 5460 23716 6750
rect 23996 6690 24052 6702
rect 23996 6638 23998 6690
rect 24050 6638 24052 6690
rect 23996 6580 24052 6638
rect 23996 6514 24052 6524
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24220 6132 24276 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24332 11620 24388 11630
rect 24332 9716 24388 11564
rect 24444 10612 24500 10622
rect 24444 10518 24500 10556
rect 25004 10612 25060 10622
rect 25004 10518 25060 10556
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 24332 9650 24388 9660
rect 24332 9380 24388 9390
rect 24332 8818 24388 9324
rect 25116 9268 25172 14476
rect 25228 14308 25284 14318
rect 25228 13748 25284 14252
rect 25228 12516 25284 13692
rect 25228 12450 25284 12460
rect 25228 12292 25284 12302
rect 25228 11394 25284 12236
rect 25228 11342 25230 11394
rect 25282 11342 25284 11394
rect 25228 11330 25284 11342
rect 24332 8766 24334 8818
rect 24386 8766 24388 8818
rect 24332 8596 24388 8766
rect 24892 9212 25172 9268
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24332 8530 24388 8540
rect 24332 8260 24388 8270
rect 24332 6916 24388 8204
rect 24668 7700 24724 7710
rect 24668 7586 24724 7644
rect 24668 7534 24670 7586
rect 24722 7534 24724 7586
rect 24668 7364 24724 7534
rect 24668 7298 24724 7308
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 24892 6916 24948 9212
rect 24332 6860 24500 6916
rect 24332 6692 24388 6702
rect 24332 6356 24388 6636
rect 24332 6290 24388 6300
rect 24444 6244 24500 6860
rect 24780 6860 24948 6916
rect 25004 8260 25060 8270
rect 25004 7474 25060 8204
rect 25004 7422 25006 7474
rect 25058 7422 25060 7474
rect 24444 6178 24500 6188
rect 24556 6802 24612 6814
rect 24556 6750 24558 6802
rect 24610 6750 24612 6802
rect 23660 5394 23716 5404
rect 23996 6076 24276 6132
rect 23996 5346 24052 6076
rect 24220 5908 24276 5918
rect 24220 5814 24276 5852
rect 24556 5796 24612 6750
rect 24780 6468 24836 6860
rect 24892 6692 24948 6702
rect 24892 6598 24948 6636
rect 24780 6412 24948 6468
rect 24668 6020 24724 6030
rect 24668 5926 24724 5964
rect 24556 5730 24612 5740
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23996 5294 23998 5346
rect 24050 5294 24052 5346
rect 23996 5282 24052 5294
rect 23548 4286 23550 4338
rect 23602 4286 23604 4338
rect 23548 3780 23604 4286
rect 23660 5234 23716 5246
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23660 4340 23716 5182
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24220 4676 24276 4686
rect 23660 4274 23716 4284
rect 23884 4340 23940 4350
rect 23884 4004 23940 4284
rect 23996 4116 24052 4126
rect 23996 4022 24052 4060
rect 23884 3938 23940 3948
rect 23548 3714 23604 3724
rect 24220 3556 24276 4620
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 24892 3778 24948 6412
rect 25004 5908 25060 7422
rect 25116 7028 25172 7038
rect 25116 6804 25172 6972
rect 25116 6738 25172 6748
rect 25228 6692 25284 6702
rect 25228 6356 25284 6636
rect 25004 5814 25060 5852
rect 25116 6300 25284 6356
rect 24892 3726 24894 3778
rect 24946 3726 24948 3778
rect 24892 3714 24948 3726
rect 25004 5234 25060 5246
rect 25004 5182 25006 5234
rect 25058 5182 25060 5234
rect 24220 3490 24276 3500
rect 24556 3666 24612 3678
rect 24556 3614 24558 3666
rect 24610 3614 24612 3666
rect 24556 3388 24612 3614
rect 23884 3332 23940 3342
rect 23436 3154 23492 3164
rect 23660 3330 23940 3332
rect 23660 3278 23886 3330
rect 23938 3278 23940 3330
rect 23660 3276 23940 3278
rect 23548 3108 23604 3118
rect 22764 2828 23268 2884
rect 22428 2772 22484 2782
rect 22428 2678 22484 2716
rect 22652 2660 22708 2670
rect 22988 2660 23044 2670
rect 22652 2658 23044 2660
rect 22652 2606 22654 2658
rect 22706 2606 22990 2658
rect 23042 2606 23044 2658
rect 22652 2604 23044 2606
rect 22652 2594 22708 2604
rect 22988 2594 23044 2604
rect 23100 2660 23156 2670
rect 23100 2566 23156 2604
rect 22540 2546 22596 2558
rect 22540 2494 22542 2546
rect 22594 2494 22596 2546
rect 22540 2100 22596 2494
rect 22540 2034 22596 2044
rect 22652 2212 22708 2222
rect 22652 2098 22708 2156
rect 22652 2046 22654 2098
rect 22706 2046 22708 2098
rect 22652 2034 22708 2046
rect 22316 1934 22318 1986
rect 22370 1934 22372 1986
rect 22316 1922 22372 1934
rect 23100 1988 23156 1998
rect 22092 1708 22260 1764
rect 21756 1652 21812 1662
rect 21084 1202 21252 1204
rect 21084 1150 21086 1202
rect 21138 1150 21252 1202
rect 21084 1148 21252 1150
rect 21644 1428 21700 1438
rect 21644 1202 21700 1372
rect 21644 1150 21646 1202
rect 21698 1150 21700 1202
rect 21084 1138 21140 1148
rect 21644 1138 21700 1150
rect 21308 980 21364 990
rect 21308 978 21476 980
rect 21308 926 21310 978
rect 21362 926 21476 978
rect 21308 924 21476 926
rect 21308 914 21364 924
rect 21308 756 21364 766
rect 21308 112 21364 700
rect 21420 644 21476 924
rect 21420 578 21476 588
rect 21756 112 21812 1596
rect 21980 1090 22036 1708
rect 21980 1038 21982 1090
rect 22034 1038 22036 1090
rect 21980 1026 22036 1038
rect 22204 112 22260 1708
rect 23100 1202 23156 1932
rect 23100 1150 23102 1202
rect 23154 1150 23156 1202
rect 23100 1138 23156 1150
rect 22316 1092 22372 1102
rect 22316 998 22372 1036
rect 22652 980 22708 990
rect 23100 980 23156 990
rect 22652 978 22820 980
rect 22652 926 22654 978
rect 22706 926 22820 978
rect 22652 924 22820 926
rect 22652 914 22708 924
rect 22652 756 22708 766
rect 22652 112 22708 700
rect 22764 420 22820 924
rect 22764 354 22820 364
rect 23100 112 23156 924
rect 23212 308 23268 2828
rect 23436 2660 23492 2670
rect 23436 2566 23492 2604
rect 23548 2324 23604 3052
rect 23660 2772 23716 3276
rect 23884 3266 23940 3276
rect 24220 3332 24612 3388
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24220 2996 24276 3332
rect 24108 2940 24276 2996
rect 24332 3220 24388 3230
rect 23772 2772 23828 2782
rect 23660 2770 23828 2772
rect 23660 2718 23774 2770
rect 23826 2718 23828 2770
rect 23660 2716 23828 2718
rect 23772 2706 23828 2716
rect 23884 2772 23940 2782
rect 23772 2436 23828 2446
rect 23884 2436 23940 2716
rect 24108 2548 24164 2940
rect 24332 2884 24388 3164
rect 24220 2828 24388 2884
rect 24220 2770 24276 2828
rect 24892 2772 24948 2782
rect 24220 2718 24222 2770
rect 24274 2718 24276 2770
rect 24220 2706 24276 2718
rect 24332 2770 24948 2772
rect 24332 2718 24894 2770
rect 24946 2718 24948 2770
rect 24332 2716 24948 2718
rect 24108 2482 24164 2492
rect 23828 2380 23940 2436
rect 23772 2370 23828 2380
rect 24332 2324 24388 2716
rect 24892 2706 24948 2716
rect 24444 2548 24500 2586
rect 24444 2482 24500 2492
rect 23548 2258 23604 2268
rect 23884 2268 24388 2324
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24892 2324 24948 2334
rect 23884 2210 23940 2268
rect 23884 2158 23886 2210
rect 23938 2158 23940 2210
rect 23884 2146 23940 2158
rect 24892 2210 24948 2268
rect 24892 2158 24894 2210
rect 24946 2158 24948 2210
rect 24892 2146 24948 2158
rect 24556 2100 24612 2110
rect 24220 2098 24612 2100
rect 24220 2046 24558 2098
rect 24610 2046 24612 2098
rect 24220 2044 24612 2046
rect 23548 1652 23604 1662
rect 23324 980 23380 990
rect 23324 886 23380 924
rect 23212 242 23268 252
rect 23548 112 23604 1596
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 24220 1202 24276 2044
rect 24556 2034 24612 2044
rect 24220 1150 24222 1202
rect 24274 1150 24276 1202
rect 24220 1138 24276 1150
rect 24332 1540 24388 1550
rect 24332 756 24388 1484
rect 25004 1428 25060 5182
rect 25116 5236 25172 6300
rect 25228 6132 25284 6142
rect 25228 5572 25284 6076
rect 25228 5506 25284 5516
rect 25340 5346 25396 17276
rect 25452 13748 25508 18284
rect 25900 17778 25956 17790
rect 25900 17726 25902 17778
rect 25954 17726 25956 17778
rect 25788 16884 25844 16894
rect 25788 16790 25844 16828
rect 25900 16324 25956 17726
rect 26124 17668 26180 18284
rect 26236 17668 26292 17678
rect 26124 17612 26236 17668
rect 26236 17574 26292 17612
rect 25900 16258 25956 16268
rect 26124 16548 26180 16558
rect 26124 16324 26180 16492
rect 26124 16258 26180 16268
rect 26124 15090 26180 15102
rect 26124 15038 26126 15090
rect 26178 15038 26180 15090
rect 25676 14642 25732 14654
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25564 14530 25620 14542
rect 25564 14478 25566 14530
rect 25618 14478 25620 14530
rect 25564 14158 25620 14478
rect 25676 14532 25732 14590
rect 26124 14642 26180 15038
rect 26124 14590 26126 14642
rect 26178 14590 26180 14642
rect 26124 14578 26180 14590
rect 25676 14466 25732 14476
rect 25900 14420 25956 14430
rect 25564 14102 25844 14158
rect 25452 13692 25732 13748
rect 25452 13524 25508 13534
rect 25452 13430 25508 13468
rect 25564 12516 25620 12526
rect 25452 12180 25508 12190
rect 25452 11844 25508 12124
rect 25564 12178 25620 12460
rect 25564 12126 25566 12178
rect 25618 12126 25620 12178
rect 25564 12114 25620 12126
rect 25564 11844 25620 11854
rect 25452 11788 25564 11844
rect 25564 11506 25620 11788
rect 25564 11454 25566 11506
rect 25618 11454 25620 11506
rect 25564 11442 25620 11454
rect 25452 11396 25508 11406
rect 25452 10724 25508 11340
rect 25452 10658 25508 10668
rect 25676 10612 25732 13692
rect 25788 13412 25844 14102
rect 25900 13746 25956 14364
rect 25900 13694 25902 13746
rect 25954 13694 25956 13746
rect 25900 13636 25956 13694
rect 25900 13570 25956 13580
rect 26236 13636 26292 13646
rect 25788 13346 25844 13356
rect 26124 13524 26180 13534
rect 25788 13188 25844 13198
rect 25788 13094 25844 13132
rect 25900 12628 25956 12638
rect 25676 10546 25732 10556
rect 25788 11172 25844 11182
rect 25788 10388 25844 11116
rect 25452 8818 25508 8830
rect 25452 8766 25454 8818
rect 25506 8766 25508 8818
rect 25452 8372 25508 8766
rect 25452 8306 25508 8316
rect 25452 8148 25508 8158
rect 25452 7812 25508 8092
rect 25676 8146 25732 8158
rect 25676 8094 25678 8146
rect 25730 8094 25732 8146
rect 25676 8036 25732 8094
rect 25676 7970 25732 7980
rect 25452 7474 25508 7756
rect 25452 7422 25454 7474
rect 25506 7422 25508 7474
rect 25452 7410 25508 7422
rect 25676 7250 25732 7262
rect 25676 7198 25678 7250
rect 25730 7198 25732 7250
rect 25564 6804 25620 6814
rect 25676 6804 25732 7198
rect 25564 6802 25732 6804
rect 25564 6750 25566 6802
rect 25618 6750 25732 6802
rect 25564 6748 25732 6750
rect 25564 6738 25620 6748
rect 25452 6468 25508 6478
rect 25452 5906 25508 6412
rect 25788 6244 25844 10332
rect 25900 8036 25956 12572
rect 26124 12516 26180 13468
rect 26236 12852 26292 13580
rect 26236 12758 26292 12796
rect 26012 10948 26068 10958
rect 26012 10610 26068 10892
rect 26012 10558 26014 10610
rect 26066 10558 26068 10610
rect 26012 10388 26068 10558
rect 26012 10322 26068 10332
rect 26124 8932 26180 12460
rect 26348 12180 26404 18732
rect 26460 17220 26516 17230
rect 26460 14084 26516 17164
rect 26460 14018 26516 14028
rect 26572 12404 26628 19852
rect 26684 20132 26740 20142
rect 26684 18338 26740 20076
rect 26796 18788 26852 21980
rect 26908 23492 26964 23502
rect 26908 19346 26964 23436
rect 27020 21810 27076 23886
rect 27020 21758 27022 21810
rect 27074 21758 27076 21810
rect 27020 21746 27076 21758
rect 26908 19294 26910 19346
rect 26962 19294 26964 19346
rect 26908 19282 26964 19294
rect 26796 18722 26852 18732
rect 26684 18286 26686 18338
rect 26738 18286 26740 18338
rect 26684 18274 26740 18286
rect 26796 18228 26852 18238
rect 26796 16882 26852 18172
rect 26796 16830 26798 16882
rect 26850 16830 26852 16882
rect 26684 16324 26740 16334
rect 26684 16098 26740 16268
rect 26796 16212 26852 16830
rect 26796 16146 26852 16156
rect 26684 16046 26686 16098
rect 26738 16046 26740 16098
rect 26684 15988 26740 16046
rect 26684 15922 26740 15932
rect 26908 15988 26964 15998
rect 26908 14980 26964 15932
rect 26796 14924 26964 14980
rect 26796 14530 26852 14924
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26796 14466 26852 14478
rect 26348 12114 26404 12124
rect 26460 12348 26628 12404
rect 26460 11060 26516 12348
rect 26572 12178 26628 12190
rect 26572 12126 26574 12178
rect 26626 12126 26628 12178
rect 26572 11732 26628 12126
rect 26572 11284 26628 11676
rect 26572 11218 26628 11228
rect 26684 12180 26740 12190
rect 26684 11172 26740 12124
rect 26796 11396 26852 11406
rect 26796 11302 26852 11340
rect 26684 11116 26852 11172
rect 26460 11004 26740 11060
rect 26348 10836 26404 10846
rect 26124 8876 26292 8932
rect 26124 8372 26180 8382
rect 26012 8260 26068 8270
rect 26012 8166 26068 8204
rect 25900 7970 25956 7980
rect 26124 7700 26180 8316
rect 26124 7474 26180 7644
rect 26124 7422 26126 7474
rect 26178 7422 26180 7474
rect 25900 6692 25956 6702
rect 25900 6598 25956 6636
rect 25900 6468 25956 6478
rect 25900 6466 26068 6468
rect 25900 6414 25902 6466
rect 25954 6414 26068 6466
rect 25900 6412 26068 6414
rect 25900 6402 25956 6412
rect 25788 6188 25956 6244
rect 25452 5854 25454 5906
rect 25506 5854 25508 5906
rect 25452 5842 25508 5854
rect 25676 5684 25732 5694
rect 25676 5682 25844 5684
rect 25676 5630 25678 5682
rect 25730 5630 25844 5682
rect 25676 5628 25844 5630
rect 25676 5618 25732 5628
rect 25340 5294 25342 5346
rect 25394 5294 25396 5346
rect 25340 5282 25396 5294
rect 25564 5572 25620 5582
rect 25116 4562 25172 5180
rect 25116 4510 25118 4562
rect 25170 4510 25172 4562
rect 25116 4498 25172 4510
rect 25564 3778 25620 5516
rect 25788 4564 25844 5628
rect 25900 5460 25956 6188
rect 25900 5394 25956 5404
rect 26012 5348 26068 6412
rect 26124 5906 26180 7422
rect 26236 6804 26292 8876
rect 26348 8372 26404 10780
rect 26572 10836 26628 10846
rect 26348 8306 26404 8316
rect 26460 10612 26516 10622
rect 26460 8258 26516 10556
rect 26572 10500 26628 10780
rect 26572 10434 26628 10444
rect 26684 8708 26740 11004
rect 26684 8642 26740 8652
rect 26684 8372 26740 8382
rect 26460 8206 26462 8258
rect 26514 8206 26516 8258
rect 26460 8194 26516 8206
rect 26572 8370 26740 8372
rect 26572 8318 26686 8370
rect 26738 8318 26740 8370
rect 26572 8316 26740 8318
rect 26460 7140 26516 7150
rect 26236 6748 26404 6804
rect 26236 6578 26292 6590
rect 26236 6526 26238 6578
rect 26290 6526 26292 6578
rect 26236 6468 26292 6526
rect 26236 6402 26292 6412
rect 26348 6020 26404 6748
rect 26460 6468 26516 7084
rect 26460 6402 26516 6412
rect 26348 5954 26404 5964
rect 26124 5854 26126 5906
rect 26178 5854 26180 5906
rect 26124 5842 26180 5854
rect 26572 5796 26628 8316
rect 26684 8306 26740 8316
rect 26684 7700 26740 7710
rect 26684 6690 26740 7644
rect 26796 7474 26852 11116
rect 26796 7422 26798 7474
rect 26850 7422 26852 7474
rect 26796 7410 26852 7422
rect 26908 7476 26964 14924
rect 27020 14196 27076 14206
rect 27020 12852 27076 14140
rect 27020 12786 27076 12796
rect 27020 11732 27076 11742
rect 27020 7812 27076 11676
rect 27132 9380 27188 27468
rect 27244 19460 27300 30044
rect 27804 29650 27860 30156
rect 27804 29598 27806 29650
rect 27858 29598 27860 29650
rect 27804 29586 27860 29598
rect 27916 30100 27972 30110
rect 27916 29540 27972 30044
rect 27916 29474 27972 29484
rect 27580 28756 27636 28766
rect 27580 28662 27636 28700
rect 28028 28754 28084 30940
rect 28028 28702 28030 28754
rect 28082 28702 28084 28754
rect 28028 28690 28084 28702
rect 27580 28084 27636 28094
rect 27580 27298 27636 28028
rect 28140 28084 28196 32396
rect 28140 28018 28196 28028
rect 27580 27246 27582 27298
rect 27634 27246 27636 27298
rect 27580 27234 27636 27246
rect 27692 27858 27748 27870
rect 27692 27806 27694 27858
rect 27746 27806 27748 27858
rect 27356 27062 27412 27074
rect 27692 27064 27748 27806
rect 27916 27748 27972 27758
rect 27916 27654 27972 27692
rect 28028 27076 28084 27086
rect 27356 27010 27358 27062
rect 27410 27010 27412 27062
rect 27356 26964 27412 27010
rect 27636 27008 27748 27064
rect 27916 27074 28084 27076
rect 27916 27022 28030 27074
rect 28082 27022 28084 27074
rect 27916 27020 28084 27022
rect 27636 26964 27692 27008
rect 27356 24612 27412 26908
rect 27356 24546 27412 24556
rect 27468 26908 27692 26964
rect 27468 20804 27524 26908
rect 27804 26292 27860 26302
rect 27804 26198 27860 26236
rect 27692 25732 27748 25742
rect 27916 25732 27972 27020
rect 28028 27010 28084 27020
rect 27692 25730 27972 25732
rect 27692 25678 27694 25730
rect 27746 25678 27972 25730
rect 27692 25676 27972 25678
rect 28028 25844 28084 25854
rect 27692 25666 27748 25676
rect 27916 24724 27972 24734
rect 27804 24612 27860 24622
rect 27804 24518 27860 24556
rect 27916 24500 27972 24668
rect 27692 24388 27748 24398
rect 27748 24332 27860 24388
rect 27692 24322 27748 24332
rect 27692 23940 27748 23950
rect 27692 23846 27748 23884
rect 27692 22596 27748 22606
rect 27692 22502 27748 22540
rect 27804 21924 27860 24332
rect 27916 23940 27972 24444
rect 27916 23874 27972 23884
rect 27804 21858 27860 21868
rect 27804 21700 27860 21710
rect 27692 21476 27748 21486
rect 27580 20804 27636 20814
rect 27468 20802 27636 20804
rect 27468 20750 27582 20802
rect 27634 20750 27636 20802
rect 27468 20748 27636 20750
rect 27468 20356 27524 20366
rect 27244 19404 27412 19460
rect 27244 19236 27300 19246
rect 27244 19142 27300 19180
rect 27356 18116 27412 19404
rect 27356 18050 27412 18060
rect 27356 17668 27412 17678
rect 27244 16548 27300 16558
rect 27244 16212 27300 16492
rect 27244 16118 27300 16156
rect 27244 15204 27300 15214
rect 27244 14532 27300 15148
rect 27244 14466 27300 14476
rect 27356 14196 27412 17612
rect 27244 12852 27300 12862
rect 27356 12852 27412 14140
rect 27244 12850 27412 12852
rect 27244 12798 27246 12850
rect 27298 12798 27412 12850
rect 27244 12796 27412 12798
rect 27244 12786 27300 12796
rect 27244 11282 27300 11294
rect 27244 11230 27246 11282
rect 27298 11230 27300 11282
rect 27244 11172 27300 11230
rect 27244 11106 27300 11116
rect 27356 10052 27412 12796
rect 27356 9986 27412 9996
rect 27468 9828 27524 20300
rect 27580 12068 27636 20748
rect 27692 19572 27748 21420
rect 27804 20692 27860 21644
rect 27804 20626 27860 20636
rect 27692 19506 27748 19516
rect 27916 19684 27972 19694
rect 27916 19458 27972 19628
rect 27916 19406 27918 19458
rect 27970 19406 27972 19458
rect 27916 19394 27972 19406
rect 27692 19234 27748 19246
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 18564 27748 19182
rect 27804 19236 27860 19246
rect 27804 18674 27860 19180
rect 27804 18622 27806 18674
rect 27858 18622 27860 18674
rect 27804 18610 27860 18622
rect 27692 18498 27748 18508
rect 28028 17780 28084 25788
rect 28140 22484 28196 22494
rect 28140 22390 28196 22428
rect 28252 21700 28308 32620
rect 28364 31108 28420 37212
rect 28588 34804 28644 38780
rect 28700 38770 28756 38780
rect 28700 38052 28756 38062
rect 28756 37996 28868 38052
rect 28700 37958 28756 37996
rect 28812 37266 28868 37996
rect 28812 37214 28814 37266
rect 28866 37214 28868 37266
rect 28812 37202 28868 37214
rect 28700 35700 28756 35710
rect 28700 35698 28868 35700
rect 28700 35646 28702 35698
rect 28754 35646 28868 35698
rect 28700 35644 28868 35646
rect 28700 35634 28756 35644
rect 28700 35476 28756 35486
rect 28700 35026 28756 35420
rect 28812 35140 28868 35644
rect 28812 35074 28868 35084
rect 28700 34974 28702 35026
rect 28754 34974 28756 35026
rect 28700 34962 28756 34974
rect 28924 34916 28980 39004
rect 29036 38052 29092 38062
rect 29036 37958 29092 37996
rect 28588 34748 28756 34804
rect 28476 33684 28532 33694
rect 28476 33348 28532 33628
rect 28588 33348 28644 33358
rect 28476 33346 28644 33348
rect 28476 33294 28590 33346
rect 28642 33294 28644 33346
rect 28476 33292 28644 33294
rect 28588 31778 28644 33292
rect 28588 31726 28590 31778
rect 28642 31726 28644 31778
rect 28588 31714 28644 31726
rect 28364 30322 28420 31052
rect 28700 30548 28756 34748
rect 28812 34020 28868 34030
rect 28812 32674 28868 33964
rect 28924 33684 28980 34860
rect 28924 33618 28980 33628
rect 29036 37156 29092 37166
rect 28812 32622 28814 32674
rect 28866 32622 28868 32674
rect 28812 32004 28868 32622
rect 28924 32340 28980 32350
rect 28924 32246 28980 32284
rect 28812 31938 28868 31948
rect 28924 31780 28980 31790
rect 28924 31106 28980 31724
rect 29036 31444 29092 37100
rect 29148 36932 29204 39228
rect 29484 39172 29540 39566
rect 29708 39284 29764 44604
rect 29820 43428 29876 44942
rect 29932 44322 29988 45836
rect 30156 45668 30212 48300
rect 30268 48242 30324 48254
rect 30268 48190 30270 48242
rect 30322 48190 30324 48242
rect 30268 47348 30324 48190
rect 30380 47572 30436 47582
rect 30380 47478 30436 47516
rect 30268 47292 30436 47348
rect 30268 46676 30324 46686
rect 30380 46676 30436 47292
rect 30492 47012 30548 48748
rect 30716 48692 30772 48702
rect 30716 48130 30772 48636
rect 30716 48078 30718 48130
rect 30770 48078 30772 48130
rect 30716 47908 30772 48078
rect 30716 47842 30772 47852
rect 30716 47572 30772 47582
rect 30716 47458 30772 47516
rect 30716 47406 30718 47458
rect 30770 47406 30772 47458
rect 30716 47394 30772 47406
rect 30828 47460 30884 47470
rect 30716 47236 30772 47246
rect 30716 47142 30772 47180
rect 30492 46946 30548 46956
rect 30268 46674 30436 46676
rect 30268 46622 30270 46674
rect 30322 46622 30436 46674
rect 30268 46620 30436 46622
rect 30268 46610 30324 46620
rect 30156 45602 30212 45612
rect 30044 45444 30100 45454
rect 30044 44884 30100 45388
rect 30156 45108 30212 45118
rect 30156 45014 30212 45052
rect 30380 45108 30436 46620
rect 30604 46676 30660 46686
rect 30660 46620 30772 46676
rect 30604 46610 30660 46620
rect 30716 46562 30772 46620
rect 30716 46510 30718 46562
rect 30770 46510 30772 46562
rect 30716 46498 30772 46510
rect 30604 46452 30660 46462
rect 30604 46004 30660 46396
rect 30604 46002 30772 46004
rect 30604 45950 30606 46002
rect 30658 45950 30772 46002
rect 30604 45948 30772 45950
rect 30604 45938 30660 45948
rect 30380 45042 30436 45052
rect 30492 45892 30548 45902
rect 30044 44818 30100 44828
rect 29932 44270 29934 44322
rect 29986 44270 29988 44322
rect 29932 43540 29988 44270
rect 29932 43474 29988 43484
rect 30492 44322 30548 45836
rect 30604 45668 30660 45678
rect 30604 45574 30660 45612
rect 30716 45444 30772 45948
rect 30828 45892 30884 47404
rect 30828 45826 30884 45836
rect 30716 45378 30772 45388
rect 30940 45332 30996 49420
rect 31388 49250 31444 49644
rect 31388 49198 31390 49250
rect 31442 49198 31444 49250
rect 31388 49186 31444 49198
rect 31164 49026 31220 49038
rect 31164 48974 31166 49026
rect 31218 48974 31220 49026
rect 31164 47460 31220 48974
rect 31500 49028 31556 50372
rect 31724 50148 31780 50542
rect 31836 50484 31892 52222
rect 32172 51828 32228 51838
rect 32172 51378 32228 51772
rect 32172 51326 32174 51378
rect 32226 51326 32228 51378
rect 32172 51314 32228 51326
rect 31836 50418 31892 50428
rect 31948 51156 32004 51166
rect 31948 50260 32004 51100
rect 32172 51156 32228 51166
rect 31724 50082 31780 50092
rect 31836 50204 32116 50260
rect 31500 48962 31556 48972
rect 31612 49700 31668 49710
rect 31276 48916 31332 48926
rect 31276 48822 31332 48860
rect 31612 48914 31668 49644
rect 31836 49698 31892 50204
rect 31836 49646 31838 49698
rect 31890 49646 31892 49698
rect 31836 49634 31892 49646
rect 31948 49700 32004 49710
rect 31612 48862 31614 48914
rect 31666 48862 31668 48914
rect 31612 48850 31668 48862
rect 31500 48804 31556 48814
rect 31388 47684 31444 47694
rect 31388 47590 31444 47628
rect 30940 45266 30996 45276
rect 31052 47458 31220 47460
rect 31052 47406 31166 47458
rect 31218 47406 31220 47458
rect 31052 47404 31220 47406
rect 31052 46340 31108 47404
rect 31164 47394 31220 47404
rect 31276 47460 31332 47470
rect 31276 47366 31332 47404
rect 30940 45108 30996 45118
rect 30940 45014 30996 45052
rect 30716 44772 30772 44782
rect 30604 44436 30660 44446
rect 30604 44342 30660 44380
rect 30492 44270 30494 44322
rect 30546 44270 30548 44322
rect 29820 41748 29876 43372
rect 30268 43316 30324 43326
rect 30268 43222 30324 43260
rect 29820 41682 29876 41692
rect 30044 42756 30100 42766
rect 29372 39116 29540 39172
rect 29596 39228 29764 39284
rect 29820 41412 29876 41422
rect 29260 38724 29316 38762
rect 29260 38658 29316 38668
rect 29260 38276 29316 38286
rect 29260 38182 29316 38220
rect 29372 37492 29428 39116
rect 29148 36866 29204 36876
rect 29260 37436 29428 37492
rect 29484 38948 29540 38958
rect 29148 35476 29204 35486
rect 29148 35382 29204 35420
rect 29260 34804 29316 37436
rect 29372 37266 29428 37278
rect 29372 37214 29374 37266
rect 29426 37214 29428 37266
rect 29372 37156 29428 37214
rect 29372 37090 29428 37100
rect 29484 37154 29540 38892
rect 29484 37102 29486 37154
rect 29538 37102 29540 37154
rect 29484 37090 29540 37102
rect 29484 36484 29540 36494
rect 29484 34916 29540 36428
rect 29596 35252 29652 39228
rect 29820 38724 29876 41356
rect 30044 41186 30100 42700
rect 30492 41748 30548 44270
rect 30604 44100 30660 44110
rect 30604 44006 30660 44044
rect 30716 43876 30772 44716
rect 30940 44772 30996 44782
rect 30940 44100 30996 44716
rect 31052 44436 31108 46284
rect 31164 47124 31220 47134
rect 31164 46114 31220 47068
rect 31164 46062 31166 46114
rect 31218 46062 31220 46114
rect 31164 44772 31220 46062
rect 31276 46116 31332 46126
rect 31276 46022 31332 46060
rect 31388 45892 31444 45902
rect 31388 45798 31444 45836
rect 31164 44706 31220 44716
rect 31388 44882 31444 44894
rect 31388 44830 31390 44882
rect 31442 44830 31444 44882
rect 31388 44772 31444 44830
rect 31388 44706 31444 44716
rect 31276 44660 31332 44670
rect 31276 44546 31332 44604
rect 31276 44494 31278 44546
rect 31330 44494 31332 44546
rect 31276 44482 31332 44494
rect 31388 44548 31444 44558
rect 31388 44454 31444 44492
rect 31164 44436 31220 44446
rect 31052 44380 31164 44436
rect 31164 44342 31220 44380
rect 31388 44324 31444 44334
rect 30940 44034 30996 44044
rect 31276 44212 31332 44222
rect 30604 43820 30772 43876
rect 30604 42082 30660 43820
rect 30828 43314 30884 43326
rect 30828 43262 30830 43314
rect 30882 43262 30884 43314
rect 30604 42030 30606 42082
rect 30658 42030 30660 42082
rect 30604 42018 30660 42030
rect 30716 42866 30772 42878
rect 30716 42814 30718 42866
rect 30770 42814 30772 42866
rect 30716 41860 30772 42814
rect 30828 42754 30884 43262
rect 30828 42702 30830 42754
rect 30882 42702 30884 42754
rect 30828 42690 30884 42702
rect 30940 43092 30996 43102
rect 30716 41794 30772 41804
rect 30492 41692 30660 41748
rect 30044 41134 30046 41186
rect 30098 41134 30100 41186
rect 29820 38658 29876 38668
rect 29932 40964 29988 40974
rect 29708 38612 29764 38622
rect 29708 38162 29764 38556
rect 29932 38276 29988 40908
rect 29708 38110 29710 38162
rect 29762 38110 29764 38162
rect 29708 38098 29764 38110
rect 29820 38220 29988 38276
rect 29820 37940 29876 38220
rect 29596 35186 29652 35196
rect 29708 37884 29876 37940
rect 29932 38050 29988 38062
rect 29932 37998 29934 38050
rect 29986 37998 29988 38050
rect 29484 34850 29540 34860
rect 29260 34738 29316 34748
rect 29372 34468 29428 34478
rect 29372 32676 29428 34412
rect 29372 32610 29428 32620
rect 29484 33684 29540 33694
rect 29260 32450 29316 32462
rect 29260 32398 29262 32450
rect 29314 32398 29316 32450
rect 29036 31378 29092 31388
rect 29148 32340 29204 32350
rect 28924 31054 28926 31106
rect 28978 31054 28980 31106
rect 28924 31042 28980 31054
rect 29148 30996 29204 32284
rect 29260 31220 29316 32398
rect 29372 32340 29428 32350
rect 29372 32246 29428 32284
rect 29484 32116 29540 33628
rect 29708 33346 29764 37884
rect 29932 37266 29988 37998
rect 29932 37214 29934 37266
rect 29986 37214 29988 37266
rect 29932 37202 29988 37214
rect 30044 36484 30100 41134
rect 30268 41524 30324 41534
rect 30156 39730 30212 39742
rect 30156 39678 30158 39730
rect 30210 39678 30212 39730
rect 30156 38948 30212 39678
rect 30156 38882 30212 38892
rect 30156 38500 30212 38510
rect 30156 36594 30212 38444
rect 30268 37268 30324 41468
rect 30492 41524 30548 41534
rect 30492 40626 30548 41468
rect 30492 40574 30494 40626
rect 30546 40574 30548 40626
rect 30492 40562 30548 40574
rect 30492 40180 30548 40190
rect 30380 39618 30436 39630
rect 30380 39566 30382 39618
rect 30434 39566 30436 39618
rect 30380 39058 30436 39566
rect 30380 39006 30382 39058
rect 30434 39006 30436 39058
rect 30380 38994 30436 39006
rect 30492 38052 30548 40124
rect 30604 39620 30660 41692
rect 30716 41188 30772 41198
rect 30940 41188 30996 43036
rect 31276 42308 31332 44156
rect 31388 43876 31444 44268
rect 31388 43810 31444 43820
rect 31388 42532 31444 42542
rect 31388 42438 31444 42476
rect 31276 42252 31444 42308
rect 31052 41972 31108 41982
rect 31052 41970 31332 41972
rect 31052 41918 31054 41970
rect 31106 41918 31332 41970
rect 31052 41916 31332 41918
rect 31052 41906 31108 41916
rect 30772 41132 30884 41188
rect 30716 41122 30772 41132
rect 30604 39554 30660 39564
rect 30828 39956 30884 41132
rect 30940 41122 30996 41132
rect 31276 41524 31332 41916
rect 30940 40964 30996 40974
rect 30940 40514 30996 40908
rect 30940 40462 30942 40514
rect 30994 40462 30996 40514
rect 30940 40450 30996 40462
rect 31276 40402 31332 41468
rect 31276 40350 31278 40402
rect 31330 40350 31332 40402
rect 31276 40338 31332 40350
rect 31388 40292 31444 42252
rect 31388 40226 31444 40236
rect 31500 41970 31556 48748
rect 31836 48804 31892 48814
rect 31836 48710 31892 48748
rect 31612 48244 31668 48254
rect 31612 47458 31668 48188
rect 31612 47406 31614 47458
rect 31666 47406 31668 47458
rect 31612 47124 31668 47406
rect 31836 48018 31892 48030
rect 31836 47966 31838 48018
rect 31890 47966 31892 48018
rect 31836 47458 31892 47966
rect 31836 47406 31838 47458
rect 31890 47406 31892 47458
rect 31836 47394 31892 47406
rect 31948 47124 32004 49644
rect 31612 47058 31668 47068
rect 31724 47068 32004 47124
rect 31612 45892 31668 45902
rect 31724 45892 31780 47068
rect 31612 45890 31780 45892
rect 31612 45838 31614 45890
rect 31666 45838 31780 45890
rect 31612 45836 31780 45838
rect 31948 46450 32004 46462
rect 31948 46398 31950 46450
rect 32002 46398 32004 46450
rect 31612 45826 31668 45836
rect 31612 45668 31668 45678
rect 31612 44322 31668 45612
rect 31836 45668 31892 45678
rect 31836 45574 31892 45612
rect 31612 44270 31614 44322
rect 31666 44270 31668 44322
rect 31612 44258 31668 44270
rect 31724 44772 31780 44782
rect 31612 43540 31668 43550
rect 31612 42532 31668 43484
rect 31724 42756 31780 44716
rect 31948 44548 32004 46398
rect 32060 46004 32116 50204
rect 32060 45938 32116 45948
rect 31948 44482 32004 44492
rect 32060 44996 32116 45006
rect 31836 44324 31892 44334
rect 31836 44230 31892 44268
rect 31948 44212 32004 44222
rect 31948 43988 32004 44156
rect 31948 43922 32004 43932
rect 32060 43426 32116 44940
rect 32060 43374 32062 43426
rect 32114 43374 32116 43426
rect 31724 42700 31892 42756
rect 31724 42532 31780 42542
rect 31612 42530 31780 42532
rect 31612 42478 31726 42530
rect 31778 42478 31780 42530
rect 31612 42476 31780 42478
rect 31724 42466 31780 42476
rect 31500 41918 31502 41970
rect 31554 41918 31556 41970
rect 30492 38050 30772 38052
rect 30492 37998 30494 38050
rect 30546 37998 30772 38050
rect 30492 37996 30772 37998
rect 30492 37986 30548 37996
rect 30604 37380 30660 37390
rect 30492 37268 30548 37278
rect 30268 37266 30548 37268
rect 30268 37214 30494 37266
rect 30546 37214 30548 37266
rect 30268 37212 30548 37214
rect 30156 36542 30158 36594
rect 30210 36542 30212 36594
rect 30156 36530 30212 36542
rect 30044 36418 30100 36428
rect 29820 36370 29876 36382
rect 29820 36318 29822 36370
rect 29874 36318 29876 36370
rect 29820 35140 29876 36318
rect 29820 35074 29876 35084
rect 30044 36036 30100 36046
rect 29820 34580 29876 34590
rect 29820 34242 29876 34524
rect 29820 34190 29822 34242
rect 29874 34190 29876 34242
rect 29820 34178 29876 34190
rect 29708 33294 29710 33346
rect 29762 33294 29764 33346
rect 29260 31154 29316 31164
rect 29372 32060 29540 32116
rect 29596 32338 29652 32350
rect 29596 32286 29598 32338
rect 29650 32286 29652 32338
rect 29148 30930 29204 30940
rect 28812 30772 28868 30782
rect 28812 30678 28868 30716
rect 29036 30770 29092 30782
rect 29036 30718 29038 30770
rect 29090 30718 29092 30770
rect 28700 30492 28868 30548
rect 28364 30270 28366 30322
rect 28418 30270 28420 30322
rect 28364 29988 28420 30270
rect 28364 29922 28420 29932
rect 28588 29540 28644 29550
rect 28364 28756 28420 28766
rect 28364 28642 28420 28700
rect 28364 28590 28366 28642
rect 28418 28590 28420 28642
rect 28364 28578 28420 28590
rect 28476 28532 28532 28542
rect 28588 28532 28644 29484
rect 28532 28476 28644 28532
rect 28700 29426 28756 29438
rect 28700 29374 28702 29426
rect 28754 29374 28756 29426
rect 28476 28466 28532 28476
rect 28252 21364 28308 21644
rect 28252 21298 28308 21308
rect 28364 28420 28420 28430
rect 28364 24612 28420 28364
rect 28700 28196 28756 29374
rect 28812 28420 28868 30492
rect 29036 30212 29092 30718
rect 29260 30772 29316 30782
rect 29260 30678 29316 30716
rect 29036 30146 29092 30156
rect 29260 30324 29316 30334
rect 29260 29652 29316 30268
rect 29260 29586 29316 29596
rect 29148 29202 29204 29214
rect 29148 29150 29150 29202
rect 29202 29150 29204 29202
rect 29148 28980 29204 29150
rect 29148 28914 29204 28924
rect 29036 28868 29092 28878
rect 29036 28774 29092 28812
rect 28924 28756 28980 28766
rect 28924 28642 28980 28700
rect 28924 28590 28926 28642
rect 28978 28590 28980 28642
rect 28924 28578 28980 28590
rect 28812 28364 29092 28420
rect 28756 28140 28868 28196
rect 28700 28130 28756 28140
rect 28700 27188 28756 27198
rect 28588 27074 28644 27086
rect 28588 27022 28590 27074
rect 28642 27022 28644 27074
rect 28476 26740 28532 26750
rect 28588 26740 28644 27022
rect 28532 26684 28644 26740
rect 28476 26674 28532 26684
rect 28588 25956 28644 26684
rect 28700 26740 28756 27132
rect 28700 26402 28756 26684
rect 28700 26350 28702 26402
rect 28754 26350 28756 26402
rect 28700 26338 28756 26350
rect 28588 25890 28644 25900
rect 28588 25508 28644 25518
rect 28476 24612 28532 24622
rect 28364 24610 28532 24612
rect 28364 24558 28478 24610
rect 28530 24558 28532 24610
rect 28364 24556 28532 24558
rect 28364 21252 28420 24556
rect 28476 24546 28532 24556
rect 28588 23156 28644 25452
rect 28812 25506 28868 28140
rect 28812 25454 28814 25506
rect 28866 25454 28868 25506
rect 28812 25442 28868 25454
rect 28924 27860 28980 27870
rect 28812 24722 28868 24734
rect 28812 24670 28814 24722
rect 28866 24670 28868 24722
rect 28700 24276 28756 24286
rect 28700 23940 28756 24220
rect 28700 23846 28756 23884
rect 28588 23090 28644 23100
rect 28700 23268 28756 23278
rect 28588 22370 28644 22382
rect 28588 22318 28590 22370
rect 28642 22318 28644 22370
rect 28476 21700 28532 21710
rect 28476 21606 28532 21644
rect 28588 21588 28644 22318
rect 28588 21522 28644 21532
rect 28588 21364 28644 21374
rect 28364 21196 28532 21252
rect 28364 20692 28420 20702
rect 28364 20598 28420 20636
rect 28364 19236 28420 19246
rect 28364 19142 28420 19180
rect 27916 17724 28084 17780
rect 27804 14532 27860 14542
rect 27916 14532 27972 17724
rect 28364 17666 28420 17678
rect 28364 17614 28366 17666
rect 28418 17614 28420 17666
rect 28028 17556 28084 17566
rect 28028 17462 28084 17500
rect 28364 16322 28420 17614
rect 28364 16270 28366 16322
rect 28418 16270 28420 16322
rect 28364 16258 28420 16270
rect 28476 15148 28532 21196
rect 28588 17444 28644 21308
rect 28700 20914 28756 23212
rect 28812 22596 28868 24670
rect 28812 22530 28868 22540
rect 28924 22370 28980 27804
rect 29036 26628 29092 28364
rect 29036 26562 29092 26572
rect 29036 26292 29092 26302
rect 29036 26198 29092 26236
rect 29260 25732 29316 25742
rect 29260 25638 29316 25676
rect 29260 24724 29316 24734
rect 29372 24724 29428 32060
rect 29596 32004 29652 32286
rect 29596 31938 29652 31948
rect 29596 31780 29652 31790
rect 29708 31780 29764 33294
rect 29596 31778 29764 31780
rect 29596 31726 29598 31778
rect 29650 31726 29764 31778
rect 29596 31724 29764 31726
rect 29932 32562 29988 32574
rect 29932 32510 29934 32562
rect 29986 32510 29988 32562
rect 29484 31668 29540 31678
rect 29484 30436 29540 31612
rect 29596 31332 29652 31724
rect 29596 31266 29652 31276
rect 29932 31108 29988 32510
rect 30044 32340 30100 35980
rect 30268 35476 30324 35486
rect 30268 35382 30324 35420
rect 30044 32274 30100 32284
rect 30156 34916 30212 34926
rect 30156 31444 30212 34860
rect 30380 34916 30436 34926
rect 30380 34822 30436 34860
rect 30268 34132 30324 34142
rect 30268 34038 30324 34076
rect 30492 33908 30548 37212
rect 30604 35810 30660 37324
rect 30604 35758 30606 35810
rect 30658 35758 30660 35810
rect 30604 34468 30660 35758
rect 30604 34402 30660 34412
rect 30380 33852 30548 33908
rect 30604 34130 30660 34142
rect 30604 34078 30606 34130
rect 30658 34078 30660 34130
rect 30380 32788 30436 33852
rect 30380 32722 30436 32732
rect 30492 33684 30548 33694
rect 30492 32452 30548 33628
rect 30604 33572 30660 34078
rect 30604 33506 30660 33516
rect 30380 32450 30548 32452
rect 30380 32398 30494 32450
rect 30546 32398 30548 32450
rect 30380 32396 30548 32398
rect 30380 32116 30436 32396
rect 30492 32386 30548 32396
rect 30604 32788 30660 32798
rect 30380 32050 30436 32060
rect 30492 32004 30548 32014
rect 30156 31388 30324 31444
rect 30156 31220 30212 31230
rect 29932 31106 30100 31108
rect 29932 31054 29934 31106
rect 29986 31054 30100 31106
rect 29932 31052 30100 31054
rect 29932 31042 29988 31052
rect 29820 30996 29876 31006
rect 29820 30436 29876 30940
rect 30044 30996 30100 31052
rect 30044 30930 30100 30940
rect 30044 30772 30100 30782
rect 29932 30436 29988 30446
rect 29820 30434 29988 30436
rect 29820 30382 29934 30434
rect 29986 30382 29988 30434
rect 29820 30380 29988 30382
rect 29484 30370 29540 30380
rect 29932 30370 29988 30380
rect 30044 30434 30100 30716
rect 30044 30382 30046 30434
rect 30098 30382 30100 30434
rect 30044 30370 30100 30382
rect 30156 30434 30212 31164
rect 30156 30382 30158 30434
rect 30210 30382 30212 30434
rect 30156 30370 30212 30382
rect 29484 30212 29540 30222
rect 30268 30212 30324 31388
rect 30380 31108 30436 31118
rect 30380 30882 30436 31052
rect 30380 30830 30382 30882
rect 30434 30830 30436 30882
rect 30380 30818 30436 30830
rect 30492 30322 30548 31948
rect 30492 30270 30494 30322
rect 30546 30270 30548 30322
rect 30492 30258 30548 30270
rect 29484 30118 29540 30156
rect 30156 30156 30324 30212
rect 30380 30212 30436 30222
rect 30044 30100 30100 30110
rect 29708 28644 29764 28654
rect 29708 28550 29764 28588
rect 30044 28642 30100 30044
rect 30044 28590 30046 28642
rect 30098 28590 30100 28642
rect 30044 28578 30100 28590
rect 30156 27858 30212 30156
rect 30380 30118 30436 30156
rect 30604 30100 30660 32732
rect 30492 30044 30660 30100
rect 30268 29202 30324 29214
rect 30268 29150 30270 29202
rect 30322 29150 30324 29202
rect 30268 28644 30324 29150
rect 30268 28578 30324 28588
rect 30156 27806 30158 27858
rect 30210 27806 30212 27858
rect 29596 27636 29652 27646
rect 29596 27076 29652 27580
rect 29596 26982 29652 27020
rect 29708 26964 29764 26974
rect 29708 26628 29764 26908
rect 29708 26516 29764 26572
rect 29596 26460 29764 26516
rect 29820 26516 29876 26526
rect 29596 26290 29652 26460
rect 29596 26238 29598 26290
rect 29650 26238 29652 26290
rect 29596 26226 29652 26238
rect 29708 26292 29764 26302
rect 29708 26178 29764 26236
rect 29708 26126 29710 26178
rect 29762 26126 29764 26178
rect 29708 26114 29764 26126
rect 29260 24722 29428 24724
rect 29260 24670 29262 24722
rect 29314 24670 29428 24722
rect 29260 24668 29428 24670
rect 29036 24388 29092 24398
rect 29036 23604 29092 24332
rect 29036 23538 29092 23548
rect 29260 23548 29316 24668
rect 29484 24498 29540 24510
rect 29484 24446 29486 24498
rect 29538 24446 29540 24498
rect 29484 24388 29540 24446
rect 29484 24322 29540 24332
rect 29708 23940 29764 23950
rect 29484 23938 29764 23940
rect 29484 23886 29710 23938
rect 29762 23886 29764 23938
rect 29484 23884 29764 23886
rect 29484 23548 29540 23884
rect 29708 23874 29764 23884
rect 29260 23492 29428 23548
rect 29484 23492 29764 23548
rect 28924 22318 28926 22370
rect 28978 22318 28980 22370
rect 28812 21588 28868 21626
rect 28812 21522 28868 21532
rect 28924 21252 28980 22318
rect 29036 23154 29092 23166
rect 29036 23102 29038 23154
rect 29090 23102 29092 23154
rect 29036 22820 29092 23102
rect 29036 21364 29092 22764
rect 29148 22484 29204 22494
rect 29148 22390 29204 22428
rect 29036 21298 29092 21308
rect 29148 21812 29204 21822
rect 29148 21588 29204 21756
rect 29260 21588 29316 21598
rect 29148 21586 29316 21588
rect 29148 21534 29262 21586
rect 29314 21534 29316 21586
rect 29148 21532 29316 21534
rect 28700 20862 28702 20914
rect 28754 20862 28756 20914
rect 28700 20850 28756 20862
rect 28812 21196 28980 21252
rect 28700 20692 28756 20702
rect 28700 20018 28756 20636
rect 28700 19966 28702 20018
rect 28754 19966 28756 20018
rect 28700 19124 28756 19966
rect 28700 19058 28756 19068
rect 28700 18564 28756 18574
rect 28700 18470 28756 18508
rect 28588 17388 28756 17444
rect 28700 16994 28756 17388
rect 28700 16942 28702 16994
rect 28754 16942 28756 16994
rect 27804 14530 27972 14532
rect 27804 14478 27806 14530
rect 27858 14478 27972 14530
rect 27804 14476 27972 14478
rect 28364 15092 28532 15148
rect 28588 16884 28644 16894
rect 27692 13076 27748 13086
rect 27692 12982 27748 13020
rect 27804 12516 27860 14476
rect 28252 13524 28308 13534
rect 27804 12450 27860 12460
rect 28140 13412 28196 13422
rect 27580 12012 27860 12068
rect 27692 11844 27748 11854
rect 27580 11396 27636 11406
rect 27580 11302 27636 11340
rect 27468 9734 27524 9772
rect 27132 9324 27636 9380
rect 27020 7746 27076 7756
rect 27132 8258 27188 8270
rect 27132 8206 27134 8258
rect 27186 8206 27188 8258
rect 27132 7700 27188 8206
rect 27132 7634 27188 7644
rect 27468 8260 27524 8270
rect 26908 7420 27412 7476
rect 27244 6802 27300 6814
rect 27244 6750 27246 6802
rect 27298 6750 27300 6802
rect 26684 6638 26686 6690
rect 26738 6638 26740 6690
rect 26684 6626 26740 6638
rect 27132 6692 27188 6702
rect 27132 6598 27188 6636
rect 27244 6132 27300 6750
rect 27244 6066 27300 6076
rect 26684 6020 26740 6030
rect 26684 5906 26740 5964
rect 26684 5854 26686 5906
rect 26738 5854 26740 5906
rect 26684 5842 26740 5854
rect 26012 5282 26068 5292
rect 26236 5740 26628 5796
rect 25900 5124 25956 5134
rect 25900 5030 25956 5068
rect 26124 5010 26180 5022
rect 26124 4958 26126 5010
rect 26178 4958 26180 5010
rect 26124 4676 26180 4958
rect 26236 5010 26292 5740
rect 26796 5348 26852 5358
rect 26796 5122 26852 5292
rect 27244 5348 27300 5358
rect 27244 5254 27300 5292
rect 27356 5346 27412 7420
rect 27468 6020 27524 8204
rect 27468 5954 27524 5964
rect 27356 5294 27358 5346
rect 27410 5294 27412 5346
rect 27356 5282 27412 5294
rect 27580 5236 27636 9324
rect 27692 6692 27748 11788
rect 27804 10388 27860 12012
rect 28140 11508 28196 13356
rect 28252 11732 28308 13468
rect 28252 11666 28308 11676
rect 28252 11508 28308 11518
rect 28140 11506 28308 11508
rect 28140 11454 28254 11506
rect 28306 11454 28308 11506
rect 28140 11452 28308 11454
rect 28252 11442 28308 11452
rect 28028 11396 28084 11406
rect 28028 10724 28084 11340
rect 28028 10658 28084 10668
rect 27804 10332 28196 10388
rect 27916 9940 27972 9950
rect 27916 9044 27972 9884
rect 27916 8978 27972 8988
rect 27916 8260 27972 8270
rect 27916 8166 27972 8204
rect 27804 7812 27860 7822
rect 27804 7588 27860 7756
rect 27804 7474 27860 7532
rect 27804 7422 27806 7474
rect 27858 7422 27860 7474
rect 27804 7410 27860 7422
rect 27692 6626 27748 6636
rect 27804 6690 27860 6702
rect 27804 6638 27806 6690
rect 27858 6638 27860 6690
rect 27692 5906 27748 5918
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5460 27748 5854
rect 27804 5908 27860 6638
rect 27804 5842 27860 5852
rect 27692 5394 27748 5404
rect 28028 5684 28084 5694
rect 28028 5236 28084 5628
rect 26796 5070 26798 5122
rect 26850 5070 26852 5122
rect 26796 5058 26852 5070
rect 26908 5180 27188 5236
rect 27580 5180 27860 5236
rect 26236 4958 26238 5010
rect 26290 4958 26292 5010
rect 26236 4946 26292 4958
rect 26572 4900 26628 4910
rect 26348 4898 26628 4900
rect 26348 4846 26574 4898
rect 26626 4846 26628 4898
rect 26348 4844 26628 4846
rect 26348 4676 26404 4844
rect 26572 4834 26628 4844
rect 26124 4620 26404 4676
rect 25788 4508 26852 4564
rect 26796 4338 26852 4508
rect 26908 4450 26964 5180
rect 27132 5124 27188 5180
rect 27468 5124 27524 5134
rect 27132 5122 27524 5124
rect 27132 5070 27470 5122
rect 27522 5070 27524 5122
rect 27132 5068 27524 5070
rect 27468 5058 27524 5068
rect 27020 5012 27076 5022
rect 27020 5010 27300 5012
rect 27020 4958 27022 5010
rect 27074 4958 27300 5010
rect 27020 4956 27300 4958
rect 27020 4946 27076 4956
rect 26908 4398 26910 4450
rect 26962 4398 26964 4450
rect 26908 4386 26964 4398
rect 27020 4788 27076 4798
rect 26796 4286 26798 4338
rect 26850 4286 26852 4338
rect 26796 4274 26852 4286
rect 27020 4338 27076 4732
rect 27020 4286 27022 4338
rect 27074 4286 27076 4338
rect 27020 4274 27076 4286
rect 27244 4226 27300 4956
rect 27244 4174 27246 4226
rect 27298 4174 27300 4226
rect 27244 4162 27300 4174
rect 27468 4338 27524 4350
rect 27468 4286 27470 4338
rect 27522 4286 27524 4338
rect 26124 4116 26180 4126
rect 26124 4114 26292 4116
rect 26124 4062 26126 4114
rect 26178 4062 26292 4114
rect 26124 4060 26292 4062
rect 26124 4050 26180 4060
rect 25564 3726 25566 3778
rect 25618 3726 25620 3778
rect 25564 3714 25620 3726
rect 26012 3780 26068 3790
rect 25228 3666 25284 3678
rect 25228 3614 25230 3666
rect 25282 3614 25284 3666
rect 25228 3388 25284 3614
rect 25116 3332 25284 3388
rect 25116 1988 25172 3332
rect 25452 3220 25508 3230
rect 25228 2212 25284 2222
rect 25228 2118 25284 2156
rect 25116 1922 25172 1932
rect 25004 1362 25060 1372
rect 24668 1204 24724 1214
rect 24444 1092 24500 1102
rect 24444 998 24500 1036
rect 24668 980 24724 1148
rect 24892 1204 24948 1214
rect 24892 1110 24948 1148
rect 25452 1202 25508 3164
rect 25676 3220 25732 3230
rect 25676 2884 25732 3164
rect 25676 2770 25732 2828
rect 25676 2718 25678 2770
rect 25730 2718 25732 2770
rect 25676 2706 25732 2718
rect 25564 2100 25620 2110
rect 25564 2098 25956 2100
rect 25564 2046 25566 2098
rect 25618 2046 25956 2098
rect 25564 2044 25956 2046
rect 25564 2034 25620 2044
rect 25452 1150 25454 1202
rect 25506 1150 25508 1202
rect 25452 1138 25508 1150
rect 25676 1764 25732 1774
rect 24668 924 24948 980
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24892 756 24948 924
rect 24332 690 24388 700
rect 24892 690 24948 700
rect 25116 978 25172 990
rect 25116 926 25118 978
rect 25170 926 25172 978
rect 24892 532 24948 542
rect 24444 308 24500 318
rect 23996 252 24276 308
rect 23996 112 24052 252
rect 13468 18 13524 28
rect 13664 0 13776 112
rect 14112 0 14224 112
rect 14560 0 14672 112
rect 15008 0 15120 112
rect 15456 0 15568 112
rect 15904 0 16016 112
rect 16352 0 16464 112
rect 16800 0 16912 112
rect 17248 0 17360 112
rect 17696 0 17808 112
rect 18144 0 18256 112
rect 18592 0 18704 112
rect 19040 0 19152 112
rect 19488 0 19600 112
rect 19936 0 20048 112
rect 20384 0 20496 112
rect 20832 0 20944 112
rect 21280 0 21392 112
rect 21728 0 21840 112
rect 22176 0 22288 112
rect 22624 0 22736 112
rect 23072 0 23184 112
rect 23520 0 23632 112
rect 23968 0 24080 112
rect 24220 94 24276 252
rect 24444 112 24500 252
rect 24892 112 24948 476
rect 25116 532 25172 926
rect 25116 466 25172 476
rect 25340 644 25396 654
rect 25340 112 25396 588
rect 25676 532 25732 1708
rect 25900 1540 25956 2044
rect 26012 1986 26068 3724
rect 26124 3556 26180 3566
rect 26124 3462 26180 3500
rect 26012 1934 26014 1986
rect 26066 1934 26068 1986
rect 26012 1922 26068 1934
rect 25900 1484 26180 1540
rect 25788 1428 25844 1438
rect 25788 1090 25844 1372
rect 26124 1202 26180 1484
rect 26124 1150 26126 1202
rect 26178 1150 26180 1202
rect 26124 1138 26180 1150
rect 26236 1204 26292 4060
rect 26460 4114 26516 4126
rect 26460 4062 26462 4114
rect 26514 4062 26516 4114
rect 26460 3444 26516 4062
rect 26572 3780 26628 3790
rect 26572 3686 26628 3724
rect 26460 3378 26516 3388
rect 27468 3332 27524 4286
rect 27692 3780 27748 3790
rect 27692 3686 27748 3724
rect 27804 3388 27860 5180
rect 28028 5142 28084 5180
rect 27916 5124 27972 5134
rect 27916 5030 27972 5068
rect 28140 5012 28196 10332
rect 28364 6692 28420 15092
rect 28588 14420 28644 16828
rect 28700 16324 28756 16942
rect 28700 16258 28756 16268
rect 28812 15540 28868 21196
rect 29036 21140 29092 21150
rect 28924 19236 28980 19246
rect 28924 19142 28980 19180
rect 29036 18338 29092 21084
rect 29148 20692 29204 21532
rect 29260 21522 29316 21532
rect 29372 21364 29428 23492
rect 29484 23156 29540 23166
rect 29484 23044 29540 23100
rect 29484 23042 29652 23044
rect 29484 22990 29486 23042
rect 29538 22990 29652 23042
rect 29484 22988 29652 22990
rect 29484 22978 29540 22988
rect 29148 20626 29204 20636
rect 29260 21308 29428 21364
rect 29484 21362 29540 21374
rect 29484 21310 29486 21362
rect 29538 21310 29540 21362
rect 29148 19908 29204 19918
rect 29148 19814 29204 19852
rect 29036 18286 29038 18338
rect 29090 18286 29092 18338
rect 29036 18274 29092 18286
rect 29036 17778 29092 17790
rect 29036 17726 29038 17778
rect 29090 17726 29092 17778
rect 28924 17666 28980 17678
rect 28924 17614 28926 17666
rect 28978 17614 28980 17666
rect 28924 16548 28980 17614
rect 29036 17220 29092 17726
rect 29036 17154 29092 17164
rect 29148 16660 29204 16670
rect 29148 16566 29204 16604
rect 28924 16482 28980 16492
rect 28588 14326 28644 14364
rect 28700 15484 28868 15540
rect 28700 14196 28756 15484
rect 28924 14532 28980 14542
rect 28364 6626 28420 6636
rect 28476 14140 28756 14196
rect 28812 14530 28980 14532
rect 28812 14478 28926 14530
rect 28978 14478 28980 14530
rect 28812 14476 28980 14478
rect 29260 14532 29316 21308
rect 29484 20804 29540 21310
rect 29484 20738 29540 20748
rect 29596 19908 29652 22988
rect 29708 22820 29764 23492
rect 29708 22754 29764 22764
rect 29820 22596 29876 26460
rect 30156 26292 30212 27806
rect 30380 27634 30436 27646
rect 30380 27582 30382 27634
rect 30434 27582 30436 27634
rect 30044 26236 30212 26292
rect 30268 27524 30324 27534
rect 30044 26180 30100 26236
rect 30044 25060 30100 26124
rect 30156 26068 30212 26078
rect 30156 25172 30212 26012
rect 30156 25106 30212 25116
rect 30044 24994 30100 25004
rect 29932 24612 29988 24622
rect 29932 24518 29988 24556
rect 30268 24162 30324 27468
rect 30380 27300 30436 27582
rect 30380 27234 30436 27244
rect 30380 26290 30436 26302
rect 30380 26238 30382 26290
rect 30434 26238 30436 26290
rect 30380 25730 30436 26238
rect 30380 25678 30382 25730
rect 30434 25678 30436 25730
rect 30380 25666 30436 25678
rect 30492 24612 30548 30044
rect 30268 24110 30270 24162
rect 30322 24110 30324 24162
rect 30268 23940 30324 24110
rect 29596 19842 29652 19852
rect 29708 22540 29876 22596
rect 30156 23604 30212 23614
rect 29708 19796 29764 22540
rect 29820 22370 29876 22382
rect 29820 22318 29822 22370
rect 29874 22318 29876 22370
rect 29820 21588 29876 22318
rect 30156 22036 30212 23548
rect 30268 23268 30324 23884
rect 30268 23202 30324 23212
rect 30380 24556 30548 24612
rect 30604 28532 30660 28542
rect 30156 21970 30212 21980
rect 30268 22372 30324 22382
rect 29932 21588 29988 21598
rect 29820 21586 29988 21588
rect 29820 21534 29934 21586
rect 29986 21534 29988 21586
rect 29820 21532 29988 21534
rect 29932 21026 29988 21532
rect 30268 21476 30324 22316
rect 30380 22370 30436 24556
rect 30604 23380 30660 28476
rect 30716 26908 30772 37996
rect 30828 34018 30884 39900
rect 30940 39394 30996 39406
rect 30940 39342 30942 39394
rect 30994 39342 30996 39394
rect 30940 38276 30996 39342
rect 31276 39396 31332 39406
rect 31276 39302 31332 39340
rect 31388 38948 31444 38958
rect 31388 38854 31444 38892
rect 31164 38724 31220 38734
rect 30940 38210 30996 38220
rect 31052 38388 31108 38398
rect 30940 38052 30996 38062
rect 30940 36820 30996 37996
rect 31052 37268 31108 38332
rect 31052 37202 31108 37212
rect 30940 34132 30996 36764
rect 31052 35700 31108 35710
rect 31052 35606 31108 35644
rect 31164 35588 31220 38668
rect 31276 38612 31332 38622
rect 31276 38050 31332 38556
rect 31276 37998 31278 38050
rect 31330 37998 31332 38050
rect 31276 37986 31332 37998
rect 31388 38164 31444 38174
rect 31388 37261 31444 38108
rect 31388 37209 31390 37261
rect 31442 37209 31444 37261
rect 31388 37197 31444 37209
rect 31388 36258 31444 36270
rect 31388 36206 31390 36258
rect 31442 36206 31444 36258
rect 31388 36036 31444 36206
rect 31388 35970 31444 35980
rect 31164 35522 31220 35532
rect 31276 35476 31332 35486
rect 31164 34804 31220 34814
rect 30940 34066 30996 34076
rect 31052 34468 31108 34478
rect 30828 33966 30830 34018
rect 30882 33966 30884 34018
rect 30828 33954 30884 33966
rect 31052 33236 31108 34412
rect 31052 33170 31108 33180
rect 31164 32788 31220 34748
rect 31276 34130 31332 35420
rect 31276 34078 31278 34130
rect 31330 34078 31332 34130
rect 31276 34066 31332 34078
rect 31500 33572 31556 41918
rect 31612 41860 31668 41870
rect 31612 41766 31668 41804
rect 31836 41748 31892 42700
rect 31724 41692 31892 41748
rect 31948 42532 32004 42542
rect 31724 41636 31780 41692
rect 31500 33506 31556 33516
rect 31612 41580 31780 41636
rect 31052 32732 31220 32788
rect 30940 32116 30996 32126
rect 30828 29428 30884 29438
rect 30828 29334 30884 29372
rect 30828 27860 30884 27870
rect 30828 27766 30884 27804
rect 30940 27188 30996 32060
rect 31052 29764 31108 32732
rect 31612 32564 31668 41580
rect 31724 40402 31780 40414
rect 31724 40350 31726 40402
rect 31778 40350 31780 40402
rect 31724 37604 31780 40350
rect 31948 40290 32004 42476
rect 31948 40238 31950 40290
rect 32002 40238 32004 40290
rect 31948 40226 32004 40238
rect 32060 38668 32116 43374
rect 31836 38612 31892 38622
rect 31836 38518 31892 38556
rect 31948 38612 32116 38668
rect 31724 37548 31892 37604
rect 31836 35588 31892 37548
rect 31836 35522 31892 35532
rect 31836 35364 31892 35374
rect 31836 34468 31892 35308
rect 31836 34402 31892 34412
rect 31388 32508 31668 32564
rect 31836 33908 31892 33918
rect 31052 29698 31108 29708
rect 31164 30996 31220 31006
rect 31052 29204 31108 29214
rect 31052 28642 31108 29148
rect 31052 28590 31054 28642
rect 31106 28590 31108 28642
rect 31052 28578 31108 28590
rect 30940 27122 30996 27132
rect 31052 28084 31108 28094
rect 30716 26852 30884 26908
rect 30716 25060 30772 25070
rect 30716 24722 30772 25004
rect 30716 24670 30718 24722
rect 30770 24670 30772 24722
rect 30716 24658 30772 24670
rect 30380 22318 30382 22370
rect 30434 22318 30436 22370
rect 30380 22306 30436 22318
rect 30492 23324 30660 23380
rect 30268 21410 30324 21420
rect 30492 21028 30548 23324
rect 30604 23156 30660 23166
rect 30604 23062 30660 23100
rect 29932 20974 29934 21026
rect 29986 20974 29988 21026
rect 29932 20962 29988 20974
rect 30380 20972 30548 21028
rect 30604 22484 30660 22494
rect 29484 19348 29540 19358
rect 29372 18452 29428 18462
rect 29372 14980 29428 18396
rect 29484 17780 29540 19292
rect 29484 17714 29540 17724
rect 29596 19236 29652 19246
rect 29372 14756 29428 14924
rect 29372 14690 29428 14700
rect 29484 16548 29540 16558
rect 29260 14476 29428 14532
rect 28476 6690 28532 14140
rect 28812 13186 28868 14476
rect 28924 14466 28980 14476
rect 29036 14420 29092 14430
rect 28924 14196 28980 14206
rect 28924 13858 28980 14140
rect 28924 13806 28926 13858
rect 28978 13806 28980 13858
rect 28924 13794 28980 13806
rect 29036 13636 29092 14364
rect 28812 13134 28814 13186
rect 28866 13134 28868 13186
rect 28812 13122 28868 13134
rect 28924 13580 29092 13636
rect 29148 14308 29204 14318
rect 28588 11954 28644 11966
rect 28588 11902 28590 11954
rect 28642 11902 28644 11954
rect 28588 11508 28644 11902
rect 28700 11508 28756 11518
rect 28588 11506 28756 11508
rect 28588 11454 28702 11506
rect 28754 11454 28756 11506
rect 28588 11452 28756 11454
rect 28700 11442 28756 11452
rect 28812 11396 28868 11406
rect 28700 11172 28756 11182
rect 28700 9268 28756 11116
rect 28812 9716 28868 11340
rect 28924 9828 28980 13580
rect 29036 10388 29092 10398
rect 29036 10050 29092 10332
rect 29036 9998 29038 10050
rect 29090 9998 29092 10050
rect 29036 9986 29092 9998
rect 28924 9772 29092 9828
rect 28812 9660 28980 9716
rect 28812 9268 28868 9278
rect 28700 9212 28812 9268
rect 28588 8484 28644 8494
rect 28588 8036 28644 8428
rect 28812 8258 28868 9212
rect 28812 8206 28814 8258
rect 28866 8206 28868 8258
rect 28812 8194 28868 8206
rect 28588 7970 28644 7980
rect 28476 6638 28478 6690
rect 28530 6638 28532 6690
rect 28476 6626 28532 6638
rect 28476 6132 28532 6142
rect 28476 6038 28532 6076
rect 28588 5682 28644 5694
rect 28588 5630 28590 5682
rect 28642 5630 28644 5682
rect 28588 5348 28644 5630
rect 28700 5684 28756 5694
rect 28700 5590 28756 5628
rect 28588 5282 28644 5292
rect 28028 4956 28196 5012
rect 27804 3332 27972 3388
rect 27468 3276 27748 3332
rect 26460 2884 26516 2894
rect 26460 2770 26516 2828
rect 26460 2718 26462 2770
rect 26514 2718 26516 2770
rect 26460 2706 26516 2718
rect 27580 2548 27636 2558
rect 26908 2546 27636 2548
rect 26908 2494 27582 2546
rect 27634 2494 27636 2546
rect 26908 2492 27636 2494
rect 26572 2212 26628 2222
rect 26572 2118 26628 2156
rect 26236 1138 26292 1148
rect 26908 1202 26964 2492
rect 27580 2482 27636 2492
rect 27692 2210 27748 3276
rect 27804 2772 27860 2782
rect 27804 2678 27860 2716
rect 27916 2548 27972 3332
rect 28028 3220 28084 4956
rect 28476 4116 28532 4126
rect 28252 4114 28532 4116
rect 28252 4062 28478 4114
rect 28530 4062 28532 4114
rect 28252 4060 28532 4062
rect 28140 3668 28196 3678
rect 28140 3574 28196 3612
rect 28028 3154 28084 3164
rect 27916 2482 27972 2492
rect 27692 2158 27694 2210
rect 27746 2158 27748 2210
rect 27692 2146 27748 2158
rect 26908 1150 26910 1202
rect 26962 1150 26964 1202
rect 26908 1138 26964 1150
rect 28028 1316 28084 1326
rect 28028 1202 28084 1260
rect 28028 1150 28030 1202
rect 28082 1150 28084 1202
rect 28028 1138 28084 1150
rect 25788 1038 25790 1090
rect 25842 1038 25844 1090
rect 25788 1026 25844 1038
rect 27020 1092 27076 1102
rect 26460 978 26516 990
rect 26460 926 26462 978
rect 26514 926 26516 978
rect 25676 476 25844 532
rect 25788 112 25844 476
rect 26236 420 26292 430
rect 26236 112 26292 364
rect 26460 308 26516 926
rect 26460 242 26516 252
rect 26684 980 26740 990
rect 26684 112 26740 924
rect 27020 532 27076 1036
rect 27132 980 27188 990
rect 27132 886 27188 924
rect 28252 756 28308 4060
rect 28476 4050 28532 4060
rect 28812 4114 28868 4126
rect 28812 4062 28814 4114
rect 28866 4062 28868 4114
rect 28476 3780 28532 3790
rect 28476 3554 28532 3724
rect 28812 3668 28868 4062
rect 28924 3780 28980 9660
rect 29036 4788 29092 9772
rect 29036 4722 29092 4732
rect 29148 4676 29204 14252
rect 29260 13636 29316 13646
rect 29260 10948 29316 13580
rect 29372 11172 29428 14476
rect 29484 14530 29540 16492
rect 29596 16324 29652 19180
rect 29708 18564 29764 19740
rect 29708 18498 29764 18508
rect 29820 20132 29876 20142
rect 29708 17666 29764 17678
rect 29708 17614 29710 17666
rect 29762 17614 29764 17666
rect 29708 17108 29764 17614
rect 29708 17042 29764 17052
rect 29596 16258 29652 16268
rect 29596 14756 29652 14766
rect 29596 14662 29652 14700
rect 29484 14478 29486 14530
rect 29538 14478 29540 14530
rect 29484 14308 29540 14478
rect 29484 14242 29540 14252
rect 29820 12066 29876 20076
rect 30380 20132 30436 20972
rect 30604 20914 30660 22428
rect 30716 21588 30772 21598
rect 30828 21588 30884 26852
rect 30940 26290 30996 26302
rect 30940 26238 30942 26290
rect 30994 26238 30996 26290
rect 30940 26068 30996 26238
rect 30940 26002 30996 26012
rect 31052 23604 31108 28028
rect 31052 23538 31108 23548
rect 31164 23154 31220 30940
rect 31276 30098 31332 30110
rect 31276 30046 31278 30098
rect 31330 30046 31332 30098
rect 31276 29540 31332 30046
rect 31276 29474 31332 29484
rect 31388 27746 31444 32508
rect 31612 32338 31668 32350
rect 31612 32286 31614 32338
rect 31666 32286 31668 32338
rect 31612 32004 31668 32286
rect 31612 31938 31668 31948
rect 31500 30772 31556 30782
rect 31500 30678 31556 30716
rect 31500 30212 31556 30222
rect 31836 30212 31892 33852
rect 31948 33124 32004 38612
rect 32172 35698 32228 51100
rect 32284 50148 32340 55804
rect 32396 55858 32452 55870
rect 32396 55806 32398 55858
rect 32450 55806 32452 55858
rect 32396 55412 32452 55806
rect 32956 55524 33012 57344
rect 33180 56308 33236 56318
rect 33180 56082 33236 56252
rect 33180 56030 33182 56082
rect 33234 56030 33236 56082
rect 33180 56018 33236 56030
rect 33404 56084 33460 57344
rect 33404 56018 33460 56028
rect 32396 55346 32452 55356
rect 32620 55468 33012 55524
rect 33404 55858 33460 55870
rect 33404 55806 33406 55858
rect 33458 55806 33460 55858
rect 32508 55300 32564 55310
rect 32508 55206 32564 55244
rect 32396 55074 32452 55086
rect 32396 55022 32398 55074
rect 32450 55022 32452 55074
rect 32396 54740 32452 55022
rect 32396 54684 32564 54740
rect 32396 54514 32452 54526
rect 32396 54462 32398 54514
rect 32450 54462 32452 54514
rect 32396 54068 32452 54462
rect 32396 54002 32452 54012
rect 32508 53956 32564 54684
rect 32508 53862 32564 53900
rect 32396 53842 32452 53854
rect 32396 53790 32398 53842
rect 32450 53790 32452 53842
rect 32396 53732 32452 53790
rect 32396 53666 32452 53676
rect 32620 52948 32676 55468
rect 33180 55410 33236 55422
rect 33180 55358 33182 55410
rect 33234 55358 33236 55410
rect 32956 55298 33012 55310
rect 32956 55246 32958 55298
rect 33010 55246 33012 55298
rect 32844 54292 32900 54302
rect 32844 54198 32900 54236
rect 32844 54068 32900 54078
rect 32732 53732 32788 53742
rect 32732 53638 32788 53676
rect 32844 53508 32900 54012
rect 32844 53284 32900 53452
rect 32732 53228 32900 53284
rect 32732 53058 32788 53228
rect 32732 53006 32734 53058
rect 32786 53006 32788 53058
rect 32732 52994 32788 53006
rect 32508 52164 32564 52174
rect 32508 52070 32564 52108
rect 32620 51156 32676 52892
rect 32620 51090 32676 51100
rect 32956 50428 33012 55246
rect 33180 54628 33236 55358
rect 33404 55188 33460 55806
rect 33740 55860 33796 55870
rect 33740 55766 33796 55804
rect 33404 55122 33460 55132
rect 33516 55748 33572 55758
rect 33516 54964 33572 55692
rect 33852 55748 33908 57344
rect 33852 55682 33908 55692
rect 34076 55858 34132 55870
rect 34076 55806 34078 55858
rect 34130 55806 34132 55858
rect 33852 55412 33908 55422
rect 33852 55318 33908 55356
rect 33628 55300 33684 55310
rect 33628 55206 33684 55244
rect 34076 55188 34132 55806
rect 34300 55524 34356 57344
rect 34524 57204 34580 57214
rect 34524 56082 34580 57148
rect 34524 56030 34526 56082
rect 34578 56030 34580 56082
rect 34524 56018 34580 56030
rect 34748 56084 34804 57344
rect 34748 56018 34804 56028
rect 34748 55860 34804 55870
rect 34300 55458 34356 55468
rect 34412 55858 34804 55860
rect 34412 55806 34750 55858
rect 34802 55806 34804 55858
rect 34412 55804 34804 55806
rect 34412 55300 34468 55804
rect 34748 55794 34804 55804
rect 33516 54898 33572 54908
rect 33852 55132 34132 55188
rect 34300 55244 34468 55300
rect 34524 55412 34580 55422
rect 34524 55298 34580 55356
rect 34524 55246 34526 55298
rect 34578 55246 34580 55298
rect 33180 54562 33236 54572
rect 33068 53506 33124 53518
rect 33068 53454 33070 53506
rect 33122 53454 33124 53506
rect 33068 53172 33124 53454
rect 33068 53106 33124 53116
rect 33628 53060 33684 53070
rect 33068 52948 33124 52958
rect 33068 52724 33124 52892
rect 33068 52658 33124 52668
rect 33180 52722 33236 52734
rect 33180 52670 33182 52722
rect 33234 52670 33236 52722
rect 32508 50372 32564 50382
rect 32508 50278 32564 50316
rect 32732 50372 32788 50382
rect 32284 50082 32340 50092
rect 32396 50036 32452 50046
rect 32284 49924 32340 49934
rect 32284 49830 32340 49868
rect 32396 48580 32452 49980
rect 32732 49924 32788 50316
rect 32732 49858 32788 49868
rect 32844 50372 33012 50428
rect 33068 52500 33124 52510
rect 33068 51490 33124 52444
rect 33180 52164 33236 52670
rect 33180 52098 33236 52108
rect 33628 52052 33684 53004
rect 33852 52612 33908 55132
rect 34188 55076 34244 55086
rect 33964 55074 34244 55076
rect 33964 55022 34190 55074
rect 34242 55022 34244 55074
rect 33964 55020 34244 55022
rect 33964 54738 34020 55020
rect 34188 55010 34244 55020
rect 33964 54686 33966 54738
rect 34018 54686 34020 54738
rect 33964 54674 34020 54686
rect 34188 53956 34244 53966
rect 34188 53862 34244 53900
rect 34300 53732 34356 55244
rect 34524 55234 34580 55246
rect 34636 55298 34692 55310
rect 34636 55246 34638 55298
rect 34690 55246 34692 55298
rect 34636 53844 34692 55246
rect 34748 55298 34804 55310
rect 34748 55246 34750 55298
rect 34802 55246 34804 55298
rect 34748 54514 34804 55246
rect 34748 54462 34750 54514
rect 34802 54462 34804 54514
rect 34748 54450 34804 54462
rect 34860 55298 34916 55310
rect 34860 55246 34862 55298
rect 34914 55246 34916 55298
rect 33964 53676 34356 53732
rect 34524 53788 34692 53844
rect 33964 53172 34020 53676
rect 33964 53106 34020 53116
rect 34076 53508 34132 53518
rect 33852 52546 33908 52556
rect 33740 52276 33796 52286
rect 33740 52182 33796 52220
rect 33068 51438 33070 51490
rect 33122 51438 33124 51490
rect 33068 50372 33124 51438
rect 32508 48804 32564 48814
rect 32508 48710 32564 48748
rect 32396 48524 32564 48580
rect 32396 48018 32452 48030
rect 32396 47966 32398 48018
rect 32450 47966 32452 48018
rect 32396 47684 32452 47966
rect 32396 47618 32452 47628
rect 32284 47124 32340 47134
rect 32284 43316 32340 47068
rect 32396 45892 32452 45902
rect 32508 45892 32564 48524
rect 32732 47348 32788 47358
rect 32620 46562 32676 46574
rect 32620 46510 32622 46562
rect 32674 46510 32676 46562
rect 32620 46116 32676 46510
rect 32732 46452 32788 47292
rect 32844 47124 32900 50372
rect 33068 50306 33124 50316
rect 33180 51828 33236 51838
rect 32956 49812 33012 49822
rect 32956 49718 33012 49756
rect 32844 47058 32900 47068
rect 33068 47570 33124 47582
rect 33068 47518 33070 47570
rect 33122 47518 33124 47570
rect 33068 47124 33124 47518
rect 33068 47058 33124 47068
rect 33180 47460 33236 51772
rect 33628 51716 33684 51996
rect 34076 52162 34132 53452
rect 34524 53284 34580 53788
rect 34860 53732 34916 55246
rect 35196 55300 35252 57344
rect 35532 56420 35588 56430
rect 35532 56082 35588 56364
rect 35532 56030 35534 56082
rect 35586 56030 35588 56082
rect 35532 56018 35588 56030
rect 35196 55234 35252 55244
rect 35308 55636 35364 55646
rect 35644 55636 35700 57344
rect 36092 56308 36148 57344
rect 36540 56420 36596 57344
rect 36540 56354 36596 56364
rect 35980 56252 36148 56308
rect 34860 53666 34916 53676
rect 34972 54514 35028 54526
rect 34972 54462 34974 54514
rect 35026 54462 35028 54514
rect 34636 53618 34692 53630
rect 34636 53566 34638 53618
rect 34690 53566 34692 53618
rect 34636 53508 34692 53566
rect 34972 53620 35028 54462
rect 35084 54404 35140 54414
rect 35084 54290 35140 54348
rect 35084 54238 35086 54290
rect 35138 54238 35140 54290
rect 35084 54226 35140 54238
rect 35196 54402 35252 54414
rect 35196 54350 35198 54402
rect 35250 54350 35252 54402
rect 35196 53844 35252 54350
rect 35308 53956 35364 55580
rect 35420 55580 35700 55636
rect 35756 55858 35812 55870
rect 35756 55806 35758 55858
rect 35810 55806 35812 55858
rect 35420 55298 35476 55580
rect 35756 55524 35812 55806
rect 35756 55458 35812 55468
rect 35420 55246 35422 55298
rect 35474 55246 35476 55298
rect 35420 55234 35476 55246
rect 35644 55410 35700 55422
rect 35644 55358 35646 55410
rect 35698 55358 35700 55410
rect 35420 54404 35476 54414
rect 35420 54402 35588 54404
rect 35420 54350 35422 54402
rect 35474 54350 35588 54402
rect 35420 54348 35588 54350
rect 35420 54338 35476 54348
rect 35308 53890 35364 53900
rect 35196 53778 35252 53788
rect 34972 53554 35028 53564
rect 35420 53620 35476 53630
rect 35420 53526 35476 53564
rect 34636 53442 34692 53452
rect 34300 53228 34580 53284
rect 34300 53170 34356 53228
rect 34300 53118 34302 53170
rect 34354 53118 34356 53170
rect 34300 53106 34356 53118
rect 34860 53116 35252 53172
rect 34748 52948 34804 52958
rect 34076 52110 34078 52162
rect 34130 52110 34132 52162
rect 34076 52052 34132 52110
rect 34076 51986 34132 51996
rect 34524 52946 34804 52948
rect 34524 52894 34750 52946
rect 34802 52894 34804 52946
rect 34524 52892 34804 52894
rect 33628 51660 33796 51716
rect 33516 51156 33572 51166
rect 33516 51062 33572 51100
rect 33740 50706 33796 51660
rect 34524 51604 34580 52892
rect 34748 52882 34804 52892
rect 34636 52388 34692 52398
rect 34636 52274 34692 52332
rect 34636 52222 34638 52274
rect 34690 52222 34692 52274
rect 34636 52210 34692 52222
rect 34748 52276 34804 52286
rect 34748 52182 34804 52220
rect 34748 51938 34804 51950
rect 34748 51886 34750 51938
rect 34802 51886 34804 51938
rect 34636 51604 34692 51614
rect 34524 51602 34692 51604
rect 34524 51550 34638 51602
rect 34690 51550 34692 51602
rect 34524 51548 34692 51550
rect 34636 51538 34692 51548
rect 34748 51156 34804 51886
rect 33740 50654 33742 50706
rect 33794 50654 33796 50706
rect 33740 50642 33796 50654
rect 34412 51100 34804 51156
rect 34076 50596 34132 50606
rect 33964 50594 34132 50596
rect 33964 50542 34078 50594
rect 34130 50542 34132 50594
rect 33964 50540 34132 50542
rect 33964 50372 34020 50540
rect 34076 50530 34132 50540
rect 33628 49138 33684 49150
rect 33628 49086 33630 49138
rect 33682 49086 33684 49138
rect 33516 49028 33572 49038
rect 32956 46788 33012 46798
rect 32956 46694 33012 46732
rect 32732 46386 32788 46396
rect 32844 46450 32900 46462
rect 32844 46398 32846 46450
rect 32898 46398 32900 46450
rect 32620 46050 32676 46060
rect 32508 45836 32676 45892
rect 32396 44100 32452 45836
rect 32508 45668 32564 45678
rect 32508 45574 32564 45612
rect 32508 44882 32564 44894
rect 32508 44830 32510 44882
rect 32562 44830 32564 44882
rect 32508 44324 32564 44830
rect 32508 44258 32564 44268
rect 32508 44100 32564 44110
rect 32396 44098 32564 44100
rect 32396 44046 32510 44098
rect 32562 44046 32564 44098
rect 32396 44044 32564 44046
rect 32508 44034 32564 44044
rect 32284 43250 32340 43260
rect 32508 43540 32564 43550
rect 32620 43540 32676 45836
rect 32844 44660 32900 46398
rect 33180 46116 33236 47404
rect 33292 48804 33348 48814
rect 33292 46676 33348 48748
rect 33516 48692 33572 48972
rect 33516 48626 33572 48636
rect 33516 48020 33572 48030
rect 33516 47926 33572 47964
rect 33628 47684 33684 49086
rect 33964 48804 34020 50316
rect 34412 49812 34468 51100
rect 34860 50428 34916 53116
rect 35084 52946 35140 52958
rect 35084 52894 35086 52946
rect 35138 52894 35140 52946
rect 34748 50372 34916 50428
rect 34972 51828 35028 51838
rect 34412 49746 34468 49756
rect 34524 49810 34580 49822
rect 34524 49758 34526 49810
rect 34578 49758 34580 49810
rect 34076 49586 34132 49598
rect 34076 49534 34078 49586
rect 34130 49534 34132 49586
rect 34076 49364 34132 49534
rect 34076 49298 34132 49308
rect 34524 49252 34580 49758
rect 33964 48354 34020 48748
rect 34188 49026 34244 49038
rect 34188 48974 34190 49026
rect 34242 48974 34244 49026
rect 34188 48804 34244 48974
rect 34188 48738 34244 48748
rect 34524 48804 34580 49196
rect 34524 48738 34580 48748
rect 34636 49700 34692 49710
rect 33964 48302 33966 48354
rect 34018 48302 34020 48354
rect 33964 48290 34020 48302
rect 34076 48692 34132 48702
rect 33516 47628 33684 47684
rect 34076 47638 34132 48636
rect 33404 47570 33460 47582
rect 33404 47518 33406 47570
rect 33458 47518 33460 47570
rect 33404 47012 33460 47518
rect 33516 47236 33572 47628
rect 33964 47582 34132 47638
rect 34412 48580 34468 48590
rect 33740 47572 33796 47582
rect 33628 47516 33740 47572
rect 33628 47458 33684 47516
rect 33740 47506 33796 47516
rect 33964 47570 34020 47582
rect 33964 47518 33966 47570
rect 34018 47518 34020 47570
rect 33964 47506 34020 47518
rect 33628 47406 33630 47458
rect 33682 47406 33684 47458
rect 33628 47394 33684 47406
rect 33516 47180 33684 47236
rect 33404 46946 33460 46956
rect 33628 46900 33684 47180
rect 33628 46834 33684 46844
rect 33404 46676 33460 46686
rect 33292 46674 33460 46676
rect 33292 46622 33406 46674
rect 33458 46622 33460 46674
rect 33292 46620 33460 46622
rect 32844 44594 32900 44604
rect 33068 46060 33236 46116
rect 32508 43538 32676 43540
rect 32508 43486 32510 43538
rect 32562 43486 32676 43538
rect 32508 43484 32676 43486
rect 32732 43764 32788 43774
rect 32508 43092 32564 43484
rect 32508 43026 32564 43036
rect 32508 42532 32564 42542
rect 32284 42530 32564 42532
rect 32284 42478 32510 42530
rect 32562 42478 32564 42530
rect 32284 42476 32564 42478
rect 32284 41970 32340 42476
rect 32508 42466 32564 42476
rect 32284 41918 32286 41970
rect 32338 41918 32340 41970
rect 32284 40404 32340 41918
rect 32620 41972 32676 41982
rect 32620 41878 32676 41916
rect 32396 40404 32452 40414
rect 32284 40402 32452 40404
rect 32284 40350 32398 40402
rect 32450 40350 32452 40402
rect 32284 40348 32452 40350
rect 32396 40338 32452 40348
rect 32732 40180 32788 43708
rect 32956 42980 33012 42990
rect 32956 41300 33012 42924
rect 32956 41186 33012 41244
rect 32956 41134 32958 41186
rect 33010 41134 33012 41186
rect 32956 41122 33012 41134
rect 32956 40516 33012 40526
rect 32956 40402 33012 40460
rect 32956 40350 32958 40402
rect 33010 40350 33012 40402
rect 32956 40338 33012 40350
rect 32732 40114 32788 40124
rect 32172 35646 32174 35698
rect 32226 35646 32228 35698
rect 32172 35634 32228 35646
rect 32284 40068 32340 40078
rect 32284 35308 32340 40012
rect 33068 40068 33124 46060
rect 33404 46004 33460 46620
rect 33852 46562 33908 46574
rect 33852 46510 33854 46562
rect 33906 46510 33908 46562
rect 33180 45948 33460 46004
rect 33628 46002 33684 46014
rect 33628 45950 33630 46002
rect 33682 45950 33684 46002
rect 33180 45108 33236 45948
rect 33628 45892 33684 45950
rect 33628 45826 33684 45836
rect 33180 44324 33236 45052
rect 33180 44258 33236 44268
rect 33292 45780 33348 45790
rect 33180 43652 33236 43662
rect 33292 43652 33348 45724
rect 33852 45444 33908 46510
rect 34076 45780 34132 45790
rect 34076 45686 34132 45724
rect 33852 45378 33908 45388
rect 33964 45556 34020 45566
rect 33516 44996 33572 45006
rect 33180 43650 33348 43652
rect 33180 43598 33182 43650
rect 33234 43598 33348 43650
rect 33180 43596 33348 43598
rect 33404 44994 33572 44996
rect 33404 44942 33518 44994
rect 33570 44942 33572 44994
rect 33404 44940 33572 44942
rect 33180 43586 33236 43596
rect 33068 40002 33124 40012
rect 33180 43316 33236 43326
rect 32508 39394 32564 39406
rect 32508 39342 32510 39394
rect 32562 39342 32564 39394
rect 32508 38668 32564 39342
rect 33180 38724 33236 43260
rect 33292 41748 33348 41758
rect 33292 40516 33348 41692
rect 33404 41412 33460 44940
rect 33516 44930 33572 44940
rect 33628 44434 33684 44446
rect 33628 44382 33630 44434
rect 33682 44382 33684 44434
rect 33516 43428 33572 43438
rect 33516 43334 33572 43372
rect 33628 43092 33684 44382
rect 33964 43764 34020 45500
rect 34188 45220 34244 45230
rect 34076 44324 34132 44334
rect 34076 44230 34132 44268
rect 33964 43698 34020 43708
rect 33516 43036 33684 43092
rect 33740 43428 33796 43438
rect 33516 41748 33572 43036
rect 33628 42868 33684 42878
rect 33628 42774 33684 42812
rect 33628 41972 33684 41982
rect 33628 41878 33684 41916
rect 33516 41692 33684 41748
rect 33404 41318 33460 41356
rect 33292 40450 33348 40460
rect 33628 40404 33684 41692
rect 32508 38612 32900 38668
rect 33180 38658 33236 38668
rect 33292 40292 33348 40302
rect 32620 37940 32676 37950
rect 32508 37938 32676 37940
rect 32508 37886 32622 37938
rect 32674 37886 32676 37938
rect 32508 37884 32676 37886
rect 32508 37154 32564 37884
rect 32620 37874 32676 37884
rect 32844 37266 32900 38612
rect 32956 38610 33012 38622
rect 32956 38558 32958 38610
rect 33010 38558 33012 38610
rect 32956 38050 33012 38558
rect 32956 37998 32958 38050
rect 33010 37998 33012 38050
rect 32956 37986 33012 37998
rect 32844 37214 32846 37266
rect 32898 37214 32900 37266
rect 32844 37202 32900 37214
rect 32508 37102 32510 37154
rect 32562 37102 32564 37154
rect 32508 37044 32564 37102
rect 32508 36978 32564 36988
rect 33068 37156 33124 37166
rect 32844 36820 32900 36830
rect 32172 35252 32340 35308
rect 32508 35698 32564 35710
rect 32508 35646 32510 35698
rect 32562 35646 32564 35698
rect 32060 34132 32116 34142
rect 32060 34038 32116 34076
rect 31948 33058 32004 33068
rect 32060 31892 32116 31902
rect 32060 31668 32116 31836
rect 32060 31602 32116 31612
rect 31948 30884 32004 30894
rect 32172 30884 32228 35252
rect 32508 35138 32564 35646
rect 32508 35086 32510 35138
rect 32562 35086 32564 35138
rect 32508 35074 32564 35086
rect 32284 34916 32340 34926
rect 32284 34244 32340 34860
rect 32844 34804 32900 36764
rect 32844 34738 32900 34748
rect 32956 36484 33012 36494
rect 32284 34178 32340 34188
rect 32508 34244 32564 34254
rect 32508 33346 32564 34188
rect 32844 34130 32900 34142
rect 32844 34078 32846 34130
rect 32898 34078 32900 34130
rect 32844 33908 32900 34078
rect 32844 33842 32900 33852
rect 32956 33684 33012 36428
rect 33068 33908 33124 37100
rect 33180 37044 33236 37054
rect 33180 36484 33236 36988
rect 33180 36390 33236 36428
rect 33292 36148 33348 40236
rect 33628 39842 33684 40348
rect 33628 39790 33630 39842
rect 33682 39790 33684 39842
rect 33628 39778 33684 39790
rect 33628 39620 33684 39630
rect 33516 38612 33572 38622
rect 33516 38518 33572 38556
rect 33628 38274 33684 39564
rect 33628 38222 33630 38274
rect 33682 38222 33684 38274
rect 33628 38210 33684 38222
rect 33292 36082 33348 36092
rect 33404 38050 33460 38062
rect 33740 38052 33796 43372
rect 33852 43092 33908 43102
rect 33852 42532 33908 43036
rect 34076 42642 34132 42654
rect 34076 42590 34078 42642
rect 34130 42590 34132 42642
rect 34076 42532 34132 42590
rect 33852 42476 34132 42532
rect 33852 40964 33908 42476
rect 33852 40404 33908 40908
rect 34076 41300 34132 41310
rect 33852 40338 33908 40348
rect 33964 40402 34020 40414
rect 33964 40350 33966 40402
rect 34018 40350 34020 40402
rect 33404 37998 33406 38050
rect 33458 37998 33460 38050
rect 33404 37266 33460 37998
rect 33404 37214 33406 37266
rect 33458 37214 33460 37266
rect 33292 35700 33348 35710
rect 33292 35606 33348 35644
rect 33180 35588 33236 35598
rect 33180 35494 33236 35532
rect 33068 33842 33124 33852
rect 33180 34804 33236 34814
rect 32508 33294 32510 33346
rect 32562 33294 32564 33346
rect 32284 32562 32340 32574
rect 32284 32510 32286 32562
rect 32338 32510 32340 32562
rect 32284 30996 32340 32510
rect 32284 30930 32340 30940
rect 32396 32004 32452 32014
rect 32396 31108 32452 31948
rect 32396 30994 32452 31052
rect 32396 30942 32398 30994
rect 32450 30942 32452 30994
rect 32396 30930 32452 30942
rect 32508 31778 32564 33294
rect 32508 31726 32510 31778
rect 32562 31726 32564 31778
rect 31948 30882 32228 30884
rect 31948 30830 31950 30882
rect 32002 30830 32228 30882
rect 31948 30828 32228 30830
rect 31948 30818 32004 30828
rect 31836 30156 32004 30212
rect 31500 30118 31556 30156
rect 31836 29986 31892 29998
rect 31836 29934 31838 29986
rect 31890 29934 31892 29986
rect 31836 29652 31892 29934
rect 31836 29586 31892 29596
rect 31836 29428 31892 29438
rect 31948 29428 32004 30156
rect 31836 29426 32004 29428
rect 31836 29374 31838 29426
rect 31890 29374 32004 29426
rect 31836 29372 32004 29374
rect 31836 29362 31892 29372
rect 31724 28868 31780 28878
rect 31724 28774 31780 28812
rect 31612 28756 31668 28766
rect 31612 28662 31668 28700
rect 31948 28644 32004 28654
rect 31724 28418 31780 28430
rect 31724 28366 31726 28418
rect 31778 28366 31780 28418
rect 31724 27860 31780 28366
rect 31724 27794 31780 27804
rect 31388 27694 31390 27746
rect 31442 27694 31444 27746
rect 31388 27524 31444 27694
rect 31388 27458 31444 27468
rect 31836 27636 31892 27646
rect 31836 27298 31892 27580
rect 31836 27246 31838 27298
rect 31890 27246 31892 27298
rect 31836 27234 31892 27246
rect 31724 27188 31780 27198
rect 31724 27094 31780 27132
rect 31836 27076 31892 27086
rect 31164 23102 31166 23154
rect 31218 23102 31220 23154
rect 31164 23044 31220 23102
rect 31276 26962 31332 26974
rect 31276 26910 31278 26962
rect 31330 26910 31332 26962
rect 31276 26740 31332 26910
rect 31388 26964 31444 27002
rect 31388 26898 31444 26908
rect 31276 23044 31332 26684
rect 31500 26740 31556 26750
rect 31500 25844 31556 26684
rect 31500 25778 31556 25788
rect 31612 26628 31668 26638
rect 31612 25618 31668 26572
rect 31836 26290 31892 27020
rect 31836 26238 31838 26290
rect 31890 26238 31892 26290
rect 31612 25566 31614 25618
rect 31666 25566 31668 25618
rect 31612 25554 31668 25566
rect 31724 25618 31780 25630
rect 31724 25566 31726 25618
rect 31778 25566 31780 25618
rect 31724 25508 31780 25566
rect 31724 25442 31780 25452
rect 31836 25396 31892 26238
rect 31836 25330 31892 25340
rect 31724 25284 31780 25294
rect 31724 25190 31780 25228
rect 31500 24724 31556 24734
rect 31500 24630 31556 24668
rect 31724 24276 31780 24286
rect 31500 24052 31556 24062
rect 31388 23714 31444 23726
rect 31388 23662 31390 23714
rect 31442 23662 31444 23714
rect 31388 23268 31444 23662
rect 31388 23202 31444 23212
rect 31276 22988 31444 23044
rect 31164 22978 31220 22988
rect 31052 22820 31108 22830
rect 30716 21586 30884 21588
rect 30716 21534 30718 21586
rect 30770 21534 30884 21586
rect 30716 21532 30884 21534
rect 30940 22036 30996 22046
rect 30716 21522 30772 21532
rect 30604 20862 30606 20914
rect 30658 20862 30660 20914
rect 30604 20850 30660 20862
rect 30716 21364 30772 21374
rect 30380 20066 30436 20076
rect 30492 20802 30548 20814
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30268 19908 30324 19918
rect 30492 19908 30548 20750
rect 30268 19906 30548 19908
rect 30268 19854 30270 19906
rect 30322 19854 30548 19906
rect 30268 19852 30548 19854
rect 30268 19842 30324 19852
rect 30716 19346 30772 21308
rect 30716 19294 30718 19346
rect 30770 19294 30772 19346
rect 30716 19282 30772 19294
rect 30828 19346 30884 19358
rect 30828 19294 30830 19346
rect 30882 19294 30884 19346
rect 29932 19236 29988 19246
rect 29932 19142 29988 19180
rect 30716 19124 30772 19134
rect 30044 18564 30100 18574
rect 29932 16212 29988 16222
rect 29932 13300 29988 16156
rect 29932 13234 29988 13244
rect 30044 16098 30100 18508
rect 30268 18452 30324 18462
rect 30268 18358 30324 18396
rect 30156 17668 30212 17678
rect 30156 17574 30212 17612
rect 30268 17108 30324 17118
rect 30268 17014 30324 17052
rect 30604 16324 30660 16334
rect 30604 16230 30660 16268
rect 30044 16046 30046 16098
rect 30098 16046 30100 16098
rect 30044 14308 30100 16046
rect 30604 16100 30660 16110
rect 30604 15764 30660 16044
rect 30268 15204 30324 15214
rect 30268 14868 30324 15148
rect 30268 14802 30324 14812
rect 30268 14532 30324 14542
rect 30268 14530 30548 14532
rect 30268 14478 30270 14530
rect 30322 14478 30548 14530
rect 30268 14476 30548 14478
rect 30268 14466 30324 14476
rect 29820 12014 29822 12066
rect 29874 12014 29876 12066
rect 29820 12002 29876 12014
rect 29484 11396 29540 11406
rect 29484 11302 29540 11340
rect 29372 11116 29540 11172
rect 29260 10892 29428 10948
rect 29260 10724 29316 10734
rect 29260 10630 29316 10668
rect 29372 6916 29428 10892
rect 29260 6860 29428 6916
rect 29260 5684 29316 6860
rect 29372 6692 29428 6702
rect 29372 6598 29428 6636
rect 29484 6580 29540 11116
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29596 10388 29652 10558
rect 29596 10322 29652 10332
rect 30044 10164 30100 14252
rect 30268 14084 30324 14094
rect 30156 13076 30212 13086
rect 30156 12290 30212 13020
rect 30156 12238 30158 12290
rect 30210 12238 30212 12290
rect 30156 12226 30212 12238
rect 30156 11844 30212 11854
rect 30268 11844 30324 14028
rect 30492 13970 30548 14476
rect 30604 14530 30660 15708
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14466 30660 14478
rect 30492 13918 30494 13970
rect 30546 13918 30548 13970
rect 30492 13906 30548 13918
rect 30716 12628 30772 19068
rect 30828 18788 30884 19294
rect 30828 18722 30884 18732
rect 30828 18450 30884 18462
rect 30828 18398 30830 18450
rect 30882 18398 30884 18450
rect 30828 18228 30884 18398
rect 30828 18162 30884 18172
rect 30716 12562 30772 12572
rect 30828 18004 30884 18014
rect 30212 11788 30324 11844
rect 30380 11956 30436 11966
rect 30156 11778 30212 11788
rect 30268 11508 30324 11518
rect 30156 11396 30212 11406
rect 30156 10610 30212 11340
rect 30268 11394 30324 11452
rect 30268 11342 30270 11394
rect 30322 11342 30324 11394
rect 30268 11330 30324 11342
rect 30380 10948 30436 11900
rect 30380 10882 30436 10892
rect 30156 10558 30158 10610
rect 30210 10558 30212 10610
rect 30156 10500 30212 10558
rect 30156 10434 30212 10444
rect 30268 10388 30324 10398
rect 30268 10294 30324 10332
rect 29820 10108 30100 10164
rect 29596 9828 29652 9838
rect 29596 9734 29652 9772
rect 29484 6514 29540 6524
rect 29260 5618 29316 5628
rect 29484 5908 29540 5918
rect 29820 5908 29876 10108
rect 30044 9938 30100 9950
rect 30044 9886 30046 9938
rect 30098 9886 30100 9938
rect 30044 9380 30100 9886
rect 30044 9314 30100 9324
rect 30380 8708 30436 8718
rect 30156 8148 30212 8158
rect 30156 8146 30324 8148
rect 30156 8094 30158 8146
rect 30210 8094 30324 8146
rect 30156 8092 30324 8094
rect 30156 8082 30212 8092
rect 29484 5906 29876 5908
rect 29484 5854 29486 5906
rect 29538 5854 29876 5906
rect 29484 5852 29876 5854
rect 30156 7924 30212 7934
rect 30156 6578 30212 7868
rect 30268 7474 30324 8092
rect 30380 7812 30436 8652
rect 30604 8596 30660 8606
rect 30380 7746 30436 7756
rect 30492 8484 30548 8494
rect 30268 7422 30270 7474
rect 30322 7422 30324 7474
rect 30268 7364 30324 7422
rect 30268 7028 30324 7308
rect 30268 6962 30324 6972
rect 30492 6804 30548 8428
rect 30604 8370 30660 8540
rect 30604 8318 30606 8370
rect 30658 8318 30660 8370
rect 30604 8306 30660 8318
rect 30492 6710 30548 6748
rect 30716 7924 30772 7934
rect 30716 7362 30772 7868
rect 30716 7310 30718 7362
rect 30770 7310 30772 7362
rect 30156 6526 30158 6578
rect 30210 6526 30212 6578
rect 29484 5460 29540 5852
rect 29932 5796 29988 5806
rect 29932 5702 29988 5740
rect 30156 5796 30212 6526
rect 30156 5730 30212 5740
rect 29148 4610 29204 4620
rect 29260 5404 29540 5460
rect 29148 3780 29204 3818
rect 28924 3724 29092 3780
rect 28812 3612 28980 3668
rect 28476 3502 28478 3554
rect 28530 3502 28532 3554
rect 28476 3490 28532 3502
rect 28700 3556 28756 3566
rect 28588 3108 28644 3118
rect 28588 2210 28644 3052
rect 28700 2882 28756 3500
rect 28700 2830 28702 2882
rect 28754 2830 28756 2882
rect 28700 2818 28756 2830
rect 28924 2548 28980 3612
rect 29036 3554 29092 3724
rect 29148 3714 29204 3724
rect 29036 3502 29038 3554
rect 29090 3502 29092 3554
rect 29036 3490 29092 3502
rect 29260 3388 29316 5404
rect 29148 3332 29316 3388
rect 29372 4788 29428 4798
rect 29372 3556 29428 4732
rect 30380 4788 30436 4798
rect 30156 4340 30212 4350
rect 29036 2660 29092 2670
rect 29036 2566 29092 2604
rect 28588 2158 28590 2210
rect 28642 2158 28644 2210
rect 28588 2146 28644 2158
rect 28812 2492 28980 2548
rect 28812 1428 28868 2492
rect 28924 2324 28980 2334
rect 28924 2210 28980 2268
rect 28924 2158 28926 2210
rect 28978 2158 28980 2210
rect 28924 2146 28980 2158
rect 28812 1362 28868 1372
rect 29148 1428 29204 3332
rect 29260 3220 29316 3230
rect 29260 2210 29316 3164
rect 29260 2158 29262 2210
rect 29314 2158 29316 2210
rect 29260 2146 29316 2158
rect 29148 1362 29204 1372
rect 28700 1316 28756 1326
rect 28700 1202 28756 1260
rect 28700 1150 28702 1202
rect 28754 1150 28756 1202
rect 28700 1138 28756 1150
rect 29372 1202 29428 3500
rect 29484 4338 30212 4340
rect 29484 4286 30158 4338
rect 30210 4286 30212 4338
rect 29484 4284 30212 4286
rect 29484 1876 29540 4284
rect 30156 4274 30212 4284
rect 29932 4116 29988 4126
rect 29708 4114 29988 4116
rect 29708 4062 29934 4114
rect 29986 4062 29988 4114
rect 29708 4060 29988 4062
rect 29596 2100 29652 2110
rect 29708 2100 29764 4060
rect 29932 4050 29988 4060
rect 29820 3554 29876 3566
rect 29820 3502 29822 3554
rect 29874 3502 29876 3554
rect 29820 3388 29876 3502
rect 30156 3556 30212 3566
rect 30156 3462 30212 3500
rect 29820 3332 30100 3388
rect 29932 3108 29988 3118
rect 30044 3108 30100 3332
rect 30044 3052 30324 3108
rect 29708 2044 29876 2100
rect 29596 2006 29652 2044
rect 29484 1820 29764 1876
rect 29372 1150 29374 1202
rect 29426 1150 29428 1202
rect 29372 1138 29428 1150
rect 29036 1092 29092 1102
rect 29036 998 29092 1036
rect 29708 1090 29764 1820
rect 29708 1038 29710 1090
rect 29762 1038 29764 1090
rect 29708 1026 29764 1038
rect 28028 700 28308 756
rect 28364 978 28420 990
rect 28364 926 28366 978
rect 28418 926 28420 978
rect 27580 532 27636 542
rect 27020 476 27188 532
rect 27132 112 27188 476
rect 27580 112 27636 476
rect 28028 112 28084 700
rect 28364 532 28420 926
rect 28364 466 28420 476
rect 28924 980 28980 990
rect 28476 308 28532 318
rect 28476 112 28532 252
rect 28924 112 28980 924
rect 29372 532 29428 542
rect 29372 112 29428 476
rect 29820 112 29876 2044
rect 29932 1540 29988 3052
rect 30268 2994 30324 3052
rect 30268 2942 30270 2994
rect 30322 2942 30324 2994
rect 30268 2930 30324 2942
rect 30268 2436 30324 2446
rect 29932 1474 29988 1484
rect 30044 1986 30100 1998
rect 30044 1934 30046 1986
rect 30098 1934 30100 1986
rect 30044 1428 30100 1934
rect 30268 1652 30324 2380
rect 30380 1988 30436 4732
rect 30604 4452 30660 4462
rect 30604 4358 30660 4396
rect 30716 3388 30772 7310
rect 30828 4340 30884 17948
rect 30940 17108 30996 21980
rect 31052 20020 31108 22764
rect 31164 22372 31220 22382
rect 31164 22278 31220 22316
rect 31276 20804 31332 20814
rect 31276 20710 31332 20748
rect 31052 19926 31108 19964
rect 31276 20132 31332 20142
rect 31052 19346 31108 19358
rect 31052 19294 31054 19346
rect 31106 19294 31108 19346
rect 31052 19236 31108 19294
rect 31164 19236 31220 19246
rect 31052 19234 31220 19236
rect 31052 19182 31166 19234
rect 31218 19182 31220 19234
rect 31052 19180 31220 19182
rect 31164 19170 31220 19180
rect 31276 19012 31332 20076
rect 31164 18956 31332 19012
rect 31052 17668 31108 17678
rect 31052 17574 31108 17612
rect 30940 17042 30996 17052
rect 31164 15988 31220 18956
rect 31164 15922 31220 15932
rect 31276 18340 31332 18350
rect 31164 13076 31220 13086
rect 31164 12290 31220 13020
rect 31164 12238 31166 12290
rect 31218 12238 31220 12290
rect 31164 12226 31220 12238
rect 31276 12180 31332 18284
rect 31388 16436 31444 22988
rect 31500 20020 31556 23996
rect 31724 21700 31780 24220
rect 31724 21634 31780 21644
rect 31612 21586 31668 21598
rect 31612 21534 31614 21586
rect 31666 21534 31668 21586
rect 31612 21252 31668 21534
rect 31948 21252 32004 28588
rect 32060 24612 32116 30828
rect 32508 30772 32564 31726
rect 32844 33628 33012 33684
rect 32732 30996 32788 31006
rect 32732 30902 32788 30940
rect 32060 24546 32116 24556
rect 32172 30716 32564 30772
rect 32732 30772 32788 30782
rect 32060 23492 32116 23502
rect 32060 23154 32116 23436
rect 32060 23102 32062 23154
rect 32114 23102 32116 23154
rect 32060 23090 32116 23102
rect 31612 21196 32004 21252
rect 31612 20580 31668 20590
rect 31612 20486 31668 20524
rect 31500 19954 31556 19964
rect 31500 19796 31556 19806
rect 31500 19702 31556 19740
rect 31612 19234 31668 19246
rect 31612 19182 31614 19234
rect 31666 19182 31668 19234
rect 31612 18788 31668 19182
rect 31836 19234 31892 19246
rect 31836 19182 31838 19234
rect 31890 19182 31892 19234
rect 31388 16370 31444 16380
rect 31500 18340 31556 18350
rect 31500 17668 31556 18284
rect 31612 17892 31668 18732
rect 31724 19122 31780 19134
rect 31724 19070 31726 19122
rect 31778 19070 31780 19122
rect 31724 18676 31780 19070
rect 31836 19124 31892 19182
rect 31836 19058 31892 19068
rect 31724 18620 31892 18676
rect 31724 18450 31780 18462
rect 31724 18398 31726 18450
rect 31778 18398 31780 18450
rect 31724 18116 31780 18398
rect 31724 18050 31780 18060
rect 31724 17892 31780 17902
rect 31612 17890 31780 17892
rect 31612 17838 31726 17890
rect 31778 17838 31780 17890
rect 31612 17836 31780 17838
rect 31724 17826 31780 17836
rect 31612 17668 31668 17678
rect 31500 17666 31668 17668
rect 31500 17614 31614 17666
rect 31666 17614 31668 17666
rect 31500 17612 31668 17614
rect 31276 12114 31332 12124
rect 31388 15876 31444 15886
rect 30940 10612 30996 10622
rect 31276 10612 31332 10622
rect 30940 10610 31220 10612
rect 30940 10558 30942 10610
rect 30994 10558 31220 10610
rect 30940 10556 31220 10558
rect 30940 10546 30996 10556
rect 31164 10052 31220 10556
rect 31276 10518 31332 10556
rect 31276 10052 31332 10062
rect 31164 10050 31332 10052
rect 31164 9998 31278 10050
rect 31330 9998 31332 10050
rect 31164 9996 31332 9998
rect 31276 9986 31332 9996
rect 31388 6692 31444 15820
rect 31500 15316 31556 17612
rect 31612 17602 31668 17612
rect 31724 17668 31780 17678
rect 31724 17442 31780 17612
rect 31724 17390 31726 17442
rect 31778 17390 31780 17442
rect 31724 17378 31780 17390
rect 31836 16884 31892 18620
rect 31836 16818 31892 16828
rect 31948 16548 32004 21196
rect 31948 16482 32004 16492
rect 32060 22596 32116 22606
rect 31500 15250 31556 15260
rect 31612 15988 31668 15998
rect 31612 15204 31668 15932
rect 31724 15874 31780 15886
rect 31724 15822 31726 15874
rect 31778 15822 31780 15874
rect 31724 15316 31780 15822
rect 31948 15652 32004 15662
rect 31948 15426 32004 15596
rect 31948 15374 31950 15426
rect 32002 15374 32004 15426
rect 31948 15362 32004 15374
rect 31724 15250 31780 15260
rect 31164 5682 31220 5694
rect 31164 5630 31166 5682
rect 31218 5630 31220 5682
rect 30828 4274 30884 4284
rect 31052 4340 31108 4350
rect 31164 4340 31220 5630
rect 31052 4338 31220 4340
rect 31052 4286 31054 4338
rect 31106 4286 31220 4338
rect 31052 4284 31220 4286
rect 31276 4452 31332 4462
rect 30716 3332 30884 3388
rect 30380 1922 30436 1932
rect 30492 3220 30548 3230
rect 30268 1586 30324 1596
rect 30044 1362 30100 1372
rect 30156 1204 30212 1214
rect 30156 1110 30212 1148
rect 30380 980 30436 990
rect 30380 886 30436 924
rect 30268 308 30324 318
rect 30268 112 30324 252
rect 30492 196 30548 3164
rect 30716 2658 30772 2670
rect 30716 2606 30718 2658
rect 30770 2606 30772 2658
rect 30716 2548 30772 2606
rect 30716 2482 30772 2492
rect 30604 2212 30660 2222
rect 30828 2212 30884 3332
rect 31052 2770 31108 4284
rect 31164 3556 31220 3566
rect 31164 3462 31220 3500
rect 31052 2718 31054 2770
rect 31106 2718 31108 2770
rect 31052 2706 31108 2718
rect 30604 2210 30884 2212
rect 30604 2158 30606 2210
rect 30658 2158 30884 2210
rect 30604 2156 30884 2158
rect 30604 2146 30660 2156
rect 31164 1764 31220 1774
rect 30492 130 30548 140
rect 30716 756 30772 766
rect 30716 112 30772 700
rect 31164 112 31220 1708
rect 31276 1204 31332 4396
rect 31388 4338 31444 6636
rect 31388 4286 31390 4338
rect 31442 4286 31444 4338
rect 31388 4274 31444 4286
rect 31500 15092 31668 15148
rect 31500 2770 31556 15092
rect 31612 14532 31668 14542
rect 31612 14438 31668 14476
rect 31836 14196 31892 14206
rect 31836 13860 31892 14140
rect 31836 13794 31892 13804
rect 31836 12852 31892 12862
rect 31724 12180 31780 12190
rect 31612 12068 31668 12078
rect 31612 11974 31668 12012
rect 31724 9604 31780 12124
rect 31836 11844 31892 12796
rect 31836 11778 31892 11788
rect 31724 9538 31780 9548
rect 32060 8930 32116 22540
rect 32172 22484 32228 30716
rect 32732 30212 32788 30716
rect 32508 30210 32788 30212
rect 32508 30158 32734 30210
rect 32786 30158 32788 30210
rect 32508 30156 32788 30158
rect 32396 30100 32452 30110
rect 32396 30006 32452 30044
rect 32508 29426 32564 30156
rect 32732 30146 32788 30156
rect 32508 29374 32510 29426
rect 32562 29374 32564 29426
rect 32508 29362 32564 29374
rect 32620 29540 32676 29550
rect 32396 29316 32452 29326
rect 32396 28754 32452 29260
rect 32396 28702 32398 28754
rect 32450 28702 32452 28754
rect 32396 28690 32452 28702
rect 32508 28084 32564 28094
rect 32620 28084 32676 29484
rect 32732 29092 32788 29102
rect 32732 28642 32788 29036
rect 32732 28590 32734 28642
rect 32786 28590 32788 28642
rect 32732 28578 32788 28590
rect 32508 28082 32676 28084
rect 32508 28030 32510 28082
rect 32562 28030 32676 28082
rect 32508 28028 32676 28030
rect 32508 27188 32564 28028
rect 32508 27122 32564 27132
rect 32732 26964 32788 26974
rect 32844 26964 32900 33628
rect 33068 33572 33124 33582
rect 33068 33478 33124 33516
rect 32956 33458 33012 33470
rect 32956 33406 32958 33458
rect 33010 33406 33012 33458
rect 32956 32452 33012 33406
rect 33068 32564 33124 32574
rect 33068 32470 33124 32508
rect 32956 32386 33012 32396
rect 33180 32340 33236 34748
rect 33068 32284 33236 32340
rect 33292 34132 33348 34142
rect 33068 31892 33124 32284
rect 33068 31798 33124 31836
rect 33180 32116 33236 32126
rect 33180 31668 33236 32060
rect 33068 31612 33236 31668
rect 32956 30770 33012 30782
rect 32956 30718 32958 30770
rect 33010 30718 33012 30770
rect 32956 30324 33012 30718
rect 32956 30258 33012 30268
rect 32956 29764 33012 29774
rect 33068 29764 33124 31612
rect 33180 30210 33236 30222
rect 33180 30158 33182 30210
rect 33234 30158 33236 30210
rect 33180 29988 33236 30158
rect 33180 29922 33236 29932
rect 33068 29708 33236 29764
rect 32956 29652 33012 29708
rect 32956 29596 33124 29652
rect 33068 29426 33124 29596
rect 33068 29374 33070 29426
rect 33122 29374 33124 29426
rect 32956 29316 33012 29326
rect 32956 29222 33012 29260
rect 33068 29092 33124 29374
rect 32956 29036 33124 29092
rect 32956 27188 33012 29036
rect 33068 28868 33124 28878
rect 33068 28082 33124 28812
rect 33180 28644 33236 29708
rect 33180 28550 33236 28588
rect 33068 28030 33070 28082
rect 33122 28030 33124 28082
rect 33068 28018 33124 28030
rect 32956 27122 33012 27132
rect 32788 26908 32900 26964
rect 32508 26852 32564 26862
rect 32508 26850 32676 26852
rect 32508 26798 32510 26850
rect 32562 26798 32676 26850
rect 32508 26796 32676 26798
rect 32508 26786 32564 26796
rect 32396 26292 32452 26302
rect 32396 25620 32452 26236
rect 32396 25554 32452 25564
rect 32620 25508 32676 26796
rect 32732 26292 32788 26908
rect 33292 26292 33348 34076
rect 33404 32452 33460 37214
rect 33516 37996 33796 38052
rect 33852 40180 33908 40190
rect 33516 37154 33572 37996
rect 33516 37102 33518 37154
rect 33570 37102 33572 37154
rect 33516 37090 33572 37102
rect 33628 37268 33684 37278
rect 33516 36594 33572 36606
rect 33516 36542 33518 36594
rect 33570 36542 33572 36594
rect 33516 33572 33572 36542
rect 33628 35140 33684 37212
rect 33852 37044 33908 40124
rect 33964 40068 34020 40350
rect 33964 40002 34020 40012
rect 34076 39620 34132 41244
rect 34188 41076 34244 45164
rect 34412 43428 34468 48524
rect 34524 47572 34580 47582
rect 34524 47478 34580 47516
rect 34636 47068 34692 49644
rect 34748 49250 34804 50372
rect 34748 49198 34750 49250
rect 34802 49198 34804 49250
rect 34748 49186 34804 49198
rect 34524 47012 34692 47068
rect 34748 48804 34804 48814
rect 34524 43876 34580 47012
rect 34748 46900 34804 48748
rect 34972 48580 35028 51772
rect 35084 51378 35140 52894
rect 35196 52946 35252 53116
rect 35196 52894 35198 52946
rect 35250 52894 35252 52946
rect 35196 52882 35252 52894
rect 35308 52722 35364 52734
rect 35308 52670 35310 52722
rect 35362 52670 35364 52722
rect 35308 52388 35364 52670
rect 35196 52332 35364 52388
rect 35420 52722 35476 52734
rect 35420 52670 35422 52722
rect 35474 52670 35476 52722
rect 35196 51828 35252 52332
rect 35420 52276 35476 52670
rect 35196 51762 35252 51772
rect 35308 52220 35476 52276
rect 35084 51326 35086 51378
rect 35138 51326 35140 51378
rect 35084 51314 35140 51326
rect 35196 51156 35252 51166
rect 35196 51062 35252 51100
rect 35084 50708 35140 50718
rect 35084 50706 35252 50708
rect 35084 50654 35086 50706
rect 35138 50654 35252 50706
rect 35084 50652 35252 50654
rect 35084 50642 35140 50652
rect 35084 50036 35140 50046
rect 35084 49942 35140 49980
rect 34972 48514 35028 48524
rect 35084 48356 35140 48366
rect 35084 48262 35140 48300
rect 34860 48244 34916 48254
rect 34860 48242 35028 48244
rect 34860 48190 34862 48242
rect 34914 48190 35028 48242
rect 34860 48188 35028 48190
rect 34860 48178 34916 48188
rect 34860 47236 34916 47246
rect 34860 47142 34916 47180
rect 34524 43810 34580 43820
rect 34636 46844 34804 46900
rect 34972 46900 35028 48188
rect 35196 48020 35252 50652
rect 35308 49364 35364 52220
rect 35420 52052 35476 52062
rect 35420 51958 35476 51996
rect 35532 51492 35588 54348
rect 35644 54068 35700 55358
rect 35980 55410 36036 56252
rect 36876 56196 36932 56206
rect 36428 56084 36484 56094
rect 36428 55990 36484 56028
rect 36876 56082 36932 56140
rect 36876 56030 36878 56082
rect 36930 56030 36932 56082
rect 36876 56018 36932 56030
rect 36988 56084 37044 57344
rect 36988 56018 37044 56028
rect 37324 56868 37380 56878
rect 36092 55860 36148 55870
rect 36092 55766 36148 55804
rect 37100 55860 37156 55870
rect 37100 55766 37156 55804
rect 35980 55358 35982 55410
rect 36034 55358 36036 55410
rect 35980 55346 36036 55358
rect 36316 55412 36372 55422
rect 36316 55318 36372 55356
rect 37212 55410 37268 55422
rect 37212 55358 37214 55410
rect 37266 55358 37268 55410
rect 35644 54002 35700 54012
rect 36540 54514 36596 54526
rect 36540 54462 36542 54514
rect 36594 54462 36596 54514
rect 35756 53844 35812 53854
rect 35756 53750 35812 53788
rect 36540 53620 36596 54462
rect 36876 54402 36932 54414
rect 36876 54350 36878 54402
rect 36930 54350 36932 54402
rect 36876 53844 36932 54350
rect 36876 53778 36932 53788
rect 36540 53554 36596 53564
rect 36988 53506 37044 53518
rect 36988 53454 36990 53506
rect 37042 53454 37044 53506
rect 36988 53060 37044 53454
rect 37100 53060 37156 53070
rect 36988 53058 37156 53060
rect 36988 53006 37102 53058
rect 37154 53006 37156 53058
rect 36988 53004 37156 53006
rect 37100 52994 37156 53004
rect 36540 52836 36596 52846
rect 35644 52724 35700 52734
rect 35644 51828 35700 52668
rect 36428 52722 36484 52734
rect 36428 52670 36430 52722
rect 36482 52670 36484 52722
rect 35868 52276 35924 52286
rect 35868 52182 35924 52220
rect 36428 52164 36484 52670
rect 36428 52098 36484 52108
rect 35644 51762 35700 51772
rect 36540 51604 36596 52780
rect 36764 52722 36820 52734
rect 36764 52670 36766 52722
rect 36818 52670 36820 52722
rect 36764 52388 36820 52670
rect 36764 52322 36820 52332
rect 36876 52724 36932 52734
rect 36540 51538 36596 51548
rect 36428 51492 36484 51502
rect 35532 51490 36484 51492
rect 35532 51438 36430 51490
rect 36482 51438 36484 51490
rect 35532 51436 36484 51438
rect 35420 51380 35476 51390
rect 35532 51380 35588 51436
rect 36428 51426 36484 51436
rect 36652 51490 36708 51502
rect 36652 51438 36654 51490
rect 36706 51438 36708 51490
rect 35420 51378 35588 51380
rect 35420 51326 35422 51378
rect 35474 51326 35588 51378
rect 35420 51324 35588 51326
rect 36540 51380 36596 51390
rect 35420 51314 35476 51324
rect 36316 51268 36372 51278
rect 36204 51266 36372 51268
rect 36204 51214 36318 51266
rect 36370 51214 36372 51266
rect 36204 51212 36372 51214
rect 35420 51156 35476 51166
rect 35420 50706 35476 51100
rect 35420 50654 35422 50706
rect 35474 50654 35476 50706
rect 35420 50642 35476 50654
rect 35532 51154 35588 51166
rect 35532 51102 35534 51154
rect 35586 51102 35588 51154
rect 35420 50036 35476 50046
rect 35532 50036 35588 51102
rect 35644 51156 35700 51166
rect 35644 51154 36148 51156
rect 35644 51102 35646 51154
rect 35698 51102 36148 51154
rect 35644 51100 36148 51102
rect 35644 51090 35700 51100
rect 35980 50820 36036 50830
rect 35980 50726 36036 50764
rect 35644 50596 35700 50606
rect 35644 50502 35700 50540
rect 35420 50034 35588 50036
rect 35420 49982 35422 50034
rect 35474 49982 35588 50034
rect 35420 49980 35588 49982
rect 35868 50484 35924 50494
rect 35420 49970 35476 49980
rect 35644 49812 35700 49822
rect 35308 49308 35588 49364
rect 35308 49140 35364 49150
rect 35308 48468 35364 49084
rect 35308 48402 35364 48412
rect 35532 48244 35588 49308
rect 35532 48150 35588 48188
rect 35196 47954 35252 47964
rect 35308 48018 35364 48030
rect 35308 47966 35310 48018
rect 35362 47966 35364 48018
rect 35308 47684 35364 47966
rect 35420 48020 35476 48030
rect 35644 48020 35700 49756
rect 35868 49250 35924 50428
rect 35868 49198 35870 49250
rect 35922 49198 35924 49250
rect 35868 49186 35924 49198
rect 35980 49028 36036 49038
rect 35980 48132 36036 48972
rect 36092 48244 36148 51100
rect 36204 50932 36260 51212
rect 36316 51202 36372 51212
rect 36540 51266 36596 51324
rect 36540 51214 36542 51266
rect 36594 51214 36596 51266
rect 36540 51202 36596 51214
rect 36204 50708 36260 50876
rect 36204 50642 36260 50652
rect 36428 50708 36484 50718
rect 36428 50614 36484 50652
rect 36428 50036 36484 50046
rect 36428 49942 36484 49980
rect 36316 49252 36372 49262
rect 36316 48914 36372 49196
rect 36316 48862 36318 48914
rect 36370 48862 36372 48914
rect 36316 48804 36372 48862
rect 36316 48738 36372 48748
rect 36540 48916 36596 48926
rect 36428 48244 36484 48254
rect 36092 48242 36484 48244
rect 36092 48190 36430 48242
rect 36482 48190 36484 48242
rect 36092 48188 36484 48190
rect 35980 48076 36260 48132
rect 35420 48018 35588 48020
rect 35420 47966 35422 48018
rect 35474 47966 35588 48018
rect 35420 47964 35588 47966
rect 35644 47964 36148 48020
rect 35420 47954 35476 47964
rect 35308 47628 35476 47684
rect 35308 47458 35364 47470
rect 35308 47406 35310 47458
rect 35362 47406 35364 47458
rect 35308 47012 35364 47406
rect 35308 46946 35364 46956
rect 35084 46900 35140 46910
rect 34972 46898 35140 46900
rect 34972 46846 35086 46898
rect 35138 46846 35140 46898
rect 34972 46844 35140 46846
rect 34412 43362 34468 43372
rect 34636 42980 34692 46844
rect 35084 46834 35140 46844
rect 34748 46676 34804 46686
rect 34748 46114 34804 46620
rect 35420 46676 35476 47628
rect 35420 46610 35476 46620
rect 35420 46450 35476 46462
rect 35420 46398 35422 46450
rect 35474 46398 35476 46450
rect 34748 46062 34750 46114
rect 34802 46062 34804 46114
rect 34748 46050 34804 46062
rect 34860 46228 34916 46238
rect 34748 44884 34804 44894
rect 34748 44790 34804 44828
rect 34860 44322 34916 46172
rect 34860 44270 34862 44322
rect 34914 44270 34916 44322
rect 34748 43652 34804 43662
rect 34748 43558 34804 43596
rect 34748 43092 34804 43102
rect 34860 43092 34916 44270
rect 35084 46004 35140 46014
rect 35084 44436 35140 45948
rect 35308 46004 35364 46014
rect 35308 45556 35364 45948
rect 35252 45500 35364 45556
rect 35252 45342 35308 45500
rect 35252 45330 35364 45342
rect 35252 45278 35310 45330
rect 35362 45278 35364 45330
rect 35252 45276 35364 45278
rect 35308 45266 35364 45276
rect 35196 44436 35252 44446
rect 35084 44434 35252 44436
rect 35084 44382 35198 44434
rect 35250 44382 35252 44434
rect 35084 44380 35252 44382
rect 34804 43036 34916 43092
rect 34748 43026 34804 43036
rect 34636 42914 34692 42924
rect 34860 42754 34916 43036
rect 34860 42702 34862 42754
rect 34914 42702 34916 42754
rect 34860 42690 34916 42702
rect 34972 43092 35028 43102
rect 34972 42196 35028 43036
rect 35084 42756 35140 44380
rect 35196 44370 35252 44380
rect 35308 43988 35364 43998
rect 35196 43538 35252 43550
rect 35196 43486 35198 43538
rect 35250 43486 35252 43538
rect 35196 43092 35252 43486
rect 35196 43026 35252 43036
rect 35308 42978 35364 43932
rect 35308 42926 35310 42978
rect 35362 42926 35364 42978
rect 35308 42914 35364 42926
rect 35084 42700 35364 42756
rect 34972 42140 35140 42196
rect 35084 42084 35140 42140
rect 35084 42018 35140 42028
rect 34524 41972 34580 41982
rect 34972 41972 35028 41982
rect 34412 41858 34468 41870
rect 34412 41806 34414 41858
rect 34466 41806 34468 41858
rect 34412 41300 34468 41806
rect 34524 41858 34580 41916
rect 34524 41806 34526 41858
rect 34578 41806 34580 41858
rect 34524 41794 34580 41806
rect 34636 41970 35028 41972
rect 34636 41918 34974 41970
rect 35026 41918 35028 41970
rect 34636 41916 35028 41918
rect 34412 41234 34468 41244
rect 34636 41412 34692 41916
rect 34972 41906 35028 41916
rect 35196 41860 35252 41870
rect 34748 41748 34804 41786
rect 35196 41766 35252 41804
rect 34748 41682 34804 41692
rect 35308 41636 35364 42700
rect 35420 41970 35476 46398
rect 35532 46004 35588 47964
rect 35644 47572 35700 47582
rect 35644 47478 35700 47516
rect 35756 46564 35812 46574
rect 35756 46562 36036 46564
rect 35756 46510 35758 46562
rect 35810 46510 36036 46562
rect 35756 46508 36036 46510
rect 35756 46498 35812 46508
rect 35532 45938 35588 45948
rect 35644 46450 35700 46462
rect 35644 46398 35646 46450
rect 35698 46398 35700 46450
rect 35644 45780 35700 46398
rect 35868 46004 35924 46014
rect 35868 45910 35924 45948
rect 35644 45724 35812 45780
rect 35644 45556 35700 45566
rect 35644 45330 35700 45500
rect 35644 45278 35646 45330
rect 35698 45278 35700 45330
rect 35644 45266 35700 45278
rect 35532 44882 35588 44894
rect 35532 44830 35534 44882
rect 35586 44830 35588 44882
rect 35532 44548 35588 44830
rect 35532 44482 35588 44492
rect 35756 43652 35812 45724
rect 35420 41918 35422 41970
rect 35474 41918 35476 41970
rect 35420 41906 35476 41918
rect 35532 43596 35812 43652
rect 35532 43538 35588 43596
rect 35532 43486 35534 43538
rect 35586 43486 35588 43538
rect 35532 42980 35588 43486
rect 35644 43428 35700 43438
rect 35644 43334 35700 43372
rect 35756 43316 35812 43326
rect 35756 43314 35924 43316
rect 35756 43262 35758 43314
rect 35810 43262 35924 43314
rect 35756 43260 35924 43262
rect 35756 43250 35812 43260
rect 35532 41860 35588 42924
rect 35644 43092 35700 43102
rect 35644 41970 35700 43036
rect 35756 42868 35812 42878
rect 35756 42082 35812 42812
rect 35756 42030 35758 42082
rect 35810 42030 35812 42082
rect 35756 42018 35812 42030
rect 35644 41918 35646 41970
rect 35698 41918 35700 41970
rect 35644 41906 35700 41918
rect 35532 41794 35588 41804
rect 35308 41580 35812 41636
rect 34188 41020 34468 41076
rect 34300 40740 34356 40750
rect 34076 38948 34132 39564
rect 34076 38882 34132 38892
rect 34188 39732 34244 39742
rect 33852 36978 33908 36988
rect 33964 38724 34020 38734
rect 33964 36820 34020 38668
rect 34076 38612 34132 38622
rect 34076 38162 34132 38556
rect 34076 38110 34078 38162
rect 34130 38110 34132 38162
rect 34076 38098 34132 38110
rect 33852 36764 34020 36820
rect 34076 37380 34132 37390
rect 34076 36820 34132 37324
rect 34188 37266 34244 39676
rect 34188 37214 34190 37266
rect 34242 37214 34244 37266
rect 34188 37202 34244 37214
rect 34076 36764 34244 36820
rect 33740 36036 33796 36046
rect 33740 35698 33796 35980
rect 33740 35646 33742 35698
rect 33794 35646 33796 35698
rect 33740 35634 33796 35646
rect 33628 35046 33684 35084
rect 33628 34804 33684 34814
rect 33628 34244 33684 34748
rect 33628 34150 33684 34188
rect 33740 34468 33796 34478
rect 33740 34132 33796 34412
rect 33740 34066 33796 34076
rect 33516 33506 33572 33516
rect 33628 33908 33684 33918
rect 33516 33348 33572 33358
rect 33516 32676 33572 33292
rect 33516 32610 33572 32620
rect 33404 32386 33460 32396
rect 33628 31220 33684 33852
rect 33852 33348 33908 36764
rect 33964 36596 34020 36606
rect 33964 36036 34020 36540
rect 33964 35970 34020 35980
rect 34188 35586 34244 36764
rect 34188 35534 34190 35586
rect 34242 35534 34244 35586
rect 34188 35476 34244 35534
rect 34188 35410 34244 35420
rect 33852 33282 33908 33292
rect 33964 35028 34020 35038
rect 33964 34804 34020 34972
rect 34076 34804 34132 34814
rect 33964 34802 34132 34804
rect 33964 34750 34078 34802
rect 34130 34750 34132 34802
rect 33964 34748 34132 34750
rect 33964 33124 34020 34748
rect 34076 34738 34132 34748
rect 34300 34244 34356 40684
rect 33740 33068 34020 33124
rect 34076 34020 34132 34030
rect 34300 34020 34356 34188
rect 34076 34018 34356 34020
rect 34076 33966 34078 34018
rect 34130 33966 34356 34018
rect 34076 33964 34356 33966
rect 33740 31332 33796 33068
rect 34076 32788 34132 33964
rect 34412 33572 34468 41020
rect 34524 40962 34580 40974
rect 34524 40910 34526 40962
rect 34578 40910 34580 40962
rect 34524 39732 34580 40910
rect 34636 40852 34692 41356
rect 34636 40786 34692 40796
rect 34748 41524 34804 41534
rect 34524 39666 34580 39676
rect 34636 38724 34692 38762
rect 34636 38658 34692 38668
rect 34748 38276 34804 41468
rect 35308 41300 35364 41310
rect 35084 41188 35140 41198
rect 34524 38220 34804 38276
rect 34860 41186 35140 41188
rect 34860 41134 35086 41186
rect 35138 41134 35140 41186
rect 34860 41132 35140 41134
rect 34860 39618 34916 41132
rect 35084 41122 35140 41132
rect 35196 40740 35252 40750
rect 35084 40404 35140 40414
rect 35084 40310 35140 40348
rect 34860 39566 34862 39618
rect 34914 39566 34916 39618
rect 34524 34804 34580 38220
rect 34860 38164 34916 39566
rect 34636 38050 34692 38062
rect 34636 37998 34638 38050
rect 34690 37998 34692 38050
rect 34636 37266 34692 37998
rect 34860 37492 34916 38108
rect 34636 37214 34638 37266
rect 34690 37214 34692 37266
rect 34636 35308 34692 37214
rect 34748 37436 34916 37492
rect 34972 40292 35028 40302
rect 34748 37156 34804 37436
rect 34748 37090 34804 37100
rect 34860 37268 34916 37278
rect 34748 36484 34804 36494
rect 34748 36390 34804 36428
rect 34636 35252 34804 35308
rect 34636 34804 34692 34814
rect 34524 34802 34692 34804
rect 34524 34750 34638 34802
rect 34690 34750 34692 34802
rect 34524 34748 34692 34750
rect 34636 34468 34692 34748
rect 34636 34402 34692 34412
rect 34188 33124 34244 33134
rect 34188 33030 34244 33068
rect 34076 32722 34132 32732
rect 34412 32562 34468 33516
rect 34412 32510 34414 32562
rect 34466 32510 34468 32562
rect 34412 32498 34468 32510
rect 34524 34132 34580 34142
rect 33852 32452 33908 32462
rect 34300 32452 34356 32462
rect 33852 32450 34244 32452
rect 33852 32398 33854 32450
rect 33906 32398 34244 32450
rect 33852 32396 34244 32398
rect 33852 32386 33908 32396
rect 34188 32002 34244 32396
rect 34300 32358 34356 32396
rect 34188 31950 34190 32002
rect 34242 31950 34244 32002
rect 34188 31938 34244 31950
rect 33740 31266 33796 31276
rect 34076 31444 34132 31454
rect 33628 31154 33684 31164
rect 33964 31108 34020 31118
rect 33404 30882 33460 30894
rect 33404 30830 33406 30882
rect 33458 30830 33460 30882
rect 33404 30772 33460 30830
rect 33404 30706 33460 30716
rect 33404 30322 33460 30334
rect 33404 30270 33406 30322
rect 33458 30270 33460 30322
rect 33404 30212 33460 30270
rect 33404 30146 33460 30156
rect 33628 30212 33684 30222
rect 33628 29428 33684 30156
rect 33964 30212 34020 31052
rect 34076 30994 34132 31388
rect 34076 30942 34078 30994
rect 34130 30942 34132 30994
rect 34076 30930 34132 30942
rect 34412 30884 34468 30894
rect 33964 30118 34020 30156
rect 34076 30772 34132 30782
rect 33964 29876 34020 29886
rect 33964 29538 34020 29820
rect 33964 29486 33966 29538
rect 34018 29486 34020 29538
rect 33964 29474 34020 29486
rect 33516 29426 33684 29428
rect 33516 29374 33630 29426
rect 33682 29374 33684 29426
rect 33516 29372 33684 29374
rect 33516 29092 33572 29372
rect 33628 29362 33684 29372
rect 33516 29026 33572 29036
rect 33964 29092 34020 29102
rect 33404 28754 33460 28766
rect 33404 28702 33406 28754
rect 33458 28702 33460 28754
rect 33404 28644 33460 28702
rect 33964 28644 34020 29036
rect 33404 28578 33460 28588
rect 33852 28588 34020 28644
rect 34076 28642 34132 30716
rect 34188 30548 34244 30558
rect 34188 29876 34244 30492
rect 34188 29810 34244 29820
rect 34300 29316 34356 29326
rect 34300 29222 34356 29260
rect 34076 28590 34078 28642
rect 34130 28590 34132 28642
rect 33740 27524 33796 27534
rect 33740 27188 33796 27468
rect 32732 26226 32788 26236
rect 33180 26236 33348 26292
rect 33404 27186 33796 27188
rect 33404 27134 33742 27186
rect 33794 27134 33796 27186
rect 33404 27132 33796 27134
rect 32956 26066 33012 26078
rect 32956 26014 32958 26066
rect 33010 26014 33012 26066
rect 32956 25620 33012 26014
rect 32956 25554 33012 25564
rect 33068 26068 33124 26078
rect 32620 25442 32676 25452
rect 32620 25282 32676 25294
rect 32620 25230 32622 25282
rect 32674 25230 32676 25282
rect 32284 25060 32340 25070
rect 32284 23044 32340 25004
rect 32620 24724 32676 25230
rect 32956 25284 33012 25294
rect 33068 25284 33124 26012
rect 32956 25282 33124 25284
rect 32956 25230 32958 25282
rect 33010 25230 33124 25282
rect 32956 25228 33124 25230
rect 32956 25218 33012 25228
rect 32956 25060 33012 25070
rect 32732 24724 32788 24734
rect 32620 24722 32788 24724
rect 32620 24670 32734 24722
rect 32786 24670 32788 24722
rect 32620 24668 32788 24670
rect 32732 24658 32788 24668
rect 32956 24722 33012 25004
rect 32956 24670 32958 24722
rect 33010 24670 33012 24722
rect 32956 24658 33012 24670
rect 32844 24498 32900 24510
rect 32844 24446 32846 24498
rect 32898 24446 32900 24498
rect 32508 24388 32564 24398
rect 32284 22978 32340 22988
rect 32396 24164 32452 24174
rect 32172 22418 32228 22428
rect 32396 21698 32452 24108
rect 32508 24162 32564 24332
rect 32508 24110 32510 24162
rect 32562 24110 32564 24162
rect 32508 24098 32564 24110
rect 32844 24164 32900 24446
rect 32844 24098 32900 24108
rect 33068 24052 33124 25228
rect 33068 23986 33124 23996
rect 33180 23828 33236 26236
rect 33292 26068 33348 26078
rect 33292 24722 33348 26012
rect 33292 24670 33294 24722
rect 33346 24670 33348 24722
rect 33292 24658 33348 24670
rect 32844 23772 33236 23828
rect 33292 24388 33348 24398
rect 32508 23492 32564 23502
rect 32508 22036 32564 23436
rect 32732 23492 32788 23502
rect 32620 23156 32676 23166
rect 32620 23062 32676 23100
rect 32508 21810 32564 21980
rect 32508 21758 32510 21810
rect 32562 21758 32564 21810
rect 32508 21746 32564 21758
rect 32396 21646 32398 21698
rect 32450 21646 32452 21698
rect 32396 21364 32452 21646
rect 32396 21298 32452 21308
rect 32620 21364 32676 21374
rect 32620 21028 32676 21308
rect 32732 21028 32788 23436
rect 32844 22482 32900 23772
rect 33292 23548 33348 24332
rect 32844 22430 32846 22482
rect 32898 22430 32900 22482
rect 32844 22418 32900 22430
rect 32956 23492 33012 23502
rect 32956 21586 33012 23436
rect 33180 23492 33348 23548
rect 33404 23604 33460 27132
rect 33740 27122 33796 27132
rect 33852 26516 33908 28588
rect 34076 28578 34132 28590
rect 34412 28642 34468 30828
rect 34524 30210 34580 34076
rect 34748 32676 34804 35252
rect 34860 34804 34916 37212
rect 34860 34738 34916 34748
rect 34748 32610 34804 32620
rect 34860 33124 34916 33134
rect 34860 32562 34916 33068
rect 34972 32788 35028 40236
rect 35196 39730 35252 40684
rect 35308 40068 35364 41244
rect 35644 41298 35700 41310
rect 35644 41246 35646 41298
rect 35698 41246 35700 41298
rect 35420 40964 35476 40974
rect 35420 40290 35476 40908
rect 35644 40516 35700 41246
rect 35756 41300 35812 41580
rect 35868 41524 35924 43260
rect 35868 41458 35924 41468
rect 35980 41300 36036 46508
rect 36092 44324 36148 47964
rect 36092 44258 36148 44268
rect 36204 43988 36260 48076
rect 36316 47348 36372 47358
rect 36428 47348 36484 48188
rect 36540 47796 36596 48860
rect 36652 48466 36708 51438
rect 36764 51380 36820 51390
rect 36764 50594 36820 51324
rect 36764 50542 36766 50594
rect 36818 50542 36820 50594
rect 36764 50530 36820 50542
rect 36876 50484 36932 52668
rect 36988 51938 37044 51950
rect 36988 51886 36990 51938
rect 37042 51886 37044 51938
rect 36988 50708 37044 51886
rect 37212 50820 37268 55358
rect 37212 50754 37268 50764
rect 36988 50642 37044 50652
rect 36876 50418 36932 50428
rect 37212 50594 37268 50606
rect 37212 50542 37214 50594
rect 37266 50542 37268 50594
rect 37212 50036 37268 50542
rect 37324 50484 37380 56812
rect 37436 56196 37492 57344
rect 37436 56130 37492 56140
rect 37548 56084 37604 56094
rect 37884 56084 37940 57344
rect 37548 56082 37940 56084
rect 37548 56030 37550 56082
rect 37602 56030 37940 56082
rect 37548 56028 37940 56030
rect 37548 56018 37604 56028
rect 37772 55858 37828 55870
rect 37772 55806 37774 55858
rect 37826 55806 37828 55858
rect 37772 55524 37828 55806
rect 38108 55860 38164 55870
rect 38108 55766 38164 55804
rect 38332 55524 38388 57344
rect 38780 56756 38836 57344
rect 38444 56700 38836 56756
rect 38444 56082 38500 56700
rect 38444 56030 38446 56082
rect 38498 56030 38500 56082
rect 38444 56018 38500 56030
rect 38780 56532 38836 56542
rect 38668 55748 38724 55758
rect 38556 55524 38612 55534
rect 38332 55522 38612 55524
rect 38332 55470 38558 55522
rect 38610 55470 38612 55522
rect 38332 55468 38612 55470
rect 37772 55458 37828 55468
rect 38556 55458 38612 55468
rect 37548 55412 37604 55422
rect 37548 55318 37604 55356
rect 38668 55188 38724 55692
rect 38668 55122 38724 55132
rect 37772 55074 37828 55086
rect 37772 55022 37774 55074
rect 37826 55022 37828 55074
rect 37548 54740 37604 54750
rect 37436 52946 37492 52958
rect 37436 52894 37438 52946
rect 37490 52894 37492 52946
rect 37436 51380 37492 52894
rect 37436 51314 37492 51324
rect 37436 50706 37492 50718
rect 37436 50654 37438 50706
rect 37490 50654 37492 50706
rect 37436 50596 37492 50654
rect 37436 50530 37492 50540
rect 37324 50418 37380 50428
rect 37212 49970 37268 49980
rect 37324 49924 37380 49934
rect 37100 49812 37156 49822
rect 37100 49028 37156 49756
rect 36652 48414 36654 48466
rect 36706 48414 36708 48466
rect 36652 48402 36708 48414
rect 36988 49026 37156 49028
rect 36988 48974 37102 49026
rect 37154 48974 37156 49026
rect 36988 48972 37156 48974
rect 36876 48130 36932 48142
rect 36876 48078 36878 48130
rect 36930 48078 36932 48130
rect 36540 47740 36820 47796
rect 36652 47570 36708 47582
rect 36652 47518 36654 47570
rect 36706 47518 36708 47570
rect 36428 47292 36596 47348
rect 36316 45780 36372 47292
rect 36428 47124 36484 47134
rect 36428 46898 36484 47068
rect 36428 46846 36430 46898
rect 36482 46846 36484 46898
rect 36428 46834 36484 46846
rect 36316 45686 36372 45724
rect 36540 45444 36596 47292
rect 36652 46228 36708 47518
rect 36764 47460 36820 47740
rect 36764 47394 36820 47404
rect 36876 47012 36932 48078
rect 36988 47348 37044 48972
rect 37100 48962 37156 48972
rect 36988 47282 37044 47292
rect 37100 48242 37156 48254
rect 37100 48190 37102 48242
rect 37154 48190 37156 48242
rect 36764 46788 36820 46798
rect 36764 46694 36820 46732
rect 36876 46564 36932 46956
rect 36988 46564 37044 46574
rect 36876 46562 37044 46564
rect 36876 46510 36990 46562
rect 37042 46510 37044 46562
rect 36876 46508 37044 46510
rect 36988 46498 37044 46508
rect 36652 46162 36708 46172
rect 36988 46340 37044 46350
rect 36988 45890 37044 46284
rect 37100 46004 37156 48190
rect 37212 48132 37268 48142
rect 37212 48038 37268 48076
rect 37324 47348 37380 49868
rect 37548 49924 37604 54684
rect 37772 54740 37828 55022
rect 38108 55074 38164 55086
rect 38108 55022 38110 55074
rect 38162 55022 38164 55074
rect 38108 54852 38164 55022
rect 38108 54786 38164 54796
rect 37772 54674 37828 54684
rect 38668 54740 38724 54750
rect 38668 54646 38724 54684
rect 38108 54290 38164 54302
rect 38108 54238 38110 54290
rect 38162 54238 38164 54290
rect 37772 53620 37828 53630
rect 37772 52052 37828 53564
rect 37996 52948 38052 52958
rect 38108 52948 38164 54238
rect 37996 52946 38164 52948
rect 37996 52894 37998 52946
rect 38050 52894 38164 52946
rect 37996 52892 38164 52894
rect 38220 53842 38276 53854
rect 38220 53790 38222 53842
rect 38274 53790 38276 53842
rect 37996 52882 38052 52892
rect 38108 52724 38164 52734
rect 38108 52630 38164 52668
rect 37996 52052 38052 52062
rect 37660 52050 38052 52052
rect 37660 51998 37998 52050
rect 38050 51998 38052 52050
rect 37660 51996 38052 51998
rect 37660 51490 37716 51996
rect 37660 51438 37662 51490
rect 37714 51438 37716 51490
rect 37660 51426 37716 51438
rect 37772 51380 37828 51390
rect 37548 49858 37604 49868
rect 37660 50708 37716 50718
rect 37660 49698 37716 50652
rect 37660 49646 37662 49698
rect 37714 49646 37716 49698
rect 37660 49634 37716 49646
rect 37324 47282 37380 47292
rect 37436 49364 37492 49374
rect 37436 49138 37492 49308
rect 37436 49086 37438 49138
rect 37490 49086 37492 49138
rect 37436 46788 37492 49086
rect 37436 46722 37492 46732
rect 37548 49252 37604 49262
rect 37772 49252 37828 51324
rect 37884 50932 37940 50942
rect 37884 50706 37940 50876
rect 37884 50654 37886 50706
rect 37938 50654 37940 50706
rect 37884 50596 37940 50654
rect 37884 50530 37940 50540
rect 37996 50036 38052 51996
rect 38108 52052 38164 52062
rect 38108 51268 38164 51996
rect 38108 51174 38164 51212
rect 38108 50036 38164 50046
rect 37996 49980 38108 50036
rect 38108 49812 38164 49980
rect 38108 49718 38164 49756
rect 37772 49196 38164 49252
rect 37324 46562 37380 46574
rect 37324 46510 37326 46562
rect 37378 46510 37380 46562
rect 37100 45948 37268 46004
rect 36988 45838 36990 45890
rect 37042 45838 37044 45890
rect 36988 45826 37044 45838
rect 36540 45378 36596 45388
rect 37212 45108 37268 45948
rect 37324 45556 37380 46510
rect 37548 46452 37604 49196
rect 37996 49028 38052 49038
rect 37996 48804 38052 48972
rect 37660 48132 37716 48142
rect 37660 48130 37940 48132
rect 37660 48078 37662 48130
rect 37714 48078 37940 48130
rect 37660 48076 37940 48078
rect 37660 48066 37716 48076
rect 37548 46386 37604 46396
rect 37772 47684 37828 47694
rect 37772 46452 37828 47628
rect 37884 47682 37940 48076
rect 37884 47630 37886 47682
rect 37938 47630 37940 47682
rect 37884 47618 37940 47630
rect 37772 46386 37828 46396
rect 37996 46340 38052 48748
rect 37996 46274 38052 46284
rect 38108 48242 38164 49196
rect 38108 48190 38110 48242
rect 38162 48190 38164 48242
rect 37436 46228 37492 46238
rect 37436 46002 37492 46172
rect 37436 45950 37438 46002
rect 37490 45950 37492 46002
rect 37436 45938 37492 45950
rect 37324 45490 37380 45500
rect 37436 45780 37492 45790
rect 37212 45042 37268 45052
rect 37436 45108 37492 45724
rect 37436 45106 37604 45108
rect 37436 45054 37438 45106
rect 37490 45054 37604 45106
rect 37436 45052 37604 45054
rect 37436 45042 37492 45052
rect 36652 44882 36708 44894
rect 36652 44830 36654 44882
rect 36706 44830 36708 44882
rect 36204 43922 36260 43932
rect 36428 44098 36484 44110
rect 36428 44046 36430 44098
rect 36482 44046 36484 44098
rect 36428 43540 36484 44046
rect 36652 43988 36708 44830
rect 36988 44884 37044 44894
rect 37324 44884 37380 44894
rect 36988 44882 37268 44884
rect 36988 44830 36990 44882
rect 37042 44830 37268 44882
rect 36988 44828 37268 44830
rect 36988 44818 37044 44828
rect 37100 44324 37156 44334
rect 37100 44230 37156 44268
rect 36652 43922 36708 43932
rect 36764 44212 36820 44222
rect 36092 43484 36484 43540
rect 36652 43764 36708 43774
rect 36092 43092 36148 43484
rect 36428 43316 36484 43326
rect 36092 43026 36148 43036
rect 36204 43314 36484 43316
rect 36204 43262 36430 43314
rect 36482 43262 36484 43314
rect 36204 43260 36484 43262
rect 35756 41244 35924 41300
rect 35644 40450 35700 40460
rect 35420 40238 35422 40290
rect 35474 40238 35476 40290
rect 35420 40226 35476 40238
rect 35756 40292 35812 40302
rect 35756 40198 35812 40236
rect 35532 40178 35588 40190
rect 35532 40126 35534 40178
rect 35586 40126 35588 40178
rect 35308 40012 35476 40068
rect 35196 39678 35198 39730
rect 35250 39678 35252 39730
rect 35196 39666 35252 39678
rect 35084 39620 35140 39630
rect 35084 38946 35140 39564
rect 35084 38894 35086 38946
rect 35138 38894 35140 38946
rect 35084 38882 35140 38894
rect 35308 39508 35364 39518
rect 35196 36932 35252 36942
rect 35196 36596 35252 36876
rect 35196 36502 35252 36540
rect 35308 36820 35364 39452
rect 35084 34914 35140 34926
rect 35084 34862 35086 34914
rect 35138 34862 35140 34914
rect 35084 34356 35140 34862
rect 35308 34916 35364 36764
rect 35420 36260 35476 40012
rect 35532 39060 35588 40126
rect 35644 40178 35700 40190
rect 35644 40126 35646 40178
rect 35698 40126 35700 40178
rect 35644 39508 35700 40126
rect 35868 39844 35924 41244
rect 35980 41234 36036 41244
rect 35868 39778 35924 39788
rect 35980 41076 36036 41086
rect 35644 39442 35700 39452
rect 35868 39172 35924 39182
rect 35644 39060 35700 39070
rect 35532 39058 35700 39060
rect 35532 39006 35646 39058
rect 35698 39006 35700 39058
rect 35532 39004 35700 39006
rect 35644 38994 35700 39004
rect 35756 38948 35812 38958
rect 35756 38854 35812 38892
rect 35868 38668 35924 39116
rect 35756 38612 35924 38668
rect 35644 38050 35700 38062
rect 35644 37998 35646 38050
rect 35698 37998 35700 38050
rect 35644 37266 35700 37998
rect 35644 37214 35646 37266
rect 35698 37214 35700 37266
rect 35644 37156 35700 37214
rect 35644 37090 35700 37100
rect 35532 36484 35588 36494
rect 35532 36390 35588 36428
rect 35420 36204 35700 36260
rect 35644 35138 35700 36204
rect 35644 35086 35646 35138
rect 35698 35086 35700 35138
rect 35644 35074 35700 35086
rect 35420 34916 35476 34926
rect 35308 34914 35476 34916
rect 35308 34862 35422 34914
rect 35474 34862 35476 34914
rect 35308 34860 35476 34862
rect 35420 34850 35476 34860
rect 35532 34804 35588 34814
rect 35420 34468 35476 34478
rect 35196 34356 35252 34366
rect 35084 34354 35252 34356
rect 35084 34302 35198 34354
rect 35250 34302 35252 34354
rect 35084 34300 35252 34302
rect 35196 34290 35252 34300
rect 35308 34244 35364 34254
rect 35308 32788 35364 34188
rect 35420 33346 35476 34412
rect 35532 33460 35588 34748
rect 35532 33394 35588 33404
rect 35644 34244 35700 34254
rect 35420 33294 35422 33346
rect 35474 33294 35476 33346
rect 35420 33282 35476 33294
rect 34972 32732 35140 32788
rect 34860 32510 34862 32562
rect 34914 32510 34916 32562
rect 34860 32498 34916 32510
rect 34860 32228 34916 32238
rect 34748 31890 34804 31902
rect 34748 31838 34750 31890
rect 34802 31838 34804 31890
rect 34636 31780 34692 31790
rect 34636 30548 34692 31724
rect 34748 31444 34804 31838
rect 34748 31378 34804 31388
rect 34636 30482 34692 30492
rect 34860 30324 34916 32172
rect 34972 31892 35028 31902
rect 34972 31798 35028 31836
rect 35084 31220 35140 32732
rect 35308 32722 35364 32732
rect 35084 31154 35140 31164
rect 35196 32676 35252 32686
rect 35196 31778 35252 32620
rect 35308 32452 35364 32462
rect 35308 32358 35364 32396
rect 35644 32116 35700 34188
rect 35644 32050 35700 32060
rect 35420 31890 35476 31902
rect 35420 31838 35422 31890
rect 35474 31838 35476 31890
rect 35196 31726 35198 31778
rect 35250 31726 35252 31778
rect 34860 30258 34916 30268
rect 34972 30994 35028 31006
rect 34972 30942 34974 30994
rect 35026 30942 35028 30994
rect 34524 30158 34526 30210
rect 34578 30158 34580 30210
rect 34524 30146 34580 30158
rect 34748 29652 34804 29662
rect 34748 29558 34804 29596
rect 34860 29426 34916 29438
rect 34860 29374 34862 29426
rect 34914 29374 34916 29426
rect 34412 28590 34414 28642
rect 34466 28590 34468 28642
rect 34412 28532 34468 28590
rect 34412 28466 34468 28476
rect 34524 29314 34580 29326
rect 34524 29262 34526 29314
rect 34578 29262 34580 29314
rect 33852 26450 33908 26460
rect 33964 28420 34020 28430
rect 33628 25618 33684 25630
rect 33628 25566 33630 25618
rect 33682 25566 33684 25618
rect 33628 25396 33684 25566
rect 33740 25508 33796 25518
rect 33740 25414 33796 25452
rect 33628 25330 33684 25340
rect 33740 24724 33796 24734
rect 33404 23538 33460 23548
rect 33516 24612 33572 24622
rect 32956 21534 32958 21586
rect 33010 21534 33012 21586
rect 32732 20972 32900 21028
rect 32620 20962 32676 20972
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32396 20692 32452 20750
rect 32732 20802 32788 20814
rect 32732 20750 32734 20802
rect 32786 20750 32788 20802
rect 32396 20636 32564 20692
rect 32508 20468 32564 20636
rect 32508 20402 32564 20412
rect 32620 20244 32676 20254
rect 32732 20244 32788 20750
rect 32620 20242 32788 20244
rect 32620 20190 32622 20242
rect 32674 20190 32788 20242
rect 32620 20188 32788 20190
rect 32620 20178 32676 20188
rect 32284 20020 32340 20030
rect 32284 15876 32340 19964
rect 32844 19796 32900 20972
rect 32844 19730 32900 19740
rect 32620 19124 32676 19134
rect 32956 19124 33012 21534
rect 33068 23044 33124 23054
rect 33068 19458 33124 22988
rect 33180 22370 33236 23492
rect 33180 22318 33182 22370
rect 33234 22318 33236 22370
rect 33180 22306 33236 22318
rect 33292 23156 33348 23166
rect 33292 22930 33348 23100
rect 33292 22878 33294 22930
rect 33346 22878 33348 22930
rect 33180 21252 33236 21262
rect 33292 21252 33348 22878
rect 33404 23154 33460 23166
rect 33404 23102 33406 23154
rect 33458 23102 33460 23154
rect 33404 22932 33460 23102
rect 33404 22484 33460 22876
rect 33404 22418 33460 22428
rect 33516 21474 33572 24556
rect 33628 24164 33684 24174
rect 33628 24070 33684 24108
rect 33628 22370 33684 22382
rect 33628 22318 33630 22370
rect 33682 22318 33684 22370
rect 33628 22148 33684 22318
rect 33628 22082 33684 22092
rect 33516 21422 33518 21474
rect 33570 21422 33572 21474
rect 33516 21410 33572 21422
rect 33236 21196 33348 21252
rect 33404 21252 33460 21262
rect 33180 21186 33236 21196
rect 33404 21026 33460 21196
rect 33404 20974 33406 21026
rect 33458 20974 33460 21026
rect 33404 20962 33460 20974
rect 33292 20802 33348 20814
rect 33292 20750 33294 20802
rect 33346 20750 33348 20802
rect 33180 20580 33236 20590
rect 33180 20242 33236 20524
rect 33180 20190 33182 20242
rect 33234 20190 33236 20242
rect 33180 20178 33236 20190
rect 33292 20132 33348 20750
rect 33348 20076 33460 20132
rect 33292 20066 33348 20076
rect 33068 19406 33070 19458
rect 33122 19406 33124 19458
rect 33068 19394 33124 19406
rect 33292 19796 33348 19806
rect 32620 19122 33012 19124
rect 32620 19070 32622 19122
rect 32674 19070 33012 19122
rect 32620 19068 33012 19070
rect 33068 19236 33124 19246
rect 32508 18788 32564 18798
rect 32508 18450 32564 18732
rect 32508 18398 32510 18450
rect 32562 18398 32564 18450
rect 32508 18386 32564 18398
rect 32620 17554 32676 19068
rect 32620 17502 32622 17554
rect 32674 17502 32676 17554
rect 32508 16884 32564 16894
rect 32508 16770 32564 16828
rect 32508 16718 32510 16770
rect 32562 16718 32564 16770
rect 32508 16706 32564 16718
rect 32284 15810 32340 15820
rect 32508 16436 32564 16446
rect 32284 15316 32340 15326
rect 32284 15222 32340 15260
rect 32284 13860 32340 13870
rect 32284 13766 32340 13804
rect 32284 11732 32340 11742
rect 32284 10610 32340 11676
rect 32284 10558 32286 10610
rect 32338 10558 32340 10610
rect 32284 10546 32340 10558
rect 32396 9714 32452 9726
rect 32396 9662 32398 9714
rect 32450 9662 32452 9714
rect 32396 9604 32452 9662
rect 32396 9538 32452 9548
rect 32060 8878 32062 8930
rect 32114 8878 32116 8930
rect 31612 8540 32004 8596
rect 31612 8372 31668 8540
rect 31612 8306 31668 8316
rect 31836 8372 31892 8382
rect 31724 8036 31780 8046
rect 31724 7942 31780 7980
rect 31836 7698 31892 8316
rect 31948 8148 32004 8540
rect 31948 8082 32004 8092
rect 32060 7812 32116 8878
rect 32396 9042 32452 9054
rect 32396 8990 32398 9042
rect 32450 8990 32452 9042
rect 32396 8372 32452 8990
rect 32396 8306 32452 8316
rect 32284 8260 32340 8270
rect 32284 8148 32340 8204
rect 32396 8148 32452 8158
rect 32284 8146 32452 8148
rect 32284 8094 32398 8146
rect 32450 8094 32452 8146
rect 32284 8092 32452 8094
rect 32284 7924 32340 8092
rect 32396 8082 32452 8092
rect 32508 7924 32564 16380
rect 32620 16100 32676 17502
rect 32732 18452 32788 18462
rect 32732 16770 32788 18396
rect 33068 18450 33124 19180
rect 33068 18398 33070 18450
rect 33122 18398 33124 18450
rect 33068 18386 33124 18398
rect 33180 18564 33236 18574
rect 32956 18226 33012 18238
rect 32956 18174 32958 18226
rect 33010 18174 33012 18226
rect 32956 17780 33012 18174
rect 33068 18004 33124 18014
rect 33068 17890 33124 17948
rect 33068 17838 33070 17890
rect 33122 17838 33124 17890
rect 33068 17826 33124 17838
rect 32956 17714 33012 17724
rect 32844 16996 32900 17034
rect 32844 16930 32900 16940
rect 32956 16884 33012 16894
rect 33180 16884 33236 18508
rect 33292 18004 33348 19740
rect 33404 19684 33460 20076
rect 33404 19618 33460 19628
rect 33516 18452 33572 18462
rect 33516 18358 33572 18396
rect 33292 17938 33348 17948
rect 32956 16882 33236 16884
rect 32956 16830 32958 16882
rect 33010 16830 33236 16882
rect 32956 16828 33236 16830
rect 33292 16884 33348 16894
rect 32956 16818 33012 16828
rect 33292 16790 33348 16828
rect 32732 16718 32734 16770
rect 32786 16718 32788 16770
rect 32732 16706 32788 16718
rect 33180 16548 33236 16558
rect 33068 16436 33124 16446
rect 32956 16212 33012 16222
rect 32956 16118 33012 16156
rect 32844 16100 32900 16110
rect 32620 16098 32844 16100
rect 32620 16046 32622 16098
rect 32674 16046 32844 16098
rect 32620 16044 32844 16046
rect 32620 16034 32676 16044
rect 32732 15876 32788 15886
rect 32732 15314 32788 15820
rect 32732 15262 32734 15314
rect 32786 15262 32788 15314
rect 32732 14868 32788 15262
rect 32732 14802 32788 14812
rect 32844 14308 32900 16044
rect 32844 14242 32900 14252
rect 32956 15090 33012 15102
rect 32956 15038 32958 15090
rect 33010 15038 33012 15090
rect 32844 14084 32900 14094
rect 32732 13746 32788 13758
rect 32732 13694 32734 13746
rect 32786 13694 32788 13746
rect 32620 13076 32676 13086
rect 32620 12962 32676 13020
rect 32620 12910 32622 12962
rect 32674 12910 32676 12962
rect 32620 12898 32676 12910
rect 32732 12402 32788 13694
rect 32732 12350 32734 12402
rect 32786 12350 32788 12402
rect 32732 12338 32788 12350
rect 32620 11060 32676 11070
rect 32620 8484 32676 11004
rect 32732 9826 32788 9838
rect 32732 9774 32734 9826
rect 32786 9774 32788 9826
rect 32732 8484 32788 9774
rect 32844 9268 32900 14028
rect 32956 13860 33012 15038
rect 32956 13794 33012 13804
rect 33068 13748 33124 16380
rect 33180 15148 33236 16492
rect 33628 15876 33684 15886
rect 33628 15314 33684 15820
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33628 15250 33684 15262
rect 33740 15204 33796 24668
rect 33852 23268 33908 23278
rect 33852 23154 33908 23212
rect 33852 23102 33854 23154
rect 33906 23102 33908 23154
rect 33852 23090 33908 23102
rect 33852 22482 33908 22494
rect 33852 22430 33854 22482
rect 33906 22430 33908 22482
rect 33852 22372 33908 22430
rect 33852 22306 33908 22316
rect 33964 22148 34020 28364
rect 34076 28308 34132 28318
rect 34076 27748 34132 28252
rect 34300 28196 34356 28206
rect 34188 27748 34244 27758
rect 34076 27746 34244 27748
rect 34076 27694 34190 27746
rect 34242 27694 34244 27746
rect 34076 27692 34244 27694
rect 34188 27682 34244 27692
rect 34188 27188 34244 27198
rect 34076 26964 34132 27002
rect 34076 26898 34132 26908
rect 34076 26066 34132 26078
rect 34076 26014 34078 26066
rect 34130 26014 34132 26066
rect 34076 25060 34132 26014
rect 34076 24994 34132 25004
rect 34076 24836 34132 24846
rect 34076 24742 34132 24780
rect 34076 23826 34132 23838
rect 34076 23774 34078 23826
rect 34130 23774 34132 23826
rect 34076 23492 34132 23774
rect 34076 23426 34132 23436
rect 34188 22820 34244 27132
rect 34300 23940 34356 28140
rect 34524 27636 34580 29262
rect 34748 28980 34804 28990
rect 34524 27570 34580 27580
rect 34636 27858 34692 27870
rect 34636 27806 34638 27858
rect 34690 27806 34692 27858
rect 34412 26964 34468 26974
rect 34412 26292 34468 26908
rect 34636 26628 34692 27806
rect 34748 27074 34804 28924
rect 34860 28868 34916 29374
rect 34860 28802 34916 28812
rect 34972 28308 35028 30942
rect 35084 29202 35140 29214
rect 35084 29150 35086 29202
rect 35138 29150 35140 29202
rect 35084 28378 35140 29150
rect 35196 29092 35252 31726
rect 35308 31780 35364 31790
rect 35308 31686 35364 31724
rect 35420 31444 35476 31838
rect 35532 31892 35588 31902
rect 35532 31798 35588 31836
rect 35420 31378 35476 31388
rect 35644 31444 35700 31454
rect 35308 31332 35364 31342
rect 35308 31220 35364 31276
rect 35308 31164 35476 31220
rect 35196 29026 35252 29036
rect 35308 29202 35364 29214
rect 35308 29150 35310 29202
rect 35362 29150 35364 29202
rect 35308 28756 35364 29150
rect 35308 28690 35364 28700
rect 35420 28420 35476 31164
rect 35532 30882 35588 30894
rect 35532 30830 35534 30882
rect 35586 30830 35588 30882
rect 35532 30436 35588 30830
rect 35644 30882 35700 31388
rect 35756 31332 35812 38612
rect 35868 37156 35924 37166
rect 35868 36708 35924 37100
rect 35980 36932 36036 41020
rect 36204 40180 36260 43260
rect 36428 43250 36484 43260
rect 36428 42980 36484 42990
rect 36428 42886 36484 42924
rect 36316 42756 36372 42766
rect 36316 40402 36372 42700
rect 36652 42644 36708 43708
rect 36764 43426 36820 44156
rect 36876 44098 36932 44110
rect 36876 44046 36878 44098
rect 36930 44046 36932 44098
rect 36876 43652 36932 44046
rect 36876 43586 36932 43596
rect 36764 43374 36766 43426
rect 36818 43374 36820 43426
rect 36764 43362 36820 43374
rect 37100 43316 37156 43326
rect 37100 42756 37156 43260
rect 37100 42662 37156 42700
rect 36652 42196 36708 42588
rect 37212 42532 37268 44828
rect 37324 44546 37380 44828
rect 37548 44660 37604 45052
rect 37884 44996 37940 45006
rect 37884 44902 37940 44940
rect 37548 44594 37604 44604
rect 37660 44772 37716 44782
rect 37324 44494 37326 44546
rect 37378 44494 37380 44546
rect 37324 44482 37380 44494
rect 37436 44548 37492 44558
rect 37436 44454 37492 44492
rect 37660 44548 37716 44716
rect 37660 44482 37716 44492
rect 37548 44436 37604 44446
rect 37548 44342 37604 44380
rect 38108 44436 38164 48190
rect 38220 46900 38276 53790
rect 38668 52946 38724 52958
rect 38668 52894 38670 52946
rect 38722 52894 38724 52946
rect 38332 52274 38388 52286
rect 38332 52222 38334 52274
rect 38386 52222 38388 52274
rect 38332 49252 38388 52222
rect 38668 51380 38724 52894
rect 38780 52500 38836 56476
rect 39116 55860 39172 55870
rect 39116 55766 39172 55804
rect 39228 55522 39284 57344
rect 39676 56644 39732 57344
rect 39452 56588 39732 56644
rect 39452 56082 39508 56588
rect 39452 56030 39454 56082
rect 39506 56030 39508 56082
rect 39452 56018 39508 56030
rect 39228 55470 39230 55522
rect 39282 55470 39284 55522
rect 39228 55458 39284 55470
rect 40012 55858 40068 55870
rect 40012 55806 40014 55858
rect 40066 55806 40068 55858
rect 38892 55412 38948 55422
rect 38892 55318 38948 55356
rect 39564 55410 39620 55422
rect 39564 55358 39566 55410
rect 39618 55358 39620 55410
rect 39564 54628 39620 55358
rect 40012 55300 40068 55806
rect 40124 55524 40180 57344
rect 40348 55858 40404 55870
rect 40348 55806 40350 55858
rect 40402 55806 40404 55858
rect 40236 55524 40292 55534
rect 40124 55522 40292 55524
rect 40124 55470 40238 55522
rect 40290 55470 40292 55522
rect 40124 55468 40292 55470
rect 40236 55458 40292 55468
rect 40012 55234 40068 55244
rect 39564 54562 39620 54572
rect 39004 54514 39060 54526
rect 39004 54462 39006 54514
rect 39058 54462 39060 54514
rect 39004 52724 39060 54462
rect 39004 52658 39060 52668
rect 39228 54402 39284 54414
rect 39228 54350 39230 54402
rect 39282 54350 39284 54402
rect 38780 52444 39060 52500
rect 38556 51324 38724 51380
rect 38892 51380 38948 51390
rect 38556 50596 38612 51324
rect 38556 50530 38612 50540
rect 38668 51156 38724 51166
rect 38668 50594 38724 51100
rect 38668 50542 38670 50594
rect 38722 50542 38724 50594
rect 38668 50530 38724 50542
rect 38556 49700 38612 49710
rect 38332 49186 38388 49196
rect 38444 49698 38612 49700
rect 38444 49646 38558 49698
rect 38610 49646 38612 49698
rect 38444 49644 38612 49646
rect 38332 48580 38388 48590
rect 38332 47570 38388 48524
rect 38444 47796 38500 49644
rect 38556 49634 38612 49644
rect 38668 49588 38724 49598
rect 38668 49586 38836 49588
rect 38668 49534 38670 49586
rect 38722 49534 38836 49586
rect 38668 49532 38836 49534
rect 38668 49522 38724 49532
rect 38668 48802 38724 48814
rect 38668 48750 38670 48802
rect 38722 48750 38724 48802
rect 38556 48244 38612 48254
rect 38668 48244 38724 48750
rect 38556 48242 38724 48244
rect 38556 48190 38558 48242
rect 38610 48190 38724 48242
rect 38556 48188 38724 48190
rect 38556 48178 38612 48188
rect 38668 48020 38724 48030
rect 38668 47926 38724 47964
rect 38444 47740 38724 47796
rect 38332 47518 38334 47570
rect 38386 47518 38388 47570
rect 38332 47506 38388 47518
rect 38444 47572 38500 47582
rect 38444 47478 38500 47516
rect 38556 47570 38612 47582
rect 38556 47518 38558 47570
rect 38610 47518 38612 47570
rect 38556 47460 38612 47518
rect 38556 47394 38612 47404
rect 38444 47236 38500 47246
rect 38220 46844 38388 46900
rect 38220 46674 38276 46686
rect 38220 46622 38222 46674
rect 38274 46622 38276 46674
rect 38220 45780 38276 46622
rect 38220 45714 38276 45724
rect 38108 44370 38164 44380
rect 38220 45332 38276 45342
rect 37660 44324 37716 44334
rect 37436 44100 37492 44110
rect 37324 43538 37380 43550
rect 37324 43486 37326 43538
rect 37378 43486 37380 43538
rect 37324 43316 37380 43486
rect 37324 43250 37380 43260
rect 37212 42466 37268 42476
rect 36764 42196 36820 42206
rect 36652 42194 36820 42196
rect 36652 42142 36766 42194
rect 36818 42142 36820 42194
rect 36652 42140 36820 42142
rect 36764 42130 36820 42140
rect 37100 42084 37156 42094
rect 36988 41858 37044 41870
rect 36988 41806 36990 41858
rect 37042 41806 37044 41858
rect 36428 41748 36484 41758
rect 36428 41746 36932 41748
rect 36428 41694 36430 41746
rect 36482 41694 36932 41746
rect 36428 41692 36932 41694
rect 36428 41682 36484 41692
rect 36764 40964 36820 40974
rect 36316 40350 36318 40402
rect 36370 40350 36372 40402
rect 36316 40338 36372 40350
rect 36652 40404 36708 40414
rect 36652 40310 36708 40348
rect 36428 40292 36484 40302
rect 36204 40124 36372 40180
rect 36204 39508 36260 39518
rect 36092 38836 36148 38846
rect 36092 37156 36148 38780
rect 36204 38834 36260 39452
rect 36204 38782 36206 38834
rect 36258 38782 36260 38834
rect 36204 38770 36260 38782
rect 36316 38052 36372 40124
rect 36428 39842 36484 40236
rect 36764 39956 36820 40908
rect 36428 39790 36430 39842
rect 36482 39790 36484 39842
rect 36428 39778 36484 39790
rect 36652 39900 36820 39956
rect 36652 38834 36708 39900
rect 36764 38948 36820 38958
rect 36764 38854 36820 38892
rect 36652 38782 36654 38834
rect 36706 38782 36708 38834
rect 36652 38770 36708 38782
rect 36876 38834 36932 41692
rect 36988 40292 37044 41806
rect 37100 41410 37156 42028
rect 37436 42084 37492 44044
rect 37436 42018 37492 42028
rect 37548 42980 37604 42990
rect 37100 41358 37102 41410
rect 37154 41358 37156 41410
rect 37100 41346 37156 41358
rect 37212 41860 37268 41870
rect 37212 41412 37268 41804
rect 37436 41860 37492 41870
rect 37436 41766 37492 41804
rect 37324 41412 37380 41422
rect 37212 41410 37380 41412
rect 37212 41358 37326 41410
rect 37378 41358 37380 41410
rect 37212 41356 37380 41358
rect 37324 41346 37380 41356
rect 37436 41186 37492 41198
rect 37436 41134 37438 41186
rect 37490 41134 37492 41186
rect 36988 40226 37044 40236
rect 37212 40402 37268 40414
rect 37212 40350 37214 40402
rect 37266 40350 37268 40402
rect 37212 40180 37268 40350
rect 37436 40292 37492 41134
rect 37548 41076 37604 42924
rect 37548 41010 37604 41020
rect 37436 40226 37492 40236
rect 37548 40852 37604 40862
rect 37548 40290 37604 40796
rect 37660 40628 37716 44268
rect 38108 44212 38164 44222
rect 38220 44212 38276 45276
rect 38108 44210 38276 44212
rect 38108 44158 38110 44210
rect 38162 44158 38276 44210
rect 38108 44156 38276 44158
rect 38108 44146 38164 44156
rect 37996 44098 38052 44110
rect 37996 44046 37998 44098
rect 38050 44046 38052 44098
rect 37996 43876 38052 44046
rect 37996 43810 38052 43820
rect 37772 43316 37828 43326
rect 37772 43222 37828 43260
rect 37884 42980 37940 42990
rect 37884 42756 37940 42924
rect 37772 42084 37828 42094
rect 37772 40852 37828 42028
rect 37772 40786 37828 40796
rect 37884 41186 37940 42700
rect 38220 42756 38276 42766
rect 38108 42084 38164 42094
rect 38108 41990 38164 42028
rect 38220 41972 38276 42700
rect 38220 41878 38276 41916
rect 37996 41748 38052 41758
rect 37996 41746 38164 41748
rect 37996 41694 37998 41746
rect 38050 41694 38164 41746
rect 37996 41692 38164 41694
rect 37996 41682 38052 41692
rect 38108 41524 38164 41692
rect 38108 41458 38164 41468
rect 37884 41134 37886 41186
rect 37938 41134 37940 41186
rect 37660 40562 37716 40572
rect 37548 40238 37550 40290
rect 37602 40238 37604 40290
rect 37212 39620 37268 40124
rect 37324 39620 37380 39630
rect 37212 39618 37380 39620
rect 37212 39566 37326 39618
rect 37378 39566 37380 39618
rect 37212 39564 37380 39566
rect 37324 39172 37380 39564
rect 36876 38782 36878 38834
rect 36930 38782 36932 38834
rect 36876 38770 36932 38782
rect 36988 38948 37044 38958
rect 36316 37986 36372 37996
rect 36316 37828 36372 37838
rect 36316 37826 36708 37828
rect 36316 37774 36318 37826
rect 36370 37774 36708 37826
rect 36316 37772 36708 37774
rect 36316 37762 36372 37772
rect 36092 37090 36148 37100
rect 36540 37268 36596 37278
rect 35980 36876 36372 36932
rect 36204 36708 36260 36718
rect 35868 36706 36260 36708
rect 35868 36654 36206 36706
rect 36258 36654 36260 36706
rect 35868 36652 36260 36654
rect 36204 36642 36260 36652
rect 35980 36482 36036 36494
rect 35980 36430 35982 36482
rect 36034 36430 36036 36482
rect 35980 36372 36036 36430
rect 35868 36148 35924 36158
rect 35868 34244 35924 36092
rect 35980 35028 36036 36316
rect 36316 35140 36372 36876
rect 36540 36372 36596 37212
rect 36652 36594 36708 37772
rect 36764 37268 36820 37278
rect 36764 37174 36820 37212
rect 36652 36542 36654 36594
rect 36706 36542 36708 36594
rect 36652 36530 36708 36542
rect 36764 37044 36820 37054
rect 36540 36306 36596 36316
rect 36764 36260 36820 36988
rect 36652 36204 36820 36260
rect 35980 34962 36036 34972
rect 36204 35084 36372 35140
rect 36428 35474 36484 35486
rect 36428 35422 36430 35474
rect 36482 35422 36484 35474
rect 36092 34244 36148 34254
rect 35868 34178 35924 34188
rect 35980 34188 36092 34244
rect 35868 33458 35924 33470
rect 35868 33406 35870 33458
rect 35922 33406 35924 33458
rect 35868 32676 35924 33406
rect 35868 32610 35924 32620
rect 35868 32452 35924 32462
rect 35868 31778 35924 32396
rect 35868 31726 35870 31778
rect 35922 31726 35924 31778
rect 35868 31714 35924 31726
rect 35756 31266 35812 31276
rect 35868 30996 35924 31006
rect 35980 30996 36036 34188
rect 36092 34178 36148 34188
rect 35868 30994 36036 30996
rect 35868 30942 35870 30994
rect 35922 30942 36036 30994
rect 35868 30940 36036 30942
rect 36092 33908 36148 33918
rect 35868 30930 35924 30940
rect 35644 30830 35646 30882
rect 35698 30830 35700 30882
rect 35644 30818 35700 30830
rect 35532 30380 35812 30436
rect 35532 30210 35588 30222
rect 35532 30158 35534 30210
rect 35586 30158 35588 30210
rect 35532 29988 35588 30158
rect 35532 29922 35588 29932
rect 35644 30212 35700 30222
rect 35532 29540 35588 29550
rect 35532 29314 35588 29484
rect 35644 29426 35700 30156
rect 35644 29374 35646 29426
rect 35698 29374 35700 29426
rect 35644 29362 35700 29374
rect 35532 29262 35534 29314
rect 35586 29262 35588 29314
rect 35532 29250 35588 29262
rect 35756 29316 35812 30380
rect 36092 30212 36148 33852
rect 36204 30772 36260 35084
rect 36316 34916 36372 34926
rect 36428 34916 36484 35422
rect 36316 34914 36484 34916
rect 36316 34862 36318 34914
rect 36370 34862 36484 34914
rect 36316 34860 36484 34862
rect 36540 35476 36596 35486
rect 36316 34850 36372 34860
rect 36540 34468 36596 35420
rect 36316 34020 36372 34030
rect 36316 32116 36372 33964
rect 36540 32676 36596 34412
rect 36652 33124 36708 36204
rect 36876 34914 36932 34926
rect 36876 34862 36878 34914
rect 36930 34862 36932 34914
rect 36876 34692 36932 34862
rect 36876 34626 36932 34636
rect 36764 34244 36820 34254
rect 36764 34130 36820 34188
rect 36764 34078 36766 34130
rect 36818 34078 36820 34130
rect 36764 34066 36820 34078
rect 36876 33908 36932 33918
rect 36876 33460 36932 33852
rect 36988 33572 37044 38892
rect 37324 38834 37380 39116
rect 37324 38782 37326 38834
rect 37378 38782 37380 38834
rect 37324 38770 37380 38782
rect 37548 38388 37604 40238
rect 37884 40180 37940 41134
rect 37884 40114 37940 40124
rect 38220 41188 38276 41198
rect 37772 39732 37828 39742
rect 37100 38332 37604 38388
rect 37660 39730 37828 39732
rect 37660 39678 37774 39730
rect 37826 39678 37828 39730
rect 37660 39676 37828 39678
rect 37660 39284 37716 39676
rect 37772 39666 37828 39676
rect 37100 33684 37156 38332
rect 37548 38164 37604 38174
rect 37660 38164 37716 39228
rect 37884 38948 37940 38958
rect 37884 38722 37940 38892
rect 37884 38670 37886 38722
rect 37938 38670 37940 38722
rect 37884 38658 37940 38670
rect 38220 38668 38276 41132
rect 37996 38612 38276 38668
rect 38332 38668 38388 46844
rect 38444 44434 38500 47180
rect 38444 44382 38446 44434
rect 38498 44382 38500 44434
rect 38444 44370 38500 44382
rect 38556 46562 38612 46574
rect 38556 46510 38558 46562
rect 38610 46510 38612 46562
rect 38556 46452 38612 46510
rect 38556 44212 38612 46396
rect 38668 45892 38724 47740
rect 38780 46452 38836 49532
rect 38780 46386 38836 46396
rect 38892 45892 38948 51324
rect 39004 48468 39060 52444
rect 39228 51380 39284 54350
rect 39564 54404 39620 54414
rect 39564 54310 39620 54348
rect 39452 53844 39508 53854
rect 39340 53506 39396 53518
rect 39340 53454 39342 53506
rect 39394 53454 39396 53506
rect 39340 52946 39396 53454
rect 39340 52894 39342 52946
rect 39394 52894 39396 52946
rect 39340 52882 39396 52894
rect 39452 52164 39508 53788
rect 40124 52948 40180 52958
rect 39564 52946 40180 52948
rect 39564 52894 40126 52946
rect 40178 52894 40180 52946
rect 39564 52892 40180 52894
rect 39564 52386 39620 52892
rect 40124 52882 40180 52892
rect 39564 52334 39566 52386
rect 39618 52334 39620 52386
rect 39564 52322 39620 52334
rect 39900 52612 39956 52622
rect 39452 52108 39844 52164
rect 39228 51314 39284 51324
rect 39340 51716 39396 51726
rect 39116 51268 39172 51278
rect 39116 50932 39172 51212
rect 39228 51156 39284 51166
rect 39228 51062 39284 51100
rect 39116 50876 39284 50932
rect 39004 48402 39060 48412
rect 39116 50596 39172 50606
rect 39116 48132 39172 50540
rect 39228 50036 39284 50876
rect 39228 49922 39284 49980
rect 39228 49870 39230 49922
rect 39282 49870 39284 49922
rect 39228 49858 39284 49870
rect 39340 49700 39396 51660
rect 39788 51266 39844 52108
rect 39788 51214 39790 51266
rect 39842 51214 39844 51266
rect 39788 51202 39844 51214
rect 39564 50596 39620 50606
rect 39564 50502 39620 50540
rect 39340 49634 39396 49644
rect 39676 49588 39732 49598
rect 39676 49494 39732 49532
rect 39676 49252 39732 49262
rect 39676 49158 39732 49196
rect 39004 48130 39172 48132
rect 39004 48078 39118 48130
rect 39170 48078 39172 48130
rect 39004 48076 39172 48078
rect 39004 47236 39060 48076
rect 39116 48066 39172 48076
rect 39452 49026 39508 49038
rect 39452 48974 39454 49026
rect 39506 48974 39508 49026
rect 39452 47684 39508 48974
rect 39900 48356 39956 52556
rect 40236 52164 40292 52174
rect 40124 51156 40180 51166
rect 40124 51062 40180 51100
rect 40236 50820 40292 52108
rect 40348 50820 40404 55806
rect 40572 55636 40628 57344
rect 40796 57092 40852 57102
rect 40460 55580 40628 55636
rect 40684 55858 40740 55870
rect 40684 55806 40686 55858
rect 40738 55806 40740 55858
rect 40460 54628 40516 55580
rect 40572 55412 40628 55422
rect 40572 55318 40628 55356
rect 40460 54562 40516 54572
rect 40460 54292 40516 54302
rect 40460 54198 40516 54236
rect 40684 53732 40740 55806
rect 40796 54402 40852 57036
rect 41020 56980 41076 57344
rect 41020 56914 41076 56924
rect 41020 56532 41076 56542
rect 41020 55970 41076 56476
rect 41020 55918 41022 55970
rect 41074 55918 41076 55970
rect 41020 55906 41076 55918
rect 41132 55860 41188 55870
rect 41356 55860 41412 55870
rect 41132 55636 41188 55804
rect 41020 55580 41188 55636
rect 41244 55858 41412 55860
rect 41244 55806 41358 55858
rect 41410 55806 41412 55858
rect 41244 55804 41412 55806
rect 41020 54516 41076 55580
rect 41132 55412 41188 55422
rect 41132 55318 41188 55356
rect 41244 54740 41300 55804
rect 41356 55794 41412 55804
rect 41468 55636 41524 57344
rect 41692 57316 41748 57326
rect 41692 56084 41748 57260
rect 41692 56028 41860 56084
rect 41468 55570 41524 55580
rect 41692 55858 41748 55870
rect 41692 55806 41694 55858
rect 41746 55806 41748 55858
rect 41468 55412 41524 55422
rect 41244 54674 41300 54684
rect 41356 55410 41524 55412
rect 41356 55358 41470 55410
rect 41522 55358 41524 55410
rect 41356 55356 41524 55358
rect 41132 54516 41188 54526
rect 41020 54514 41188 54516
rect 41020 54462 41134 54514
rect 41186 54462 41188 54514
rect 41020 54460 41188 54462
rect 41132 54450 41188 54460
rect 40796 54350 40798 54402
rect 40850 54350 40852 54402
rect 40796 54338 40852 54350
rect 40572 53676 40740 53732
rect 40908 54068 40964 54078
rect 40460 53508 40516 53518
rect 40460 52162 40516 53452
rect 40460 52110 40462 52162
rect 40514 52110 40516 52162
rect 40460 51380 40516 52110
rect 40460 51314 40516 51324
rect 40348 50764 40516 50820
rect 40236 50754 40292 50764
rect 40348 50596 40404 50606
rect 40348 50502 40404 50540
rect 40460 49588 40516 50764
rect 40460 49522 40516 49532
rect 40572 49252 40628 53676
rect 40684 53506 40740 53518
rect 40684 53454 40686 53506
rect 40738 53454 40740 53506
rect 40684 52052 40740 53454
rect 40908 52836 40964 54012
rect 41020 53508 41076 53518
rect 41020 53506 41188 53508
rect 41020 53454 41022 53506
rect 41074 53454 41188 53506
rect 41020 53452 41188 53454
rect 41020 53442 41076 53452
rect 41132 53396 41188 53452
rect 41020 52836 41076 52846
rect 40908 52834 41076 52836
rect 40908 52782 41022 52834
rect 41074 52782 41076 52834
rect 40908 52780 41076 52782
rect 41020 52770 41076 52780
rect 40908 52276 40964 52286
rect 40908 52182 40964 52220
rect 41132 52052 41188 53340
rect 41356 53060 41412 55356
rect 41468 55346 41524 55356
rect 41580 54852 41636 54862
rect 41244 53004 41412 53060
rect 41468 54290 41524 54302
rect 41468 54238 41470 54290
rect 41522 54238 41524 54290
rect 41244 52276 41300 53004
rect 41244 52210 41300 52220
rect 41356 52722 41412 52734
rect 41356 52670 41358 52722
rect 41410 52670 41412 52722
rect 41244 52052 41300 52062
rect 41132 51996 41244 52052
rect 40684 51986 40740 51996
rect 41244 51986 41300 51996
rect 40684 51378 40740 51390
rect 40684 51326 40686 51378
rect 40738 51326 40740 51378
rect 40684 51156 40740 51326
rect 41132 51268 41188 51278
rect 41132 51174 41188 51212
rect 40684 51090 40740 51100
rect 41244 51156 41300 51166
rect 40572 49186 40628 49196
rect 40796 49586 40852 49598
rect 40796 49534 40798 49586
rect 40850 49534 40852 49586
rect 40348 49028 40404 49038
rect 40348 48934 40404 48972
rect 39900 48290 39956 48300
rect 40460 48692 40516 48702
rect 39788 48242 39844 48254
rect 39788 48190 39790 48242
rect 39842 48190 39844 48242
rect 39452 47618 39508 47628
rect 39676 48132 39732 48142
rect 39004 47170 39060 47180
rect 39116 47458 39172 47470
rect 39116 47406 39118 47458
rect 39170 47406 39172 47458
rect 39116 46340 39172 47406
rect 39452 47458 39508 47470
rect 39452 47406 39454 47458
rect 39506 47406 39508 47458
rect 39004 46284 39172 46340
rect 39228 47346 39284 47358
rect 39228 47294 39230 47346
rect 39282 47294 39284 47346
rect 39004 46116 39060 46284
rect 39004 46050 39060 46060
rect 39116 46116 39172 46126
rect 39228 46116 39284 47294
rect 39116 46114 39284 46116
rect 39116 46062 39118 46114
rect 39170 46062 39284 46114
rect 39116 46060 39284 46062
rect 39340 46452 39396 46462
rect 39116 46050 39172 46060
rect 39228 45892 39284 45902
rect 38668 45836 38836 45892
rect 38892 45890 39284 45892
rect 38892 45838 39230 45890
rect 39282 45838 39284 45890
rect 38892 45836 39284 45838
rect 38780 45780 38836 45836
rect 39228 45826 39284 45836
rect 39340 45890 39396 46396
rect 39340 45838 39342 45890
rect 39394 45838 39396 45890
rect 38780 45724 39172 45780
rect 38668 45666 38724 45678
rect 38668 45614 38670 45666
rect 38722 45614 38724 45666
rect 38668 44772 38724 45614
rect 38668 44706 38724 44716
rect 38780 45332 38836 45342
rect 38780 44546 38836 45276
rect 39116 45330 39172 45724
rect 39340 45444 39396 45838
rect 39340 45378 39396 45388
rect 39116 45278 39118 45330
rect 39170 45278 39172 45330
rect 39116 45266 39172 45278
rect 38780 44494 38782 44546
rect 38834 44494 38836 44546
rect 38780 44482 38836 44494
rect 38892 45220 38948 45230
rect 38668 44436 38724 44446
rect 38668 44342 38724 44380
rect 38892 44322 38948 45164
rect 39452 45108 39508 47406
rect 39564 47460 39620 47470
rect 39564 45892 39620 47404
rect 39564 45826 39620 45836
rect 39676 45556 39732 48076
rect 39788 46898 39844 48190
rect 39788 46846 39790 46898
rect 39842 46846 39844 46898
rect 39788 46834 39844 46846
rect 40124 47684 40180 47694
rect 39788 45892 39844 45902
rect 39788 45798 39844 45836
rect 39676 45490 39732 45500
rect 39900 45332 39956 45342
rect 39340 45052 39508 45108
rect 39788 45108 39844 45118
rect 38892 44270 38894 44322
rect 38946 44270 38948 44322
rect 38892 44258 38948 44270
rect 39116 44884 39172 44894
rect 38444 44156 38612 44212
rect 39116 44210 39172 44828
rect 39116 44158 39118 44210
rect 39170 44158 39172 44210
rect 38444 41410 38500 44156
rect 39004 43876 39060 43886
rect 38892 43316 38948 43326
rect 38892 43222 38948 43260
rect 38556 43204 38612 43214
rect 38780 43204 38836 43214
rect 38612 43148 38780 43204
rect 38556 43138 38612 43148
rect 38780 43138 38836 43148
rect 38668 42756 38724 42766
rect 38668 42308 38724 42700
rect 38668 42242 38724 42252
rect 38556 41972 38612 41982
rect 38556 41878 38612 41916
rect 38444 41358 38446 41410
rect 38498 41358 38500 41410
rect 38444 41076 38500 41358
rect 38444 40068 38500 41020
rect 38780 41748 38836 41758
rect 38780 40740 38836 41692
rect 38444 40002 38500 40012
rect 38668 40684 38836 40740
rect 38668 39732 38724 40684
rect 38780 40404 38836 40414
rect 38780 40310 38836 40348
rect 39004 40180 39060 43820
rect 39116 42978 39172 44158
rect 39340 44322 39396 45052
rect 39676 44996 39732 45006
rect 39340 44270 39342 44322
rect 39394 44270 39396 44322
rect 39228 44100 39284 44110
rect 39228 43204 39284 44044
rect 39340 43876 39396 44270
rect 39340 43810 39396 43820
rect 39452 44994 39732 44996
rect 39452 44942 39678 44994
rect 39730 44942 39732 44994
rect 39452 44940 39732 44942
rect 39340 43428 39396 43438
rect 39340 43334 39396 43372
rect 39228 43148 39396 43204
rect 39116 42926 39118 42978
rect 39170 42926 39172 42978
rect 39116 42914 39172 42926
rect 39228 42980 39284 42990
rect 39228 42082 39284 42924
rect 39228 42030 39230 42082
rect 39282 42030 39284 42082
rect 39228 42018 39284 42030
rect 39340 41860 39396 43148
rect 39004 40114 39060 40124
rect 39116 41804 39396 41860
rect 39452 42754 39508 44940
rect 39676 44930 39732 44940
rect 39788 44100 39844 45052
rect 39900 44994 39956 45276
rect 40012 45220 40068 45230
rect 40012 45126 40068 45164
rect 40124 45108 40180 47628
rect 40236 47460 40292 47470
rect 40236 47366 40292 47404
rect 40348 47348 40404 47358
rect 40348 47254 40404 47292
rect 40460 47068 40516 48636
rect 40796 48242 40852 49534
rect 40908 49476 40964 49486
rect 40908 49250 40964 49420
rect 40908 49198 40910 49250
rect 40962 49198 40964 49250
rect 40908 49186 40964 49198
rect 40796 48190 40798 48242
rect 40850 48190 40852 48242
rect 40796 48178 40852 48190
rect 40908 48916 40964 48926
rect 40796 47460 40852 47470
rect 40796 47366 40852 47404
rect 40124 45042 40180 45052
rect 40236 47012 40516 47068
rect 39900 44942 39902 44994
rect 39954 44942 39956 44994
rect 39900 44930 39956 44942
rect 40012 44884 40068 44894
rect 39676 43876 39732 43886
rect 39676 43650 39732 43820
rect 39676 43598 39678 43650
rect 39730 43598 39732 43650
rect 39676 43586 39732 43598
rect 39676 43426 39732 43438
rect 39676 43374 39678 43426
rect 39730 43374 39732 43426
rect 39564 43314 39620 43326
rect 39564 43262 39566 43314
rect 39618 43262 39620 43314
rect 39564 43092 39620 43262
rect 39564 43026 39620 43036
rect 39676 42868 39732 43374
rect 39788 43426 39844 44044
rect 39788 43374 39790 43426
rect 39842 43374 39844 43426
rect 39788 43362 39844 43374
rect 39900 44436 39956 44446
rect 39676 42802 39732 42812
rect 39788 42980 39844 42990
rect 39452 42702 39454 42754
rect 39506 42702 39508 42754
rect 39116 39956 39172 41804
rect 39452 40852 39508 42702
rect 39676 42644 39732 42654
rect 39788 42644 39844 42924
rect 39676 42642 39844 42644
rect 39676 42590 39678 42642
rect 39730 42590 39844 42642
rect 39676 42588 39844 42590
rect 39676 42420 39732 42588
rect 39676 42354 39732 42364
rect 39564 42308 39620 42318
rect 39564 41188 39620 42252
rect 39788 41972 39844 41982
rect 39676 41748 39732 41786
rect 39676 41682 39732 41692
rect 39564 41132 39732 41188
rect 39564 40964 39620 40974
rect 39564 40870 39620 40908
rect 39452 40786 39508 40796
rect 39564 40404 39620 40414
rect 39564 40310 39620 40348
rect 38668 39666 38724 39676
rect 38892 39900 39172 39956
rect 39228 40290 39284 40302
rect 39228 40238 39230 40290
rect 39282 40238 39284 40290
rect 39228 40068 39284 40238
rect 38556 39284 38612 39294
rect 38444 38948 38500 38958
rect 38556 38948 38612 39228
rect 38500 38892 38612 38948
rect 38444 38882 38500 38892
rect 38444 38724 38500 38734
rect 38332 38612 38500 38668
rect 37548 38162 37716 38164
rect 37548 38110 37550 38162
rect 37602 38110 37716 38162
rect 37548 38108 37716 38110
rect 37884 38164 37940 38174
rect 37548 38098 37604 38108
rect 37884 38050 37940 38108
rect 37884 37998 37886 38050
rect 37938 37998 37940 38050
rect 37884 37986 37940 37998
rect 37548 37380 37604 37390
rect 37212 37268 37268 37278
rect 37212 37154 37268 37212
rect 37212 37102 37214 37154
rect 37266 37102 37268 37154
rect 37212 37090 37268 37102
rect 37436 36484 37492 36494
rect 37436 36390 37492 36428
rect 37548 35586 37604 37324
rect 37548 35534 37550 35586
rect 37602 35534 37604 35586
rect 37548 35476 37604 35534
rect 37548 35410 37604 35420
rect 37660 37268 37716 37278
rect 37324 34468 37380 34478
rect 37324 34242 37380 34412
rect 37324 34190 37326 34242
rect 37378 34190 37380 34242
rect 37324 34178 37380 34190
rect 37436 34020 37492 34030
rect 37436 33926 37492 33964
rect 37212 33908 37268 33918
rect 37212 33814 37268 33852
rect 37324 33684 37380 33694
rect 37100 33628 37268 33684
rect 36988 33516 37156 33572
rect 36876 33404 37044 33460
rect 36988 33346 37044 33404
rect 36988 33294 36990 33346
rect 37042 33294 37044 33346
rect 36988 33282 37044 33294
rect 36652 33058 36708 33068
rect 37100 32788 37156 33516
rect 36988 32732 37156 32788
rect 36652 32676 36708 32686
rect 36540 32620 36652 32676
rect 36652 32610 36708 32620
rect 36876 32676 36932 32686
rect 36764 32452 36820 32462
rect 36428 32338 36484 32350
rect 36428 32286 36430 32338
rect 36482 32286 36484 32338
rect 36428 32228 36484 32286
rect 36764 32228 36820 32396
rect 36428 32172 36820 32228
rect 36316 32060 36484 32116
rect 36316 31668 36372 31678
rect 36316 31574 36372 31612
rect 36428 31444 36484 32060
rect 36764 31778 36820 32172
rect 36764 31726 36766 31778
rect 36818 31726 36820 31778
rect 36764 31714 36820 31726
rect 36204 30706 36260 30716
rect 36316 31388 36484 31444
rect 36092 30146 36148 30156
rect 36316 30212 36372 31388
rect 36540 31108 36596 31118
rect 36876 31108 36932 32620
rect 36540 31106 36932 31108
rect 36540 31054 36542 31106
rect 36594 31054 36932 31106
rect 36540 31052 36932 31054
rect 36316 30146 36372 30156
rect 36428 30324 36484 30334
rect 36204 30098 36260 30110
rect 36204 30046 36206 30098
rect 36258 30046 36260 30098
rect 36204 29540 36260 30046
rect 36428 29650 36484 30268
rect 36428 29598 36430 29650
rect 36482 29598 36484 29650
rect 36428 29586 36484 29598
rect 36540 29652 36596 31052
rect 36988 30996 37044 32732
rect 36876 30940 37044 30996
rect 37100 31778 37156 31790
rect 37100 31726 37102 31778
rect 37154 31726 37156 31778
rect 37100 30996 37156 31726
rect 36652 30884 36708 30894
rect 36652 30436 36708 30828
rect 36876 30548 36932 30940
rect 37100 30930 37156 30940
rect 36988 30772 37044 30782
rect 37212 30772 37268 33628
rect 37324 32116 37380 33628
rect 37660 33460 37716 37212
rect 37884 36372 37940 36382
rect 37884 35700 37940 36316
rect 37996 36148 38052 38612
rect 38332 37268 38388 38612
rect 38108 37212 38388 37268
rect 38108 36260 38164 37212
rect 38332 37042 38388 37054
rect 38332 36990 38334 37042
rect 38386 36990 38388 37042
rect 38220 36596 38276 36606
rect 38220 36482 38276 36540
rect 38220 36430 38222 36482
rect 38274 36430 38276 36482
rect 38220 36418 38276 36430
rect 38108 36204 38276 36260
rect 37996 36082 38052 36092
rect 37996 35700 38052 35710
rect 37884 35698 38052 35700
rect 37884 35646 37998 35698
rect 38050 35646 38052 35698
rect 37884 35644 38052 35646
rect 37884 35308 37940 35644
rect 37996 35634 38052 35644
rect 37884 35252 38052 35308
rect 37772 34914 37828 34926
rect 37772 34862 37774 34914
rect 37826 34862 37828 34914
rect 37772 34244 37828 34862
rect 37772 34178 37828 34188
rect 37884 33908 37940 33918
rect 37324 32050 37380 32060
rect 37436 32564 37492 32574
rect 37324 31890 37380 31902
rect 37324 31838 37326 31890
rect 37378 31838 37380 31890
rect 37324 30996 37380 31838
rect 37436 31220 37492 32508
rect 37548 32340 37604 32350
rect 37548 32246 37604 32284
rect 37660 32116 37716 33404
rect 37436 31154 37492 31164
rect 37548 32060 37716 32116
rect 37772 33684 37828 33694
rect 37324 30930 37380 30940
rect 37212 30716 37492 30772
rect 36988 30678 37044 30716
rect 36876 30492 37044 30548
rect 36652 30434 36932 30436
rect 36652 30382 36654 30434
rect 36706 30382 36932 30434
rect 36652 30380 36932 30382
rect 36652 30370 36708 30380
rect 36540 29586 36596 29596
rect 36204 29474 36260 29484
rect 36316 29316 36372 29326
rect 35756 29314 36484 29316
rect 35756 29262 36318 29314
rect 36370 29262 36484 29314
rect 35756 29260 36484 29262
rect 36316 29250 36372 29260
rect 35868 28868 35924 28878
rect 35532 28644 35588 28654
rect 35532 28550 35588 28588
rect 35084 28322 35252 28378
rect 35420 28354 35476 28364
rect 35756 28532 35812 28542
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 26964 34804 27022
rect 34748 26898 34804 26908
rect 34860 28252 35028 28308
rect 34860 26852 34916 28252
rect 35196 28084 35252 28322
rect 35196 28018 35252 28028
rect 35196 27860 35252 27870
rect 35196 27766 35252 27804
rect 35756 27858 35812 28476
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35756 27794 35812 27806
rect 35420 27746 35476 27758
rect 35420 27694 35422 27746
rect 35474 27694 35476 27746
rect 35420 27636 35476 27694
rect 35420 27570 35476 27580
rect 35644 27634 35700 27646
rect 35644 27582 35646 27634
rect 35698 27582 35700 27634
rect 35532 27412 35588 27422
rect 35196 27188 35252 27198
rect 35196 27094 35252 27132
rect 35532 26852 35588 27356
rect 35644 27300 35700 27582
rect 35868 27524 35924 28812
rect 36092 28754 36148 28766
rect 36092 28702 36094 28754
rect 36146 28702 36148 28754
rect 35868 27458 35924 27468
rect 35980 28642 36036 28654
rect 35980 28590 35982 28642
rect 36034 28590 36036 28642
rect 35644 27244 35924 27300
rect 35756 26964 35812 26974
rect 35644 26852 35700 26862
rect 35532 26796 35644 26852
rect 34860 26786 34916 26796
rect 34636 26572 34916 26628
rect 34412 25506 34468 26236
rect 34412 25454 34414 25506
rect 34466 25454 34468 25506
rect 34412 25442 34468 25454
rect 34524 26290 34580 26302
rect 34524 26238 34526 26290
rect 34578 26238 34580 26290
rect 34524 25284 34580 26238
rect 34860 25844 34916 26572
rect 35420 26516 35476 26526
rect 35308 26292 35364 26302
rect 34524 25218 34580 25228
rect 34636 25788 34916 25844
rect 34972 26178 35028 26190
rect 34972 26126 34974 26178
rect 35026 26126 35028 26178
rect 34636 25060 34692 25788
rect 34860 25620 34916 25658
rect 34860 25554 34916 25564
rect 34524 25004 34692 25060
rect 34860 25396 34916 25406
rect 34412 24612 34468 24622
rect 34412 24518 34468 24556
rect 34300 23874 34356 23884
rect 34412 24388 34468 24398
rect 34300 23042 34356 23054
rect 34300 22990 34302 23042
rect 34354 22990 34356 23042
rect 34300 22932 34356 22990
rect 34300 22866 34356 22876
rect 33964 22082 34020 22092
rect 34076 22764 34244 22820
rect 33964 21812 34020 21822
rect 33852 20802 33908 20814
rect 33852 20750 33854 20802
rect 33906 20750 33908 20802
rect 33852 20580 33908 20750
rect 33852 20514 33908 20524
rect 33964 18450 34020 21756
rect 33964 18398 33966 18450
rect 34018 18398 34020 18450
rect 33964 18386 34020 18398
rect 33852 17108 33908 17118
rect 33852 16884 33908 17052
rect 34076 17108 34132 22764
rect 34412 22708 34468 24332
rect 34188 22652 34468 22708
rect 34524 23268 34580 25004
rect 34748 24724 34804 24734
rect 34188 19236 34244 22652
rect 34524 22596 34580 23212
rect 34636 23604 34692 23614
rect 34636 22820 34692 23548
rect 34636 22754 34692 22764
rect 34748 22596 34804 24668
rect 34860 24050 34916 25340
rect 34972 25060 35028 26126
rect 35084 26066 35140 26078
rect 35084 26014 35086 26066
rect 35138 26014 35140 26066
rect 35084 25508 35140 26014
rect 35196 26068 35252 26078
rect 35196 25974 35252 26012
rect 35308 26066 35364 26236
rect 35308 26014 35310 26066
rect 35362 26014 35364 26066
rect 35084 25442 35140 25452
rect 35196 25844 35252 25854
rect 35196 25284 35252 25788
rect 35308 25732 35364 26014
rect 35308 25666 35364 25676
rect 35420 25620 35476 26460
rect 35644 26402 35700 26796
rect 35756 26514 35812 26908
rect 35756 26462 35758 26514
rect 35810 26462 35812 26514
rect 35756 26450 35812 26462
rect 35644 26350 35646 26402
rect 35698 26350 35700 26402
rect 35644 26338 35700 26350
rect 35420 25554 35476 25564
rect 35868 25284 35924 27244
rect 35980 26404 36036 28590
rect 36092 26628 36148 28702
rect 36316 28642 36372 28654
rect 36316 28590 36318 28642
rect 36370 28590 36372 28642
rect 36316 28308 36372 28590
rect 36316 28242 36372 28252
rect 36428 27748 36484 29260
rect 36764 29314 36820 29326
rect 36764 29262 36766 29314
rect 36818 29262 36820 29314
rect 36764 29204 36820 29262
rect 36764 29138 36820 29148
rect 36652 28980 36708 28990
rect 36652 28642 36708 28924
rect 36876 28980 36932 30380
rect 36876 28914 36932 28924
rect 36652 28590 36654 28642
rect 36706 28590 36708 28642
rect 36092 26562 36148 26572
rect 36204 27692 36484 27748
rect 36540 27860 36596 27870
rect 36652 27860 36708 28590
rect 36988 28532 37044 30492
rect 37212 29988 37268 29998
rect 37212 29426 37268 29932
rect 37212 29374 37214 29426
rect 37266 29374 37268 29426
rect 37212 29362 37268 29374
rect 37324 29652 37380 29662
rect 37212 28756 37268 28766
rect 37212 28662 37268 28700
rect 36988 28476 37268 28532
rect 36540 27858 36708 27860
rect 36540 27806 36542 27858
rect 36594 27806 36708 27858
rect 36540 27804 36708 27806
rect 36764 28308 36820 28318
rect 35980 26348 36148 26404
rect 34972 24994 35028 25004
rect 35084 25228 35252 25284
rect 35308 25228 35924 25284
rect 35980 26180 36036 26190
rect 35980 25282 36036 26124
rect 36092 25844 36148 26348
rect 36092 25778 36148 25788
rect 35980 25230 35982 25282
rect 36034 25230 36036 25282
rect 34860 23998 34862 24050
rect 34914 23998 34916 24050
rect 34860 23986 34916 23998
rect 35084 23938 35140 25228
rect 35084 23886 35086 23938
rect 35138 23886 35140 23938
rect 35084 23874 35140 23886
rect 35196 24724 35252 24734
rect 35196 23154 35252 24668
rect 35196 23102 35198 23154
rect 35250 23102 35252 23154
rect 35196 23090 35252 23102
rect 35308 23156 35364 25228
rect 35980 25060 36036 25230
rect 35308 23090 35364 23100
rect 35420 25004 36036 25060
rect 35420 23044 35476 25004
rect 36204 24948 36260 27692
rect 36540 27412 36596 27804
rect 36540 27346 36596 27356
rect 36428 26852 36484 26862
rect 36316 26850 36484 26852
rect 36316 26798 36430 26850
rect 36482 26798 36484 26850
rect 36316 26796 36484 26798
rect 36316 26066 36372 26796
rect 36428 26786 36484 26796
rect 36540 26292 36596 26302
rect 36540 26178 36596 26236
rect 36540 26126 36542 26178
rect 36594 26126 36596 26178
rect 36540 26114 36596 26126
rect 36652 26180 36708 26190
rect 36652 26086 36708 26124
rect 36764 26178 36820 28252
rect 36988 28308 37044 28318
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 36764 26114 36820 26126
rect 36876 28084 36932 28094
rect 36316 26014 36318 26066
rect 36370 26014 36372 26066
rect 36316 25844 36372 26014
rect 36316 25778 36372 25788
rect 36428 26066 36484 26078
rect 36428 26014 36430 26066
rect 36482 26014 36484 26066
rect 36428 25620 36484 26014
rect 36540 25732 36596 25770
rect 36540 25666 36596 25676
rect 35532 24892 36260 24948
rect 36316 25564 36484 25620
rect 36764 25620 36820 25630
rect 35532 23268 35588 24892
rect 36316 24724 36372 25564
rect 36540 25508 36596 25518
rect 36428 25396 36484 25406
rect 36428 25302 36484 25340
rect 36540 24836 36596 25452
rect 36540 24742 36596 24780
rect 36764 24836 36820 25564
rect 36764 24770 36820 24780
rect 36316 24658 36372 24668
rect 35644 24500 35700 24510
rect 35644 24498 36372 24500
rect 35644 24446 35646 24498
rect 35698 24446 36372 24498
rect 35644 24444 36372 24446
rect 35644 24434 35700 24444
rect 36204 24276 36260 24286
rect 36316 24276 36372 24444
rect 36316 24220 36820 24276
rect 35644 24052 35700 24062
rect 35644 23938 35700 23996
rect 35644 23886 35646 23938
rect 35698 23886 35700 23938
rect 35644 23874 35700 23886
rect 35980 23716 36036 23726
rect 35756 23714 36036 23716
rect 35756 23662 35982 23714
rect 36034 23662 36036 23714
rect 35756 23660 36036 23662
rect 35644 23268 35700 23278
rect 35532 23266 35700 23268
rect 35532 23214 35646 23266
rect 35698 23214 35700 23266
rect 35532 23212 35700 23214
rect 35644 23202 35700 23212
rect 35756 23154 35812 23660
rect 35980 23650 36036 23660
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 35756 23090 35812 23102
rect 35532 23044 35588 23054
rect 35420 23042 35588 23044
rect 35420 22990 35534 23042
rect 35586 22990 35588 23042
rect 35420 22988 35588 22990
rect 35532 22978 35588 22988
rect 35308 22932 35364 22942
rect 35196 22820 35252 22830
rect 34524 22540 34692 22596
rect 34748 22540 35140 22596
rect 34524 22370 34580 22382
rect 34524 22318 34526 22370
rect 34578 22318 34580 22370
rect 34524 21812 34580 22318
rect 34636 22036 34692 22540
rect 34860 22372 34916 22382
rect 34636 21980 34804 22036
rect 34636 21812 34692 21822
rect 34524 21810 34692 21812
rect 34524 21758 34638 21810
rect 34690 21758 34692 21810
rect 34524 21756 34692 21758
rect 34636 21746 34692 21756
rect 34412 20804 34468 20814
rect 34412 20710 34468 20748
rect 34300 20356 34356 20366
rect 34300 19796 34356 20300
rect 34748 20132 34804 21980
rect 34860 20804 34916 22316
rect 34860 20738 34916 20748
rect 34748 20130 35028 20132
rect 34748 20078 34750 20130
rect 34802 20078 35028 20130
rect 34748 20076 35028 20078
rect 34748 20066 34804 20076
rect 34300 19702 34356 19740
rect 34972 19908 35028 20076
rect 34188 19170 34244 19180
rect 34860 19122 34916 19134
rect 34860 19070 34862 19122
rect 34914 19070 34916 19122
rect 34188 19010 34244 19022
rect 34188 18958 34190 19010
rect 34242 18958 34244 19010
rect 34188 18788 34244 18958
rect 34860 19012 34916 19070
rect 34860 18946 34916 18956
rect 34188 18722 34244 18732
rect 34860 18788 34916 18798
rect 34300 18564 34356 18574
rect 34300 18470 34356 18508
rect 34412 18452 34468 18462
rect 34636 18452 34692 18462
rect 34412 18358 34468 18396
rect 34524 18450 34692 18452
rect 34524 18398 34638 18450
rect 34690 18398 34692 18450
rect 34524 18396 34692 18398
rect 34524 18116 34580 18396
rect 34636 18386 34692 18396
rect 34860 18338 34916 18732
rect 34860 18286 34862 18338
rect 34914 18286 34916 18338
rect 34860 18274 34916 18286
rect 34972 18228 35028 19852
rect 35084 18450 35140 22540
rect 35196 19346 35252 22764
rect 35308 20468 35364 22876
rect 35980 22372 36036 22382
rect 35980 22370 36148 22372
rect 35980 22318 35982 22370
rect 36034 22318 36148 22370
rect 35980 22316 36148 22318
rect 35980 22306 36036 22316
rect 35420 21924 35476 21934
rect 35420 20802 35476 21868
rect 35420 20750 35422 20802
rect 35474 20750 35476 20802
rect 35420 20738 35476 20750
rect 35532 21812 35588 21822
rect 35308 20132 35364 20412
rect 35308 20066 35364 20076
rect 35532 19796 35588 21756
rect 35532 19730 35588 19740
rect 35980 20804 36036 20814
rect 35196 19294 35198 19346
rect 35250 19294 35252 19346
rect 35196 19282 35252 19294
rect 35308 19348 35364 19358
rect 35084 18398 35086 18450
rect 35138 18398 35140 18450
rect 35084 18386 35140 18398
rect 34972 18172 35252 18228
rect 34188 18060 34580 18116
rect 34188 17892 34244 18060
rect 35196 18004 35252 18172
rect 34524 17948 35028 18004
rect 34524 17892 34580 17948
rect 34188 17826 34244 17836
rect 34300 17836 34580 17892
rect 34972 17890 35028 17948
rect 35196 17938 35252 17948
rect 34972 17838 34974 17890
rect 35026 17838 35028 17890
rect 34076 17042 34132 17052
rect 34188 17444 34244 17454
rect 34300 17444 34356 17836
rect 34972 17826 35028 17838
rect 35084 17892 35140 17902
rect 35084 17798 35140 17836
rect 34636 17780 34692 17790
rect 34524 17666 34580 17678
rect 34524 17614 34526 17666
rect 34578 17614 34580 17666
rect 34188 17442 34356 17444
rect 34188 17390 34190 17442
rect 34242 17390 34356 17442
rect 34188 17388 34356 17390
rect 34412 17556 34468 17566
rect 34188 16884 34244 17388
rect 33852 16882 34020 16884
rect 33852 16830 33854 16882
rect 33906 16830 34020 16882
rect 33852 16828 34020 16830
rect 33852 16818 33908 16828
rect 33180 15092 33348 15148
rect 33740 15138 33796 15148
rect 33852 16212 33908 16222
rect 33292 14084 33348 15092
rect 33852 14308 33908 16156
rect 33964 14532 34020 16828
rect 34188 16818 34244 16828
rect 34300 16660 34356 16670
rect 34300 16212 34356 16604
rect 34300 16146 34356 16156
rect 34188 15876 34244 15886
rect 34188 15782 34244 15820
rect 34188 15316 34244 15326
rect 34412 15316 34468 17500
rect 34524 16996 34580 17614
rect 34636 17668 34692 17724
rect 35196 17668 35252 17678
rect 34636 17666 35252 17668
rect 34636 17614 35198 17666
rect 35250 17614 35252 17666
rect 34636 17612 35252 17614
rect 35196 17602 35252 17612
rect 34524 16930 34580 16940
rect 34972 16996 35028 17006
rect 34972 16098 35028 16940
rect 34972 16046 34974 16098
rect 35026 16046 35028 16098
rect 34972 16034 35028 16046
rect 34188 15314 34468 15316
rect 34188 15262 34190 15314
rect 34242 15262 34468 15314
rect 34188 15260 34468 15262
rect 34972 15876 35028 15886
rect 34972 15316 35028 15820
rect 34972 15314 35252 15316
rect 34972 15262 34974 15314
rect 35026 15262 35252 15314
rect 34972 15260 35252 15262
rect 34188 15250 34244 15260
rect 34972 15250 35028 15260
rect 33964 14466 34020 14476
rect 34748 15204 34804 15214
rect 33852 14242 33908 14252
rect 33292 14018 33348 14028
rect 33068 13654 33124 13692
rect 33180 13860 33236 13870
rect 33068 13074 33124 13086
rect 33068 13022 33070 13074
rect 33122 13022 33124 13074
rect 33068 12964 33124 13022
rect 33068 12898 33124 12908
rect 33068 12740 33124 12750
rect 32956 12180 33012 12190
rect 32956 10610 33012 12124
rect 32956 10558 32958 10610
rect 33010 10558 33012 10610
rect 32956 10546 33012 10558
rect 33068 9828 33124 12684
rect 33180 10164 33236 13804
rect 33292 13748 33348 13758
rect 33292 13634 33348 13692
rect 33964 13748 34020 13758
rect 33964 13746 34244 13748
rect 33964 13694 33966 13746
rect 34018 13694 34244 13746
rect 33964 13692 34244 13694
rect 33964 13682 34020 13692
rect 33292 13582 33294 13634
rect 33346 13582 33348 13634
rect 33292 13570 33348 13582
rect 34188 13186 34244 13692
rect 34412 13746 34468 13758
rect 34412 13694 34414 13746
rect 34466 13694 34468 13746
rect 34412 13636 34468 13694
rect 34412 13570 34468 13580
rect 34636 13636 34692 13646
rect 34188 13134 34190 13186
rect 34242 13134 34244 13186
rect 34188 13122 34244 13134
rect 33852 12292 33908 12302
rect 33180 10098 33236 10108
rect 33292 10388 33348 10398
rect 33180 9828 33236 9838
rect 33068 9826 33236 9828
rect 33068 9774 33182 9826
rect 33234 9774 33236 9826
rect 33068 9772 33236 9774
rect 33068 9492 33124 9772
rect 33180 9762 33236 9772
rect 33068 9426 33124 9436
rect 33292 9492 33348 10332
rect 33516 10388 33572 10398
rect 33516 10294 33572 10332
rect 33292 9426 33348 9436
rect 33404 9938 33460 9950
rect 33404 9886 33406 9938
rect 33458 9886 33460 9938
rect 32844 9212 33348 9268
rect 32844 9044 32900 9054
rect 32844 8950 32900 8988
rect 33068 8820 33124 8830
rect 32956 8818 33124 8820
rect 32956 8766 33070 8818
rect 33122 8766 33124 8818
rect 32956 8764 33124 8766
rect 32732 8428 32900 8484
rect 32620 8418 32676 8428
rect 32732 8260 32788 8270
rect 32732 8166 32788 8204
rect 32284 7858 32340 7868
rect 32396 7868 32564 7924
rect 32844 8036 32900 8428
rect 32060 7746 32116 7756
rect 31836 7646 31838 7698
rect 31890 7646 31892 7698
rect 31836 7634 31892 7646
rect 31948 7364 32004 7374
rect 31724 6468 31780 6478
rect 31724 6374 31780 6412
rect 31724 4900 31780 4910
rect 31724 4676 31780 4844
rect 31948 4900 32004 7308
rect 31948 4834 32004 4844
rect 32284 5124 32340 5134
rect 32172 4788 32228 4798
rect 32060 4732 32172 4788
rect 32060 4676 32116 4732
rect 32172 4722 32228 4732
rect 31724 4620 32116 4676
rect 32172 4338 32228 4350
rect 32172 4286 32174 4338
rect 32226 4286 32228 4338
rect 31612 4116 31668 4126
rect 31612 4022 31668 4060
rect 32060 3780 32116 3790
rect 31948 2772 32004 2782
rect 31500 2718 31502 2770
rect 31554 2718 31556 2770
rect 31500 2706 31556 2718
rect 31836 2716 31948 2772
rect 31724 2548 31780 2558
rect 31724 2454 31780 2492
rect 31724 2212 31780 2222
rect 31836 2212 31892 2716
rect 31948 2706 32004 2716
rect 31724 2210 31892 2212
rect 31724 2158 31726 2210
rect 31778 2158 31892 2210
rect 31724 2156 31892 2158
rect 31724 2146 31780 2156
rect 31276 1138 31332 1148
rect 31612 1652 31668 1662
rect 31612 112 31668 1596
rect 31724 1428 31780 1438
rect 31724 1314 31780 1372
rect 31724 1262 31726 1314
rect 31778 1262 31780 1314
rect 31724 1250 31780 1262
rect 32060 1090 32116 3724
rect 32172 2772 32228 4286
rect 32284 4228 32340 5068
rect 32284 4162 32340 4172
rect 32396 3778 32452 7868
rect 32508 7588 32564 7598
rect 32508 7140 32564 7532
rect 32844 7474 32900 7980
rect 32844 7422 32846 7474
rect 32898 7422 32900 7474
rect 32844 7410 32900 7422
rect 32508 7074 32564 7084
rect 32508 6578 32564 6590
rect 32508 6526 32510 6578
rect 32562 6526 32564 6578
rect 32508 6468 32564 6526
rect 32508 6402 32564 6412
rect 32620 6468 32676 6478
rect 32620 6466 32900 6468
rect 32620 6414 32622 6466
rect 32674 6414 32900 6466
rect 32620 6412 32900 6414
rect 32620 6402 32676 6412
rect 32620 5906 32676 5918
rect 32620 5854 32622 5906
rect 32674 5854 32676 5906
rect 32620 5796 32676 5854
rect 32620 5730 32676 5740
rect 32732 5684 32788 5694
rect 32620 4340 32676 4350
rect 32620 4246 32676 4284
rect 32732 4228 32788 5628
rect 32844 5348 32900 6412
rect 32956 6356 33012 8764
rect 33068 8754 33124 8764
rect 33180 8258 33236 8270
rect 33180 8206 33182 8258
rect 33234 8206 33236 8258
rect 33180 8148 33236 8206
rect 33180 7364 33236 8092
rect 33292 7474 33348 9212
rect 33404 8596 33460 9886
rect 33404 8530 33460 8540
rect 33740 9042 33796 9054
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33516 8484 33572 8494
rect 33292 7422 33294 7474
rect 33346 7422 33348 7474
rect 33292 7410 33348 7422
rect 33404 8370 33460 8382
rect 33404 8318 33406 8370
rect 33458 8318 33460 8370
rect 33180 7298 33236 7308
rect 33068 6804 33124 6814
rect 33068 6710 33124 6748
rect 33292 6690 33348 6702
rect 33292 6638 33294 6690
rect 33346 6638 33348 6690
rect 33180 6580 33236 6590
rect 33180 6486 33236 6524
rect 33292 6356 33348 6638
rect 32956 6300 33236 6356
rect 32844 5122 32900 5292
rect 32844 5070 32846 5122
rect 32898 5070 32900 5122
rect 32844 5058 32900 5070
rect 32956 6132 33012 6142
rect 32732 4162 32788 4172
rect 32396 3726 32398 3778
rect 32450 3726 32452 3778
rect 32396 3714 32452 3726
rect 32508 4116 32564 4126
rect 32172 2678 32228 2716
rect 32284 3668 32340 3678
rect 32284 2436 32340 3612
rect 32284 2370 32340 2380
rect 32508 2098 32564 4060
rect 32732 3668 32788 3678
rect 32732 3574 32788 3612
rect 32956 2996 33012 6076
rect 33068 5684 33124 5722
rect 33068 5618 33124 5628
rect 33068 5460 33124 5470
rect 33068 5346 33124 5404
rect 33068 5294 33070 5346
rect 33122 5294 33124 5346
rect 33068 5282 33124 5294
rect 33180 5010 33236 6300
rect 33292 5460 33348 6300
rect 33292 5394 33348 5404
rect 33404 5348 33460 8318
rect 33516 7588 33572 8428
rect 33740 8260 33796 8990
rect 33852 9044 33908 12236
rect 33964 12180 34020 12190
rect 33964 12086 34020 12124
rect 34524 12068 34580 12078
rect 34636 12068 34692 13580
rect 34524 12066 34692 12068
rect 34524 12014 34526 12066
rect 34578 12014 34692 12066
rect 34524 12012 34692 12014
rect 34412 11394 34468 11406
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 34300 10164 34356 10174
rect 34076 9828 34132 9838
rect 34076 9826 34244 9828
rect 34076 9774 34078 9826
rect 34130 9774 34244 9826
rect 34076 9772 34244 9774
rect 34076 9762 34132 9772
rect 34076 9044 34132 9054
rect 33852 9042 34132 9044
rect 33852 8990 34078 9042
rect 34130 8990 34132 9042
rect 33852 8988 34132 8990
rect 34076 8978 34132 8988
rect 34188 8372 34244 9772
rect 33852 8260 33908 8270
rect 33740 8258 33908 8260
rect 33740 8206 33854 8258
rect 33906 8206 33908 8258
rect 33740 8204 33908 8206
rect 33852 8036 33908 8204
rect 33852 7970 33908 7980
rect 33516 7522 33572 7532
rect 34188 7474 34244 8316
rect 34188 7422 34190 7474
rect 34242 7422 34244 7474
rect 34188 7410 34244 7422
rect 33516 7250 33572 7262
rect 33516 7198 33518 7250
rect 33570 7198 33572 7250
rect 33516 7028 33572 7198
rect 33516 6962 33572 6972
rect 33516 6580 33572 6590
rect 33516 6486 33572 6524
rect 34188 6580 34244 6590
rect 34188 6486 34244 6524
rect 33740 6468 33796 6478
rect 34076 6468 34132 6478
rect 33740 6466 34132 6468
rect 33740 6414 33742 6466
rect 33794 6414 34078 6466
rect 34130 6414 34132 6466
rect 33740 6412 34132 6414
rect 33740 6402 33796 6412
rect 33852 6020 33908 6412
rect 34076 6402 34132 6412
rect 34188 6132 34244 6142
rect 34188 6038 34244 6076
rect 33628 5964 33908 6020
rect 33516 5348 33572 5358
rect 33404 5346 33572 5348
rect 33404 5294 33518 5346
rect 33570 5294 33572 5346
rect 33404 5292 33572 5294
rect 33516 5282 33572 5292
rect 33628 5346 33684 5964
rect 34300 5684 34356 10108
rect 34412 10052 34468 11342
rect 34524 11172 34580 12012
rect 34524 11106 34580 11116
rect 34748 11508 34804 15148
rect 34636 10388 34692 10398
rect 34412 9716 34468 9996
rect 34412 9650 34468 9660
rect 34524 10386 34692 10388
rect 34524 10334 34638 10386
rect 34690 10334 34692 10386
rect 34524 10332 34692 10334
rect 34524 10164 34580 10332
rect 34636 10322 34692 10332
rect 34412 8260 34468 8270
rect 34412 8166 34468 8204
rect 34524 8036 34580 10108
rect 34636 9828 34692 9838
rect 34636 9734 34692 9772
rect 34412 7980 34580 8036
rect 34636 8596 34692 8606
rect 34412 6802 34468 7980
rect 34412 6750 34414 6802
rect 34466 6750 34468 6802
rect 34412 6738 34468 6750
rect 34524 7028 34580 7038
rect 34524 6580 34580 6972
rect 34300 5618 34356 5628
rect 34412 6524 34580 6580
rect 34412 5460 34468 6524
rect 34076 5404 34468 5460
rect 34524 6132 34580 6142
rect 33628 5294 33630 5346
rect 33682 5294 33684 5346
rect 33628 5282 33684 5294
rect 33740 5348 33796 5358
rect 33740 5254 33796 5292
rect 33180 4958 33182 5010
rect 33234 4958 33236 5010
rect 33180 4946 33236 4958
rect 34076 4900 34132 5404
rect 34412 5236 34468 5246
rect 34188 5234 34468 5236
rect 34188 5182 34414 5234
rect 34466 5182 34468 5234
rect 34188 5180 34468 5182
rect 34188 5122 34244 5180
rect 34412 5170 34468 5180
rect 34524 5234 34580 6076
rect 34636 6130 34692 8540
rect 34748 7474 34804 11452
rect 34748 7422 34750 7474
rect 34802 7422 34804 7474
rect 34748 7410 34804 7422
rect 34860 14532 34916 14542
rect 34860 12964 34916 14476
rect 34972 14418 35028 14430
rect 34972 14366 34974 14418
rect 35026 14366 35028 14418
rect 34972 14308 35028 14366
rect 34972 14242 35028 14252
rect 34972 12964 35028 12974
rect 34860 12962 35028 12964
rect 34860 12910 34974 12962
rect 35026 12910 35028 12962
rect 34860 12908 35028 12910
rect 34860 7476 34916 12908
rect 34972 12898 35028 12908
rect 35084 12628 35140 12638
rect 34972 12292 35028 12302
rect 34972 11956 35028 12236
rect 34972 9044 35028 11900
rect 35084 9828 35140 12572
rect 35196 11396 35252 15260
rect 35308 14084 35364 19292
rect 35980 18564 36036 20748
rect 35980 18498 36036 18508
rect 35420 18340 35476 18350
rect 35420 18246 35476 18284
rect 35532 18340 35588 18350
rect 35756 18340 35812 18350
rect 35532 18338 35756 18340
rect 35532 18286 35534 18338
rect 35586 18286 35756 18338
rect 35532 18284 35756 18286
rect 35532 18274 35588 18284
rect 35756 18274 35812 18284
rect 35532 16996 35588 17006
rect 35420 16658 35476 16670
rect 35420 16606 35422 16658
rect 35474 16606 35476 16658
rect 35420 14530 35476 16606
rect 35532 16322 35588 16940
rect 35532 16270 35534 16322
rect 35586 16270 35588 16322
rect 35532 16258 35588 16270
rect 35756 15876 35812 15886
rect 35756 15092 35812 15820
rect 36092 15148 36148 22316
rect 36204 21588 36260 24220
rect 36764 23938 36820 24220
rect 36764 23886 36766 23938
rect 36818 23886 36820 23938
rect 36764 23874 36820 23886
rect 36428 23828 36484 23838
rect 36652 23828 36708 23838
rect 36428 23734 36484 23772
rect 36540 23772 36652 23828
rect 36316 23268 36372 23278
rect 36316 23174 36372 23212
rect 36428 22932 36484 22942
rect 36428 22838 36484 22876
rect 36540 22708 36596 23772
rect 36652 23762 36708 23772
rect 36764 23716 36820 23726
rect 36652 23156 36708 23166
rect 36652 23062 36708 23100
rect 36204 21522 36260 21532
rect 36316 22652 36596 22708
rect 36204 20692 36260 20702
rect 36204 20598 36260 20636
rect 36316 20468 36372 22652
rect 36540 22370 36596 22382
rect 36540 22318 36542 22370
rect 36594 22318 36596 22370
rect 36428 21586 36484 21598
rect 36428 21534 36430 21586
rect 36482 21534 36484 21586
rect 36428 21140 36484 21534
rect 36428 21074 36484 21084
rect 36540 20692 36596 22318
rect 36764 22036 36820 23660
rect 36876 23268 36932 28028
rect 36988 27746 37044 28252
rect 36988 27694 36990 27746
rect 37042 27694 37044 27746
rect 36988 27682 37044 27694
rect 37100 27412 37156 27422
rect 37100 27074 37156 27356
rect 37100 27022 37102 27074
rect 37154 27022 37156 27074
rect 36988 25508 37044 25518
rect 36988 25414 37044 25452
rect 36988 24498 37044 24510
rect 36988 24446 36990 24498
rect 37042 24446 37044 24498
rect 36988 24164 37044 24446
rect 36988 24098 37044 24108
rect 36876 23156 36932 23212
rect 37100 23268 37156 27022
rect 37212 26292 37268 28476
rect 37212 26226 37268 26236
rect 37324 25508 37380 29596
rect 37436 26908 37492 30716
rect 37548 27298 37604 32060
rect 37772 30212 37828 33628
rect 37884 31778 37940 33852
rect 37996 33346 38052 35252
rect 38220 35028 38276 36204
rect 38220 34962 38276 34972
rect 38220 34468 38276 34478
rect 38108 34244 38164 34254
rect 38108 34130 38164 34188
rect 38108 34078 38110 34130
rect 38162 34078 38164 34130
rect 38108 33796 38164 34078
rect 38108 33730 38164 33740
rect 37996 33294 37998 33346
rect 38050 33294 38052 33346
rect 37996 32900 38052 33294
rect 38220 33124 38276 34412
rect 38332 34244 38388 36990
rect 38444 35140 38500 35150
rect 38556 35140 38612 38892
rect 38668 38948 38724 38958
rect 38668 35252 38724 38892
rect 38892 37940 38948 39900
rect 39228 39732 39284 40012
rect 39228 39666 39284 39676
rect 39452 40292 39508 40302
rect 39452 39730 39508 40236
rect 39564 39844 39620 39854
rect 39676 39844 39732 41132
rect 39564 39842 39732 39844
rect 39564 39790 39566 39842
rect 39618 39790 39732 39842
rect 39564 39788 39732 39790
rect 39788 39842 39844 41916
rect 39788 39790 39790 39842
rect 39842 39790 39844 39842
rect 39564 39778 39620 39788
rect 39788 39778 39844 39790
rect 39452 39678 39454 39730
rect 39506 39678 39508 39730
rect 39004 39396 39060 39406
rect 39004 39394 39284 39396
rect 39004 39342 39006 39394
rect 39058 39342 39284 39394
rect 39004 39340 39284 39342
rect 39004 39330 39060 39340
rect 39004 38612 39060 38622
rect 39004 38610 39172 38612
rect 39004 38558 39006 38610
rect 39058 38558 39172 38610
rect 39004 38556 39172 38558
rect 39004 38546 39060 38556
rect 38892 37874 38948 37884
rect 39116 37266 39172 38556
rect 39116 37214 39118 37266
rect 39170 37214 39172 37266
rect 39116 37202 39172 37214
rect 38780 37154 38836 37166
rect 38780 37102 38782 37154
rect 38834 37102 38836 37154
rect 38780 35812 38836 37102
rect 38892 35812 38948 35822
rect 38780 35810 38948 35812
rect 38780 35758 38894 35810
rect 38946 35758 38948 35810
rect 38780 35756 38948 35758
rect 38780 35588 38836 35756
rect 38892 35746 38948 35756
rect 38780 35522 38836 35532
rect 39116 35700 39172 35710
rect 38668 35186 38724 35196
rect 38500 35084 38612 35140
rect 38444 35074 38500 35084
rect 38332 34178 38388 34188
rect 38556 34804 38612 35084
rect 38780 34804 38836 34814
rect 38556 34748 38780 34804
rect 38444 33796 38500 33806
rect 38556 33796 38612 34748
rect 38780 34738 38836 34748
rect 38500 33740 38612 33796
rect 38892 34580 38948 34590
rect 38892 33796 38948 34524
rect 39004 34132 39060 34142
rect 39004 33908 39060 34076
rect 39004 33842 39060 33852
rect 38444 33570 38500 33740
rect 38892 33730 38948 33740
rect 38444 33518 38446 33570
rect 38498 33518 38500 33570
rect 38444 33506 38500 33518
rect 38220 33068 38612 33124
rect 37996 32844 38164 32900
rect 37996 32676 38052 32686
rect 37996 32582 38052 32620
rect 37884 31726 37886 31778
rect 37938 31726 37940 31778
rect 37884 31444 37940 31726
rect 37884 31378 37940 31388
rect 37996 31780 38052 31790
rect 37884 31220 37940 31230
rect 37884 30436 37940 31164
rect 37884 30370 37940 30380
rect 37772 30156 37940 30212
rect 37772 29988 37828 29998
rect 37772 29894 37828 29932
rect 37660 29426 37716 29438
rect 37660 29374 37662 29426
rect 37714 29374 37716 29426
rect 37660 29092 37716 29374
rect 37772 29316 37828 29326
rect 37884 29316 37940 30156
rect 37772 29314 37940 29316
rect 37772 29262 37774 29314
rect 37826 29262 37940 29314
rect 37772 29260 37940 29262
rect 37772 29250 37828 29260
rect 37716 29036 37828 29092
rect 37660 29026 37716 29036
rect 37548 27246 37550 27298
rect 37602 27246 37604 27298
rect 37548 27234 37604 27246
rect 37436 26852 37716 26908
rect 37324 25442 37380 25452
rect 37548 25620 37604 25630
rect 37324 24724 37380 24734
rect 37212 23938 37268 23950
rect 37212 23886 37214 23938
rect 37266 23886 37268 23938
rect 37212 23492 37268 23886
rect 37212 23426 37268 23436
rect 37100 23202 37156 23212
rect 36988 23156 37044 23166
rect 36876 23154 37044 23156
rect 36876 23102 36990 23154
rect 37042 23102 37044 23154
rect 36876 23100 37044 23102
rect 36988 23090 37044 23100
rect 37212 23156 37268 23166
rect 37212 23062 37268 23100
rect 37100 22930 37156 22942
rect 37100 22878 37102 22930
rect 37154 22878 37156 22930
rect 37100 22708 37156 22878
rect 37100 22642 37156 22652
rect 37100 22484 37156 22494
rect 37324 22484 37380 24668
rect 37436 24050 37492 24062
rect 37436 23998 37438 24050
rect 37490 23998 37492 24050
rect 37436 23940 37492 23998
rect 37436 23874 37492 23884
rect 37100 22482 37380 22484
rect 37100 22430 37102 22482
rect 37154 22430 37380 22482
rect 37100 22428 37380 22430
rect 37100 22418 37156 22428
rect 37548 22372 37604 25564
rect 37660 24724 37716 26852
rect 37660 24658 37716 24668
rect 37660 24388 37716 24398
rect 37660 23828 37716 24332
rect 37660 23762 37716 23772
rect 37548 22306 37604 22316
rect 37660 23154 37716 23166
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 37436 22148 37492 22158
rect 36764 21980 36932 22036
rect 36764 21812 36820 21822
rect 36652 21028 36708 21038
rect 36652 20934 36708 20972
rect 36540 20626 36596 20636
rect 36204 20412 36372 20468
rect 36204 16772 36260 20412
rect 36428 19012 36484 19022
rect 36428 19010 36708 19012
rect 36428 18958 36430 19010
rect 36482 18958 36708 19010
rect 36428 18956 36708 18958
rect 36428 18946 36484 18956
rect 36540 18564 36596 18574
rect 36316 18340 36372 18350
rect 36316 17778 36372 18284
rect 36316 17726 36318 17778
rect 36370 17726 36372 17778
rect 36316 17714 36372 17726
rect 36204 16706 36260 16716
rect 36316 17444 36372 17454
rect 35756 15026 35812 15036
rect 35980 15092 36036 15102
rect 36092 15092 36260 15148
rect 35980 14754 36036 15036
rect 35980 14702 35982 14754
rect 36034 14702 36036 14754
rect 35980 14690 36036 14702
rect 36092 14868 36148 14878
rect 35420 14478 35422 14530
rect 35474 14478 35476 14530
rect 35420 14466 35476 14478
rect 35532 14532 35588 14542
rect 35308 14018 35364 14028
rect 35420 14308 35476 14318
rect 35308 13746 35364 13758
rect 35308 13694 35310 13746
rect 35362 13694 35364 13746
rect 35308 11620 35364 13694
rect 35308 11554 35364 11564
rect 35308 11396 35364 11406
rect 35196 11394 35364 11396
rect 35196 11342 35310 11394
rect 35362 11342 35364 11394
rect 35196 11340 35364 11342
rect 35308 11330 35364 11340
rect 35420 10948 35476 14252
rect 35532 13300 35588 14476
rect 35532 13186 35588 13244
rect 35532 13134 35534 13186
rect 35586 13134 35588 13186
rect 35532 13122 35588 13134
rect 35868 14530 35924 14542
rect 35868 14478 35870 14530
rect 35922 14478 35924 14530
rect 35644 11956 35700 11966
rect 35644 11954 35812 11956
rect 35644 11902 35646 11954
rect 35698 11902 35812 11954
rect 35644 11900 35812 11902
rect 35644 11890 35700 11900
rect 35644 11620 35700 11630
rect 35084 9762 35140 9772
rect 35308 10892 35476 10948
rect 35532 11394 35588 11406
rect 35532 11342 35534 11394
rect 35586 11342 35588 11394
rect 35084 9044 35140 9054
rect 34972 9042 35140 9044
rect 34972 8990 35086 9042
rect 35138 8990 35140 9042
rect 34972 8988 35140 8990
rect 35084 8978 35140 8988
rect 34860 7410 34916 7420
rect 34748 6804 34804 6842
rect 34748 6738 34804 6748
rect 35196 6804 35252 6814
rect 34972 6690 35028 6702
rect 34972 6638 34974 6690
rect 35026 6638 35028 6690
rect 34972 6468 35028 6638
rect 34748 6412 35028 6468
rect 35084 6578 35140 6590
rect 35084 6526 35086 6578
rect 35138 6526 35140 6578
rect 34748 6356 34804 6412
rect 34748 6290 34804 6300
rect 35084 6238 35140 6526
rect 35196 6468 35252 6748
rect 35308 6468 35364 10892
rect 35532 10724 35588 11342
rect 35644 10948 35700 11564
rect 35756 11396 35812 11900
rect 35868 11620 35924 14478
rect 36092 12292 36148 14812
rect 36204 12852 36260 15092
rect 36316 13636 36372 17388
rect 36540 16882 36596 18508
rect 36652 18450 36708 18956
rect 36652 18398 36654 18450
rect 36706 18398 36708 18450
rect 36652 18386 36708 18398
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 36540 16100 36596 16830
rect 36652 17666 36708 17678
rect 36652 17614 36654 17666
rect 36706 17614 36708 17666
rect 36652 16322 36708 17614
rect 36652 16270 36654 16322
rect 36706 16270 36708 16322
rect 36652 16258 36708 16270
rect 36540 16044 36708 16100
rect 36316 13570 36372 13580
rect 36540 15428 36596 15438
rect 36540 13412 36596 15372
rect 36652 14980 36708 16044
rect 36764 15148 36820 21756
rect 36876 21588 36932 21980
rect 37324 21588 37380 21598
rect 36876 21586 37380 21588
rect 36876 21534 37326 21586
rect 37378 21534 37380 21586
rect 36876 21532 37380 21534
rect 37100 20020 37156 20030
rect 37100 19926 37156 19964
rect 36988 19236 37044 19246
rect 36988 18564 37044 19180
rect 37324 18564 37380 21532
rect 37436 19236 37492 22092
rect 37660 21028 37716 23102
rect 37772 21812 37828 29036
rect 37884 28756 37940 28766
rect 37884 26404 37940 28700
rect 37884 26310 37940 26348
rect 37884 24836 37940 24846
rect 37884 23492 37940 24780
rect 37996 24388 38052 31724
rect 38108 31444 38164 32844
rect 38220 32564 38276 32574
rect 38220 32228 38276 32508
rect 38556 32562 38612 33068
rect 39116 32788 39172 35644
rect 39228 35698 39284 39340
rect 39452 38668 39508 39678
rect 39900 39620 39956 44380
rect 39228 35646 39230 35698
rect 39282 35646 39284 35698
rect 39228 35634 39284 35646
rect 39340 38612 39508 38668
rect 39564 39564 39956 39620
rect 39228 35364 39284 35374
rect 39228 32900 39284 35308
rect 39340 33684 39396 38612
rect 39564 35308 39620 39564
rect 39788 39172 39844 39182
rect 39676 38948 39732 38958
rect 39676 38854 39732 38892
rect 39788 38164 39844 39116
rect 40012 39060 40068 44828
rect 40236 44436 40292 47012
rect 40684 46674 40740 46686
rect 40684 46622 40686 46674
rect 40738 46622 40740 46674
rect 40348 46340 40404 46350
rect 40348 44772 40404 46284
rect 40460 45780 40516 45790
rect 40684 45780 40740 46622
rect 40460 45778 40740 45780
rect 40460 45726 40462 45778
rect 40514 45726 40740 45778
rect 40460 45724 40740 45726
rect 40460 45714 40516 45724
rect 40684 45556 40740 45724
rect 40572 45108 40628 45118
rect 40684 45108 40740 45500
rect 40572 45106 40740 45108
rect 40572 45054 40574 45106
rect 40626 45054 40740 45106
rect 40572 45052 40740 45054
rect 40572 45042 40628 45052
rect 40348 44716 40628 44772
rect 40236 44370 40292 44380
rect 40348 43876 40404 43886
rect 40236 43428 40292 43438
rect 40236 41412 40292 43372
rect 40348 41972 40404 43820
rect 40460 43428 40516 43438
rect 40460 43334 40516 43372
rect 40572 43092 40628 44716
rect 40684 44322 40740 45052
rect 40796 46002 40852 46014
rect 40796 45950 40798 46002
rect 40850 45950 40852 46002
rect 40796 44884 40852 45950
rect 40796 44818 40852 44828
rect 40908 44436 40964 48860
rect 41244 48692 41300 51100
rect 41356 48916 41412 52670
rect 41468 50596 41524 54238
rect 41580 53842 41636 54796
rect 41580 53790 41582 53842
rect 41634 53790 41636 53842
rect 41580 53396 41636 53790
rect 41580 53330 41636 53340
rect 41580 52276 41636 52286
rect 41580 52052 41636 52220
rect 41692 52164 41748 55806
rect 41804 54964 41860 56028
rect 41916 55524 41972 57344
rect 42140 56644 42196 56654
rect 42140 56082 42196 56588
rect 42140 56030 42142 56082
rect 42194 56030 42196 56082
rect 42140 56018 42196 56030
rect 42364 56084 42420 57344
rect 42364 56018 42420 56028
rect 41916 55458 41972 55468
rect 42364 55858 42420 55870
rect 42364 55806 42366 55858
rect 42418 55806 42420 55858
rect 42140 55410 42196 55422
rect 42140 55358 42142 55410
rect 42194 55358 42196 55410
rect 41804 54898 41860 54908
rect 41916 55298 41972 55310
rect 41916 55246 41918 55298
rect 41970 55246 41972 55298
rect 41916 54404 41972 55246
rect 42028 54852 42084 54862
rect 42028 54404 42084 54796
rect 42140 54628 42196 55358
rect 42364 54964 42420 55806
rect 42812 55636 42868 57344
rect 43260 56420 43316 57344
rect 43708 57316 43764 57344
rect 43708 57250 43764 57260
rect 43260 56354 43316 56364
rect 43484 56980 43540 56990
rect 42812 55570 42868 55580
rect 43260 56082 43316 56094
rect 43260 56030 43262 56082
rect 43314 56030 43316 56082
rect 42812 55412 42868 55422
rect 42812 55410 42980 55412
rect 42812 55358 42814 55410
rect 42866 55358 42980 55410
rect 42812 55356 42980 55358
rect 42812 55346 42868 55356
rect 42588 55298 42644 55310
rect 42588 55246 42590 55298
rect 42642 55246 42644 55298
rect 42588 55188 42644 55246
rect 42588 55122 42644 55132
rect 42364 54898 42420 54908
rect 42140 54562 42196 54572
rect 42476 54516 42532 54526
rect 42252 54514 42532 54516
rect 42252 54462 42478 54514
rect 42530 54462 42532 54514
rect 42252 54460 42532 54462
rect 42140 54404 42196 54414
rect 42028 54402 42196 54404
rect 42028 54350 42142 54402
rect 42194 54350 42196 54402
rect 42028 54348 42196 54350
rect 41916 54338 41972 54348
rect 42140 54338 42196 54348
rect 41804 54292 41860 54302
rect 41804 54198 41860 54236
rect 41804 53730 41860 53742
rect 41804 53678 41806 53730
rect 41858 53678 41860 53730
rect 41804 53284 41860 53678
rect 42140 53732 42196 53742
rect 41804 53228 42084 53284
rect 41804 52948 41860 52958
rect 41804 52724 41860 52892
rect 41804 52630 41860 52668
rect 42028 52386 42084 53228
rect 42028 52334 42030 52386
rect 42082 52334 42084 52386
rect 42028 52322 42084 52334
rect 41692 52108 42084 52164
rect 41580 51996 41860 52052
rect 41580 51044 41636 51054
rect 41580 50706 41636 50988
rect 41580 50654 41582 50706
rect 41634 50654 41636 50706
rect 41580 50642 41636 50654
rect 41468 50530 41524 50540
rect 41692 49810 41748 49822
rect 41692 49758 41694 49810
rect 41746 49758 41748 49810
rect 41692 49028 41748 49758
rect 41804 49252 41860 51996
rect 41916 51380 41972 51390
rect 41916 50594 41972 51324
rect 41916 50542 41918 50594
rect 41970 50542 41972 50594
rect 41916 50530 41972 50542
rect 41804 49186 41860 49196
rect 42028 49028 42084 52108
rect 42140 51492 42196 53676
rect 42252 51602 42308 54460
rect 42476 54450 42532 54460
rect 42700 54516 42756 54526
rect 42700 54422 42756 54460
rect 42812 54180 42868 54190
rect 42700 53618 42756 53630
rect 42700 53566 42702 53618
rect 42754 53566 42756 53618
rect 42700 53508 42756 53566
rect 42700 53442 42756 53452
rect 42252 51550 42254 51602
rect 42306 51550 42308 51602
rect 42252 51538 42308 51550
rect 42588 52162 42644 52174
rect 42588 52110 42590 52162
rect 42642 52110 42644 52162
rect 42140 50428 42196 51436
rect 42476 51380 42532 51390
rect 42476 50932 42532 51324
rect 42588 51044 42644 52110
rect 42700 51604 42756 51614
rect 42700 51510 42756 51548
rect 42812 51378 42868 54124
rect 42924 53284 42980 55356
rect 43148 55298 43204 55310
rect 43148 55246 43150 55298
rect 43202 55246 43204 55298
rect 43036 54290 43092 54302
rect 43036 54238 43038 54290
rect 43090 54238 43092 54290
rect 43036 54180 43092 54238
rect 43036 54114 43092 54124
rect 43148 54068 43204 55246
rect 43260 55076 43316 56030
rect 43484 55970 43540 56924
rect 44156 56644 44212 57344
rect 44380 56644 44436 56654
rect 44156 56588 44380 56644
rect 44380 56578 44436 56588
rect 43484 55918 43486 55970
rect 43538 55918 43540 55970
rect 43484 55906 43540 55918
rect 43596 56532 43652 56542
rect 44604 56532 44660 57344
rect 45052 56868 45108 57344
rect 45052 56802 45108 56812
rect 45276 56868 45332 56878
rect 45164 56756 45220 56766
rect 43596 55636 43652 56476
rect 43804 56476 44068 56486
rect 44604 56476 44996 56532
rect 43860 56420 43908 56476
rect 43964 56420 44012 56476
rect 43804 56410 44068 56420
rect 44156 56420 44212 56430
rect 43820 56308 43876 56318
rect 43820 56082 43876 56252
rect 43820 56030 43822 56082
rect 43874 56030 43876 56082
rect 43820 56018 43876 56030
rect 44156 55970 44212 56364
rect 44716 56308 44772 56318
rect 44268 56252 44716 56308
rect 44268 56196 44324 56252
rect 44716 56242 44772 56252
rect 44268 56130 44324 56140
rect 44156 55918 44158 55970
rect 44210 55918 44212 55970
rect 44156 55906 44212 55918
rect 44492 55860 44548 55898
rect 44492 55794 44548 55804
rect 44828 55860 44884 55870
rect 44828 55766 44884 55804
rect 44464 55692 44728 55702
rect 43596 55570 43652 55580
rect 44268 55636 44324 55646
rect 44520 55636 44568 55692
rect 44624 55636 44672 55692
rect 44464 55626 44728 55636
rect 44940 55636 44996 56476
rect 45164 56082 45220 56700
rect 45276 56196 45332 56812
rect 45276 56130 45332 56140
rect 45500 56196 45556 57344
rect 45500 56130 45556 56140
rect 45164 56030 45166 56082
rect 45218 56030 45220 56082
rect 45164 56018 45220 56030
rect 45836 56084 45892 56094
rect 45836 55990 45892 56028
rect 45500 55860 45556 55870
rect 45500 55858 45668 55860
rect 45500 55806 45502 55858
rect 45554 55806 45668 55858
rect 45500 55804 45668 55806
rect 45500 55794 45556 55804
rect 43484 55524 43540 55534
rect 43484 55430 43540 55468
rect 44268 55468 44324 55580
rect 44940 55570 44996 55580
rect 43820 55410 43876 55422
rect 44268 55412 44436 55468
rect 43820 55358 43822 55410
rect 43874 55358 43876 55410
rect 43820 55300 43876 55358
rect 43820 55234 43876 55244
rect 44156 55300 44212 55310
rect 44156 55206 44212 55244
rect 44380 55300 44436 55412
rect 44492 55412 44548 55422
rect 45164 55412 45220 55422
rect 44492 55318 44548 55356
rect 44940 55410 45220 55412
rect 44940 55358 45166 55410
rect 45218 55358 45220 55410
rect 44940 55356 45220 55358
rect 45612 55412 45668 55804
rect 45948 55636 46004 57344
rect 46172 57316 46228 57326
rect 46172 55970 46228 57260
rect 46172 55918 46174 55970
rect 46226 55918 46228 55970
rect 46172 55906 46228 55918
rect 46284 56532 46340 56542
rect 45948 55570 46004 55580
rect 45612 55356 46004 55412
rect 44380 55234 44436 55244
rect 44828 55298 44884 55310
rect 44828 55246 44830 55298
rect 44882 55246 44884 55298
rect 43260 55010 43316 55020
rect 43596 55020 44212 55076
rect 43596 54964 43652 55020
rect 44156 54964 44212 55020
rect 43596 54898 43652 54908
rect 43804 54908 44068 54918
rect 43860 54852 43908 54908
rect 43964 54852 44012 54908
rect 44156 54898 44212 54908
rect 43804 54842 44068 54852
rect 44268 54852 44324 54862
rect 44156 54516 44212 54526
rect 43372 54514 44212 54516
rect 43372 54462 44158 54514
rect 44210 54462 44212 54514
rect 43372 54460 44212 54462
rect 43372 54402 43428 54460
rect 43372 54350 43374 54402
rect 43426 54350 43428 54402
rect 43148 54012 43316 54068
rect 43148 53844 43204 53854
rect 43148 53750 43204 53788
rect 43260 53620 43316 54012
rect 43372 53732 43428 54350
rect 43372 53666 43428 53676
rect 43484 54290 43540 54302
rect 43708 54292 43764 54302
rect 43484 54238 43486 54290
rect 43538 54238 43540 54290
rect 43260 53554 43316 53564
rect 42924 53228 43092 53284
rect 42924 53060 42980 53070
rect 42924 52834 42980 53004
rect 42924 52782 42926 52834
rect 42978 52782 42980 52834
rect 42924 52770 42980 52782
rect 42924 52274 42980 52286
rect 42924 52222 42926 52274
rect 42978 52222 42980 52274
rect 42924 51492 42980 52222
rect 43036 52276 43092 53228
rect 43372 52946 43428 52958
rect 43372 52894 43374 52946
rect 43426 52894 43428 52946
rect 43372 52724 43428 52894
rect 43372 52658 43428 52668
rect 43484 52388 43540 54238
rect 43036 52210 43092 52220
rect 43372 52332 43540 52388
rect 43596 54290 43764 54292
rect 43596 54238 43710 54290
rect 43762 54238 43764 54290
rect 43596 54236 43764 54238
rect 43596 52388 43652 54236
rect 43708 54226 43764 54236
rect 44156 53732 44212 54460
rect 44268 54402 44324 54796
rect 44492 54516 44548 54526
rect 44492 54422 44548 54460
rect 44268 54350 44270 54402
rect 44322 54350 44324 54402
rect 44268 54338 44324 54350
rect 44716 54292 44772 54330
rect 44716 54226 44772 54236
rect 44464 54124 44728 54134
rect 44520 54068 44568 54124
rect 44624 54068 44672 54124
rect 44464 54058 44728 54068
rect 44828 53956 44884 55246
rect 44940 54740 44996 55356
rect 45164 55346 45220 55356
rect 45388 55298 45444 55310
rect 45388 55246 45390 55298
rect 45442 55246 45444 55298
rect 45388 54852 45444 55246
rect 45388 54786 45444 54796
rect 45724 54964 45780 54974
rect 45724 54740 45780 54908
rect 45948 54964 46004 55356
rect 46060 55410 46116 55422
rect 46060 55358 46062 55410
rect 46114 55358 46116 55410
rect 46060 55188 46116 55358
rect 46060 55122 46116 55132
rect 45948 54898 46004 54908
rect 46060 54740 46116 54750
rect 45724 54684 46060 54740
rect 44940 54674 44996 54684
rect 46060 54674 46116 54684
rect 45612 54514 45668 54526
rect 45612 54462 45614 54514
rect 45666 54462 45668 54514
rect 45388 54404 45444 54414
rect 45388 54310 45444 54348
rect 44604 53900 44884 53956
rect 45052 54290 45108 54302
rect 45052 54238 45054 54290
rect 45106 54238 45108 54290
rect 44604 53732 44660 53900
rect 44156 53676 44548 53732
rect 44268 53508 44324 53518
rect 44492 53508 44548 53676
rect 44604 53666 44660 53676
rect 44716 53788 44996 53844
rect 44716 53730 44772 53788
rect 44716 53678 44718 53730
rect 44770 53678 44772 53730
rect 44716 53666 44772 53678
rect 44268 53506 44436 53508
rect 44268 53454 44270 53506
rect 44322 53454 44436 53506
rect 44268 53452 44436 53454
rect 44268 53442 44324 53452
rect 44380 53396 44436 53452
rect 43804 53340 44068 53350
rect 43860 53284 43908 53340
rect 43964 53284 44012 53340
rect 44380 53330 44436 53340
rect 43804 53274 44068 53284
rect 43820 53172 43876 53182
rect 43820 52724 43876 53116
rect 44044 53116 44436 53172
rect 44044 53060 44100 53116
rect 43932 53004 44100 53060
rect 43932 52948 43988 53004
rect 43932 52882 43988 52892
rect 44156 52946 44212 52958
rect 44156 52894 44158 52946
rect 44210 52894 44212 52946
rect 44156 52724 44212 52894
rect 44380 52946 44436 53116
rect 44492 53060 44548 53452
rect 44828 53618 44884 53630
rect 44828 53566 44830 53618
rect 44882 53566 44884 53618
rect 44828 53172 44884 53566
rect 44828 53106 44884 53116
rect 44492 53004 44772 53060
rect 44380 52894 44382 52946
rect 44434 52894 44436 52946
rect 44380 52882 44436 52894
rect 44716 52946 44772 53004
rect 44716 52894 44718 52946
rect 44770 52894 44772 52946
rect 44716 52882 44772 52894
rect 43820 52668 44212 52724
rect 44604 52724 44660 52734
rect 44604 52722 44884 52724
rect 44604 52670 44606 52722
rect 44658 52670 44884 52722
rect 44604 52668 44884 52670
rect 44604 52658 44660 52668
rect 44464 52556 44728 52566
rect 44156 52500 44212 52510
rect 44520 52500 44568 52556
rect 44624 52500 44672 52556
rect 44212 52444 44324 52500
rect 44464 52490 44728 52500
rect 44156 52434 44212 52444
rect 43260 52052 43316 52062
rect 43260 51958 43316 51996
rect 43260 51604 43316 51614
rect 43260 51510 43316 51548
rect 43148 51492 43204 51502
rect 42924 51436 43092 51492
rect 42812 51326 42814 51378
rect 42866 51326 42868 51378
rect 42812 51314 42868 51326
rect 42588 50988 42756 51044
rect 42476 50876 42644 50932
rect 42140 50372 42420 50428
rect 42364 49812 42420 50372
rect 42364 49746 42420 49756
rect 42140 49700 42196 49710
rect 42140 49606 42196 49644
rect 42476 49028 42532 49038
rect 41692 48962 41748 48972
rect 41916 48972 42084 49028
rect 42364 49026 42532 49028
rect 42364 48974 42478 49026
rect 42530 48974 42532 49026
rect 42364 48972 42532 48974
rect 41356 48850 41412 48860
rect 41580 48916 41636 48926
rect 41244 48636 41412 48692
rect 41244 48244 41300 48254
rect 41020 48132 41076 48142
rect 41020 47682 41076 48076
rect 41020 47630 41022 47682
rect 41074 47630 41076 47682
rect 41020 47618 41076 47630
rect 41132 46452 41188 46462
rect 41132 46358 41188 46396
rect 41244 46116 41300 48188
rect 41356 48244 41412 48636
rect 41356 48242 41524 48244
rect 41356 48190 41358 48242
rect 41410 48190 41524 48242
rect 41356 48188 41524 48190
rect 41356 48178 41412 48188
rect 41356 47684 41412 47694
rect 41356 47590 41412 47628
rect 41244 46050 41300 46060
rect 41356 45108 41412 45118
rect 41020 44884 41076 44894
rect 41020 44790 41076 44828
rect 41244 44660 41300 44670
rect 40908 44370 40964 44380
rect 41132 44434 41188 44446
rect 41132 44382 41134 44434
rect 41186 44382 41188 44434
rect 40684 44270 40686 44322
rect 40738 44270 40740 44322
rect 40684 44258 40740 44270
rect 41020 43764 41076 43774
rect 40796 43426 40852 43438
rect 40796 43374 40798 43426
rect 40850 43374 40852 43426
rect 40348 41906 40404 41916
rect 40460 43036 40628 43092
rect 40684 43314 40740 43326
rect 40684 43262 40686 43314
rect 40738 43262 40740 43314
rect 40236 41346 40292 41356
rect 40348 41186 40404 41198
rect 40348 41134 40350 41186
rect 40402 41134 40404 41186
rect 40236 40852 40292 40862
rect 40124 40396 40180 40408
rect 40124 40344 40126 40396
rect 40178 40344 40180 40396
rect 40124 40068 40180 40344
rect 40236 40290 40292 40796
rect 40236 40238 40238 40290
rect 40290 40238 40292 40290
rect 40236 40226 40292 40238
rect 40124 40002 40180 40012
rect 40236 39732 40292 39742
rect 40236 39638 40292 39676
rect 39788 38098 39844 38108
rect 39900 39004 40068 39060
rect 39676 37266 39732 37278
rect 39676 37214 39678 37266
rect 39730 37214 39732 37266
rect 39676 35700 39732 37214
rect 39788 37268 39844 37278
rect 39788 37154 39844 37212
rect 39788 37102 39790 37154
rect 39842 37102 39844 37154
rect 39788 37090 39844 37102
rect 39788 35700 39844 35710
rect 39676 35644 39788 35700
rect 39900 35700 39956 39004
rect 40348 38948 40404 41134
rect 40348 38882 40404 38892
rect 40012 38724 40068 38762
rect 40012 38658 40068 38668
rect 40348 37826 40404 37838
rect 40348 37774 40350 37826
rect 40402 37774 40404 37826
rect 40124 37380 40180 37390
rect 39900 35644 40068 35700
rect 39788 35606 39844 35644
rect 39900 35476 39956 35486
rect 39900 35382 39956 35420
rect 39340 33618 39396 33628
rect 39452 35252 39620 35308
rect 40012 35252 40068 35644
rect 39228 32834 39284 32844
rect 39116 32722 39172 32732
rect 38556 32510 38558 32562
rect 38610 32510 38612 32562
rect 38556 32498 38612 32510
rect 39228 32562 39284 32574
rect 39228 32510 39230 32562
rect 39282 32510 39284 32562
rect 38780 32452 38836 32462
rect 38780 32358 38836 32396
rect 38892 32450 38948 32462
rect 38892 32398 38894 32450
rect 38946 32398 38948 32450
rect 38220 32162 38276 32172
rect 38668 32338 38724 32350
rect 38668 32286 38670 32338
rect 38722 32286 38724 32338
rect 38108 31378 38164 31388
rect 38444 31778 38500 31790
rect 38444 31726 38446 31778
rect 38498 31726 38500 31778
rect 38444 31332 38500 31726
rect 38444 31266 38500 31276
rect 38220 30996 38276 31006
rect 38108 30772 38164 30782
rect 38108 30678 38164 30716
rect 38220 30322 38276 30940
rect 38444 30772 38500 30782
rect 38444 30434 38500 30716
rect 38444 30382 38446 30434
rect 38498 30382 38500 30434
rect 38444 30370 38500 30382
rect 38668 30434 38724 32286
rect 38892 31892 38948 32398
rect 38892 31826 38948 31836
rect 39116 32228 39172 32238
rect 38668 30382 38670 30434
rect 38722 30382 38724 30434
rect 38668 30370 38724 30382
rect 38780 31444 38836 31454
rect 38780 31106 38836 31388
rect 38780 31054 38782 31106
rect 38834 31054 38836 31106
rect 38220 30270 38222 30322
rect 38274 30270 38276 30322
rect 38220 30258 38276 30270
rect 38332 30098 38388 30110
rect 38332 30046 38334 30098
rect 38386 30046 38388 30098
rect 38332 29988 38388 30046
rect 38332 29922 38388 29932
rect 38780 29764 38836 31054
rect 39116 30882 39172 32172
rect 39116 30830 39118 30882
rect 39170 30830 39172 30882
rect 39116 30818 39172 30830
rect 39228 30772 39284 32510
rect 39340 31780 39396 31790
rect 39340 31686 39396 31724
rect 39228 30706 39284 30716
rect 38668 29708 38780 29764
rect 38332 29426 38388 29438
rect 38332 29374 38334 29426
rect 38386 29374 38388 29426
rect 38332 28866 38388 29374
rect 38332 28814 38334 28866
rect 38386 28814 38388 28866
rect 38332 28802 38388 28814
rect 38668 28756 38724 29708
rect 38780 29698 38836 29708
rect 38892 30492 39396 30548
rect 38780 29428 38836 29438
rect 38780 29334 38836 29372
rect 38668 28690 38724 28700
rect 38780 28868 38836 28878
rect 38892 28868 38948 30492
rect 39340 30378 39396 30492
rect 39228 30322 39284 30334
rect 39228 30270 39230 30322
rect 39282 30270 39284 30322
rect 39340 30326 39342 30378
rect 39394 30326 39396 30378
rect 39340 30314 39396 30326
rect 39228 30212 39284 30270
rect 39228 30156 39396 30212
rect 38780 28866 38948 28868
rect 38780 28814 38782 28866
rect 38834 28814 38948 28866
rect 38780 28812 38948 28814
rect 39228 29986 39284 29998
rect 39228 29934 39230 29986
rect 39282 29934 39284 29986
rect 38780 28532 38836 28812
rect 39004 28642 39060 28654
rect 39004 28590 39006 28642
rect 39058 28590 39060 28642
rect 38556 28476 38780 28532
rect 38108 28084 38164 28094
rect 38556 28084 38612 28476
rect 38780 28466 38836 28476
rect 38892 28530 38948 28542
rect 38892 28478 38894 28530
rect 38946 28478 38948 28530
rect 38892 28420 38948 28478
rect 38892 28354 38948 28364
rect 39004 28196 39060 28590
rect 38108 28082 38612 28084
rect 38108 28030 38110 28082
rect 38162 28030 38612 28082
rect 38108 28028 38612 28030
rect 38108 28018 38164 28028
rect 38332 27860 38388 27870
rect 38220 27188 38276 27198
rect 38332 27188 38388 27804
rect 38556 27858 38612 28028
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 27794 38612 27806
rect 38668 28140 39060 28196
rect 38668 27524 38724 28140
rect 38892 27972 38948 27982
rect 38892 27970 39172 27972
rect 38892 27918 38894 27970
rect 38946 27918 39172 27970
rect 38892 27916 39172 27918
rect 38892 27906 38948 27916
rect 38892 27746 38948 27758
rect 38892 27694 38894 27746
rect 38946 27694 38948 27746
rect 38276 27132 38388 27188
rect 38556 27468 38724 27524
rect 38780 27634 38836 27646
rect 38780 27582 38782 27634
rect 38834 27582 38836 27634
rect 38108 26516 38164 26526
rect 38108 26180 38164 26460
rect 38108 26114 38164 26124
rect 37996 24164 38052 24332
rect 37996 24098 38052 24108
rect 38108 24498 38164 24510
rect 38108 24446 38110 24498
rect 38162 24446 38164 24498
rect 38108 23938 38164 24446
rect 38108 23886 38110 23938
rect 38162 23886 38164 23938
rect 38108 23874 38164 23886
rect 37884 23436 38052 23492
rect 37772 21746 37828 21756
rect 37996 23044 38052 23436
rect 38220 23268 38276 27132
rect 38556 26964 38612 27468
rect 38668 27300 38724 27310
rect 38668 27206 38724 27244
rect 38556 26898 38612 26908
rect 38556 26628 38612 26638
rect 38332 26180 38388 26190
rect 38332 25284 38388 26124
rect 38332 25218 38388 25228
rect 38444 23938 38500 23950
rect 38444 23886 38446 23938
rect 38498 23886 38500 23938
rect 38444 23828 38500 23886
rect 38220 23212 38388 23268
rect 38220 23044 38276 23054
rect 37996 23042 38276 23044
rect 37996 22990 38222 23042
rect 38274 22990 38276 23042
rect 37996 22988 38276 22990
rect 37660 20962 37716 20972
rect 37772 21588 37828 21598
rect 37772 21026 37828 21532
rect 37996 21364 38052 22988
rect 38220 22978 38276 22988
rect 38220 22148 38276 22158
rect 38108 22146 38276 22148
rect 38108 22094 38222 22146
rect 38274 22094 38276 22146
rect 38108 22092 38276 22094
rect 38108 21586 38164 22092
rect 38220 22082 38276 22092
rect 38108 21534 38110 21586
rect 38162 21534 38164 21586
rect 38108 21522 38164 21534
rect 38220 21924 38276 21934
rect 37996 21308 38164 21364
rect 37772 20974 37774 21026
rect 37826 20974 37828 21026
rect 37772 20962 37828 20974
rect 37548 20356 37604 20366
rect 37548 19906 37604 20300
rect 37548 19854 37550 19906
rect 37602 19854 37604 19906
rect 37548 19842 37604 19854
rect 37548 19460 37604 19470
rect 37548 19366 37604 19404
rect 37436 19180 37716 19236
rect 37324 18508 37492 18564
rect 36988 18498 37044 18508
rect 37100 18452 37156 18462
rect 37100 17892 37156 18396
rect 37324 18340 37380 18350
rect 37324 18246 37380 18284
rect 37100 17666 37156 17836
rect 37324 17892 37380 17902
rect 37324 17798 37380 17836
rect 37100 17614 37102 17666
rect 37154 17614 37156 17666
rect 37100 17602 37156 17614
rect 36988 16772 37044 16782
rect 36988 16678 37044 16716
rect 37324 16100 37380 16110
rect 37212 15988 37268 15998
rect 37324 15988 37380 16044
rect 37212 15986 37380 15988
rect 37212 15934 37214 15986
rect 37266 15934 37380 15986
rect 37212 15932 37380 15934
rect 37212 15922 37268 15932
rect 37436 15876 37492 18508
rect 37548 18340 37604 18350
rect 37548 16436 37604 18284
rect 37548 16370 37604 16380
rect 37324 15820 37492 15876
rect 37100 15204 37156 15214
rect 36764 15092 36932 15148
rect 36652 14924 36820 14980
rect 36540 13346 36596 13356
rect 36652 14530 36708 14542
rect 36652 14478 36654 14530
rect 36706 14478 36708 14530
rect 36652 13186 36708 14478
rect 36764 13636 36820 14924
rect 36764 13570 36820 13580
rect 36652 13134 36654 13186
rect 36706 13134 36708 13186
rect 36652 13122 36708 13134
rect 36204 12628 36260 12796
rect 36204 12562 36260 12572
rect 35868 11554 35924 11564
rect 35980 12236 36148 12292
rect 35868 11396 35924 11406
rect 35756 11394 35924 11396
rect 35756 11342 35870 11394
rect 35922 11342 35924 11394
rect 35756 11340 35924 11342
rect 35868 11330 35924 11340
rect 35644 10892 35924 10948
rect 35644 10724 35700 10734
rect 35532 10722 35700 10724
rect 35532 10670 35646 10722
rect 35698 10670 35700 10722
rect 35532 10668 35700 10670
rect 35644 10658 35700 10668
rect 35756 10612 35812 10622
rect 35756 10518 35812 10556
rect 35868 10388 35924 10892
rect 35532 10332 35924 10388
rect 35420 10276 35476 10286
rect 35420 8484 35476 10220
rect 35532 9826 35588 10332
rect 35980 10276 36036 12236
rect 36092 12124 36820 12180
rect 36092 11506 36148 12124
rect 36764 12066 36820 12124
rect 36764 12014 36766 12066
rect 36818 12014 36820 12066
rect 36316 11956 36372 11966
rect 36316 11862 36372 11900
rect 36428 11954 36484 11966
rect 36428 11902 36430 11954
rect 36482 11902 36484 11954
rect 36092 11454 36094 11506
rect 36146 11454 36148 11506
rect 36092 11442 36148 11454
rect 35532 9774 35534 9826
rect 35586 9774 35588 9826
rect 35532 9762 35588 9774
rect 35644 10220 36036 10276
rect 36316 10610 36372 10622
rect 36316 10558 36318 10610
rect 36370 10558 36372 10610
rect 35644 9716 35700 10220
rect 35868 10052 35924 10062
rect 36204 10052 36260 10062
rect 36316 10052 36372 10558
rect 35924 9996 36148 10052
rect 35868 9986 35924 9996
rect 36092 9938 36148 9996
rect 36204 10050 36372 10052
rect 36204 9998 36206 10050
rect 36258 9998 36372 10050
rect 36204 9996 36372 9998
rect 36204 9986 36260 9996
rect 36092 9886 36094 9938
rect 36146 9886 36148 9938
rect 36092 9874 36148 9886
rect 35420 8428 35588 8484
rect 35420 8258 35476 8270
rect 35420 8206 35422 8258
rect 35474 8206 35476 8258
rect 35420 8148 35476 8206
rect 35420 8082 35476 8092
rect 35532 7028 35588 8428
rect 35644 7474 35700 9660
rect 36316 9602 36372 9614
rect 36316 9550 36318 9602
rect 36370 9550 36372 9602
rect 36316 9380 36372 9550
rect 36316 9314 36372 9324
rect 35644 7422 35646 7474
rect 35698 7422 35700 7474
rect 35644 7410 35700 7422
rect 35868 7476 35924 7486
rect 35532 6972 35812 7028
rect 35420 6916 35476 6926
rect 35420 6822 35476 6860
rect 35644 6804 35700 6814
rect 35644 6710 35700 6748
rect 35532 6692 35588 6702
rect 35532 6598 35588 6636
rect 35308 6412 35700 6468
rect 35196 6402 35252 6412
rect 35252 6238 35476 6244
rect 35084 6188 35476 6238
rect 35084 6182 35308 6188
rect 34636 6078 34638 6130
rect 34690 6078 34692 6130
rect 34636 6066 34692 6078
rect 35084 5908 35140 5918
rect 34860 5852 35084 5908
rect 34860 5794 34916 5852
rect 35084 5842 35140 5852
rect 35420 5908 35476 6188
rect 35420 5842 35476 5852
rect 34860 5742 34862 5794
rect 34914 5742 34916 5794
rect 34860 5730 34916 5742
rect 34748 5682 34804 5694
rect 34748 5630 34750 5682
rect 34802 5630 34804 5682
rect 34748 5348 34804 5630
rect 34748 5282 34804 5292
rect 35084 5684 35140 5694
rect 34524 5182 34526 5234
rect 34578 5182 34580 5234
rect 34524 5170 34580 5182
rect 34188 5070 34190 5122
rect 34242 5070 34244 5122
rect 34188 5058 34244 5070
rect 34076 4844 34356 4900
rect 33740 4340 33796 4350
rect 33740 4246 33796 4284
rect 34188 4114 34244 4126
rect 34188 4062 34190 4114
rect 34242 4062 34244 4114
rect 32956 2930 33012 2940
rect 33628 4004 33684 4014
rect 32956 2772 33012 2782
rect 32956 2678 33012 2716
rect 33292 2548 33348 2558
rect 32508 2046 32510 2098
rect 32562 2046 32564 2098
rect 32508 2034 32564 2046
rect 32956 2100 33012 2110
rect 32060 1038 32062 1090
rect 32114 1038 32116 1090
rect 32060 1026 32116 1038
rect 32060 532 32116 542
rect 32060 112 32116 476
rect 32508 196 32564 206
rect 32508 112 32564 140
rect 32956 112 33012 2044
rect 33068 2098 33124 2110
rect 33068 2046 33070 2098
rect 33122 2046 33124 2098
rect 33068 1428 33124 2046
rect 33292 1986 33348 2492
rect 33628 2210 33684 3948
rect 33852 3780 33908 3790
rect 33852 3554 33908 3724
rect 33852 3502 33854 3554
rect 33906 3502 33908 3554
rect 33852 3490 33908 3502
rect 33740 2772 33796 2782
rect 33740 2678 33796 2716
rect 33628 2158 33630 2210
rect 33682 2158 33684 2210
rect 33628 2146 33684 2158
rect 33964 2324 34020 2334
rect 33292 1934 33294 1986
rect 33346 1934 33348 1986
rect 33292 1922 33348 1934
rect 33852 1876 33908 1886
rect 33292 1428 33348 1438
rect 33068 1426 33348 1428
rect 33068 1374 33294 1426
rect 33346 1374 33348 1426
rect 33068 1372 33348 1374
rect 33292 1362 33348 1372
rect 33740 980 33796 990
rect 33516 978 33796 980
rect 33516 926 33742 978
rect 33794 926 33796 978
rect 33516 924 33796 926
rect 33404 868 33460 878
rect 33404 112 33460 812
rect 33516 308 33572 924
rect 33740 914 33796 924
rect 33516 242 33572 252
rect 33852 112 33908 1820
rect 33964 1428 34020 2268
rect 34076 2098 34132 2110
rect 34076 2046 34078 2098
rect 34130 2046 34132 2098
rect 34076 1764 34132 2046
rect 34188 2100 34244 4062
rect 34300 3778 34356 4844
rect 34300 3726 34302 3778
rect 34354 3726 34356 3778
rect 34300 3714 34356 3726
rect 34524 4114 34580 4126
rect 34524 4062 34526 4114
rect 34578 4062 34580 4114
rect 34412 3668 34468 3678
rect 34300 2772 34356 2782
rect 34300 2678 34356 2716
rect 34412 2210 34468 3612
rect 34524 3388 34580 4062
rect 34524 3332 35028 3388
rect 34972 2658 35028 3332
rect 35084 2996 35140 5628
rect 35308 5348 35364 5358
rect 35308 4900 35364 5292
rect 35308 4834 35364 4844
rect 35532 5012 35588 5022
rect 35420 4116 35476 4126
rect 35084 2930 35140 2940
rect 35308 4114 35476 4116
rect 35308 4062 35422 4114
rect 35474 4062 35476 4114
rect 35308 4060 35476 4062
rect 35196 2772 35252 2782
rect 35196 2678 35252 2716
rect 34972 2606 34974 2658
rect 35026 2606 35028 2658
rect 34972 2594 35028 2606
rect 34412 2158 34414 2210
rect 34466 2158 34468 2210
rect 34412 2146 34468 2158
rect 34636 2546 34692 2558
rect 34636 2494 34638 2546
rect 34690 2494 34692 2546
rect 34188 2034 34244 2044
rect 34076 1698 34132 1708
rect 33964 1362 34020 1372
rect 34636 1204 34692 2494
rect 35084 2212 35140 2222
rect 35084 2118 35140 2156
rect 35308 2100 35364 4060
rect 35420 4050 35476 4060
rect 35532 3556 35588 4956
rect 35644 3668 35700 6412
rect 35756 4788 35812 6972
rect 35868 6916 35924 7420
rect 35868 6850 35924 6860
rect 36316 7028 36372 7038
rect 36316 6804 36372 6972
rect 36316 6738 36372 6748
rect 36428 6802 36484 11902
rect 36540 11956 36596 11966
rect 36540 11954 36708 11956
rect 36540 11902 36542 11954
rect 36594 11902 36708 11954
rect 36540 11900 36708 11902
rect 36540 11890 36596 11900
rect 36652 11732 36708 11900
rect 36652 11666 36708 11676
rect 36540 11620 36596 11630
rect 36540 11526 36596 11564
rect 36652 11396 36708 11406
rect 36652 11302 36708 11340
rect 36652 10836 36708 10846
rect 36764 10836 36820 12014
rect 36652 10834 36820 10836
rect 36652 10782 36654 10834
rect 36706 10782 36820 10834
rect 36652 10780 36820 10782
rect 36652 10770 36708 10780
rect 36764 10612 36820 10622
rect 36764 10518 36820 10556
rect 36652 10386 36708 10398
rect 36876 10388 36932 15092
rect 36652 10334 36654 10386
rect 36706 10334 36708 10386
rect 36428 6750 36430 6802
rect 36482 6750 36484 6802
rect 36428 6738 36484 6750
rect 36540 8818 36596 8830
rect 36540 8766 36542 8818
rect 36594 8766 36596 8818
rect 35980 6690 36036 6702
rect 35980 6638 35982 6690
rect 36034 6638 36036 6690
rect 35980 6132 36036 6638
rect 35980 6066 36036 6076
rect 36316 6466 36372 6478
rect 36316 6414 36318 6466
rect 36370 6414 36372 6466
rect 36316 5906 36372 6414
rect 36428 6356 36484 6366
rect 36428 6020 36484 6300
rect 36540 6244 36596 8766
rect 36652 7588 36708 10334
rect 36764 10332 36932 10388
rect 36988 15092 37156 15148
rect 36988 14530 37044 15092
rect 36988 14478 36990 14530
rect 37042 14478 37044 14530
rect 36764 9042 36820 10332
rect 36988 10276 37044 14478
rect 37100 14308 37156 14318
rect 37100 13524 37156 14252
rect 37100 13458 37156 13468
rect 37324 13300 37380 15820
rect 37324 13234 37380 13244
rect 37436 15652 37492 15662
rect 37324 12964 37380 12974
rect 37324 12870 37380 12908
rect 37100 11732 37156 11742
rect 37100 11394 37156 11676
rect 37100 11342 37102 11394
rect 37154 11342 37156 11394
rect 37100 10500 37156 11342
rect 37324 11172 37380 11182
rect 37100 10498 37268 10500
rect 37100 10446 37102 10498
rect 37154 10446 37268 10498
rect 37100 10444 37268 10446
rect 37100 10434 37156 10444
rect 36988 10220 37156 10276
rect 36764 8990 36766 9042
rect 36818 8990 36820 9042
rect 36764 8978 36820 8990
rect 36876 9828 36932 9838
rect 36764 8260 36820 8270
rect 36876 8260 36932 9772
rect 36764 8258 36932 8260
rect 36764 8206 36766 8258
rect 36818 8206 36932 8258
rect 36764 8204 36932 8206
rect 36764 8194 36820 8204
rect 36876 8148 36932 8204
rect 36876 8082 36932 8092
rect 36652 7532 36932 7588
rect 36540 6178 36596 6188
rect 36652 7028 36708 7038
rect 36428 5954 36484 5964
rect 36316 5854 36318 5906
rect 36370 5854 36372 5906
rect 36316 5842 36372 5854
rect 36540 5908 36596 5918
rect 36540 5814 36596 5852
rect 36652 5460 36708 6972
rect 36876 6692 36932 7532
rect 36876 6636 37044 6692
rect 36876 6130 36932 6142
rect 36876 6078 36878 6130
rect 36930 6078 36932 6130
rect 36764 5684 36820 5694
rect 36764 5590 36820 5628
rect 36540 5404 36708 5460
rect 36540 5012 36596 5404
rect 36876 5346 36932 6078
rect 36988 5906 37044 6636
rect 36988 5854 36990 5906
rect 37042 5854 37044 5906
rect 36988 5842 37044 5854
rect 36876 5294 36878 5346
rect 36930 5294 36932 5346
rect 36652 5236 36708 5246
rect 36652 5234 36820 5236
rect 36652 5182 36654 5234
rect 36706 5182 36820 5234
rect 36652 5180 36820 5182
rect 36652 5170 36708 5180
rect 36540 4956 36708 5012
rect 35756 4722 35812 4732
rect 35756 4340 35812 4350
rect 35756 4246 35812 4284
rect 36428 4340 36484 4350
rect 36428 4246 36484 4284
rect 36316 4226 36372 4238
rect 36316 4174 36318 4226
rect 36370 4174 36372 4226
rect 35644 3602 35700 3612
rect 35868 3668 35924 3678
rect 35868 3574 35924 3612
rect 36092 3668 36148 3678
rect 36316 3668 36372 4174
rect 36092 3666 36372 3668
rect 36092 3614 36094 3666
rect 36146 3614 36372 3666
rect 36092 3612 36372 3614
rect 36652 3780 36708 4956
rect 35532 3490 35588 3500
rect 35420 3444 35476 3482
rect 35420 3378 35476 3388
rect 36092 3444 36148 3612
rect 36092 3378 36148 3388
rect 36204 3444 36260 3454
rect 36540 3444 36596 3454
rect 36204 3442 36596 3444
rect 36204 3390 36206 3442
rect 36258 3390 36542 3442
rect 36594 3390 36596 3442
rect 36204 3388 36596 3390
rect 36204 3378 36260 3388
rect 36540 3378 36596 3388
rect 36652 3388 36708 3724
rect 36764 3778 36820 5180
rect 36876 4340 36932 5294
rect 37100 5346 37156 10220
rect 37212 10164 37268 10444
rect 37212 10098 37268 10108
rect 37324 10050 37380 11116
rect 37324 9998 37326 10050
rect 37378 9998 37380 10050
rect 37324 9986 37380 9998
rect 37212 9604 37268 9614
rect 37212 9154 37268 9548
rect 37212 9102 37214 9154
rect 37266 9102 37268 9154
rect 37212 9090 37268 9102
rect 37100 5294 37102 5346
rect 37154 5294 37156 5346
rect 37100 5282 37156 5294
rect 37212 8370 37268 8382
rect 37212 8318 37214 8370
rect 37266 8318 37268 8370
rect 37212 6916 37268 8318
rect 37324 6916 37380 6926
rect 37212 6860 37324 6916
rect 36988 5012 37044 5022
rect 36988 4918 37044 4956
rect 36876 4274 36932 4284
rect 37212 4228 37268 6860
rect 37324 6850 37380 6860
rect 37212 4162 37268 4172
rect 36764 3726 36766 3778
rect 36818 3726 36820 3778
rect 36764 3668 36820 3726
rect 36764 3602 36820 3612
rect 37212 3666 37268 3678
rect 37212 3614 37214 3666
rect 37266 3614 37268 3666
rect 36876 3444 36932 3482
rect 37212 3388 37268 3614
rect 36652 3332 36820 3388
rect 36876 3378 36932 3388
rect 36204 3220 36260 3230
rect 35756 2772 35812 2810
rect 35756 2706 35812 2716
rect 35644 2658 35700 2670
rect 35644 2606 35646 2658
rect 35698 2606 35700 2658
rect 35644 2212 35700 2606
rect 35644 2146 35700 2156
rect 35756 2548 35812 2558
rect 34636 1138 34692 1148
rect 35196 2044 35364 2100
rect 34748 1092 34804 1102
rect 34748 998 34804 1036
rect 34076 980 34132 990
rect 34076 886 34132 924
rect 34412 978 34468 990
rect 34412 926 34414 978
rect 34466 926 34468 978
rect 34412 756 34468 926
rect 34412 690 34468 700
rect 34748 420 34804 430
rect 34300 308 34356 318
rect 34300 112 34356 252
rect 34748 112 34804 364
rect 35196 112 35252 2044
rect 35308 1652 35364 1662
rect 35308 1090 35364 1596
rect 35532 1428 35588 1438
rect 35532 1202 35588 1372
rect 35532 1150 35534 1202
rect 35586 1150 35588 1202
rect 35532 1138 35588 1150
rect 35308 1038 35310 1090
rect 35362 1038 35364 1090
rect 35308 1026 35364 1038
rect 35756 756 35812 2492
rect 36204 2210 36260 3164
rect 36652 2772 36708 2782
rect 36652 2678 36708 2716
rect 36204 2158 36206 2210
rect 36258 2158 36260 2210
rect 36204 2146 36260 2158
rect 36316 2546 36372 2558
rect 36316 2494 36318 2546
rect 36370 2494 36372 2546
rect 36092 2100 36148 2110
rect 35644 700 35812 756
rect 35980 978 36036 990
rect 35980 926 35982 978
rect 36034 926 36036 978
rect 35644 112 35700 700
rect 35980 532 36036 926
rect 35980 466 36036 476
rect 36092 112 36148 2044
rect 36316 1876 36372 2494
rect 36316 1810 36372 1820
rect 36428 1988 36484 1998
rect 36316 1204 36372 1214
rect 36428 1204 36484 1932
rect 36764 1986 36820 3332
rect 37100 3332 37268 3388
rect 37436 3332 37492 15596
rect 37548 15540 37604 15550
rect 37548 15426 37604 15484
rect 37548 15374 37550 15426
rect 37602 15374 37604 15426
rect 37548 15362 37604 15374
rect 37548 13860 37604 13870
rect 37548 13766 37604 13804
rect 37548 13300 37604 13310
rect 37548 11956 37604 13244
rect 37548 11506 37604 11900
rect 37660 11844 37716 19180
rect 37996 19012 38052 19022
rect 37996 18450 38052 18956
rect 37996 18398 37998 18450
rect 38050 18398 38052 18450
rect 37996 18386 38052 18398
rect 37996 17666 38052 17678
rect 37996 17614 37998 17666
rect 38050 17614 38052 17666
rect 37996 17108 38052 17614
rect 38108 17444 38164 21308
rect 38108 17378 38164 17388
rect 38108 17108 38164 17118
rect 37996 17106 38164 17108
rect 37996 17054 38110 17106
rect 38162 17054 38164 17106
rect 37996 17052 38164 17054
rect 38108 17042 38164 17052
rect 37772 16212 37828 16222
rect 37772 13186 37828 16156
rect 37884 16100 37940 16110
rect 37884 15314 37940 16044
rect 37884 15262 37886 15314
rect 37938 15262 37940 15314
rect 37884 15250 37940 15262
rect 37996 15540 38052 15550
rect 37996 15148 38052 15484
rect 38220 15316 38276 21868
rect 38332 21700 38388 23212
rect 38444 21924 38500 23772
rect 38556 23492 38612 26572
rect 38780 25732 38836 27582
rect 38892 27300 38948 27694
rect 38892 27234 38948 27244
rect 39116 27076 39172 27916
rect 39228 27858 39284 29934
rect 39340 29092 39396 30156
rect 39340 29026 39396 29036
rect 39452 28868 39508 35252
rect 39900 35196 40068 35252
rect 39564 34130 39620 34142
rect 39564 34078 39566 34130
rect 39618 34078 39620 34130
rect 39564 33570 39620 34078
rect 39564 33518 39566 33570
rect 39618 33518 39620 33570
rect 39564 33506 39620 33518
rect 39676 34020 39732 34030
rect 39676 33348 39732 33964
rect 39228 27806 39230 27858
rect 39282 27806 39284 27858
rect 39228 27794 39284 27806
rect 39340 28812 39508 28868
rect 39564 33292 39732 33348
rect 39340 27860 39396 28812
rect 39452 28642 39508 28654
rect 39452 28590 39454 28642
rect 39506 28590 39508 28642
rect 39452 28084 39508 28590
rect 39452 28018 39508 28028
rect 39340 27804 39508 27860
rect 39452 27412 39508 27804
rect 39564 27524 39620 33292
rect 39788 29426 39844 29438
rect 39788 29374 39790 29426
rect 39842 29374 39844 29426
rect 39788 28644 39844 29374
rect 39788 28578 39844 28588
rect 39676 28532 39732 28542
rect 39676 27858 39732 28476
rect 39788 28084 39844 28094
rect 39788 27970 39844 28028
rect 39788 27918 39790 27970
rect 39842 27918 39844 27970
rect 39788 27906 39844 27918
rect 39676 27806 39678 27858
rect 39730 27806 39732 27858
rect 39676 27794 39732 27806
rect 39564 27468 39844 27524
rect 39452 27356 39732 27412
rect 38780 25666 38836 25676
rect 39004 27074 39172 27076
rect 39004 27022 39118 27074
rect 39170 27022 39172 27074
rect 39004 27020 39172 27022
rect 38556 23426 38612 23436
rect 38668 25282 38724 25294
rect 38668 25230 38670 25282
rect 38722 25230 38724 25282
rect 38668 23154 38724 25230
rect 38892 24610 38948 24622
rect 38892 24558 38894 24610
rect 38946 24558 38948 24610
rect 38892 24388 38948 24558
rect 39004 24610 39060 27020
rect 39116 27010 39172 27020
rect 39564 27076 39620 27086
rect 39676 27076 39732 27356
rect 39788 27188 39844 27468
rect 39900 27300 39956 35196
rect 40124 32452 40180 37324
rect 40348 37266 40404 37774
rect 40348 37214 40350 37266
rect 40402 37214 40404 37266
rect 40348 37202 40404 37214
rect 40236 35700 40292 35710
rect 40236 34018 40292 35644
rect 40348 34690 40404 34702
rect 40348 34638 40350 34690
rect 40402 34638 40404 34690
rect 40348 34468 40404 34638
rect 40348 34402 40404 34412
rect 40348 34132 40404 34142
rect 40348 34038 40404 34076
rect 40236 33966 40238 34018
rect 40290 33966 40292 34018
rect 40236 33954 40292 33966
rect 40012 32396 40180 32452
rect 40236 33796 40292 33806
rect 40012 28084 40068 32396
rect 40236 31444 40292 33740
rect 40460 33460 40516 43036
rect 40684 42980 40740 43262
rect 40572 42924 40740 42980
rect 40572 42308 40628 42924
rect 40796 42868 40852 43374
rect 40908 43426 40964 43438
rect 40908 43374 40910 43426
rect 40962 43374 40964 43426
rect 40908 43316 40964 43374
rect 40908 43250 40964 43260
rect 40572 42242 40628 42252
rect 40684 42812 40852 42868
rect 40908 42868 40964 42878
rect 40572 41972 40628 41982
rect 40572 41188 40628 41916
rect 40684 41860 40740 42812
rect 40796 42644 40852 42654
rect 40908 42644 40964 42812
rect 40796 42642 40964 42644
rect 40796 42590 40798 42642
rect 40850 42590 40964 42642
rect 40796 42588 40964 42590
rect 40796 42578 40852 42588
rect 40908 42420 40964 42588
rect 40908 42354 40964 42364
rect 40684 41794 40740 41804
rect 41020 42308 41076 43708
rect 40796 41746 40852 41758
rect 40796 41694 40798 41746
rect 40850 41694 40852 41746
rect 40572 41122 40628 41132
rect 40684 41636 40740 41646
rect 40572 40964 40628 40974
rect 40572 39618 40628 40908
rect 40572 39566 40574 39618
rect 40626 39566 40628 39618
rect 40572 39554 40628 39566
rect 40572 36708 40628 36718
rect 40572 35698 40628 36652
rect 40572 35646 40574 35698
rect 40626 35646 40628 35698
rect 40572 35634 40628 35646
rect 40684 34692 40740 41580
rect 40796 40402 40852 41694
rect 40908 41412 40964 41422
rect 41020 41412 41076 42252
rect 41132 41748 41188 44382
rect 41244 43876 41300 44604
rect 41244 43810 41300 43820
rect 41356 43764 41412 45052
rect 41356 43698 41412 43708
rect 41244 43650 41300 43662
rect 41244 43598 41246 43650
rect 41298 43598 41300 43650
rect 41244 43428 41300 43598
rect 41244 43362 41300 43372
rect 41468 43092 41524 48188
rect 41580 44436 41636 48860
rect 41916 48580 41972 48972
rect 41916 48514 41972 48524
rect 42028 48804 42084 48814
rect 42364 48804 42420 48972
rect 42476 48962 42532 48972
rect 42028 48802 42420 48804
rect 42028 48750 42030 48802
rect 42082 48750 42420 48802
rect 42028 48748 42420 48750
rect 42476 48802 42532 48814
rect 42476 48750 42478 48802
rect 42530 48750 42532 48802
rect 41804 48130 41860 48142
rect 41804 48078 41806 48130
rect 41858 48078 41860 48130
rect 41692 47570 41748 47582
rect 41692 47518 41694 47570
rect 41746 47518 41748 47570
rect 41692 46340 41748 47518
rect 41692 46274 41748 46284
rect 41804 46788 41860 48078
rect 42028 47570 42084 48748
rect 42028 47518 42030 47570
rect 42082 47518 42084 47570
rect 42028 47506 42084 47518
rect 42252 48020 42308 48030
rect 42140 47346 42196 47358
rect 42140 47294 42142 47346
rect 42194 47294 42196 47346
rect 42140 47124 42196 47294
rect 42140 47058 42196 47068
rect 42252 47012 42308 47964
rect 42364 47458 42420 47470
rect 42364 47406 42366 47458
rect 42418 47406 42420 47458
rect 42364 47236 42420 47406
rect 42476 47458 42532 48750
rect 42476 47406 42478 47458
rect 42530 47406 42532 47458
rect 42476 47394 42532 47406
rect 42588 47236 42644 50876
rect 42364 47180 42644 47236
rect 42252 46946 42308 46956
rect 42700 47012 42756 50988
rect 42812 50820 42868 50830
rect 42812 50726 42868 50764
rect 42924 50148 42980 50158
rect 42812 48804 42868 48814
rect 42812 48710 42868 48748
rect 42700 46946 42756 46956
rect 42812 48580 42868 48590
rect 41804 46004 41860 46732
rect 42700 46788 42756 46798
rect 42700 46694 42756 46732
rect 42812 46676 42868 48524
rect 42924 48244 42980 50092
rect 43036 48916 43092 51436
rect 43036 48850 43092 48860
rect 43148 48914 43204 51436
rect 43260 50596 43316 50606
rect 43260 49028 43316 50540
rect 43372 50372 43428 52332
rect 43596 52322 43652 52332
rect 43596 52164 43652 52174
rect 43484 52052 43540 52062
rect 43484 51602 43540 51996
rect 43484 51550 43486 51602
rect 43538 51550 43540 51602
rect 43484 51538 43540 51550
rect 43596 51154 43652 52108
rect 44268 52052 44324 52444
rect 44828 52388 44884 52668
rect 44604 52332 44884 52388
rect 44268 51996 44436 52052
rect 44380 51940 44436 51996
rect 44380 51874 44436 51884
rect 44492 51828 44548 51838
rect 43804 51772 44068 51782
rect 43860 51716 43908 51772
rect 43964 51716 44012 51772
rect 43804 51706 44068 51716
rect 44492 51380 44548 51772
rect 44604 51604 44660 52332
rect 44940 51828 44996 53788
rect 45052 53060 45108 54238
rect 45164 54180 45220 54190
rect 45164 53508 45220 54124
rect 45500 53842 45556 53854
rect 45500 53790 45502 53842
rect 45554 53790 45556 53842
rect 45276 53732 45332 53742
rect 45276 53638 45332 53676
rect 45164 53442 45220 53452
rect 45052 52994 45108 53004
rect 45276 53396 45332 53406
rect 45052 52836 45108 52846
rect 45052 52742 45108 52780
rect 45276 52834 45332 53340
rect 45500 53396 45556 53790
rect 45500 53330 45556 53340
rect 45276 52782 45278 52834
rect 45330 52782 45332 52834
rect 45276 52770 45332 52782
rect 45164 52722 45220 52734
rect 45164 52670 45166 52722
rect 45218 52670 45220 52722
rect 45164 52052 45220 52670
rect 45388 52164 45444 52174
rect 45388 52070 45444 52108
rect 45164 51986 45220 51996
rect 45612 51940 45668 54462
rect 46172 54516 46228 54526
rect 46172 54422 46228 54460
rect 46284 54068 46340 56476
rect 46396 55524 46452 57344
rect 46396 55458 46452 55468
rect 46620 57092 46676 57102
rect 46508 55412 46564 55422
rect 46396 55300 46452 55310
rect 46396 55206 46452 55244
rect 46508 54516 46564 55356
rect 46620 55300 46676 57036
rect 46732 55858 46788 55870
rect 46732 55806 46734 55858
rect 46786 55806 46788 55858
rect 46732 55636 46788 55806
rect 46732 55570 46788 55580
rect 46844 55524 46900 57344
rect 47068 56644 47124 56654
rect 47068 55970 47124 56588
rect 47068 55918 47070 55970
rect 47122 55918 47124 55970
rect 47068 55906 47124 55918
rect 46844 55458 46900 55468
rect 47292 55524 47348 57344
rect 47740 56420 47796 57344
rect 47740 56364 47908 56420
rect 47740 56196 47796 56206
rect 47740 55970 47796 56140
rect 47740 55918 47742 55970
rect 47794 55918 47796 55970
rect 47740 55906 47796 55918
rect 47404 55860 47460 55870
rect 47404 55766 47460 55804
rect 47292 55458 47348 55468
rect 47628 55636 47684 55646
rect 46620 55234 46676 55244
rect 46732 55410 46788 55422
rect 46732 55358 46734 55410
rect 46786 55358 46788 55410
rect 46732 55076 46788 55358
rect 46732 55010 46788 55020
rect 46956 55298 47012 55310
rect 46956 55246 46958 55298
rect 47010 55246 47012 55298
rect 46508 54450 46564 54460
rect 46284 54002 46340 54012
rect 46172 53842 46228 53854
rect 46172 53790 46174 53842
rect 46226 53790 46228 53842
rect 45948 53730 46004 53742
rect 45948 53678 45950 53730
rect 46002 53678 46004 53730
rect 45948 53508 46004 53678
rect 45948 53442 46004 53452
rect 46172 53172 46228 53790
rect 46508 53842 46564 53854
rect 46508 53790 46510 53842
rect 46562 53790 46564 53842
rect 46508 53620 46564 53790
rect 46508 53554 46564 53564
rect 46732 53730 46788 53742
rect 46732 53678 46734 53730
rect 46786 53678 46788 53730
rect 46172 53106 46228 53116
rect 44940 51762 44996 51772
rect 45388 51884 45668 51940
rect 46060 52946 46116 52958
rect 46060 52894 46062 52946
rect 46114 52894 46116 52946
rect 44604 51538 44660 51548
rect 44492 51286 44548 51324
rect 44716 51380 44772 51390
rect 44940 51380 44996 51390
rect 44716 51378 44884 51380
rect 44716 51326 44718 51378
rect 44770 51326 44884 51378
rect 44716 51324 44884 51326
rect 44716 51314 44772 51324
rect 43596 51102 43598 51154
rect 43650 51102 43652 51154
rect 43596 51090 43652 51102
rect 44268 51268 44324 51278
rect 44268 51154 44324 51212
rect 44268 51102 44270 51154
rect 44322 51102 44324 51154
rect 44268 50932 44324 51102
rect 44380 51156 44436 51194
rect 44380 51090 44436 51100
rect 44464 50988 44728 50998
rect 44520 50932 44568 50988
rect 44624 50932 44672 50988
rect 44464 50922 44728 50932
rect 44268 50866 44324 50876
rect 43932 50708 43988 50718
rect 43932 50614 43988 50652
rect 44380 50484 44436 50494
rect 44828 50428 44884 51324
rect 44940 51286 44996 51324
rect 45276 51378 45332 51390
rect 45276 51326 45278 51378
rect 45330 51326 45332 51378
rect 45276 51268 45332 51326
rect 45276 51202 45332 51212
rect 45164 51156 45220 51166
rect 44380 50390 44436 50428
rect 43372 50306 43428 50316
rect 44604 50372 44884 50428
rect 44940 50932 44996 50942
rect 44940 50482 44996 50876
rect 45052 50708 45108 50718
rect 45052 50614 45108 50652
rect 44940 50430 44942 50482
rect 44994 50430 44996 50482
rect 44940 50418 44996 50430
rect 43804 50204 44068 50214
rect 43860 50148 43908 50204
rect 43964 50148 44012 50204
rect 43804 50138 44068 50148
rect 44492 50148 44548 50158
rect 43372 50036 43428 50046
rect 43372 49942 43428 49980
rect 44492 49924 44548 50092
rect 43260 48962 43316 48972
rect 43820 49868 44548 49924
rect 43148 48862 43150 48914
rect 43202 48862 43204 48914
rect 43148 48850 43204 48862
rect 43820 48804 43876 49868
rect 44492 49810 44548 49868
rect 44604 49922 44660 50372
rect 45052 50148 45108 50158
rect 44604 49870 44606 49922
rect 44658 49870 44660 49922
rect 44604 49858 44660 49870
rect 44828 49924 44884 49934
rect 44492 49758 44494 49810
rect 44546 49758 44548 49810
rect 44492 49746 44548 49758
rect 44716 49812 44772 49822
rect 44716 49718 44772 49756
rect 44156 49700 44212 49710
rect 43596 48748 43876 48804
rect 43932 49698 44212 49700
rect 43932 49646 44158 49698
rect 44210 49646 44212 49698
rect 43932 49644 44212 49646
rect 43932 48804 43988 49644
rect 44156 49634 44212 49644
rect 44268 49476 44324 49486
rect 43036 48580 43092 48590
rect 43036 48466 43092 48524
rect 43596 48580 43652 48748
rect 43932 48738 43988 48748
rect 44156 49364 44212 49374
rect 44156 48804 44212 49308
rect 44268 49252 44324 49420
rect 44464 49420 44728 49430
rect 44520 49364 44568 49420
rect 44624 49364 44672 49420
rect 44464 49354 44728 49364
rect 44828 49364 44884 49868
rect 45052 49924 45108 50092
rect 45052 49858 45108 49868
rect 44828 49298 44884 49308
rect 44940 49476 44996 49486
rect 44268 49196 44660 49252
rect 44604 48916 44660 49196
rect 44604 48850 44660 48860
rect 44156 48738 44212 48748
rect 43804 48636 44068 48646
rect 43860 48580 43908 48636
rect 43964 48580 44012 48636
rect 44940 48580 44996 49420
rect 45164 49140 45220 51100
rect 45276 50596 45332 50606
rect 45276 50502 45332 50540
rect 45276 49812 45332 49822
rect 45276 49718 45332 49756
rect 45276 49140 45332 49150
rect 45164 49138 45332 49140
rect 45164 49086 45278 49138
rect 45330 49086 45332 49138
rect 45164 49084 45332 49086
rect 45276 49074 45332 49084
rect 45052 49028 45108 49038
rect 45052 48692 45108 48972
rect 45052 48626 45108 48636
rect 43804 48570 44068 48580
rect 43596 48514 43652 48524
rect 44156 48524 44996 48580
rect 44156 48468 44212 48524
rect 43036 48414 43038 48466
rect 43090 48414 43092 48466
rect 43036 48402 43092 48414
rect 43708 48412 44212 48468
rect 43596 48244 43652 48254
rect 42924 48188 43092 48244
rect 42812 46610 42868 46620
rect 42924 47348 42980 47358
rect 42924 46786 42980 47292
rect 42924 46734 42926 46786
rect 42978 46734 42980 46786
rect 42252 46452 42308 46462
rect 42252 46358 42308 46396
rect 42924 46452 42980 46734
rect 43036 46788 43092 48188
rect 43372 48242 43652 48244
rect 43372 48190 43598 48242
rect 43650 48190 43652 48242
rect 43372 48188 43652 48190
rect 43372 47908 43428 48188
rect 43596 48178 43652 48188
rect 43484 48020 43540 48030
rect 43484 47926 43540 47964
rect 43708 48020 43764 48412
rect 44380 48244 44436 48254
rect 44940 48244 44996 48254
rect 45276 48244 45332 48254
rect 44380 48242 44884 48244
rect 44380 48190 44382 48242
rect 44434 48190 44884 48242
rect 44380 48188 44884 48190
rect 44380 48178 44436 48188
rect 44828 48132 44884 48188
rect 44940 48242 45108 48244
rect 44940 48190 44942 48242
rect 44994 48190 45108 48242
rect 44940 48188 45108 48190
rect 44940 48178 44996 48188
rect 44828 48066 44884 48076
rect 43708 47954 43764 47964
rect 44044 48018 44100 48030
rect 44268 48020 44324 48030
rect 44044 47966 44046 48018
rect 44098 47966 44100 48018
rect 43372 47842 43428 47852
rect 44044 47796 44100 47966
rect 43596 47740 44100 47796
rect 44156 48018 44324 48020
rect 44156 47966 44270 48018
rect 44322 47966 44324 48018
rect 44156 47964 44324 47966
rect 43596 47460 43652 47740
rect 43596 47404 43764 47460
rect 43148 47236 43204 47246
rect 43708 47236 43764 47404
rect 44156 47348 44212 47964
rect 44268 47954 44324 47964
rect 44604 48020 44660 48030
rect 44940 48020 44996 48030
rect 44660 47964 44884 47998
rect 44604 47942 44884 47964
rect 44828 47908 44884 47942
rect 44464 47852 44728 47862
rect 44520 47796 44568 47852
rect 44624 47796 44672 47852
rect 44828 47842 44884 47852
rect 44464 47786 44728 47796
rect 44268 47684 44324 47722
rect 44940 47684 44996 47964
rect 45052 47796 45108 48188
rect 45388 48244 45444 51884
rect 45724 51380 45780 51390
rect 45724 51286 45780 51324
rect 45612 51154 45668 51166
rect 45612 51102 45614 51154
rect 45666 51102 45668 51154
rect 45500 51044 45556 51054
rect 45500 50820 45556 50988
rect 45500 50754 45556 50764
rect 45500 50148 45556 50158
rect 45500 49252 45556 50092
rect 45612 50036 45668 51102
rect 45836 51156 45892 51166
rect 45836 51062 45892 51100
rect 45836 50484 45892 50494
rect 45836 50482 46004 50484
rect 45836 50430 45838 50482
rect 45890 50430 46004 50482
rect 45836 50428 46004 50430
rect 45836 50418 45892 50428
rect 45612 49970 45668 49980
rect 45836 50260 45892 50270
rect 45500 49186 45556 49196
rect 45724 49586 45780 49598
rect 45724 49534 45726 49586
rect 45778 49534 45780 49586
rect 45612 49028 45668 49038
rect 45388 48188 45556 48244
rect 45276 48130 45332 48188
rect 45276 48078 45278 48130
rect 45330 48078 45332 48130
rect 45276 48066 45332 48078
rect 45052 47730 45108 47740
rect 44268 47618 44324 47628
rect 44492 47628 44996 47684
rect 44492 47460 44548 47628
rect 44492 47394 44548 47404
rect 44828 47458 44884 47470
rect 44828 47406 44830 47458
rect 44882 47406 44884 47458
rect 44156 47292 44436 47348
rect 43148 47234 43652 47236
rect 43148 47182 43150 47234
rect 43202 47182 43652 47234
rect 43148 47180 43652 47182
rect 43148 47170 43204 47180
rect 43036 46722 43092 46732
rect 43148 46676 43204 46686
rect 43148 46674 43540 46676
rect 43148 46622 43150 46674
rect 43202 46622 43540 46674
rect 43148 46620 43540 46622
rect 43148 46610 43204 46620
rect 42924 46386 42980 46396
rect 43260 46450 43316 46462
rect 43260 46398 43262 46450
rect 43314 46398 43316 46450
rect 43260 46228 43316 46398
rect 42588 46172 43316 46228
rect 43372 46450 43428 46462
rect 43372 46398 43374 46450
rect 43426 46398 43428 46450
rect 43372 46228 43428 46398
rect 42588 46114 42644 46172
rect 42588 46062 42590 46114
rect 42642 46062 42644 46114
rect 42588 46050 42644 46062
rect 41804 45938 41860 45948
rect 43372 46004 43428 46172
rect 43372 45938 43428 45948
rect 41580 44370 41636 44380
rect 41692 45892 41748 45902
rect 41692 43650 41748 45836
rect 42028 45724 42644 45780
rect 42028 45666 42084 45724
rect 42028 45614 42030 45666
rect 42082 45614 42084 45666
rect 42028 45602 42084 45614
rect 42588 45330 42644 45724
rect 42588 45278 42590 45330
rect 42642 45278 42644 45330
rect 42588 45266 42644 45278
rect 42700 45778 42756 45790
rect 42700 45726 42702 45778
rect 42754 45726 42756 45778
rect 41916 45108 41972 45118
rect 42140 45108 42196 45118
rect 41972 45106 42196 45108
rect 41972 45054 42142 45106
rect 42194 45054 42196 45106
rect 41972 45052 42196 45054
rect 41916 45042 41972 45052
rect 42140 45042 42196 45052
rect 42252 45108 42308 45118
rect 42140 44772 42196 44782
rect 42140 44436 42196 44716
rect 42140 44370 42196 44380
rect 41692 43598 41694 43650
rect 41746 43598 41748 43650
rect 41692 43586 41748 43598
rect 42252 43538 42308 45052
rect 42588 44772 42644 44782
rect 42588 44660 42644 44716
rect 42364 44604 42644 44660
rect 42364 44546 42420 44604
rect 42364 44494 42366 44546
rect 42418 44494 42420 44546
rect 42700 44578 42756 45726
rect 43372 45778 43428 45790
rect 43372 45726 43374 45778
rect 43426 45726 43428 45778
rect 42812 45668 42868 45678
rect 42812 45666 43204 45668
rect 42812 45614 42814 45666
rect 42866 45614 43204 45666
rect 42812 45612 43204 45614
rect 42812 45602 42868 45612
rect 43036 45332 43092 45342
rect 42924 45108 42980 45118
rect 42924 45014 42980 45052
rect 43036 45106 43092 45276
rect 43148 45218 43204 45612
rect 43372 45444 43428 45726
rect 43372 45378 43428 45388
rect 43148 45166 43150 45218
rect 43202 45166 43204 45218
rect 43148 45154 43204 45166
rect 43036 45054 43038 45106
rect 43090 45054 43092 45106
rect 43036 45042 43092 45054
rect 43372 45108 43428 45118
rect 43260 44882 43316 44894
rect 43260 44830 43262 44882
rect 43314 44830 43316 44882
rect 42700 44522 43204 44578
rect 42364 44482 42420 44494
rect 42924 44436 42980 44446
rect 42924 44342 42980 44380
rect 42812 44100 42868 44110
rect 42812 44006 42868 44044
rect 42252 43486 42254 43538
rect 42306 43486 42308 43538
rect 42252 43474 42308 43486
rect 42924 43876 42980 43886
rect 41916 43428 41972 43438
rect 41356 43036 41524 43092
rect 41580 43314 41636 43326
rect 41580 43262 41582 43314
rect 41634 43262 41636 43314
rect 41244 42868 41300 42878
rect 41244 42774 41300 42812
rect 41132 41682 41188 41692
rect 40908 41410 41076 41412
rect 40908 41358 40910 41410
rect 40962 41358 41076 41410
rect 40908 41356 41076 41358
rect 40908 41346 40964 41356
rect 41244 40404 41300 40414
rect 40796 40350 40798 40402
rect 40850 40350 40852 40402
rect 40796 40338 40852 40350
rect 41132 40402 41300 40404
rect 41132 40350 41246 40402
rect 41298 40350 41300 40402
rect 41132 40348 41300 40350
rect 41020 40068 41076 40078
rect 41020 39618 41076 40012
rect 41020 39566 41022 39618
rect 41074 39566 41076 39618
rect 41020 39554 41076 39566
rect 41132 39508 41188 40348
rect 41244 40338 41300 40348
rect 41244 40068 41300 40078
rect 41244 39842 41300 40012
rect 41244 39790 41246 39842
rect 41298 39790 41300 39842
rect 41244 39778 41300 39790
rect 40796 38948 40852 38958
rect 40796 37716 40852 38892
rect 41132 38668 41188 39452
rect 40796 35140 40852 37660
rect 41020 38612 41188 38668
rect 41356 39284 41412 43036
rect 41468 42868 41524 42878
rect 41468 40404 41524 42812
rect 41580 42084 41636 43262
rect 41804 43316 41860 43354
rect 41916 43334 41972 43372
rect 42476 43428 42532 43438
rect 41804 43250 41860 43260
rect 41580 42018 41636 42028
rect 42252 42756 42308 42766
rect 42252 42084 42308 42700
rect 42252 41990 42308 42028
rect 42364 42530 42420 42542
rect 42364 42478 42366 42530
rect 42418 42478 42420 42530
rect 41468 40338 41524 40348
rect 41580 41858 41636 41870
rect 41580 41806 41582 41858
rect 41634 41806 41636 41858
rect 40908 37266 40964 37278
rect 40908 37214 40910 37266
rect 40962 37214 40964 37266
rect 40908 35700 40964 37214
rect 40908 35606 40964 35644
rect 40796 35074 40852 35084
rect 40684 34626 40740 34636
rect 40684 34468 40740 34478
rect 40460 33404 40628 33460
rect 40460 33234 40516 33246
rect 40460 33182 40462 33234
rect 40514 33182 40516 33234
rect 40348 33012 40404 33022
rect 40348 32674 40404 32956
rect 40348 32622 40350 32674
rect 40402 32622 40404 32674
rect 40348 32610 40404 32622
rect 40236 31378 40292 31388
rect 40460 30996 40516 33182
rect 40572 32340 40628 33404
rect 40684 32562 40740 34412
rect 40796 34244 40852 34254
rect 40796 34130 40852 34188
rect 40796 34078 40798 34130
rect 40850 34078 40852 34130
rect 40796 34066 40852 34078
rect 40908 34132 40964 34142
rect 40908 33570 40964 34076
rect 40908 33518 40910 33570
rect 40962 33518 40964 33570
rect 40908 33506 40964 33518
rect 40684 32510 40686 32562
rect 40738 32510 40740 32562
rect 40684 32498 40740 32510
rect 40796 33458 40852 33470
rect 40796 33406 40798 33458
rect 40850 33406 40852 33458
rect 40572 32284 40740 32340
rect 40460 30930 40516 30940
rect 40348 30772 40404 30782
rect 40348 30770 40628 30772
rect 40348 30718 40350 30770
rect 40402 30718 40628 30770
rect 40348 30716 40628 30718
rect 40348 30706 40404 30716
rect 40236 30212 40292 30222
rect 40236 30118 40292 30156
rect 40572 30210 40628 30716
rect 40572 30158 40574 30210
rect 40626 30158 40628 30210
rect 40572 30146 40628 30158
rect 40460 29764 40516 29774
rect 40012 28018 40068 28028
rect 40236 29428 40292 29438
rect 40012 27860 40068 27870
rect 40012 27766 40068 27804
rect 40124 27858 40180 27870
rect 40124 27806 40126 27858
rect 40178 27806 40180 27858
rect 40124 27412 40180 27806
rect 40236 27860 40292 29372
rect 40460 29426 40516 29708
rect 40460 29374 40462 29426
rect 40514 29374 40516 29426
rect 40236 27794 40292 27804
rect 40348 29316 40404 29326
rect 40124 27356 40292 27412
rect 40236 27300 40292 27356
rect 39900 27244 40180 27300
rect 39788 27132 40068 27188
rect 39676 27020 39844 27076
rect 39228 26964 39284 26974
rect 39340 26964 39396 26974
rect 39284 26962 39396 26964
rect 39284 26910 39342 26962
rect 39394 26910 39396 26962
rect 39284 26908 39396 26910
rect 39116 25508 39172 25518
rect 39116 25414 39172 25452
rect 39228 25172 39284 26908
rect 39340 26898 39396 26908
rect 39452 26740 39508 26750
rect 39452 26068 39508 26684
rect 39340 26066 39508 26068
rect 39340 26014 39454 26066
rect 39506 26014 39508 26066
rect 39340 26012 39508 26014
rect 39340 25508 39396 26012
rect 39452 26002 39508 26012
rect 39340 25442 39396 25452
rect 39340 25284 39396 25294
rect 39340 25190 39396 25228
rect 39004 24558 39006 24610
rect 39058 24558 39060 24610
rect 39004 24546 39060 24558
rect 39116 25116 39284 25172
rect 39116 24388 39172 25116
rect 39564 24836 39620 27020
rect 39676 26852 39732 26862
rect 39676 26758 39732 26796
rect 39676 25844 39732 25854
rect 39676 25730 39732 25788
rect 39676 25678 39678 25730
rect 39730 25678 39732 25730
rect 39676 25666 39732 25678
rect 39788 25396 39844 27020
rect 39228 24780 39620 24836
rect 39676 25060 39732 25070
rect 39676 24834 39732 25004
rect 39676 24782 39678 24834
rect 39730 24782 39732 24834
rect 39228 24722 39284 24780
rect 39676 24770 39732 24782
rect 39228 24670 39230 24722
rect 39282 24670 39284 24722
rect 39228 24658 39284 24670
rect 39788 24612 39844 25340
rect 38892 24332 39172 24388
rect 39564 24556 39844 24612
rect 39900 26964 39956 26974
rect 39340 23940 39396 23950
rect 39116 23492 39172 23502
rect 39004 23156 39060 23166
rect 38668 23102 38670 23154
rect 38722 23102 38724 23154
rect 38668 23090 38724 23102
rect 38780 23154 39060 23156
rect 38780 23102 39006 23154
rect 39058 23102 39060 23154
rect 38780 23100 39060 23102
rect 38444 21858 38500 21868
rect 38668 21924 38724 21934
rect 38332 21644 38444 21700
rect 38388 21476 38444 21644
rect 38332 21420 38444 21476
rect 38668 21586 38724 21868
rect 38668 21534 38670 21586
rect 38722 21534 38724 21586
rect 38332 16322 38388 21420
rect 38556 21364 38612 21374
rect 38332 16270 38334 16322
rect 38386 16270 38388 16322
rect 38332 16212 38388 16270
rect 38332 16146 38388 16156
rect 38444 21362 38612 21364
rect 38444 21310 38558 21362
rect 38610 21310 38612 21362
rect 38444 21308 38612 21310
rect 38444 15652 38500 21308
rect 38556 21298 38612 21308
rect 38668 21178 38724 21534
rect 38556 21122 38724 21178
rect 38556 20356 38612 21122
rect 38556 20290 38612 20300
rect 38668 21028 38724 21038
rect 38668 20242 38724 20972
rect 38668 20190 38670 20242
rect 38722 20190 38724 20242
rect 38668 20178 38724 20190
rect 38556 19796 38612 19806
rect 38556 18676 38612 19740
rect 38668 19012 38724 19022
rect 38668 18918 38724 18956
rect 38556 18620 38724 18676
rect 38220 15250 38276 15260
rect 38332 15596 38500 15652
rect 38556 18450 38612 18462
rect 38556 18398 38558 18450
rect 38610 18398 38612 18450
rect 38556 17666 38612 18398
rect 38556 17614 38558 17666
rect 38610 17614 38612 17666
rect 37772 13134 37774 13186
rect 37826 13134 37828 13186
rect 37772 13122 37828 13134
rect 37884 15092 38052 15148
rect 37660 11778 37716 11788
rect 37548 11454 37550 11506
rect 37602 11454 37604 11506
rect 37548 11442 37604 11454
rect 37548 10164 37604 10174
rect 37548 7140 37604 10108
rect 37660 9042 37716 9054
rect 37660 8990 37662 9042
rect 37714 8990 37716 9042
rect 37660 8372 37716 8990
rect 37660 8306 37716 8316
rect 37548 7074 37604 7084
rect 37772 8260 37828 8270
rect 37548 5682 37604 5694
rect 37548 5630 37550 5682
rect 37602 5630 37604 5682
rect 37548 5124 37604 5630
rect 37548 5058 37604 5068
rect 37548 4340 37604 4350
rect 37548 3778 37604 4284
rect 37548 3726 37550 3778
rect 37602 3726 37604 3778
rect 37548 3714 37604 3726
rect 36988 2548 37044 2558
rect 36988 2454 37044 2492
rect 36764 1934 36766 1986
rect 36818 1934 36820 1986
rect 36764 1922 36820 1934
rect 36316 1202 36484 1204
rect 36316 1150 36318 1202
rect 36370 1150 36484 1202
rect 36316 1148 36484 1150
rect 36876 1204 36932 1214
rect 36316 1138 36372 1148
rect 36876 1110 36932 1148
rect 36652 980 36708 990
rect 36652 978 36820 980
rect 36652 926 36654 978
rect 36706 926 36820 978
rect 36652 924 36820 926
rect 36652 914 36708 924
rect 36540 532 36596 542
rect 36540 112 36596 476
rect 36764 196 36820 924
rect 37100 756 37156 3332
rect 37436 3266 37492 3276
rect 37660 2996 37716 3006
rect 37324 2772 37380 2782
rect 37324 2678 37380 2716
rect 37660 2770 37716 2940
rect 37660 2718 37662 2770
rect 37714 2718 37716 2770
rect 37660 2706 37716 2718
rect 37548 2212 37604 2222
rect 37548 2118 37604 2156
rect 36764 130 36820 140
rect 36988 700 37156 756
rect 37212 2098 37268 2110
rect 37212 2046 37214 2098
rect 37266 2046 37268 2098
rect 36988 112 37044 700
rect 37212 420 37268 2046
rect 37772 1876 37828 8204
rect 37884 7586 37940 15092
rect 37996 14530 38052 14542
rect 37996 14478 37998 14530
rect 38050 14478 38052 14530
rect 37996 14308 38052 14478
rect 37996 14242 38052 14252
rect 38220 14084 38276 14094
rect 37996 13636 38052 13646
rect 37996 13542 38052 13580
rect 38108 12964 38164 12974
rect 38108 11998 38164 12908
rect 38220 12178 38276 14028
rect 38220 12126 38222 12178
rect 38274 12126 38276 12178
rect 38220 12114 38276 12126
rect 38108 11942 38276 11998
rect 37996 11844 38052 11854
rect 37996 9042 38052 11788
rect 37996 8990 37998 9042
rect 38050 8990 38052 9042
rect 37996 8978 38052 8990
rect 38108 11732 38164 11742
rect 37884 7534 37886 7586
rect 37938 7534 37940 7586
rect 37884 7522 37940 7534
rect 38108 7252 38164 11676
rect 38220 10722 38276 11942
rect 38332 11732 38388 15596
rect 38444 15316 38500 15354
rect 38444 15250 38500 15260
rect 38556 15202 38612 17614
rect 38556 15150 38558 15202
rect 38610 15150 38612 15202
rect 38556 15138 38612 15150
rect 38668 14084 38724 18620
rect 38780 18452 38836 23100
rect 39004 23090 39060 23100
rect 39116 21588 39172 23436
rect 39228 22932 39284 22942
rect 39228 22838 39284 22876
rect 39340 21924 39396 23884
rect 39564 23938 39620 24556
rect 39564 23886 39566 23938
rect 39618 23886 39620 23938
rect 39564 23874 39620 23886
rect 39676 24276 39732 24286
rect 39676 23548 39732 24220
rect 39900 23828 39956 26908
rect 40012 23940 40068 27132
rect 40124 26908 40180 27244
rect 40236 27234 40292 27244
rect 40236 27076 40292 27114
rect 40236 27010 40292 27020
rect 40124 26852 40292 26908
rect 40124 26292 40180 26302
rect 40124 26198 40180 26236
rect 40124 25844 40180 25854
rect 40124 25620 40180 25788
rect 40124 25554 40180 25564
rect 40012 23874 40068 23884
rect 40124 24500 40180 24510
rect 40236 24500 40292 26852
rect 40348 25284 40404 29260
rect 40460 28642 40516 29374
rect 40460 28590 40462 28642
rect 40514 28590 40516 28642
rect 40460 28578 40516 28590
rect 40684 28084 40740 32284
rect 40796 28196 40852 33406
rect 40908 33348 40964 33358
rect 40908 29316 40964 33292
rect 41020 32004 41076 38612
rect 41244 38610 41300 38622
rect 41244 38558 41246 38610
rect 41298 38558 41300 38610
rect 41244 36708 41300 38558
rect 41244 36642 41300 36652
rect 41356 36484 41412 39228
rect 41468 38276 41524 38286
rect 41468 38182 41524 38220
rect 41468 37716 41524 37726
rect 41468 37380 41524 37660
rect 41468 37314 41524 37324
rect 41580 37044 41636 41806
rect 41916 41860 41972 41870
rect 41916 41766 41972 41804
rect 42364 41860 42420 42478
rect 42364 41794 42420 41804
rect 42364 41524 42420 41534
rect 42252 41076 42308 41086
rect 42028 40964 42084 40974
rect 41916 40962 42084 40964
rect 41916 40910 42030 40962
rect 42082 40910 42084 40962
rect 41916 40908 42084 40910
rect 41916 39618 41972 40908
rect 42028 40898 42084 40908
rect 41916 39566 41918 39618
rect 41970 39566 41972 39618
rect 41916 39554 41972 39566
rect 42028 40404 42084 40414
rect 41916 39172 41972 39182
rect 41916 38834 41972 39116
rect 41916 38782 41918 38834
rect 41970 38782 41972 38834
rect 41916 38724 41972 38782
rect 42028 38836 42084 40348
rect 42252 39844 42308 41020
rect 42364 40628 42420 41468
rect 42476 41186 42532 43372
rect 42924 43314 42980 43820
rect 43148 43652 43204 44522
rect 43260 44436 43316 44830
rect 43260 43876 43316 44380
rect 43260 43810 43316 43820
rect 43148 43596 43316 43652
rect 43036 43540 43092 43550
rect 43092 43484 43204 43540
rect 43036 43474 43092 43484
rect 43148 43426 43204 43484
rect 43148 43374 43150 43426
rect 43202 43374 43204 43426
rect 43148 43362 43204 43374
rect 42924 43262 42926 43314
rect 42978 43262 42980 43314
rect 42924 43204 42980 43262
rect 42700 43148 42980 43204
rect 43036 43314 43092 43326
rect 43036 43262 43038 43314
rect 43090 43262 43092 43314
rect 42588 41860 42644 41870
rect 42588 41766 42644 41804
rect 42588 41412 42644 41422
rect 42588 41318 42644 41356
rect 42476 41134 42478 41186
rect 42530 41134 42532 41186
rect 42476 40852 42532 41134
rect 42700 41188 42756 43148
rect 42812 42642 42868 42654
rect 42812 42590 42814 42642
rect 42866 42590 42868 42642
rect 42812 41412 42868 42590
rect 42924 42530 42980 42542
rect 42924 42478 42926 42530
rect 42978 42478 42980 42530
rect 42924 41524 42980 42478
rect 43036 42084 43092 43262
rect 43260 42194 43316 43596
rect 43372 43650 43428 45052
rect 43484 44772 43540 46620
rect 43484 44706 43540 44716
rect 43372 43598 43374 43650
rect 43426 43598 43428 43650
rect 43372 43586 43428 43598
rect 43484 44210 43540 44222
rect 43484 44158 43486 44210
rect 43538 44158 43540 44210
rect 43372 42756 43428 42766
rect 43484 42756 43540 44158
rect 43596 43650 43652 47180
rect 43708 47170 43764 47180
rect 43804 47068 44068 47078
rect 43860 47012 43908 47068
rect 43964 47012 44012 47068
rect 43804 47002 44068 47012
rect 44380 46676 44436 47292
rect 44828 47236 44884 47406
rect 44828 47170 44884 47180
rect 45164 47236 45220 47246
rect 44156 46620 44436 46676
rect 43820 46564 43876 46574
rect 43820 46114 43876 46508
rect 43820 46062 43822 46114
rect 43874 46062 43876 46114
rect 43820 45780 43876 46062
rect 43820 45714 43876 45724
rect 43804 45500 44068 45510
rect 43860 45444 43908 45500
rect 43964 45444 44012 45500
rect 43804 45434 44068 45444
rect 43820 44660 43876 44670
rect 43820 44434 43876 44604
rect 43820 44382 43822 44434
rect 43874 44382 43876 44434
rect 43820 44370 43876 44382
rect 43804 43932 44068 43942
rect 43860 43876 43908 43932
rect 43964 43876 44012 43932
rect 43804 43866 44068 43876
rect 43596 43598 43598 43650
rect 43650 43598 43652 43650
rect 43596 43586 43652 43598
rect 43708 43764 43764 43774
rect 43372 42754 43540 42756
rect 43372 42702 43374 42754
rect 43426 42702 43540 42754
rect 43372 42700 43540 42702
rect 43596 43316 43652 43326
rect 43372 42644 43428 42700
rect 43372 42420 43428 42588
rect 43372 42354 43428 42364
rect 43260 42142 43262 42194
rect 43314 42142 43316 42194
rect 43260 42130 43316 42142
rect 43484 42308 43540 42318
rect 43036 42028 43204 42084
rect 43036 41860 43092 41870
rect 43036 41766 43092 41804
rect 42924 41458 42980 41468
rect 42812 41346 42868 41356
rect 43148 41300 43204 42028
rect 43372 41860 43428 41870
rect 43260 41748 43316 41758
rect 43260 41410 43316 41692
rect 43260 41358 43262 41410
rect 43314 41358 43316 41410
rect 43260 41346 43316 41358
rect 43148 41234 43204 41244
rect 42812 41188 42868 41198
rect 43036 41188 43092 41198
rect 42700 41186 42868 41188
rect 42700 41134 42814 41186
rect 42866 41134 42868 41186
rect 42700 41132 42868 41134
rect 42812 41122 42868 41132
rect 42924 41186 43092 41188
rect 42924 41134 43038 41186
rect 43090 41134 43092 41186
rect 42924 41132 43092 41134
rect 42476 40786 42532 40796
rect 42364 40572 42532 40628
rect 42252 39778 42308 39788
rect 42364 40402 42420 40414
rect 42364 40350 42366 40402
rect 42418 40350 42420 40402
rect 42252 39618 42308 39630
rect 42252 39566 42254 39618
rect 42306 39566 42308 39618
rect 42252 39508 42308 39566
rect 42252 39442 42308 39452
rect 42364 39396 42420 40350
rect 42476 39620 42532 40572
rect 42924 40626 42980 41132
rect 43036 41122 43092 41132
rect 43372 40964 43428 41804
rect 43372 40870 43428 40908
rect 42924 40574 42926 40626
rect 42978 40574 42980 40626
rect 42924 40562 42980 40574
rect 42812 40516 42868 40526
rect 42812 40422 42868 40460
rect 43372 40404 43428 40414
rect 43484 40404 43540 42252
rect 43596 42194 43652 43260
rect 43708 42980 43764 43708
rect 43708 42914 43764 42924
rect 43932 43764 43988 43774
rect 44156 43708 44212 46620
rect 43932 42978 43988 43708
rect 43932 42926 43934 42978
rect 43986 42926 43988 42978
rect 43932 42756 43988 42926
rect 44044 43652 44212 43708
rect 44268 46450 44324 46462
rect 44268 46398 44270 46450
rect 44322 46398 44324 46450
rect 44044 42980 44100 43652
rect 44268 43540 44324 46398
rect 44464 46284 44728 46294
rect 44520 46228 44568 46284
rect 44624 46228 44672 46284
rect 44464 46218 44728 46228
rect 45052 45892 45108 45902
rect 44940 45668 44996 45678
rect 44940 45574 44996 45612
rect 44828 45444 44884 45454
rect 44380 45332 44436 45342
rect 44380 45218 44436 45276
rect 44380 45166 44382 45218
rect 44434 45166 44436 45218
rect 44380 45154 44436 45166
rect 44828 44882 44884 45388
rect 44828 44830 44830 44882
rect 44882 44830 44884 44882
rect 44464 44716 44728 44726
rect 44520 44660 44568 44716
rect 44624 44660 44672 44716
rect 44464 44650 44728 44660
rect 44828 43764 44884 44830
rect 45052 44660 45108 45836
rect 45164 45332 45220 47180
rect 45500 47012 45556 48188
rect 45500 46562 45556 46956
rect 45500 46510 45502 46562
rect 45554 46510 45556 46562
rect 45500 46498 45556 46510
rect 45164 45266 45220 45276
rect 45388 46452 45444 46462
rect 45052 44594 45108 44604
rect 44940 44436 44996 44446
rect 44940 43876 44996 44380
rect 45052 44100 45108 44110
rect 45052 44098 45332 44100
rect 45052 44046 45054 44098
rect 45106 44046 45332 44098
rect 45052 44044 45332 44046
rect 45052 44034 45108 44044
rect 44940 43820 45108 43876
rect 44828 43708 44996 43764
rect 44268 43474 44324 43484
rect 44492 43540 44548 43550
rect 44492 43446 44548 43484
rect 44828 43538 44884 43550
rect 44828 43486 44830 43538
rect 44882 43486 44884 43538
rect 44156 43428 44212 43438
rect 44156 43334 44212 43372
rect 44268 43314 44324 43326
rect 44268 43262 44270 43314
rect 44322 43262 44324 43314
rect 44268 43204 44324 43262
rect 44268 43138 44324 43148
rect 44464 43148 44728 43158
rect 44520 43092 44568 43148
rect 44624 43092 44672 43148
rect 44464 43082 44728 43092
rect 44044 42924 44212 42980
rect 43932 42690 43988 42700
rect 43804 42364 44068 42374
rect 43860 42308 43908 42364
rect 43964 42308 44012 42364
rect 43804 42298 44068 42308
rect 43596 42142 43598 42194
rect 43650 42142 43652 42194
rect 43596 42130 43652 42142
rect 43820 41412 43876 41422
rect 43820 41318 43876 41356
rect 44156 40852 44212 42924
rect 43804 40796 44068 40806
rect 43860 40740 43908 40796
rect 43964 40740 44012 40796
rect 43804 40730 44068 40740
rect 43484 40348 43764 40404
rect 43372 40310 43428 40348
rect 43596 40180 43652 40190
rect 43372 40178 43652 40180
rect 43372 40126 43598 40178
rect 43650 40126 43652 40178
rect 43372 40124 43652 40126
rect 42476 39554 42532 39564
rect 43260 39618 43316 39630
rect 43260 39566 43262 39618
rect 43314 39566 43316 39618
rect 43260 39396 43316 39566
rect 42364 39340 43316 39396
rect 42028 38770 42084 38780
rect 42588 39172 42644 39182
rect 41916 38658 41972 38668
rect 42364 38722 42420 38734
rect 42364 38670 42366 38722
rect 42418 38670 42420 38722
rect 42364 38668 42420 38670
rect 42364 38612 42532 38668
rect 42476 38546 42532 38556
rect 42028 38276 42084 38286
rect 41916 38220 42028 38276
rect 41916 37940 41972 38220
rect 42028 38210 42084 38220
rect 41804 37938 41972 37940
rect 41804 37886 41918 37938
rect 41970 37886 41972 37938
rect 41804 37884 41972 37886
rect 41804 37380 41860 37884
rect 41916 37874 41972 37884
rect 42476 37940 42532 37950
rect 42476 37846 42532 37884
rect 41804 37314 41860 37324
rect 41916 37266 41972 37278
rect 41916 37214 41918 37266
rect 41970 37214 41972 37266
rect 41916 37156 41972 37214
rect 41916 37100 42084 37156
rect 41244 36428 41412 36484
rect 41468 36988 41636 37044
rect 41132 36372 41188 36382
rect 41132 36278 41188 36316
rect 41244 35308 41300 36428
rect 41132 35252 41300 35308
rect 41356 36260 41412 36270
rect 41132 32900 41188 35252
rect 41356 34356 41412 36204
rect 41468 35476 41524 36988
rect 41804 36932 41860 36942
rect 41580 36482 41636 36494
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 35924 41636 36430
rect 41580 35858 41636 35868
rect 41692 36372 41748 36382
rect 41468 35410 41524 35420
rect 41356 34290 41412 34300
rect 41468 35140 41524 35150
rect 41244 34018 41300 34030
rect 41244 33966 41246 34018
rect 41298 33966 41300 34018
rect 41244 33796 41300 33966
rect 41244 33730 41300 33740
rect 41468 33348 41524 35084
rect 41580 35026 41636 35038
rect 41580 34974 41582 35026
rect 41634 34974 41636 35026
rect 41580 34468 41636 34974
rect 41692 34804 41748 36316
rect 41692 34738 41748 34748
rect 41580 34402 41636 34412
rect 41804 34244 41860 36876
rect 42028 36708 42084 37100
rect 42476 36932 42532 36942
rect 42140 36708 42196 36718
rect 42028 36706 42196 36708
rect 42028 36654 42142 36706
rect 42194 36654 42196 36706
rect 42028 36652 42196 36654
rect 41916 36482 41972 36494
rect 41916 36430 41918 36482
rect 41970 36430 41972 36482
rect 41916 35812 41972 36430
rect 41916 35746 41972 35756
rect 42028 35698 42084 36652
rect 42140 36642 42196 36652
rect 42252 36708 42308 36718
rect 42028 35646 42030 35698
rect 42082 35646 42084 35698
rect 42028 35634 42084 35646
rect 42028 35140 42084 35150
rect 42028 34914 42084 35084
rect 42028 34862 42030 34914
rect 42082 34862 42084 34914
rect 42028 34580 42084 34862
rect 42028 34514 42084 34524
rect 41468 33282 41524 33292
rect 41580 34188 41804 34244
rect 41132 32834 41188 32844
rect 41244 33012 41300 33022
rect 41020 31938 41076 31948
rect 41132 32562 41188 32574
rect 41132 32510 41134 32562
rect 41186 32510 41188 32562
rect 41132 31780 41188 32510
rect 41244 31890 41300 32956
rect 41356 32340 41412 32350
rect 41356 32246 41412 32284
rect 41244 31838 41246 31890
rect 41298 31838 41300 31890
rect 41244 31826 41300 31838
rect 41580 32228 41636 34188
rect 41804 34178 41860 34188
rect 41692 33906 41748 33918
rect 41692 33854 41694 33906
rect 41746 33854 41748 33906
rect 41692 32564 41748 33854
rect 42028 33124 42084 33134
rect 41916 33122 42084 33124
rect 41916 33070 42030 33122
rect 42082 33070 42084 33122
rect 41916 33068 42084 33070
rect 41804 32564 41860 32574
rect 41692 32562 41860 32564
rect 41692 32510 41806 32562
rect 41858 32510 41860 32562
rect 41692 32508 41860 32510
rect 41804 32498 41860 32508
rect 41132 31714 41188 31724
rect 41132 30996 41188 31006
rect 41132 30324 41188 30940
rect 41580 30882 41636 32172
rect 41692 31780 41748 31790
rect 41916 31780 41972 33068
rect 42028 33058 42084 33068
rect 42252 32228 42308 36652
rect 42364 35588 42420 35598
rect 42364 32788 42420 35532
rect 42476 33012 42532 36876
rect 42588 36594 42644 39116
rect 43260 38276 43316 39340
rect 43260 38210 43316 38220
rect 42812 38050 42868 38062
rect 42812 37998 42814 38050
rect 42866 37998 42868 38050
rect 42812 37380 42868 37998
rect 42812 37314 42868 37324
rect 43260 37604 43316 37614
rect 43260 37266 43316 37548
rect 43260 37214 43262 37266
rect 43314 37214 43316 37266
rect 43260 37202 43316 37214
rect 42700 37154 42756 37166
rect 42700 37102 42702 37154
rect 42754 37102 42756 37154
rect 42700 37044 42756 37102
rect 42700 36978 42756 36988
rect 42812 37042 42868 37054
rect 42812 36990 42814 37042
rect 42866 36990 42868 37042
rect 42812 36708 42868 36990
rect 43036 37044 43092 37054
rect 43036 37042 43316 37044
rect 43036 36990 43038 37042
rect 43090 36990 43316 37042
rect 43036 36988 43316 36990
rect 43036 36978 43092 36988
rect 42588 36542 42590 36594
rect 42642 36542 42644 36594
rect 42588 36530 42644 36542
rect 42700 36652 42868 36708
rect 42700 35140 42756 36652
rect 43148 36482 43204 36494
rect 43148 36430 43150 36482
rect 43202 36430 43204 36482
rect 42924 35588 42980 35598
rect 42924 35494 42980 35532
rect 43148 35588 43204 36430
rect 43148 35522 43204 35532
rect 43036 35474 43092 35486
rect 43036 35422 43038 35474
rect 43090 35422 43092 35474
rect 42700 35074 42756 35084
rect 42812 35252 42868 35262
rect 42700 34802 42756 34814
rect 42700 34750 42702 34802
rect 42754 34750 42756 34802
rect 42700 33348 42756 34750
rect 42812 34018 42868 35196
rect 42812 33966 42814 34018
rect 42866 33966 42868 34018
rect 42812 33954 42868 33966
rect 43036 34020 43092 35422
rect 43036 33954 43092 33964
rect 43148 35026 43204 35038
rect 43148 34974 43150 35026
rect 43202 34974 43204 35026
rect 42700 33282 42756 33292
rect 42476 32946 42532 32956
rect 43148 33012 43204 34974
rect 43260 34692 43316 36988
rect 43372 36708 43428 40124
rect 43596 40114 43652 40124
rect 43708 39508 43764 40348
rect 44156 40068 44212 40796
rect 44268 41746 44324 41758
rect 44268 41694 44270 41746
rect 44322 41694 44324 41746
rect 44268 40516 44324 41694
rect 44828 41748 44884 43486
rect 44940 41972 44996 43708
rect 45052 43762 45108 43820
rect 45052 43710 45054 43762
rect 45106 43710 45108 43762
rect 45052 43698 45108 43710
rect 45164 43538 45220 43550
rect 45164 43486 45166 43538
rect 45218 43486 45220 43538
rect 45052 42980 45108 42990
rect 45164 42980 45220 43486
rect 45052 42978 45220 42980
rect 45052 42926 45054 42978
rect 45106 42926 45220 42978
rect 45052 42924 45220 42926
rect 45052 42914 45108 42924
rect 45276 42868 45332 44044
rect 45388 43540 45444 46396
rect 45612 46340 45668 48972
rect 45724 48916 45780 49534
rect 45724 48850 45780 48860
rect 45724 47684 45780 47694
rect 45836 47684 45892 50204
rect 45724 47682 45892 47684
rect 45724 47630 45726 47682
rect 45778 47630 45892 47682
rect 45724 47628 45892 47630
rect 45724 47618 45780 47628
rect 45948 47236 46004 50428
rect 46060 50260 46116 52894
rect 46508 52948 46564 52958
rect 46284 52500 46340 52510
rect 46060 49812 46116 50204
rect 46060 49746 46116 49756
rect 46172 52162 46228 52174
rect 46172 52110 46174 52162
rect 46226 52110 46228 52162
rect 46172 50484 46228 52110
rect 46284 50818 46340 52444
rect 46508 52386 46564 52892
rect 46620 52724 46676 52734
rect 46620 52630 46676 52668
rect 46508 52334 46510 52386
rect 46562 52334 46564 52386
rect 46508 52322 46564 52334
rect 46620 52276 46676 52286
rect 46284 50766 46286 50818
rect 46338 50766 46340 50818
rect 46284 50754 46340 50766
rect 46396 51490 46452 51502
rect 46396 51438 46398 51490
rect 46450 51438 46452 51490
rect 46396 50820 46452 51438
rect 46620 51268 46676 52220
rect 46732 52164 46788 53678
rect 46956 53284 47012 55246
rect 47292 54292 47348 54302
rect 47180 53842 47236 53854
rect 47180 53790 47182 53842
rect 47234 53790 47236 53842
rect 47180 53732 47236 53790
rect 47180 53666 47236 53676
rect 46956 53218 47012 53228
rect 46732 52098 46788 52108
rect 46844 52274 46900 52286
rect 46844 52222 46846 52274
rect 46898 52222 46900 52274
rect 46844 52052 46900 52222
rect 47292 52162 47348 54236
rect 47516 53732 47572 53742
rect 47516 53638 47572 53676
rect 47292 52110 47294 52162
rect 47346 52110 47348 52162
rect 47292 52098 47348 52110
rect 47516 52274 47572 52286
rect 47516 52222 47518 52274
rect 47570 52222 47572 52274
rect 46844 51986 46900 51996
rect 47516 51828 47572 52222
rect 47516 51762 47572 51772
rect 46620 51202 46676 51212
rect 46060 49028 46116 49038
rect 46172 49028 46228 50428
rect 46396 49700 46452 50764
rect 47068 51044 47124 51054
rect 46844 49812 46900 49822
rect 46844 49718 46900 49756
rect 46396 49634 46452 49644
rect 46060 49026 46228 49028
rect 46060 48974 46062 49026
rect 46114 48974 46228 49026
rect 46060 48972 46228 48974
rect 46284 49196 46564 49252
rect 46060 48962 46116 48972
rect 45948 46674 46004 47180
rect 45948 46622 45950 46674
rect 46002 46622 46004 46674
rect 45948 46610 46004 46622
rect 46284 46340 46340 49196
rect 46508 49138 46564 49196
rect 46508 49086 46510 49138
rect 46562 49086 46564 49138
rect 46508 49074 46564 49086
rect 46396 49028 46452 49038
rect 46396 46674 46452 48972
rect 46620 49026 46676 49038
rect 46620 48974 46622 49026
rect 46674 48974 46676 49026
rect 46620 48916 46676 48974
rect 46620 48850 46676 48860
rect 46732 49026 46788 49038
rect 46732 48974 46734 49026
rect 46786 48974 46788 49026
rect 46732 48804 46788 48974
rect 47068 48916 47124 50988
rect 47628 51044 47684 55580
rect 47852 55412 47908 56364
rect 48188 56084 48244 57344
rect 48636 56756 48692 57344
rect 48636 56690 48692 56700
rect 49084 56532 49140 57344
rect 49532 56868 49588 57344
rect 49532 56802 49588 56812
rect 49084 56466 49140 56476
rect 49756 56532 49812 56542
rect 48188 56018 48244 56028
rect 49084 55972 49140 55982
rect 49084 55878 49140 55916
rect 49756 55970 49812 56476
rect 49756 55918 49758 55970
rect 49810 55918 49812 55970
rect 49756 55906 49812 55918
rect 47852 55346 47908 55356
rect 48076 55858 48132 55870
rect 48076 55806 48078 55858
rect 48130 55806 48132 55858
rect 48076 55188 48132 55806
rect 48412 55860 48468 55870
rect 48412 55766 48468 55804
rect 48748 55858 48804 55870
rect 48748 55806 48750 55858
rect 48802 55806 48804 55858
rect 48748 55524 48804 55806
rect 49420 55858 49476 55870
rect 49420 55806 49422 55858
rect 49474 55806 49476 55858
rect 48748 55458 48804 55468
rect 48972 55748 49028 55758
rect 48076 55122 48132 55132
rect 48860 55298 48916 55310
rect 48860 55246 48862 55298
rect 48914 55246 48916 55298
rect 48748 54740 48804 54750
rect 48636 54404 48692 54414
rect 48412 53844 48468 53854
rect 48412 53842 48580 53844
rect 48412 53790 48414 53842
rect 48466 53790 48580 53842
rect 48412 53788 48580 53790
rect 48412 53778 48468 53788
rect 48188 53732 48244 53742
rect 48188 53638 48244 53676
rect 48412 52836 48468 52846
rect 48412 52742 48468 52780
rect 47740 52724 47796 52734
rect 47740 52722 48244 52724
rect 47740 52670 47742 52722
rect 47794 52670 48244 52722
rect 47740 52668 48244 52670
rect 47740 52658 47796 52668
rect 48076 52164 48132 52174
rect 48076 51156 48132 52108
rect 48188 52162 48244 52668
rect 48188 52110 48190 52162
rect 48242 52110 48244 52162
rect 48188 52098 48244 52110
rect 48300 52388 48356 52398
rect 48300 51604 48356 52332
rect 48524 52388 48580 53788
rect 48636 53284 48692 54348
rect 48748 54180 48804 54684
rect 48860 54626 48916 55246
rect 48860 54574 48862 54626
rect 48914 54574 48916 54626
rect 48860 54562 48916 54574
rect 48748 54114 48804 54124
rect 48972 54180 49028 55692
rect 48972 54114 49028 54124
rect 49196 55748 49252 55758
rect 49084 53842 49140 53854
rect 49084 53790 49086 53842
rect 49138 53790 49140 53842
rect 49084 53732 49140 53790
rect 49196 53844 49252 55692
rect 49420 55524 49476 55806
rect 49420 55458 49476 55468
rect 49980 55524 50036 57344
rect 50428 55468 50484 57344
rect 50540 57204 50596 57214
rect 50540 55970 50596 57148
rect 50876 57092 50932 57344
rect 50876 57026 50932 57036
rect 50540 55918 50542 55970
rect 50594 55918 50596 55970
rect 50540 55906 50596 55918
rect 49980 55458 50036 55468
rect 50316 55412 50484 55468
rect 50876 55858 50932 55870
rect 50876 55806 50878 55858
rect 50930 55806 50932 55858
rect 50876 55524 50932 55806
rect 51212 55858 51268 55870
rect 51212 55806 51214 55858
rect 51266 55806 51268 55858
rect 50876 55458 50932 55468
rect 51100 55636 51156 55646
rect 50316 54964 50372 55412
rect 50428 55188 50484 55198
rect 50428 55094 50484 55132
rect 50316 54898 50372 54908
rect 50652 54852 50708 54862
rect 49980 54740 50036 54750
rect 49420 54068 49476 54078
rect 49420 53954 49476 54012
rect 49420 53902 49422 53954
rect 49474 53902 49476 53954
rect 49420 53890 49476 53902
rect 49196 53778 49252 53788
rect 49084 53666 49140 53676
rect 49868 53730 49924 53742
rect 49868 53678 49870 53730
rect 49922 53678 49924 53730
rect 48636 53218 48692 53228
rect 49868 53060 49924 53678
rect 49868 52994 49924 53004
rect 48524 52322 48580 52332
rect 48748 52722 48804 52734
rect 48748 52670 48750 52722
rect 48802 52670 48804 52722
rect 48748 52276 48804 52670
rect 49196 52724 49252 52734
rect 49196 52630 49252 52668
rect 49532 52724 49588 52734
rect 49532 52722 49812 52724
rect 49532 52670 49534 52722
rect 49586 52670 49812 52722
rect 49532 52668 49812 52670
rect 49532 52658 49588 52668
rect 48748 52210 48804 52220
rect 48860 52612 48916 52622
rect 48860 52052 48916 52556
rect 49532 52274 49588 52286
rect 49532 52222 49534 52274
rect 49586 52222 49588 52274
rect 48860 51986 48916 51996
rect 49420 52050 49476 52062
rect 49420 51998 49422 52050
rect 49474 51998 49476 52050
rect 48300 51538 48356 51548
rect 48412 51938 48468 51950
rect 48412 51886 48414 51938
rect 48466 51886 48468 51938
rect 48076 51090 48132 51100
rect 47628 50978 47684 50988
rect 47740 50932 47796 50942
rect 47180 50708 47236 50718
rect 47180 50428 47236 50652
rect 47404 50708 47460 50718
rect 47404 50614 47460 50652
rect 47516 50596 47572 50606
rect 47180 50372 47348 50428
rect 47292 49812 47348 50372
rect 47180 49810 47348 49812
rect 47180 49758 47294 49810
rect 47346 49758 47348 49810
rect 47180 49756 47348 49758
rect 47180 49250 47236 49756
rect 47292 49746 47348 49756
rect 47404 50260 47460 50270
rect 47180 49198 47182 49250
rect 47234 49198 47236 49250
rect 47180 49186 47236 49198
rect 47068 48850 47124 48860
rect 46732 48738 46788 48748
rect 46956 48354 47012 48366
rect 46956 48302 46958 48354
rect 47010 48302 47012 48354
rect 46508 48018 46564 48030
rect 46508 47966 46510 48018
rect 46562 47966 46564 48018
rect 46508 47460 46564 47966
rect 46844 47572 46900 47582
rect 46844 47478 46900 47516
rect 46508 47394 46564 47404
rect 46396 46622 46398 46674
rect 46450 46622 46452 46674
rect 46396 46610 46452 46622
rect 46732 46676 46788 46686
rect 46732 46582 46788 46620
rect 46508 46452 46564 46462
rect 46956 46452 47012 48302
rect 46508 46450 47012 46452
rect 46508 46398 46510 46450
rect 46562 46398 47012 46450
rect 46508 46396 47012 46398
rect 47068 47796 47124 47806
rect 47068 46674 47124 47740
rect 47068 46622 47070 46674
rect 47122 46622 47124 46674
rect 46508 46386 46564 46396
rect 45500 46284 45668 46340
rect 45724 46284 46340 46340
rect 45500 44548 45556 46284
rect 45612 46004 45668 46014
rect 45612 45890 45668 45948
rect 45612 45838 45614 45890
rect 45666 45838 45668 45890
rect 45612 45826 45668 45838
rect 45500 44492 45668 44548
rect 45388 43474 45444 43484
rect 45500 43426 45556 43438
rect 45500 43374 45502 43426
rect 45554 43374 45556 43426
rect 45388 43314 45444 43326
rect 45388 43262 45390 43314
rect 45442 43262 45444 43314
rect 45388 42980 45444 43262
rect 45388 42914 45444 42924
rect 45276 42802 45332 42812
rect 44940 41906 44996 41916
rect 45052 42756 45108 42766
rect 44828 41682 44884 41692
rect 44464 41580 44728 41590
rect 44520 41524 44568 41580
rect 44624 41524 44672 41580
rect 44464 41514 44728 41524
rect 44940 41298 44996 41310
rect 44940 41246 44942 41298
rect 44994 41246 44996 41298
rect 44940 41188 44996 41246
rect 44940 41122 44996 41132
rect 45052 40964 45108 42700
rect 45500 42754 45556 43374
rect 45500 42702 45502 42754
rect 45554 42702 45556 42754
rect 45164 42644 45220 42654
rect 45164 41188 45220 42588
rect 45388 41746 45444 41758
rect 45388 41694 45390 41746
rect 45442 41694 45444 41746
rect 45388 41524 45444 41694
rect 45388 41458 45444 41468
rect 45500 41748 45556 42702
rect 45388 41188 45444 41198
rect 45164 41186 45444 41188
rect 45164 41134 45390 41186
rect 45442 41134 45444 41186
rect 45164 41132 45444 41134
rect 45388 41122 45444 41132
rect 44940 40908 45108 40964
rect 45500 40964 45556 41692
rect 44492 40516 44548 40526
rect 44268 40450 44324 40460
rect 44380 40460 44492 40516
rect 44380 40402 44436 40460
rect 44492 40450 44548 40460
rect 44380 40350 44382 40402
rect 44434 40350 44436 40402
rect 44380 40180 44436 40350
rect 44156 40002 44212 40012
rect 44268 40124 44436 40180
rect 44828 40180 44884 40190
rect 43708 39442 43764 39452
rect 43932 39396 43988 39406
rect 43932 39394 44212 39396
rect 43932 39342 43934 39394
rect 43986 39342 44212 39394
rect 43932 39340 44212 39342
rect 43932 39330 43988 39340
rect 43804 39228 44068 39238
rect 43484 39172 43540 39182
rect 43860 39172 43908 39228
rect 43964 39172 44012 39228
rect 43804 39162 44068 39172
rect 43484 39058 43540 39116
rect 44156 39060 44212 39340
rect 43484 39006 43486 39058
rect 43538 39006 43540 39058
rect 43484 38994 43540 39006
rect 44044 39004 44212 39060
rect 43932 38724 43988 38734
rect 43708 38052 43764 38062
rect 43596 38050 43764 38052
rect 43596 37998 43710 38050
rect 43762 37998 43764 38050
rect 43596 37996 43764 37998
rect 43596 37604 43652 37996
rect 43708 37986 43764 37996
rect 43932 37828 43988 38668
rect 44044 38052 44100 39004
rect 44268 38388 44324 40124
rect 44828 40086 44884 40124
rect 44464 40012 44728 40022
rect 44520 39956 44568 40012
rect 44624 39956 44672 40012
rect 44464 39946 44728 39956
rect 44716 39508 44772 39518
rect 44380 39172 44436 39182
rect 44380 38946 44436 39116
rect 44380 38894 44382 38946
rect 44434 38894 44436 38946
rect 44380 38724 44436 38894
rect 44380 38658 44436 38668
rect 44716 38724 44772 39452
rect 44940 38668 44996 40908
rect 45500 40898 45556 40908
rect 45276 40852 45332 40862
rect 45164 40740 45220 40750
rect 45052 39844 45108 39854
rect 45052 39396 45108 39788
rect 45052 39330 45108 39340
rect 44716 38658 44772 38668
rect 44828 38612 44996 38668
rect 44464 38444 44728 38454
rect 44520 38388 44568 38444
rect 44624 38388 44672 38444
rect 44464 38378 44728 38388
rect 44268 38322 44324 38332
rect 44268 38052 44324 38062
rect 44044 38050 44324 38052
rect 44044 37998 44270 38050
rect 44322 37998 44324 38050
rect 44044 37996 44324 37998
rect 44268 37986 44324 37996
rect 44492 38052 44548 38062
rect 43932 37772 44212 37828
rect 44156 37716 44212 37772
rect 43372 36642 43428 36652
rect 43484 37548 43652 37604
rect 43804 37660 44068 37670
rect 43860 37604 43908 37660
rect 43964 37604 44012 37660
rect 44156 37650 44212 37660
rect 43804 37594 44068 37604
rect 44492 37604 44548 37996
rect 43372 36484 43428 36494
rect 43372 35698 43428 36428
rect 43484 36372 43540 37548
rect 44492 37538 44548 37548
rect 43596 37380 43652 37390
rect 43596 37154 43652 37324
rect 43596 37102 43598 37154
rect 43650 37102 43652 37154
rect 43596 37090 43652 37102
rect 43708 37268 43764 37278
rect 43484 36306 43540 36316
rect 43708 36372 43764 37212
rect 44492 37268 44548 37278
rect 44156 37156 44212 37166
rect 44156 37062 44212 37100
rect 44492 37154 44548 37212
rect 44492 37102 44494 37154
rect 44546 37102 44548 37154
rect 44492 37090 44548 37102
rect 44716 37156 44772 37166
rect 44716 37062 44772 37100
rect 44464 36876 44728 36886
rect 44156 36820 44212 36830
rect 44520 36820 44568 36876
rect 44624 36820 44672 36876
rect 44464 36810 44728 36820
rect 44156 36482 44212 36764
rect 44156 36430 44158 36482
rect 44210 36430 44212 36482
rect 44156 36418 44212 36430
rect 43708 36306 43764 36316
rect 43804 36092 44068 36102
rect 43860 36036 43908 36092
rect 43964 36036 44012 36092
rect 43804 36026 44068 36036
rect 44380 36036 44436 36046
rect 44268 35924 44324 35934
rect 44268 35830 44324 35868
rect 43372 35646 43374 35698
rect 43426 35646 43428 35698
rect 43372 35364 43428 35646
rect 43484 35812 43540 35822
rect 43484 35586 43540 35756
rect 43484 35534 43486 35586
rect 43538 35534 43540 35586
rect 43484 35522 43540 35534
rect 43596 35700 43652 35710
rect 44380 35700 44436 35980
rect 43372 35298 43428 35308
rect 43596 35252 43652 35644
rect 44268 35644 44436 35700
rect 43708 35588 43764 35598
rect 43708 35494 43764 35532
rect 43596 35186 43652 35196
rect 44268 34916 44324 35644
rect 44828 35364 44884 38612
rect 44940 38276 44996 38286
rect 44940 38182 44996 38220
rect 45052 38052 45108 38062
rect 45052 37958 45108 37996
rect 44464 35308 44728 35318
rect 44520 35252 44568 35308
rect 44624 35252 44672 35308
rect 44828 35298 44884 35308
rect 44940 37716 44996 37726
rect 44940 36370 44996 37660
rect 45164 37380 45220 40684
rect 45276 40180 45332 40796
rect 45276 40114 45332 40124
rect 45500 39844 45556 39854
rect 45500 39620 45556 39788
rect 45388 39618 45556 39620
rect 45388 39566 45502 39618
rect 45554 39566 45556 39618
rect 45388 39564 45556 39566
rect 45388 39172 45444 39564
rect 45500 39554 45556 39564
rect 45388 39106 45444 39116
rect 45612 39172 45668 44492
rect 45724 43316 45780 46284
rect 46060 46116 46116 46126
rect 46060 46114 46452 46116
rect 46060 46062 46062 46114
rect 46114 46062 46452 46114
rect 46060 46060 46452 46062
rect 46060 46050 46116 46060
rect 45948 45890 46004 45902
rect 45948 45838 45950 45890
rect 46002 45838 46004 45890
rect 45948 45556 46004 45838
rect 46284 45892 46340 45902
rect 46284 45798 46340 45836
rect 46172 45778 46228 45790
rect 46172 45726 46174 45778
rect 46226 45726 46228 45778
rect 45948 45500 46116 45556
rect 45948 45332 46004 45342
rect 45948 45238 46004 45276
rect 45836 44436 45892 44446
rect 45836 44322 45892 44380
rect 45836 44270 45838 44322
rect 45890 44270 45892 44322
rect 45836 44258 45892 44270
rect 45948 43540 46004 43550
rect 45724 43250 45780 43260
rect 45836 43314 45892 43326
rect 45836 43262 45838 43314
rect 45890 43262 45892 43314
rect 45724 42868 45780 42878
rect 45724 42774 45780 42812
rect 45724 42644 45780 42654
rect 45724 41972 45780 42588
rect 45836 42196 45892 43262
rect 45948 42754 46004 43484
rect 46060 42980 46116 45500
rect 46172 43652 46228 45726
rect 46396 45108 46452 46060
rect 46508 45220 46564 45230
rect 46508 45126 46564 45164
rect 46396 45014 46452 45052
rect 46620 44772 46676 46396
rect 46956 45780 47012 45790
rect 46844 45778 47012 45780
rect 46844 45726 46958 45778
rect 47010 45726 47012 45778
rect 46844 45724 47012 45726
rect 46732 45668 46788 45678
rect 46732 45574 46788 45612
rect 46620 44706 46676 44716
rect 46732 45444 46788 45454
rect 46284 44434 46340 44446
rect 46284 44382 46286 44434
rect 46338 44382 46340 44434
rect 46284 43988 46340 44382
rect 46284 43922 46340 43932
rect 46172 43596 46564 43652
rect 46172 43314 46228 43326
rect 46172 43262 46174 43314
rect 46226 43262 46228 43314
rect 46172 43204 46228 43262
rect 46172 43138 46228 43148
rect 46060 42924 46228 42980
rect 45948 42702 45950 42754
rect 46002 42702 46004 42754
rect 45948 42690 46004 42702
rect 46060 42754 46116 42766
rect 46060 42702 46062 42754
rect 46114 42702 46116 42754
rect 46060 42644 46116 42702
rect 46060 42578 46116 42588
rect 45836 42140 46116 42196
rect 45948 41972 46004 41982
rect 45724 41970 46004 41972
rect 45724 41918 45950 41970
rect 46002 41918 46004 41970
rect 45724 41916 46004 41918
rect 45724 41636 45780 41646
rect 45724 39620 45780 41580
rect 45724 39554 45780 39564
rect 45836 41524 45892 41534
rect 45612 39106 45668 39116
rect 45836 38948 45892 41468
rect 45948 40964 46004 41916
rect 46060 40964 46116 42140
rect 46172 41412 46228 42924
rect 46284 42978 46340 42990
rect 46284 42926 46286 42978
rect 46338 42926 46340 42978
rect 46284 42756 46340 42926
rect 46508 42756 46564 43596
rect 46620 43316 46676 43326
rect 46620 43222 46676 43260
rect 46620 42756 46676 42766
rect 46508 42754 46676 42756
rect 46508 42702 46622 42754
rect 46674 42702 46676 42754
rect 46508 42700 46676 42702
rect 46284 42690 46340 42700
rect 46620 42690 46676 42700
rect 46732 42532 46788 45388
rect 46844 43540 46900 45724
rect 46956 45714 47012 45724
rect 47068 45218 47124 46622
rect 47404 47458 47460 50204
rect 47404 47406 47406 47458
rect 47458 47406 47460 47458
rect 47404 46452 47460 47406
rect 47404 46386 47460 46396
rect 47516 50034 47572 50540
rect 47516 49982 47518 50034
rect 47570 49982 47572 50034
rect 47516 46228 47572 49982
rect 47628 49924 47684 49934
rect 47628 46676 47684 49868
rect 47740 47684 47796 50876
rect 48076 50932 48132 50942
rect 47852 50372 47908 50382
rect 47852 49810 47908 50316
rect 47852 49758 47854 49810
rect 47906 49758 47908 49810
rect 47852 49746 47908 49758
rect 48076 49812 48132 50876
rect 48412 50036 48468 51886
rect 48748 51940 48804 51950
rect 48524 51492 48580 51502
rect 48524 51398 48580 51436
rect 48748 51156 48804 51884
rect 48748 51090 48804 51100
rect 48972 51940 49028 51950
rect 48860 50820 48916 50830
rect 48524 50596 48580 50606
rect 48524 50502 48580 50540
rect 48860 50594 48916 50764
rect 48860 50542 48862 50594
rect 48914 50542 48916 50594
rect 48860 50530 48916 50542
rect 48972 50428 49028 51884
rect 49308 51938 49364 51950
rect 49308 51886 49310 51938
rect 49362 51886 49364 51938
rect 49308 51604 49364 51886
rect 49308 51538 49364 51548
rect 49196 51378 49252 51390
rect 49196 51326 49198 51378
rect 49250 51326 49252 51378
rect 49084 50708 49140 50718
rect 49084 50614 49140 50652
rect 49196 50484 49252 51326
rect 49420 50428 49476 51998
rect 48972 50372 49140 50428
rect 48748 50036 48804 50046
rect 48412 50034 48804 50036
rect 48412 49982 48750 50034
rect 48802 49982 48804 50034
rect 48412 49980 48804 49982
rect 48412 49924 48468 49980
rect 48748 49970 48804 49980
rect 48412 49858 48468 49868
rect 48860 49924 48916 49934
rect 48076 49810 48244 49812
rect 48076 49758 48078 49810
rect 48130 49758 48244 49810
rect 48076 49756 48244 49758
rect 48076 49746 48132 49756
rect 47964 49700 48020 49710
rect 47964 49606 48020 49644
rect 48076 48804 48132 48814
rect 47740 47618 47796 47628
rect 47852 48802 48132 48804
rect 47852 48750 48078 48802
rect 48130 48750 48132 48802
rect 47852 48748 48132 48750
rect 47852 46676 47908 48748
rect 48076 48738 48132 48748
rect 48188 48244 48244 49756
rect 48524 49700 48580 49710
rect 48412 49586 48468 49598
rect 48412 49534 48414 49586
rect 48466 49534 48468 49586
rect 48300 49028 48356 49038
rect 48412 49028 48468 49534
rect 48356 48972 48468 49028
rect 48524 49028 48580 49644
rect 48860 49252 48916 49868
rect 48972 49812 49028 49822
rect 48972 49718 49028 49756
rect 49084 49476 49140 50372
rect 49084 49410 49140 49420
rect 48748 49196 48916 49252
rect 48972 49250 49028 49262
rect 48972 49198 48974 49250
rect 49026 49198 49028 49250
rect 48636 49028 48692 49038
rect 48524 49026 48692 49028
rect 48524 48974 48638 49026
rect 48690 48974 48692 49026
rect 48524 48972 48692 48974
rect 48300 48934 48356 48972
rect 48636 48962 48692 48972
rect 47628 46620 47796 46676
rect 47628 46452 47684 46462
rect 47628 46358 47684 46396
rect 47516 46172 47684 46228
rect 47404 46004 47460 46014
rect 47404 45910 47460 45948
rect 47180 45890 47236 45902
rect 47180 45838 47182 45890
rect 47234 45838 47236 45890
rect 47180 45332 47236 45838
rect 47292 45780 47348 45790
rect 47292 45686 47348 45724
rect 47180 45266 47236 45276
rect 47068 45166 47070 45218
rect 47122 45166 47124 45218
rect 46844 43474 46900 43484
rect 46956 44884 47012 44894
rect 46844 42980 46900 42990
rect 46844 42754 46900 42924
rect 46844 42702 46846 42754
rect 46898 42702 46900 42754
rect 46844 42690 46900 42702
rect 46396 42476 46788 42532
rect 46284 41412 46340 41422
rect 46172 41410 46340 41412
rect 46172 41358 46286 41410
rect 46338 41358 46340 41410
rect 46172 41356 46340 41358
rect 46284 41346 46340 41356
rect 46060 40908 46340 40964
rect 45948 40898 46004 40908
rect 45948 40180 46004 40190
rect 45948 40178 46228 40180
rect 45948 40126 45950 40178
rect 46002 40126 46228 40178
rect 45948 40124 46228 40126
rect 45948 40114 46004 40124
rect 46172 39618 46228 40124
rect 46172 39566 46174 39618
rect 46226 39566 46228 39618
rect 46172 39554 46228 39566
rect 45388 38892 45892 38948
rect 45388 38668 45444 38892
rect 46060 38724 46116 38734
rect 46284 38668 46340 40908
rect 46396 39618 46452 42476
rect 46732 41972 46788 41982
rect 46508 41746 46564 41758
rect 46508 41694 46510 41746
rect 46562 41694 46564 41746
rect 46508 41188 46564 41694
rect 46620 41188 46676 41198
rect 46508 41186 46676 41188
rect 46508 41134 46622 41186
rect 46674 41134 46676 41186
rect 46508 41132 46676 41134
rect 46620 41122 46676 41132
rect 46620 40516 46676 40526
rect 46732 40516 46788 41916
rect 46676 40460 46788 40516
rect 46844 40852 46900 40862
rect 46620 40422 46676 40460
rect 46844 40292 46900 40796
rect 46396 39566 46398 39618
rect 46450 39566 46452 39618
rect 46396 38836 46452 39566
rect 46620 40236 46900 40292
rect 46396 38770 46452 38780
rect 46508 39396 46564 39406
rect 46508 38668 46564 39340
rect 45388 38612 45556 38668
rect 45948 38612 46004 38622
rect 45164 37314 45220 37324
rect 44940 36318 44942 36370
rect 44994 36318 44996 36370
rect 44464 35242 44728 35252
rect 44828 35140 44884 35150
rect 44268 34860 44436 34916
rect 44268 34692 44324 34702
rect 43260 34626 43316 34636
rect 44156 34690 44324 34692
rect 44156 34638 44270 34690
rect 44322 34638 44324 34690
rect 44156 34636 44324 34638
rect 43372 34580 43428 34590
rect 43148 32946 43204 32956
rect 43260 34468 43316 34478
rect 43260 33684 43316 34412
rect 43372 34130 43428 34524
rect 43804 34524 44068 34534
rect 43860 34468 43908 34524
rect 43964 34468 44012 34524
rect 43804 34458 44068 34468
rect 43372 34078 43374 34130
rect 43426 34078 43428 34130
rect 43372 33796 43428 34078
rect 43372 33730 43428 33740
rect 42364 32732 42644 32788
rect 42252 32162 42308 32172
rect 42476 32562 42532 32574
rect 42476 32510 42478 32562
rect 42530 32510 42532 32562
rect 42252 31890 42308 31902
rect 42252 31838 42254 31890
rect 42306 31838 42308 31890
rect 41692 31778 41972 31780
rect 41692 31726 41694 31778
rect 41746 31726 41972 31778
rect 41692 31724 41972 31726
rect 42028 31780 42084 31790
rect 41692 31714 41748 31724
rect 42028 31686 42084 31724
rect 42252 31220 42308 31838
rect 42252 31154 42308 31164
rect 42476 31780 42532 32510
rect 41580 30830 41582 30882
rect 41634 30830 41636 30882
rect 41580 30818 41636 30830
rect 41132 30258 41188 30268
rect 41244 30322 41300 30334
rect 41244 30270 41246 30322
rect 41298 30270 41300 30322
rect 41020 30212 41076 30222
rect 41020 30118 41076 30156
rect 41244 30212 41300 30270
rect 41244 30146 41300 30156
rect 41916 30212 41972 30222
rect 41916 30210 42196 30212
rect 41916 30158 41918 30210
rect 41970 30158 42196 30210
rect 41916 30156 42196 30158
rect 41916 30146 41972 30156
rect 42140 29650 42196 30156
rect 42140 29598 42142 29650
rect 42194 29598 42196 29650
rect 42140 29586 42196 29598
rect 42364 30210 42420 30222
rect 42364 30158 42366 30210
rect 42418 30158 42420 30210
rect 40908 29250 40964 29260
rect 41020 29202 41076 29214
rect 41020 29150 41022 29202
rect 41074 29150 41076 29202
rect 41020 28980 41076 29150
rect 41020 28914 41076 28924
rect 42140 28980 42196 28990
rect 40908 28868 40964 28878
rect 40908 28774 40964 28812
rect 40796 28130 40852 28140
rect 41916 28756 41972 28766
rect 40684 28018 40740 28028
rect 40908 27860 40964 27870
rect 40572 27858 40964 27860
rect 40572 27806 40910 27858
rect 40962 27806 40964 27858
rect 40572 27804 40964 27806
rect 40572 27188 40628 27804
rect 40908 27794 40964 27804
rect 41020 27804 41748 27860
rect 40684 27636 40740 27646
rect 40684 27542 40740 27580
rect 40796 27634 40852 27646
rect 40796 27582 40798 27634
rect 40850 27582 40852 27634
rect 40572 27074 40628 27132
rect 40572 27022 40574 27074
rect 40626 27022 40628 27074
rect 40460 26962 40516 26974
rect 40460 26910 40462 26962
rect 40514 26910 40516 26962
rect 40460 26852 40516 26910
rect 40460 26786 40516 26796
rect 40572 26740 40628 27022
rect 40572 26674 40628 26684
rect 40684 27076 40740 27086
rect 40684 26292 40740 27020
rect 40796 26516 40852 27582
rect 40908 27188 40964 27198
rect 41020 27188 41076 27804
rect 41132 27636 41188 27646
rect 41132 27634 41412 27636
rect 41132 27582 41134 27634
rect 41186 27582 41412 27634
rect 41132 27580 41412 27582
rect 41132 27570 41188 27580
rect 40908 27186 41076 27188
rect 40908 27134 40910 27186
rect 40962 27134 41076 27186
rect 40908 27132 41076 27134
rect 40908 27122 40964 27132
rect 41132 27076 41188 27086
rect 41132 26982 41188 27020
rect 41356 26628 41412 27580
rect 41692 27298 41748 27804
rect 41804 27858 41860 27870
rect 41804 27806 41806 27858
rect 41858 27806 41860 27858
rect 41804 27412 41860 27806
rect 41804 27346 41860 27356
rect 41692 27246 41694 27298
rect 41746 27246 41748 27298
rect 41692 27234 41748 27246
rect 41468 27188 41524 27198
rect 41804 27188 41860 27198
rect 41916 27188 41972 28700
rect 41524 27132 41636 27188
rect 41468 27122 41524 27132
rect 41580 27074 41636 27132
rect 41804 27186 41972 27188
rect 41804 27134 41806 27186
rect 41858 27134 41972 27186
rect 41804 27132 41972 27134
rect 42028 28418 42084 28430
rect 42028 28366 42030 28418
rect 42082 28366 42084 28418
rect 41804 27122 41860 27132
rect 41580 27022 41582 27074
rect 41634 27022 41636 27074
rect 41580 27010 41636 27022
rect 41692 27076 41748 27086
rect 41356 26572 41636 26628
rect 40796 26450 40852 26460
rect 41468 26404 41524 26414
rect 40796 26292 40852 26302
rect 40684 26290 40964 26292
rect 40684 26238 40798 26290
rect 40850 26238 40964 26290
rect 40684 26236 40964 26238
rect 40796 26226 40852 26236
rect 40572 26180 40628 26190
rect 40572 26178 40740 26180
rect 40572 26126 40574 26178
rect 40626 26126 40740 26178
rect 40572 26124 40740 26126
rect 40572 26114 40628 26124
rect 40460 26066 40516 26078
rect 40460 26014 40462 26066
rect 40514 26014 40516 26066
rect 40460 25844 40516 26014
rect 40460 25778 40516 25788
rect 40684 25732 40740 26124
rect 40684 25638 40740 25676
rect 40796 25620 40852 25630
rect 40908 25620 40964 26236
rect 41468 26290 41524 26348
rect 41468 26238 41470 26290
rect 41522 26238 41524 26290
rect 41468 26226 41524 26238
rect 41244 26180 41300 26190
rect 41244 26086 41300 26124
rect 41356 26178 41412 26190
rect 41356 26126 41358 26178
rect 41410 26126 41412 26178
rect 41020 25620 41076 25658
rect 40908 25564 41020 25620
rect 40796 25526 40852 25564
rect 41020 25554 41076 25564
rect 40460 25508 40516 25518
rect 40460 25414 40516 25452
rect 41132 25506 41188 25518
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 41020 25396 41076 25406
rect 40348 25228 40628 25284
rect 40124 24498 40292 24500
rect 40124 24446 40126 24498
rect 40178 24446 40292 24498
rect 40124 24444 40292 24446
rect 39340 21858 39396 21868
rect 39452 23492 39732 23548
rect 39788 23772 39956 23828
rect 39004 21532 39172 21588
rect 39228 21588 39284 21626
rect 38892 20804 38948 20814
rect 38892 20710 38948 20748
rect 38780 18386 38836 18396
rect 38892 19236 38948 19246
rect 38780 16884 38836 16894
rect 38780 16790 38836 16828
rect 38892 16100 38948 19180
rect 39004 17556 39060 21532
rect 39228 21522 39284 21532
rect 39228 21140 39284 21150
rect 39116 21028 39172 21038
rect 39116 20914 39172 20972
rect 39116 20862 39118 20914
rect 39170 20862 39172 20914
rect 39116 20692 39172 20862
rect 39228 20914 39284 21084
rect 39228 20862 39230 20914
rect 39282 20862 39284 20914
rect 39228 20850 39284 20862
rect 39116 20626 39172 20636
rect 39228 20690 39284 20702
rect 39228 20638 39230 20690
rect 39282 20638 39284 20690
rect 39228 20580 39284 20638
rect 39228 20514 39284 20524
rect 39340 20020 39396 20030
rect 39452 20020 39508 23492
rect 39564 21588 39620 21598
rect 39564 21494 39620 21532
rect 39788 21252 39844 23772
rect 39900 23492 39956 23502
rect 39900 23154 39956 23436
rect 39900 23102 39902 23154
rect 39954 23102 39956 23154
rect 39900 23090 39956 23102
rect 40012 21700 40068 21710
rect 40012 21586 40068 21644
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 21522 40068 21534
rect 39788 21196 39956 21252
rect 39676 20804 39732 20814
rect 39676 20710 39732 20748
rect 39396 19964 39508 20020
rect 39564 20692 39620 20702
rect 39340 19926 39396 19964
rect 39564 19458 39620 20636
rect 39564 19406 39566 19458
rect 39618 19406 39620 19458
rect 39564 19394 39620 19406
rect 39788 19908 39844 19918
rect 39788 19794 39844 19852
rect 39788 19742 39790 19794
rect 39842 19742 39844 19794
rect 39340 19010 39396 19022
rect 39340 18958 39342 19010
rect 39394 18958 39396 19010
rect 39340 18788 39396 18958
rect 39340 18450 39396 18732
rect 39676 19010 39732 19022
rect 39676 18958 39678 19010
rect 39730 18958 39732 19010
rect 39676 18676 39732 18958
rect 39676 18610 39732 18620
rect 39340 18398 39342 18450
rect 39394 18398 39396 18450
rect 39340 17666 39396 18398
rect 39340 17614 39342 17666
rect 39394 17614 39396 17666
rect 39340 17602 39396 17614
rect 39004 17490 39060 17500
rect 39228 16660 39284 16670
rect 39228 16566 39284 16604
rect 39564 16548 39620 16558
rect 38780 15204 38836 15214
rect 38780 14868 38836 15148
rect 38780 14802 38836 14812
rect 38668 14018 38724 14028
rect 38892 13860 38948 16044
rect 38892 13794 38948 13804
rect 39004 16436 39060 16446
rect 38556 13636 38612 13646
rect 38556 11732 38612 13580
rect 38892 12738 38948 12750
rect 38892 12686 38894 12738
rect 38946 12686 38948 12738
rect 38892 12180 38948 12686
rect 38892 12114 38948 12124
rect 39004 12068 39060 16380
rect 39116 15314 39172 15326
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 13970 39172 15262
rect 39564 15314 39620 16492
rect 39564 15262 39566 15314
rect 39618 15262 39620 15314
rect 39564 15204 39620 15262
rect 39564 15138 39620 15148
rect 39340 14980 39396 14990
rect 39340 14420 39396 14924
rect 39340 14354 39396 14364
rect 39788 13972 39844 19742
rect 39116 13918 39118 13970
rect 39170 13918 39172 13970
rect 39116 13906 39172 13918
rect 39676 13916 39844 13972
rect 39004 12002 39060 12012
rect 39116 13412 39172 13422
rect 38556 11676 38836 11732
rect 38332 11666 38388 11676
rect 38444 11508 38500 11518
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10658 38276 10670
rect 38332 11506 38500 11508
rect 38332 11454 38446 11506
rect 38498 11454 38500 11506
rect 38332 11452 38500 11454
rect 38220 8932 38276 8942
rect 38332 8932 38388 11452
rect 38444 11442 38500 11452
rect 38668 10500 38724 10510
rect 38780 10500 38836 11676
rect 39004 11508 39060 11518
rect 39004 11414 39060 11452
rect 39116 11396 39172 13356
rect 39228 12852 39284 12862
rect 39228 12178 39284 12796
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 12114 39284 12126
rect 39452 12740 39508 12750
rect 39116 11330 39172 11340
rect 39340 12068 39396 12078
rect 39228 11172 39284 11182
rect 38668 10498 38836 10500
rect 38668 10446 38670 10498
rect 38722 10446 38836 10498
rect 38668 10444 38836 10446
rect 38892 11170 39284 11172
rect 38892 11118 39230 11170
rect 39282 11118 39284 11170
rect 38892 11116 39284 11118
rect 38668 10434 38724 10444
rect 38220 8930 38388 8932
rect 38220 8878 38222 8930
rect 38274 8878 38388 8930
rect 38220 8876 38388 8878
rect 38444 9602 38500 9614
rect 38444 9550 38446 9602
rect 38498 9550 38500 9602
rect 38444 9044 38500 9550
rect 38780 9380 38836 9390
rect 38220 8866 38276 8876
rect 38444 8708 38500 8988
rect 38668 9044 38724 9054
rect 38668 8950 38724 8988
rect 38220 8652 38500 8708
rect 38220 7474 38276 8652
rect 38332 8372 38388 8382
rect 38388 8316 38500 8372
rect 38332 8278 38388 8316
rect 38220 7422 38222 7474
rect 38274 7422 38276 7474
rect 38220 7410 38276 7422
rect 38444 7476 38500 8316
rect 38444 7410 38500 7420
rect 38780 7474 38836 9324
rect 38780 7422 38782 7474
rect 38834 7422 38836 7474
rect 38780 7410 38836 7422
rect 38892 7362 38948 11116
rect 39228 11106 39284 11116
rect 38892 7310 38894 7362
rect 38946 7310 38948 7362
rect 38892 7298 38948 7310
rect 39004 10948 39060 10958
rect 38108 7196 38388 7252
rect 37996 6578 38052 6590
rect 37996 6526 37998 6578
rect 38050 6526 38052 6578
rect 37996 6356 38052 6526
rect 37996 6290 38052 6300
rect 38108 5908 38164 5918
rect 37884 5682 37940 5694
rect 37884 5630 37886 5682
rect 37938 5630 37940 5682
rect 37884 5124 37940 5630
rect 37884 5058 37940 5068
rect 37996 5012 38052 5022
rect 37996 4562 38052 4956
rect 37996 4510 37998 4562
rect 38050 4510 38052 4562
rect 37996 4498 38052 4510
rect 38108 4452 38164 5852
rect 38332 5124 38388 7196
rect 38444 6804 38500 6814
rect 38444 6710 38500 6748
rect 39004 6130 39060 10892
rect 39340 10388 39396 12012
rect 39340 10322 39396 10332
rect 39452 10276 39508 12684
rect 39676 12068 39732 13916
rect 39788 13746 39844 13758
rect 39788 13694 39790 13746
rect 39842 13694 39844 13746
rect 39788 12740 39844 13694
rect 39788 12674 39844 12684
rect 39676 12002 39732 12012
rect 39788 12066 39844 12078
rect 39788 12014 39790 12066
rect 39842 12014 39844 12066
rect 39564 11172 39620 11182
rect 39564 11170 39732 11172
rect 39564 11118 39566 11170
rect 39618 11118 39732 11170
rect 39564 11116 39732 11118
rect 39564 11106 39620 11116
rect 39452 10220 39620 10276
rect 39452 9604 39508 9614
rect 39452 9268 39508 9548
rect 39452 9042 39508 9212
rect 39452 8990 39454 9042
rect 39506 8990 39508 9042
rect 39452 8978 39508 8990
rect 39340 7476 39396 7486
rect 39564 7476 39620 10220
rect 39676 7588 39732 11116
rect 39788 10834 39844 12014
rect 39788 10782 39790 10834
rect 39842 10782 39844 10834
rect 39788 10770 39844 10782
rect 39900 10500 39956 21196
rect 40124 18116 40180 24444
rect 40348 23714 40404 23726
rect 40348 23662 40350 23714
rect 40402 23662 40404 23714
rect 40348 23604 40404 23662
rect 40236 23548 40404 23604
rect 40236 23492 40292 23548
rect 40236 23426 40292 23436
rect 40236 23156 40292 23166
rect 40236 23062 40292 23100
rect 40460 22484 40516 22494
rect 40460 22390 40516 22428
rect 40348 22146 40404 22158
rect 40348 22094 40350 22146
rect 40402 22094 40404 22146
rect 40348 21700 40404 22094
rect 40572 22036 40628 25228
rect 41020 24164 41076 25340
rect 41132 24948 41188 25454
rect 41244 25396 41300 25406
rect 41356 25396 41412 26126
rect 41468 25844 41524 25854
rect 41468 25506 41524 25788
rect 41468 25454 41470 25506
rect 41522 25454 41524 25506
rect 41468 25442 41524 25454
rect 41244 25394 41412 25396
rect 41244 25342 41246 25394
rect 41298 25342 41412 25394
rect 41244 25340 41412 25342
rect 41580 25396 41636 26572
rect 41692 26180 41748 27020
rect 42028 27076 42084 28366
rect 42140 27748 42196 28924
rect 42364 28308 42420 30158
rect 42476 29876 42532 31724
rect 42588 30884 42644 32732
rect 43260 32452 43316 33628
rect 43932 33572 43988 33582
rect 43932 33348 43988 33516
rect 43932 33282 43988 33292
rect 44044 33348 44100 33358
rect 44156 33348 44212 34636
rect 44268 34626 44324 34636
rect 44380 34132 44436 34860
rect 44380 34066 44436 34076
rect 44716 34804 44772 34814
rect 44716 34018 44772 34748
rect 44828 34132 44884 35084
rect 44828 34038 44884 34076
rect 44940 35140 44996 36318
rect 45276 36594 45332 36606
rect 45276 36542 45278 36594
rect 45330 36542 45332 36594
rect 45276 35700 45332 36542
rect 45276 35364 45332 35644
rect 45388 36372 45444 36382
rect 45388 35586 45444 36316
rect 45500 35812 45556 38612
rect 45836 38610 46004 38612
rect 45836 38558 45950 38610
rect 46002 38558 46004 38610
rect 45836 38556 46004 38558
rect 45612 38052 45668 38062
rect 45836 38052 45892 38556
rect 45948 38546 46004 38556
rect 45612 38050 45892 38052
rect 45612 37998 45614 38050
rect 45666 37998 45892 38050
rect 45612 37996 45892 37998
rect 45612 37986 45668 37996
rect 45948 37940 46004 37950
rect 45948 37846 46004 37884
rect 45612 37268 45668 37278
rect 45612 37266 45780 37268
rect 45612 37214 45614 37266
rect 45666 37214 45780 37266
rect 45612 37212 45780 37214
rect 45612 37202 45668 37212
rect 45500 35746 45556 35756
rect 45388 35534 45390 35586
rect 45442 35534 45444 35586
rect 45388 35522 45444 35534
rect 45500 35476 45556 35486
rect 45276 35308 45444 35364
rect 45052 35140 45108 35150
rect 44940 35084 45052 35140
rect 44716 33966 44718 34018
rect 44770 33966 44772 34018
rect 44716 33908 44772 33966
rect 44716 33852 44884 33908
rect 44044 33346 44212 33348
rect 44044 33294 44046 33346
rect 44098 33294 44212 33346
rect 44044 33292 44212 33294
rect 44268 33796 44324 33806
rect 44044 33282 44100 33292
rect 43596 33234 43652 33246
rect 43596 33182 43598 33234
rect 43650 33182 43652 33234
rect 43260 32116 43316 32396
rect 43148 32060 43316 32116
rect 43372 32900 43428 32910
rect 42812 31778 42868 31790
rect 42812 31726 42814 31778
rect 42866 31726 42868 31778
rect 42812 31218 42868 31726
rect 42812 31166 42814 31218
rect 42866 31166 42868 31218
rect 42812 31154 42868 31166
rect 42588 30818 42644 30828
rect 42476 29810 42532 29820
rect 42364 28242 42420 28252
rect 42700 29204 42756 29214
rect 42700 28530 42756 29148
rect 43148 28980 43204 32060
rect 43260 31780 43316 31790
rect 43260 31686 43316 31724
rect 43260 31444 43316 31454
rect 43260 30210 43316 31388
rect 43260 30158 43262 30210
rect 43314 30158 43316 30210
rect 43260 30146 43316 30158
rect 43148 28914 43204 28924
rect 43372 28980 43428 32844
rect 43484 32564 43540 32574
rect 43484 32470 43540 32508
rect 43596 32116 43652 33182
rect 44268 33012 44324 33740
rect 44464 33740 44728 33750
rect 44520 33684 44568 33740
rect 44624 33684 44672 33740
rect 44464 33674 44728 33684
rect 44828 33684 44884 33852
rect 44828 33618 44884 33628
rect 44604 33458 44660 33470
rect 44604 33406 44606 33458
rect 44658 33406 44660 33458
rect 44380 33348 44436 33358
rect 44380 33254 44436 33292
rect 43804 32956 44068 32966
rect 43860 32900 43908 32956
rect 43964 32900 44012 32956
rect 44268 32946 44324 32956
rect 43804 32890 44068 32900
rect 44380 32674 44436 32686
rect 44380 32622 44382 32674
rect 44434 32622 44436 32674
rect 43596 31892 43652 32060
rect 43596 31826 43652 31836
rect 44268 32564 44324 32574
rect 44380 32564 44436 32622
rect 44492 32564 44548 32574
rect 44380 32508 44492 32564
rect 44268 32340 44324 32508
rect 44492 32498 44548 32508
rect 44604 32340 44660 33406
rect 44940 32564 44996 35084
rect 45052 35074 45108 35084
rect 45276 34132 45332 34142
rect 45164 34130 45332 34132
rect 45164 34078 45278 34130
rect 45330 34078 45332 34130
rect 45164 34076 45332 34078
rect 45052 33796 45108 33806
rect 45052 33572 45108 33740
rect 45052 33506 45108 33516
rect 44940 32498 44996 32508
rect 45052 33012 45108 33022
rect 44268 32284 44660 32340
rect 44828 32338 44884 32350
rect 44828 32286 44830 32338
rect 44882 32286 44884 32338
rect 44268 31778 44324 32284
rect 44464 32172 44728 32182
rect 44520 32116 44568 32172
rect 44624 32116 44672 32172
rect 44464 32106 44728 32116
rect 44268 31726 44270 31778
rect 44322 31726 44324 31778
rect 44268 31714 44324 31726
rect 44492 31556 44548 31566
rect 43804 31388 44068 31398
rect 43860 31332 43908 31388
rect 43964 31332 44012 31388
rect 43804 31322 44068 31332
rect 43484 31220 43540 31230
rect 43484 31106 43540 31164
rect 43484 31054 43486 31106
rect 43538 31054 43540 31106
rect 43484 31042 43540 31054
rect 44156 30884 44212 30894
rect 44380 30884 44436 30894
rect 43596 30772 43652 30782
rect 43596 30678 43652 30716
rect 43804 29820 44068 29830
rect 43860 29764 43908 29820
rect 43964 29764 44012 29820
rect 43804 29754 44068 29764
rect 44156 29764 44212 30828
rect 44156 29698 44212 29708
rect 44268 30882 44436 30884
rect 44268 30830 44382 30882
rect 44434 30830 44436 30882
rect 44268 30828 44436 30830
rect 44268 30212 44324 30828
rect 44380 30818 44436 30828
rect 44492 30882 44548 31500
rect 44492 30830 44494 30882
rect 44546 30830 44548 30882
rect 44492 30818 44548 30830
rect 44716 30884 44772 30894
rect 44716 30790 44772 30828
rect 44464 30604 44728 30614
rect 44520 30548 44568 30604
rect 44624 30548 44672 30604
rect 44464 30538 44728 30548
rect 44268 29428 44324 30156
rect 44492 30324 44548 30334
rect 44492 30210 44548 30268
rect 44492 30158 44494 30210
rect 44546 30158 44548 30210
rect 44492 30146 44548 30158
rect 44268 29362 44324 29372
rect 44268 29202 44324 29214
rect 44268 29150 44270 29202
rect 44322 29150 44324 29202
rect 43372 28914 43428 28924
rect 43484 29092 43540 29102
rect 43148 28644 43204 28654
rect 43148 28642 43428 28644
rect 43148 28590 43150 28642
rect 43202 28590 43428 28642
rect 43148 28588 43428 28590
rect 43148 28578 43204 28588
rect 42700 28478 42702 28530
rect 42754 28478 42756 28530
rect 42588 28084 42644 28094
rect 42140 27746 42420 27748
rect 42140 27694 42142 27746
rect 42194 27694 42420 27746
rect 42140 27692 42420 27694
rect 42140 27682 42196 27692
rect 42252 27188 42308 27198
rect 42252 27094 42308 27132
rect 42028 27010 42084 27020
rect 42364 26908 42420 27692
rect 42140 26852 42196 26862
rect 41692 26114 41748 26124
rect 41804 26850 42196 26852
rect 41804 26798 42142 26850
rect 42194 26798 42196 26850
rect 41804 26796 42196 26798
rect 41804 25732 41860 26796
rect 42140 26786 42196 26796
rect 42252 26852 42420 26908
rect 42252 26404 42308 26852
rect 42252 26348 42420 26404
rect 41916 26180 41972 26190
rect 42252 26180 42308 26190
rect 41916 26178 42308 26180
rect 41916 26126 41918 26178
rect 41970 26126 42254 26178
rect 42306 26126 42308 26178
rect 41916 26124 42308 26126
rect 41916 26114 41972 26124
rect 42252 26114 42308 26124
rect 41916 25732 41972 25742
rect 41860 25730 41972 25732
rect 41860 25678 41918 25730
rect 41970 25678 41972 25730
rect 41860 25676 41972 25678
rect 41804 25638 41860 25676
rect 41916 25508 41972 25676
rect 42028 25732 42084 25742
rect 42028 25638 42084 25676
rect 41916 25452 42084 25508
rect 41244 25330 41300 25340
rect 41580 25330 41636 25340
rect 41804 25284 41860 25294
rect 41580 25060 41636 25070
rect 41244 24948 41300 24958
rect 41132 24946 41300 24948
rect 41132 24894 41246 24946
rect 41298 24894 41300 24946
rect 41132 24892 41300 24894
rect 41244 24882 41300 24892
rect 41020 24098 41076 24108
rect 41356 24612 41412 24622
rect 40796 23604 40852 23614
rect 40796 22482 40852 23548
rect 41356 23604 41412 24556
rect 41468 24276 41524 24286
rect 41468 24162 41524 24220
rect 41468 24110 41470 24162
rect 41522 24110 41524 24162
rect 41468 23940 41524 24110
rect 41468 23874 41524 23884
rect 41356 23154 41412 23548
rect 41356 23102 41358 23154
rect 41410 23102 41412 23154
rect 41356 23090 41412 23102
rect 41580 23044 41636 25004
rect 41692 24610 41748 24622
rect 41692 24558 41694 24610
rect 41746 24558 41748 24610
rect 41692 24500 41748 24558
rect 41692 24434 41748 24444
rect 41580 22978 41636 22988
rect 41692 24276 41748 24286
rect 41580 22708 41636 22718
rect 41692 22708 41748 24220
rect 41804 24052 41860 25228
rect 41916 24836 41972 24846
rect 41916 24742 41972 24780
rect 42028 24722 42084 25452
rect 42140 25506 42196 25518
rect 42140 25454 42142 25506
rect 42194 25454 42196 25506
rect 42140 25060 42196 25454
rect 42140 24994 42196 25004
rect 42028 24670 42030 24722
rect 42082 24670 42084 24722
rect 42028 24658 42084 24670
rect 41804 23986 41860 23996
rect 41916 24164 41972 24174
rect 41916 23826 41972 24108
rect 41916 23774 41918 23826
rect 41970 23774 41972 23826
rect 41916 23548 41972 23774
rect 41636 22652 41748 22708
rect 41804 23492 41972 23548
rect 41580 22642 41636 22652
rect 41468 22538 41524 22550
rect 40796 22430 40798 22482
rect 40850 22430 40852 22482
rect 40796 22418 40852 22430
rect 41020 22482 41076 22494
rect 41468 22486 41470 22538
rect 41522 22486 41524 22538
rect 41468 22484 41524 22486
rect 41020 22430 41022 22482
rect 41074 22430 41076 22482
rect 40460 21980 40628 22036
rect 40908 22258 40964 22270
rect 40908 22206 40910 22258
rect 40962 22206 40964 22258
rect 40460 21924 40516 21980
rect 40908 21924 40964 22206
rect 40460 21858 40516 21868
rect 40572 21868 40964 21924
rect 40572 21810 40628 21868
rect 40572 21758 40574 21810
rect 40626 21758 40628 21810
rect 40572 21746 40628 21758
rect 40348 21634 40404 21644
rect 40572 21588 40628 21598
rect 40460 21586 40628 21588
rect 40460 21534 40574 21586
rect 40626 21534 40628 21586
rect 40460 21532 40628 21534
rect 40236 21474 40292 21486
rect 40236 21422 40238 21474
rect 40290 21422 40292 21474
rect 40236 20692 40292 21422
rect 40236 20626 40292 20636
rect 40348 20916 40404 20926
rect 40460 20916 40516 21532
rect 40572 21522 40628 21532
rect 40908 21476 40964 21486
rect 40796 21362 40852 21374
rect 40796 21310 40798 21362
rect 40850 21310 40852 21362
rect 40796 21028 40852 21310
rect 40796 20962 40852 20972
rect 40348 20914 40516 20916
rect 40348 20862 40350 20914
rect 40402 20862 40516 20914
rect 40348 20860 40516 20862
rect 40684 20916 40740 20926
rect 40348 20804 40404 20860
rect 40684 20822 40740 20860
rect 40348 19796 40404 20748
rect 40572 20802 40628 20814
rect 40572 20750 40574 20802
rect 40626 20750 40628 20802
rect 40572 20692 40628 20750
rect 40796 20804 40852 20814
rect 40796 20710 40852 20748
rect 40572 20626 40628 20636
rect 40908 20580 40964 21420
rect 40908 20514 40964 20524
rect 41020 20692 41076 22430
rect 41356 22428 41524 22484
rect 41580 22484 41636 22494
rect 41804 22484 41860 23492
rect 41916 23426 41972 23436
rect 42028 23940 42084 23950
rect 41916 23156 41972 23166
rect 41916 22708 41972 23100
rect 41916 22642 41972 22652
rect 42028 22484 42084 23884
rect 41580 22482 41748 22484
rect 41580 22430 41582 22482
rect 41634 22430 41748 22482
rect 41580 22428 41748 22430
rect 41804 22428 41972 22484
rect 41356 22260 41412 22428
rect 41580 22418 41636 22428
rect 41132 22204 41412 22260
rect 41692 22260 41748 22428
rect 41692 22204 41860 22260
rect 41132 21476 41188 22204
rect 41580 22146 41636 22158
rect 41580 22094 41582 22146
rect 41634 22094 41636 22146
rect 41580 22078 41636 22094
rect 41132 21410 41188 21420
rect 41244 22022 41636 22078
rect 40908 19796 40964 19806
rect 40348 19794 40964 19796
rect 40348 19742 40910 19794
rect 40962 19742 40964 19794
rect 40348 19740 40964 19742
rect 40124 18050 40180 18060
rect 40460 19236 40516 19246
rect 40460 17892 40516 19180
rect 40572 19124 40628 19134
rect 40572 19030 40628 19068
rect 40572 18676 40628 18686
rect 40572 18582 40628 18620
rect 40572 18452 40628 18462
rect 40796 18452 40852 19740
rect 40908 19730 40964 19740
rect 41020 19572 41076 20636
rect 41132 21140 41188 21150
rect 41132 20356 41188 21084
rect 41244 21026 41300 22022
rect 41356 21812 41412 21822
rect 41356 21698 41412 21756
rect 41804 21700 41860 22204
rect 41916 21812 41972 22428
rect 42028 22418 42084 22428
rect 42140 22258 42196 22270
rect 42140 22206 42142 22258
rect 42194 22206 42196 22258
rect 42140 21924 42196 22206
rect 42140 21858 42196 21868
rect 41916 21746 41972 21756
rect 42364 21812 42420 26348
rect 42476 26178 42532 26190
rect 42476 26126 42478 26178
rect 42530 26126 42532 26178
rect 42476 25732 42532 26126
rect 42476 25666 42532 25676
rect 42476 25282 42532 25294
rect 42476 25230 42478 25282
rect 42530 25230 42532 25282
rect 42476 24836 42532 25230
rect 42476 24770 42532 24780
rect 42588 24612 42644 28028
rect 42700 26908 42756 28478
rect 43372 28082 43428 28588
rect 43372 28030 43374 28082
rect 43426 28030 43428 28082
rect 43372 28018 43428 28030
rect 43484 28642 43540 29036
rect 43708 28756 43764 28766
rect 43708 28662 43764 28700
rect 43484 28590 43486 28642
rect 43538 28590 43540 28642
rect 43484 27524 43540 28590
rect 44268 28642 44324 29150
rect 44464 29036 44728 29046
rect 44520 28980 44568 29036
rect 44624 28980 44672 29036
rect 44464 28970 44728 28980
rect 44268 28590 44270 28642
rect 44322 28590 44324 28642
rect 44268 28578 44324 28590
rect 44716 28642 44772 28654
rect 44716 28590 44718 28642
rect 44770 28590 44772 28642
rect 44604 28532 44660 28542
rect 43484 27458 43540 27468
rect 43596 28420 43652 28430
rect 43260 27188 43316 27198
rect 42812 27076 42868 27114
rect 42812 27010 42868 27020
rect 43260 26964 43316 27132
rect 42700 26852 42868 26908
rect 43260 26898 43316 26908
rect 43596 26964 43652 28364
rect 44268 28420 44324 28430
rect 43804 28252 44068 28262
rect 43860 28196 43908 28252
rect 43964 28196 44012 28252
rect 43804 28186 44068 28196
rect 43596 26898 43652 26908
rect 44156 27524 44212 27534
rect 42700 26066 42756 26078
rect 42700 26014 42702 26066
rect 42754 26014 42756 26066
rect 42700 25844 42756 26014
rect 42812 26068 42868 26852
rect 43148 26852 43204 26862
rect 43148 26514 43204 26796
rect 43804 26684 44068 26694
rect 43860 26628 43908 26684
rect 43964 26628 44012 26684
rect 43804 26618 44068 26628
rect 43148 26462 43150 26514
rect 43202 26462 43204 26514
rect 43148 26450 43204 26462
rect 43596 26516 43652 26526
rect 44156 26516 44212 27468
rect 42924 26292 42980 26302
rect 43260 26292 43316 26302
rect 42924 26290 43316 26292
rect 42924 26238 42926 26290
rect 42978 26238 43262 26290
rect 43314 26238 43316 26290
rect 42924 26236 43316 26238
rect 42924 26226 42980 26236
rect 43260 26226 43316 26236
rect 43372 26180 43428 26190
rect 43372 26086 43428 26124
rect 43260 26068 43316 26078
rect 42812 26012 42980 26068
rect 42924 25844 42980 26012
rect 43260 25956 43316 26012
rect 43484 26068 43540 26078
rect 43260 25900 43428 25956
rect 42700 25788 42868 25844
rect 42924 25788 43204 25844
rect 42700 25620 42756 25658
rect 42700 25554 42756 25564
rect 42700 25396 42756 25406
rect 42812 25396 42868 25788
rect 43148 25618 43204 25788
rect 43148 25566 43150 25618
rect 43202 25566 43204 25618
rect 43148 25554 43204 25566
rect 43036 25508 43092 25518
rect 42924 25396 42980 25406
rect 42812 25340 42924 25396
rect 42700 25302 42756 25340
rect 42924 25330 42980 25340
rect 42476 24556 42644 24612
rect 42476 22148 42532 24556
rect 42700 23826 42756 23838
rect 42700 23774 42702 23826
rect 42754 23774 42756 23826
rect 42700 23492 42756 23774
rect 42700 23426 42756 23436
rect 42924 23044 42980 23054
rect 42588 22372 42644 22382
rect 42588 22370 42868 22372
rect 42588 22318 42590 22370
rect 42642 22318 42868 22370
rect 42588 22316 42868 22318
rect 42588 22306 42644 22316
rect 42476 22092 42756 22148
rect 42364 21746 42420 21756
rect 41356 21646 41358 21698
rect 41410 21646 41412 21698
rect 41356 21634 41412 21646
rect 41580 21644 41860 21700
rect 41244 20974 41246 21026
rect 41298 20974 41300 21026
rect 41244 20962 41300 20974
rect 41356 21476 41412 21486
rect 41356 21026 41412 21420
rect 41356 20974 41358 21026
rect 41410 20974 41412 21026
rect 41356 20962 41412 20974
rect 41468 21028 41524 21038
rect 41468 20934 41524 20972
rect 41468 20804 41524 20814
rect 41132 20290 41188 20300
rect 41244 20580 41300 20590
rect 40572 18450 40852 18452
rect 40572 18398 40574 18450
rect 40626 18398 40852 18450
rect 40572 18396 40852 18398
rect 40908 19516 41076 19572
rect 41132 19908 41188 19918
rect 40908 18450 40964 19516
rect 41020 19348 41076 19358
rect 41132 19348 41188 19852
rect 41020 19346 41188 19348
rect 41020 19294 41022 19346
rect 41074 19294 41188 19346
rect 41020 19292 41188 19294
rect 41020 18788 41076 19292
rect 41020 18722 41076 18732
rect 41132 19124 41188 19134
rect 41020 18564 41076 18574
rect 41132 18564 41188 19068
rect 41244 18900 41300 20524
rect 41468 20130 41524 20748
rect 41468 20078 41470 20130
rect 41522 20078 41524 20130
rect 41468 20066 41524 20078
rect 41580 20802 41636 21644
rect 41804 21362 41860 21374
rect 41804 21310 41806 21362
rect 41858 21310 41860 21362
rect 41804 21140 41860 21310
rect 41804 21074 41860 21084
rect 41580 20750 41582 20802
rect 41634 20750 41636 20802
rect 41356 20020 41412 20030
rect 41356 19926 41412 19964
rect 41580 19460 41636 20750
rect 42364 20804 42420 20814
rect 42364 20710 42420 20748
rect 42588 20690 42644 20702
rect 42588 20638 42590 20690
rect 42642 20638 42644 20690
rect 41916 20580 41972 20590
rect 42140 20580 42196 20590
rect 42588 20580 42644 20638
rect 41916 20578 42084 20580
rect 41916 20526 41918 20578
rect 41970 20526 42084 20578
rect 41916 20524 42084 20526
rect 41916 20514 41972 20524
rect 41580 19394 41636 19404
rect 41916 20356 41972 20366
rect 41244 18834 41300 18844
rect 41804 19012 41860 19022
rect 41020 18562 41188 18564
rect 41020 18510 41022 18562
rect 41074 18510 41188 18562
rect 41020 18508 41188 18510
rect 41020 18498 41076 18508
rect 40908 18398 40910 18450
rect 40962 18398 40964 18450
rect 40572 18386 40628 18396
rect 40908 18386 40964 18398
rect 41580 18452 41636 18462
rect 41580 18358 41636 18396
rect 41132 18338 41188 18350
rect 41132 18286 41134 18338
rect 41186 18286 41188 18338
rect 40796 18004 40852 18014
rect 40460 17836 40740 17892
rect 40572 17668 40628 17678
rect 40348 17666 40628 17668
rect 40348 17614 40574 17666
rect 40626 17614 40628 17666
rect 40348 17612 40628 17614
rect 40236 17554 40292 17566
rect 40236 17502 40238 17554
rect 40290 17502 40292 17554
rect 40236 15988 40292 17502
rect 40348 17106 40404 17612
rect 40572 17602 40628 17612
rect 40348 17054 40350 17106
rect 40402 17054 40404 17106
rect 40348 17042 40404 17054
rect 40572 16324 40628 16334
rect 40684 16324 40740 17836
rect 40572 16322 40740 16324
rect 40572 16270 40574 16322
rect 40626 16270 40740 16322
rect 40572 16268 40740 16270
rect 40572 16258 40628 16268
rect 40236 15922 40292 15932
rect 40460 15988 40516 15998
rect 40460 15894 40516 15932
rect 40796 15764 40852 17948
rect 41020 17668 41076 17678
rect 41020 17220 41076 17612
rect 41020 17154 41076 17164
rect 40348 15708 40852 15764
rect 40908 16884 40964 16894
rect 40908 16100 40964 16828
rect 41020 16100 41076 16110
rect 40908 16098 41076 16100
rect 40908 16046 41022 16098
rect 41074 16046 41076 16098
rect 40908 16044 41076 16046
rect 40236 15652 40292 15662
rect 40236 13636 40292 15596
rect 40124 13634 40292 13636
rect 40124 13582 40238 13634
rect 40290 13582 40292 13634
rect 40124 13580 40292 13582
rect 40124 11172 40180 13580
rect 40236 13570 40292 13580
rect 40236 12852 40292 12862
rect 40236 12758 40292 12796
rect 40348 12178 40404 15708
rect 40460 15316 40516 15326
rect 40684 15316 40740 15326
rect 40516 15260 40628 15316
rect 40460 15250 40516 15260
rect 40572 14196 40628 15260
rect 40684 15222 40740 15260
rect 40348 12126 40350 12178
rect 40402 12126 40404 12178
rect 40236 11954 40292 11966
rect 40236 11902 40238 11954
rect 40290 11902 40292 11954
rect 40236 11284 40292 11902
rect 40348 11620 40404 12126
rect 40348 11554 40404 11564
rect 40460 13524 40516 13534
rect 40236 11218 40292 11228
rect 40124 11106 40180 11116
rect 40460 10612 40516 13468
rect 40460 10546 40516 10556
rect 39900 10434 39956 10444
rect 40124 10500 40180 10510
rect 39900 9044 39956 9054
rect 39900 8372 39956 8988
rect 39900 8306 39956 8316
rect 39676 7532 39844 7588
rect 39564 7420 39732 7476
rect 39340 7382 39396 7420
rect 39564 6692 39620 6702
rect 39564 6598 39620 6636
rect 39004 6078 39006 6130
rect 39058 6078 39060 6130
rect 39004 6066 39060 6078
rect 39676 6356 39732 7420
rect 39676 6018 39732 6300
rect 39676 5966 39678 6018
rect 39730 5966 39732 6018
rect 39676 5954 39732 5966
rect 39004 5908 39060 5918
rect 39004 5906 39284 5908
rect 39004 5854 39006 5906
rect 39058 5854 39284 5906
rect 39004 5852 39284 5854
rect 39004 5842 39060 5852
rect 38668 5794 38724 5806
rect 38668 5742 38670 5794
rect 38722 5742 38724 5794
rect 38444 5684 38500 5694
rect 38444 5346 38500 5628
rect 38444 5294 38446 5346
rect 38498 5294 38500 5346
rect 38444 5282 38500 5294
rect 38668 5348 38724 5742
rect 38668 5292 38836 5348
rect 38332 5068 38500 5124
rect 38108 4386 38164 4396
rect 38220 5010 38276 5022
rect 38220 4958 38222 5010
rect 38274 4958 38276 5010
rect 38220 4226 38276 4958
rect 38332 4452 38388 4462
rect 38332 4358 38388 4396
rect 38220 4174 38222 4226
rect 38274 4174 38276 4226
rect 37996 3780 38052 3790
rect 37996 3686 38052 3724
rect 37884 3444 37940 3482
rect 37884 3378 37940 3388
rect 38220 3220 38276 4174
rect 37884 3164 38276 3220
rect 37884 2324 37940 3164
rect 37996 2548 38052 2558
rect 37996 2454 38052 2492
rect 38332 2546 38388 2558
rect 38332 2494 38334 2546
rect 38386 2494 38388 2546
rect 37884 2258 37940 2268
rect 38220 2212 38276 2222
rect 38220 2118 38276 2156
rect 37884 2100 37940 2110
rect 37884 2006 37940 2044
rect 37772 1820 38276 1876
rect 37660 1204 37716 1214
rect 37660 1110 37716 1148
rect 37884 1148 38164 1204
rect 37324 978 37380 990
rect 37324 926 37326 978
rect 37378 926 37380 978
rect 37324 868 37380 926
rect 37324 802 37380 812
rect 37436 980 37492 990
rect 37212 354 37268 364
rect 37436 112 37492 924
rect 37884 112 37940 1148
rect 37996 978 38052 990
rect 37996 926 37998 978
rect 38050 926 38052 978
rect 37996 308 38052 926
rect 38108 980 38164 1148
rect 38220 1202 38276 1820
rect 38220 1150 38222 1202
rect 38274 1150 38276 1202
rect 38220 1138 38276 1150
rect 38332 980 38388 2494
rect 38444 2212 38500 5068
rect 38668 5122 38724 5134
rect 38668 5070 38670 5122
rect 38722 5070 38724 5122
rect 38556 5012 38612 5022
rect 38556 4918 38612 4956
rect 38668 4900 38724 5070
rect 38668 3780 38724 4844
rect 38780 4452 38836 5292
rect 39228 5346 39284 5852
rect 39228 5294 39230 5346
rect 39282 5294 39284 5346
rect 39228 5282 39284 5294
rect 39340 5684 39396 5694
rect 39340 5346 39396 5628
rect 39340 5294 39342 5346
rect 39394 5294 39396 5346
rect 39340 5282 39396 5294
rect 39116 4900 39172 4910
rect 39116 4806 39172 4844
rect 38780 4386 38836 4396
rect 39788 4338 39844 7532
rect 39900 7476 39956 7486
rect 39900 7382 39956 7420
rect 40124 5796 40180 10444
rect 40348 9714 40404 9726
rect 40348 9662 40350 9714
rect 40402 9662 40404 9714
rect 40348 9492 40404 9662
rect 40348 9426 40404 9436
rect 40460 9602 40516 9614
rect 40460 9550 40462 9602
rect 40514 9550 40516 9602
rect 40236 9042 40292 9054
rect 40236 8990 40238 9042
rect 40290 8990 40292 9042
rect 40236 8708 40292 8990
rect 40236 8642 40292 8652
rect 40460 7700 40516 9550
rect 40460 7634 40516 7644
rect 40572 7476 40628 14140
rect 40908 13748 40964 16044
rect 41020 16034 41076 16044
rect 41132 15540 41188 18286
rect 41244 17778 41300 17790
rect 41244 17726 41246 17778
rect 41298 17726 41300 17778
rect 41244 17444 41300 17726
rect 41244 17378 41300 17388
rect 41468 17780 41524 17790
rect 41468 17220 41524 17724
rect 41468 17154 41524 17164
rect 41468 16660 41524 16670
rect 41468 16658 41636 16660
rect 41468 16606 41470 16658
rect 41522 16606 41636 16658
rect 41468 16604 41636 16606
rect 41468 16594 41524 16604
rect 41468 16436 41524 16446
rect 41468 16210 41524 16380
rect 41468 16158 41470 16210
rect 41522 16158 41524 16210
rect 41468 16146 41524 16158
rect 41132 15474 41188 15484
rect 41580 15988 41636 16604
rect 41244 15090 41300 15102
rect 41244 15038 41246 15090
rect 41298 15038 41300 15090
rect 41020 14868 41076 14878
rect 41020 14642 41076 14812
rect 41020 14590 41022 14642
rect 41074 14590 41076 14642
rect 41020 14578 41076 14590
rect 41244 14532 41300 15038
rect 41356 14532 41412 14542
rect 41244 14530 41412 14532
rect 41244 14478 41358 14530
rect 41410 14478 41412 14530
rect 41244 14476 41412 14478
rect 41356 14466 41412 14476
rect 41580 14532 41636 15932
rect 41804 15428 41860 18956
rect 41916 18228 41972 20300
rect 42028 19124 42084 20524
rect 42140 20578 42644 20580
rect 42140 20526 42142 20578
rect 42194 20526 42644 20578
rect 42140 20524 42644 20526
rect 42140 20514 42196 20524
rect 42700 20468 42756 22092
rect 42812 21812 42868 22316
rect 42924 22370 42980 22988
rect 42924 22318 42926 22370
rect 42978 22318 42980 22370
rect 42924 22306 42980 22318
rect 43036 22260 43092 25452
rect 43260 25508 43316 25518
rect 43260 25060 43316 25452
rect 43260 24994 43316 25004
rect 43148 24052 43204 24062
rect 43148 22820 43204 23996
rect 43148 22754 43204 22764
rect 43036 22194 43092 22204
rect 43148 22482 43204 22494
rect 43148 22430 43150 22482
rect 43202 22430 43204 22482
rect 43036 21924 43092 21934
rect 42924 21812 42980 21822
rect 42812 21810 42980 21812
rect 42812 21758 42926 21810
rect 42978 21758 42980 21810
rect 42812 21756 42980 21758
rect 42924 21746 42980 21756
rect 42924 21252 42980 21262
rect 43036 21252 43092 21868
rect 43148 21476 43204 22430
rect 43148 21410 43204 21420
rect 43036 21196 43204 21252
rect 42812 20802 42868 20814
rect 42812 20750 42814 20802
rect 42866 20750 42868 20802
rect 42812 20692 42868 20750
rect 42812 20626 42868 20636
rect 42476 20412 42756 20468
rect 42140 19908 42196 19918
rect 42140 19906 42308 19908
rect 42140 19854 42142 19906
rect 42194 19854 42308 19906
rect 42140 19852 42308 19854
rect 42140 19842 42196 19852
rect 42140 19460 42196 19470
rect 42140 19366 42196 19404
rect 42028 19058 42084 19068
rect 42252 18452 42308 19852
rect 42364 19906 42420 19918
rect 42364 19854 42366 19906
rect 42418 19854 42420 19906
rect 42364 19460 42420 19854
rect 42364 19394 42420 19404
rect 42252 18386 42308 18396
rect 42364 19124 42420 19134
rect 41916 18162 41972 18172
rect 42140 18226 42196 18238
rect 42140 18174 42142 18226
rect 42194 18174 42196 18226
rect 42140 18116 42196 18174
rect 42140 18050 42196 18060
rect 41916 17666 41972 17678
rect 41916 17614 41918 17666
rect 41970 17614 41972 17666
rect 41916 17108 41972 17614
rect 42252 17668 42308 17678
rect 42364 17668 42420 19068
rect 42252 17666 42420 17668
rect 42252 17614 42254 17666
rect 42306 17614 42420 17666
rect 42252 17612 42420 17614
rect 42252 17578 42308 17612
rect 41916 17042 41972 17052
rect 42028 17522 42308 17578
rect 41804 15362 41860 15372
rect 41916 16100 41972 16110
rect 41580 14466 41636 14476
rect 41804 14530 41860 14542
rect 41804 14478 41806 14530
rect 41858 14478 41860 14530
rect 41804 14196 41860 14478
rect 41804 14130 41860 14140
rect 40908 13682 40964 13692
rect 41580 13748 41636 13758
rect 41468 13636 41524 13646
rect 41356 13524 41412 13534
rect 40684 13522 41412 13524
rect 40684 13470 41358 13522
rect 41410 13470 41412 13522
rect 40684 13468 41412 13470
rect 40684 12962 40740 13468
rect 41356 13458 41412 13468
rect 41244 13188 41300 13198
rect 41468 13188 41524 13580
rect 41244 13186 41524 13188
rect 41244 13134 41246 13186
rect 41298 13134 41524 13186
rect 41244 13132 41524 13134
rect 41244 13122 41300 13132
rect 40684 12910 40686 12962
rect 40738 12910 40740 12962
rect 40684 12898 40740 12910
rect 40908 13076 40964 13086
rect 40796 12180 40852 12190
rect 40796 12086 40852 12124
rect 40908 11998 40964 13020
rect 40796 11942 40964 11998
rect 41020 12964 41076 12974
rect 40796 9044 40852 11942
rect 41020 11732 41076 12908
rect 41020 11666 41076 11676
rect 41244 12066 41300 12078
rect 41244 12014 41246 12066
rect 41298 12014 41300 12066
rect 40908 11508 40964 11518
rect 40908 9266 40964 11452
rect 41132 11508 41188 11518
rect 41020 10612 41076 10622
rect 41020 9716 41076 10556
rect 41132 10276 41188 11452
rect 41132 10210 41188 10220
rect 41020 9714 41188 9716
rect 41020 9662 41022 9714
rect 41074 9662 41188 9714
rect 41020 9660 41188 9662
rect 41020 9650 41076 9660
rect 40908 9214 40910 9266
rect 40962 9214 40964 9266
rect 40908 9202 40964 9214
rect 41020 9380 41076 9390
rect 40796 8988 40964 9044
rect 40908 8596 40964 8988
rect 41020 8708 41076 9324
rect 41020 8642 41076 8652
rect 40796 8370 40852 8382
rect 40796 8318 40798 8370
rect 40850 8318 40852 8370
rect 40460 7420 40628 7476
rect 40684 8258 40740 8270
rect 40684 8206 40686 8258
rect 40738 8206 40740 8258
rect 40236 6580 40292 6590
rect 40236 6486 40292 6524
rect 40124 5702 40180 5740
rect 40348 5236 40404 5246
rect 40348 4450 40404 5180
rect 40460 5124 40516 7420
rect 40684 6916 40740 8206
rect 40796 8036 40852 8318
rect 40796 7970 40852 7980
rect 40908 7474 40964 8540
rect 41132 8596 41188 9660
rect 41132 8530 41188 8540
rect 41020 8260 41076 8270
rect 41020 8166 41076 8204
rect 40908 7422 40910 7474
rect 40962 7422 40964 7474
rect 40908 7410 40964 7422
rect 41244 7364 41300 12014
rect 41580 11788 41636 13692
rect 41692 12962 41748 12974
rect 41692 12910 41694 12962
rect 41746 12910 41748 12962
rect 41692 12402 41748 12910
rect 41692 12350 41694 12402
rect 41746 12350 41748 12402
rect 41692 12338 41748 12350
rect 41804 12516 41860 12526
rect 41580 11732 41748 11788
rect 41580 10610 41636 10622
rect 41580 10558 41582 10610
rect 41634 10558 41636 10610
rect 41468 10052 41524 10062
rect 41468 9958 41524 9996
rect 41580 8372 41636 10558
rect 41580 8306 41636 8316
rect 41356 8036 41412 8046
rect 41356 7942 41412 7980
rect 41692 7924 41748 11732
rect 41804 9940 41860 12460
rect 41804 9874 41860 9884
rect 41692 7858 41748 7868
rect 41804 8372 41860 8382
rect 41804 7474 41860 8316
rect 41804 7422 41806 7474
rect 41858 7422 41860 7474
rect 41244 7298 41300 7308
rect 41580 7364 41636 7374
rect 40684 6860 41188 6916
rect 41132 6804 41188 6860
rect 41244 6804 41300 6814
rect 41132 6802 41300 6804
rect 41132 6750 41246 6802
rect 41298 6750 41300 6802
rect 41132 6748 41300 6750
rect 40572 6692 40628 6702
rect 40572 6598 40628 6636
rect 40796 6692 40852 6702
rect 40460 5058 40516 5068
rect 40348 4398 40350 4450
rect 40402 4398 40404 4450
rect 40348 4386 40404 4398
rect 39788 4286 39790 4338
rect 39842 4286 39844 4338
rect 39788 4274 39844 4286
rect 40684 4338 40740 4350
rect 40684 4286 40686 4338
rect 40738 4286 40740 4338
rect 38668 3714 38724 3724
rect 40012 4114 40068 4126
rect 40012 4062 40014 4114
rect 40066 4062 40068 4114
rect 40012 3780 40068 4062
rect 40012 3714 40068 3724
rect 39676 3666 39732 3678
rect 39676 3614 39678 3666
rect 39730 3614 39732 3666
rect 39340 3556 39396 3566
rect 38892 3554 39396 3556
rect 38892 3502 39342 3554
rect 39394 3502 39396 3554
rect 38892 3500 39396 3502
rect 38556 2772 38612 2782
rect 38556 2678 38612 2716
rect 38556 2212 38612 2222
rect 38444 2210 38612 2212
rect 38444 2158 38558 2210
rect 38610 2158 38612 2210
rect 38444 2156 38612 2158
rect 38556 2146 38612 2156
rect 38892 2210 38948 3500
rect 39340 3490 39396 3500
rect 38892 2158 38894 2210
rect 38946 2158 38948 2210
rect 38892 2146 38948 2158
rect 39228 3332 39284 3342
rect 39228 2210 39284 3276
rect 39340 2772 39396 2782
rect 39340 2678 39396 2716
rect 39564 2548 39620 2558
rect 39228 2158 39230 2210
rect 39282 2158 39284 2210
rect 39228 2146 39284 2158
rect 39452 2546 39620 2548
rect 39452 2494 39566 2546
rect 39618 2494 39620 2546
rect 39452 2492 39620 2494
rect 39452 1540 39508 2492
rect 39564 2482 39620 2492
rect 39564 2100 39620 2110
rect 39564 2006 39620 2044
rect 39452 1474 39508 1484
rect 38108 924 38388 980
rect 38780 1428 38836 1438
rect 37996 242 38052 252
rect 38332 756 38388 766
rect 38332 112 38388 700
rect 38780 112 38836 1372
rect 39452 1204 39508 1214
rect 39452 1110 39508 1148
rect 39116 978 39172 990
rect 39116 926 39118 978
rect 39170 926 39172 978
rect 39116 532 39172 926
rect 39116 466 39172 476
rect 39228 420 39284 430
rect 39228 112 39284 364
rect 39676 112 39732 3614
rect 40572 3444 40628 3482
rect 40012 2996 40068 3006
rect 40012 2902 40068 2940
rect 40572 2772 40628 3388
rect 40684 2996 40740 4286
rect 40796 3388 40852 6636
rect 41020 6690 41076 6702
rect 41020 6638 41022 6690
rect 41074 6638 41076 6690
rect 41020 6468 41076 6638
rect 41020 6402 41076 6412
rect 41132 4900 41188 6748
rect 41244 6738 41300 6748
rect 41580 6804 41636 7308
rect 41804 7140 41860 7422
rect 41804 7074 41860 7084
rect 41580 6738 41636 6748
rect 41692 6690 41748 6702
rect 41692 6638 41694 6690
rect 41746 6638 41748 6690
rect 41244 6132 41300 6142
rect 41692 6132 41748 6638
rect 41244 6130 41748 6132
rect 41244 6078 41246 6130
rect 41298 6078 41748 6130
rect 41244 6076 41748 6078
rect 41244 6066 41300 6076
rect 41916 6020 41972 16044
rect 42028 14754 42084 17522
rect 42028 14702 42030 14754
rect 42082 14702 42084 14754
rect 42028 14690 42084 14702
rect 42140 16772 42196 16782
rect 42028 11508 42084 11518
rect 42028 11414 42084 11452
rect 42028 10500 42084 10510
rect 42028 10406 42084 10444
rect 42140 10164 42196 16716
rect 42364 16660 42420 16670
rect 42364 15316 42420 16604
rect 42364 15202 42420 15260
rect 42364 15150 42366 15202
rect 42418 15150 42420 15202
rect 42364 15138 42420 15150
rect 42476 15148 42532 20412
rect 42700 20020 42756 20030
rect 42588 19236 42644 19246
rect 42588 19142 42644 19180
rect 42700 19124 42756 19964
rect 42924 19796 42980 21196
rect 43036 20916 43092 20926
rect 43036 20822 43092 20860
rect 42924 19730 42980 19740
rect 43036 19794 43092 19806
rect 43036 19742 43038 19794
rect 43090 19742 43092 19794
rect 42700 19058 42756 19068
rect 42812 19460 42868 19470
rect 42812 18676 42868 19404
rect 43036 19460 43092 19742
rect 43036 19394 43092 19404
rect 43036 19234 43092 19246
rect 43036 19182 43038 19234
rect 43090 19182 43092 19234
rect 42588 17108 42644 17118
rect 42588 17014 42644 17052
rect 42700 16324 42756 16334
rect 42812 16324 42868 18620
rect 42924 19122 42980 19134
rect 42924 19070 42926 19122
rect 42978 19070 42980 19122
rect 42924 16882 42980 19070
rect 43036 18564 43092 19182
rect 43036 18498 43092 18508
rect 43148 18004 43204 21196
rect 43372 20020 43428 25900
rect 43484 23604 43540 26012
rect 43596 25506 43652 26460
rect 44044 26460 44212 26516
rect 43708 26180 43764 26190
rect 43708 25956 43764 26124
rect 43708 25890 43764 25900
rect 43596 25454 43598 25506
rect 43650 25454 43652 25506
rect 43596 25442 43652 25454
rect 44044 25620 44100 26460
rect 44044 25506 44100 25564
rect 44044 25454 44046 25506
rect 44098 25454 44100 25506
rect 44044 25442 44100 25454
rect 44156 25618 44212 25630
rect 44156 25566 44158 25618
rect 44210 25566 44212 25618
rect 44156 25508 44212 25566
rect 44156 25442 44212 25452
rect 44268 25284 44324 28364
rect 44492 28084 44548 28094
rect 44492 27970 44548 28028
rect 44604 28082 44660 28476
rect 44604 28030 44606 28082
rect 44658 28030 44660 28082
rect 44604 28018 44660 28030
rect 44716 28196 44772 28590
rect 44492 27918 44494 27970
rect 44546 27918 44548 27970
rect 44492 27906 44548 27918
rect 44716 27860 44772 28140
rect 44716 27794 44772 27804
rect 44464 27468 44728 27478
rect 44520 27412 44568 27468
rect 44624 27412 44672 27468
rect 44464 27402 44728 27412
rect 44380 26850 44436 26862
rect 44380 26798 44382 26850
rect 44434 26798 44436 26850
rect 44380 26516 44436 26798
rect 44380 26450 44436 26460
rect 44604 26292 44660 26302
rect 44604 26038 44660 26236
rect 44828 26292 44884 32286
rect 45052 32228 45108 32956
rect 45052 31778 45108 32172
rect 45052 31726 45054 31778
rect 45106 31726 45108 31778
rect 45052 31714 45108 31726
rect 45164 31220 45220 34076
rect 45276 34066 45332 34076
rect 45276 33346 45332 33358
rect 45276 33294 45278 33346
rect 45330 33294 45332 33346
rect 45276 32788 45332 33294
rect 45276 32722 45332 32732
rect 45388 32116 45444 35308
rect 45500 34580 45556 35420
rect 45500 34514 45556 34524
rect 45612 34356 45668 34366
rect 45612 34262 45668 34300
rect 45612 33572 45668 33582
rect 45612 33346 45668 33516
rect 45612 33294 45614 33346
rect 45666 33294 45668 33346
rect 45612 33282 45668 33294
rect 45612 33124 45668 33134
rect 45388 32060 45556 32116
rect 45388 31892 45444 31902
rect 45388 31798 45444 31836
rect 44940 31164 45220 31220
rect 44940 29988 44996 31164
rect 45164 30994 45220 31006
rect 45164 30942 45166 30994
rect 45218 30942 45220 30994
rect 44940 29922 44996 29932
rect 45052 30322 45108 30334
rect 45052 30270 45054 30322
rect 45106 30270 45108 30322
rect 44940 29204 44996 29214
rect 44940 27858 44996 29148
rect 45052 28420 45108 30270
rect 45052 28354 45108 28364
rect 45164 30324 45220 30942
rect 44940 27806 44942 27858
rect 44994 27806 44996 27858
rect 44940 26628 44996 27806
rect 45052 27860 45108 27870
rect 45052 27766 45108 27804
rect 44940 26562 44996 26572
rect 45052 27076 45108 27086
rect 45164 27076 45220 30268
rect 45276 29988 45332 29998
rect 45276 28756 45332 29932
rect 45500 29316 45556 32060
rect 45612 30996 45668 33068
rect 45612 30930 45668 30940
rect 45612 30770 45668 30782
rect 45612 30718 45614 30770
rect 45666 30718 45668 30770
rect 45612 30548 45668 30718
rect 45612 30212 45668 30492
rect 45612 30146 45668 30156
rect 45500 29314 45668 29316
rect 45500 29262 45502 29314
rect 45554 29262 45668 29314
rect 45500 29260 45668 29262
rect 45500 29250 45556 29260
rect 45276 28690 45332 28700
rect 45500 28980 45556 28990
rect 45500 27858 45556 28924
rect 45500 27806 45502 27858
rect 45554 27806 45556 27858
rect 45500 27794 45556 27806
rect 45276 27748 45332 27758
rect 45276 27746 45444 27748
rect 45276 27694 45278 27746
rect 45330 27694 45444 27746
rect 45276 27692 45444 27694
rect 45276 27682 45332 27692
rect 45052 27074 45220 27076
rect 45052 27022 45054 27074
rect 45106 27022 45220 27074
rect 45052 27020 45220 27022
rect 44828 26226 44884 26236
rect 44940 26404 44996 26414
rect 44604 25982 44884 26038
rect 44464 25900 44728 25910
rect 44520 25844 44568 25900
rect 44624 25844 44672 25900
rect 44464 25834 44728 25844
rect 44156 25228 44324 25284
rect 44604 25506 44660 25518
rect 44604 25454 44606 25506
rect 44658 25454 44660 25506
rect 43804 25116 44068 25126
rect 43860 25060 43908 25116
rect 43964 25060 44012 25116
rect 43804 25050 44068 25060
rect 44156 25060 44212 25228
rect 44156 24836 44212 25004
rect 44268 24948 44324 24958
rect 44604 24948 44660 25454
rect 44268 24946 44660 24948
rect 44268 24894 44270 24946
rect 44322 24894 44660 24946
rect 44268 24892 44660 24894
rect 44268 24882 44324 24892
rect 44156 24770 44212 24780
rect 43596 24724 43652 24734
rect 43596 24388 43652 24668
rect 43596 24322 43652 24332
rect 44464 24332 44728 24342
rect 44520 24276 44568 24332
rect 44624 24276 44672 24332
rect 44464 24266 44728 24276
rect 44380 24052 44436 24062
rect 44268 23716 44324 23726
rect 44156 23714 44324 23716
rect 44156 23662 44270 23714
rect 44322 23662 44324 23714
rect 44156 23660 44324 23662
rect 43484 23538 43540 23548
rect 43804 23548 44068 23558
rect 43860 23492 43908 23548
rect 43964 23492 44012 23548
rect 43804 23482 44068 23492
rect 43596 23156 43652 23166
rect 43484 22484 43540 22494
rect 43484 21924 43540 22428
rect 43484 21858 43540 21868
rect 43372 19954 43428 19964
rect 43484 20804 43540 20814
rect 43260 19234 43316 19246
rect 43260 19182 43262 19234
rect 43314 19182 43316 19234
rect 43260 18676 43316 19182
rect 43260 18674 43428 18676
rect 43260 18622 43262 18674
rect 43314 18622 43428 18674
rect 43260 18620 43428 18622
rect 43260 18610 43316 18620
rect 43148 17938 43204 17948
rect 43260 18452 43316 18462
rect 43260 17666 43316 18396
rect 43260 17614 43262 17666
rect 43314 17614 43316 17666
rect 43260 17332 43316 17614
rect 43260 17266 43316 17276
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42924 16818 42980 16830
rect 43372 16882 43428 18620
rect 43484 16994 43540 20748
rect 43596 20802 43652 23100
rect 44156 23044 44212 23660
rect 44268 23650 44324 23660
rect 43820 22988 44212 23044
rect 43820 22370 43876 22988
rect 44380 22932 44436 23996
rect 44268 22876 44436 22932
rect 43820 22318 43822 22370
rect 43874 22318 43876 22370
rect 43820 22306 43876 22318
rect 44156 22596 44212 22606
rect 44156 22370 44212 22540
rect 44156 22318 44158 22370
rect 44210 22318 44212 22370
rect 44156 22306 44212 22318
rect 43804 21980 44068 21990
rect 43860 21924 43908 21980
rect 43964 21924 44012 21980
rect 43804 21914 44068 21924
rect 44156 21028 44212 21038
rect 44268 21028 44324 22876
rect 44464 22764 44728 22774
rect 44520 22708 44568 22764
rect 44624 22708 44672 22764
rect 44464 22698 44728 22708
rect 44380 22596 44436 22606
rect 44380 21812 44436 22540
rect 44380 21746 44436 21756
rect 44828 21812 44884 25982
rect 44828 21746 44884 21756
rect 44940 23938 44996 26348
rect 44940 23886 44942 23938
rect 44994 23886 44996 23938
rect 44828 21364 44884 21374
rect 44464 21196 44728 21206
rect 44520 21140 44568 21196
rect 44624 21140 44672 21196
rect 44464 21130 44728 21140
rect 44156 21026 44324 21028
rect 44156 20974 44158 21026
rect 44210 20974 44324 21026
rect 44156 20972 44324 20974
rect 44156 20962 44212 20972
rect 43596 20750 43598 20802
rect 43650 20750 43652 20802
rect 43596 19796 43652 20750
rect 43804 20412 44068 20422
rect 43860 20356 43908 20412
rect 43964 20356 44012 20412
rect 43804 20346 44068 20356
rect 44268 19908 44324 19918
rect 43596 19740 43764 19796
rect 43484 16942 43486 16994
rect 43538 16942 43540 16994
rect 43484 16930 43540 16942
rect 43596 19460 43652 19470
rect 43372 16830 43374 16882
rect 43426 16830 43428 16882
rect 43372 16818 43428 16830
rect 43596 16770 43652 19404
rect 43708 19236 43764 19740
rect 43708 19170 43764 19180
rect 44156 19684 44212 19694
rect 44156 18900 44212 19628
rect 44268 19572 44324 19852
rect 44464 19628 44728 19638
rect 44520 19572 44568 19628
rect 44624 19572 44672 19628
rect 44464 19562 44728 19572
rect 44268 19346 44324 19516
rect 44268 19294 44270 19346
rect 44322 19294 44324 19346
rect 44268 19282 44324 19294
rect 44604 19236 44660 19246
rect 43804 18844 44068 18854
rect 43860 18788 43908 18844
rect 43964 18788 44012 18844
rect 44156 18834 44212 18844
rect 44380 19234 44660 19236
rect 44380 19182 44606 19234
rect 44658 19182 44660 19234
rect 44380 19180 44660 19182
rect 43804 18778 44068 18788
rect 43932 18676 43988 18686
rect 43708 18564 43764 18574
rect 43708 17890 43764 18508
rect 43708 17838 43710 17890
rect 43762 17838 43764 17890
rect 43708 17826 43764 17838
rect 43932 17890 43988 18620
rect 44268 18676 44324 18686
rect 44380 18676 44436 19180
rect 44604 19170 44660 19180
rect 44268 18674 44436 18676
rect 44268 18622 44270 18674
rect 44322 18622 44436 18674
rect 44268 18620 44436 18622
rect 44268 18610 44324 18620
rect 44828 18564 44884 21308
rect 44828 18498 44884 18508
rect 44940 20804 44996 23886
rect 45052 23156 45108 27020
rect 45388 26964 45444 27692
rect 45612 27524 45668 29260
rect 45724 28868 45780 37212
rect 46060 36708 46116 38668
rect 45948 36652 46116 36708
rect 46172 38612 46340 38668
rect 46396 38612 46564 38668
rect 46620 38946 46676 40236
rect 46620 38894 46622 38946
rect 46674 38894 46676 38946
rect 45836 35698 45892 35710
rect 45836 35646 45838 35698
rect 45890 35646 45892 35698
rect 45836 35140 45892 35646
rect 45948 35700 46004 36652
rect 45948 35634 46004 35644
rect 46060 36484 46116 36494
rect 45836 35074 45892 35084
rect 45948 35252 46004 35262
rect 45948 35026 46004 35196
rect 45948 34974 45950 35026
rect 46002 34974 46004 35026
rect 45948 34468 46004 34974
rect 45836 34412 46004 34468
rect 45836 33796 45892 34412
rect 46060 34356 46116 36428
rect 45836 33730 45892 33740
rect 45948 34300 46116 34356
rect 45836 33348 45892 33358
rect 45836 31332 45892 33292
rect 45948 33012 46004 34300
rect 46060 34132 46116 34142
rect 46060 34038 46116 34076
rect 45948 32956 46116 33012
rect 45948 32788 46004 32798
rect 45948 32694 46004 32732
rect 45836 31266 45892 31276
rect 45948 31780 46004 31790
rect 45724 28802 45780 28812
rect 45836 29426 45892 29438
rect 45836 29374 45838 29426
rect 45890 29374 45892 29426
rect 45612 27458 45668 27468
rect 45724 28644 45780 28654
rect 45500 27300 45556 27310
rect 45500 27206 45556 27244
rect 45724 27300 45780 28588
rect 45724 27234 45780 27244
rect 45276 26628 45332 26638
rect 45276 26178 45332 26572
rect 45276 26126 45278 26178
rect 45330 26126 45332 26178
rect 45276 25396 45332 26126
rect 45388 26178 45444 26908
rect 45388 26126 45390 26178
rect 45442 26126 45444 26178
rect 45388 26114 45444 26126
rect 45500 27076 45556 27086
rect 45500 26068 45556 27020
rect 45612 26292 45668 26302
rect 45612 26198 45668 26236
rect 45836 26068 45892 29374
rect 45948 28980 46004 31724
rect 46060 29204 46116 32956
rect 46172 30660 46228 38612
rect 46284 37380 46340 37390
rect 46284 37286 46340 37324
rect 46396 35364 46452 38612
rect 46396 35298 46452 35308
rect 46508 36258 46564 36270
rect 46508 36206 46510 36258
rect 46562 36206 46564 36258
rect 46284 35140 46340 35150
rect 46284 34916 46340 35084
rect 46508 35140 46564 36206
rect 46620 35700 46676 38894
rect 46732 39394 46788 39406
rect 46732 39342 46734 39394
rect 46786 39342 46788 39394
rect 46732 38164 46788 39342
rect 46732 38098 46788 38108
rect 46844 38836 46900 38846
rect 46732 37940 46788 37950
rect 46732 37846 46788 37884
rect 46620 35606 46676 35644
rect 46732 35812 46788 35822
rect 46396 34916 46452 34926
rect 46284 34914 46452 34916
rect 46284 34862 46398 34914
rect 46450 34862 46452 34914
rect 46284 34860 46452 34862
rect 46396 34850 46452 34860
rect 46508 34804 46564 35084
rect 46508 34738 46564 34748
rect 46620 34692 46676 34702
rect 46284 34244 46340 34254
rect 46508 34244 46564 34254
rect 46284 34242 46508 34244
rect 46284 34190 46286 34242
rect 46338 34190 46508 34242
rect 46284 34188 46508 34190
rect 46284 34178 46340 34188
rect 46508 34178 46564 34188
rect 46284 34020 46340 34030
rect 46284 33926 46340 33964
rect 46396 34018 46452 34030
rect 46396 33966 46398 34018
rect 46450 33966 46452 34018
rect 46396 33572 46452 33966
rect 46620 34018 46676 34636
rect 46620 33966 46622 34018
rect 46674 33966 46676 34018
rect 46620 33954 46676 33966
rect 46396 33506 46452 33516
rect 46620 33346 46676 33358
rect 46620 33294 46622 33346
rect 46674 33294 46676 33346
rect 46620 33236 46676 33294
rect 46620 33170 46676 33180
rect 46732 33012 46788 35756
rect 46508 32900 46564 32910
rect 46508 32452 46564 32844
rect 46508 32386 46564 32396
rect 46620 32562 46676 32574
rect 46620 32510 46622 32562
rect 46674 32510 46676 32562
rect 46620 32228 46676 32510
rect 46732 32452 46788 32956
rect 46732 32386 46788 32396
rect 46620 32162 46676 32172
rect 46620 31556 46676 31566
rect 46620 31462 46676 31500
rect 46172 30594 46228 30604
rect 46732 30770 46788 30782
rect 46732 30718 46734 30770
rect 46786 30718 46788 30770
rect 46284 30436 46340 30446
rect 46172 30212 46228 30222
rect 46172 30118 46228 30156
rect 46060 29138 46116 29148
rect 45948 28924 46116 28980
rect 45948 28756 46004 28766
rect 45948 26290 46004 28700
rect 46060 27748 46116 28924
rect 46172 28868 46228 28878
rect 46172 28644 46228 28812
rect 46284 28866 46340 30380
rect 46620 30212 46676 30222
rect 46620 29428 46676 30156
rect 46508 29426 46676 29428
rect 46508 29374 46622 29426
rect 46674 29374 46676 29426
rect 46508 29372 46676 29374
rect 46284 28814 46286 28866
rect 46338 28814 46340 28866
rect 46284 28802 46340 28814
rect 46396 29314 46452 29326
rect 46396 29262 46398 29314
rect 46450 29262 46452 29314
rect 46396 28866 46452 29262
rect 46396 28814 46398 28866
rect 46450 28814 46452 28866
rect 46396 28802 46452 28814
rect 46508 28866 46564 29372
rect 46620 29362 46676 29372
rect 46732 30210 46788 30718
rect 46732 30158 46734 30210
rect 46786 30158 46788 30210
rect 46508 28814 46510 28866
rect 46562 28814 46564 28866
rect 46508 28802 46564 28814
rect 46732 28866 46788 30158
rect 46844 29988 46900 38780
rect 46956 38724 47012 44828
rect 47068 44436 47124 45166
rect 47516 44884 47572 44894
rect 47516 44790 47572 44828
rect 47068 44370 47124 44380
rect 47404 44098 47460 44110
rect 47404 44046 47406 44098
rect 47458 44046 47460 44098
rect 47404 43540 47460 44046
rect 47404 43474 47460 43484
rect 47180 43316 47236 43326
rect 47068 42756 47124 42766
rect 47068 42662 47124 42700
rect 47180 41298 47236 43260
rect 47292 42868 47348 42878
rect 47292 42754 47348 42812
rect 47404 42868 47460 42878
rect 47628 42868 47684 46172
rect 47740 45444 47796 46620
rect 47852 46610 47908 46620
rect 47964 48188 48244 48244
rect 48412 48804 48468 48814
rect 47740 45378 47796 45388
rect 47852 43428 47908 43438
rect 47852 43334 47908 43372
rect 47404 42866 47684 42868
rect 47404 42814 47406 42866
rect 47458 42814 47684 42866
rect 47404 42812 47684 42814
rect 47852 42868 47908 42878
rect 47404 42802 47460 42812
rect 47292 42702 47294 42754
rect 47346 42702 47348 42754
rect 47292 42690 47348 42702
rect 47740 42532 47796 42542
rect 47180 41246 47182 41298
rect 47234 41246 47236 41298
rect 47180 41234 47236 41246
rect 47404 41972 47460 41982
rect 47404 41748 47460 41916
rect 47404 41186 47460 41692
rect 47404 41134 47406 41186
rect 47458 41134 47460 41186
rect 47404 41122 47460 41134
rect 47628 41746 47684 41758
rect 47628 41694 47630 41746
rect 47682 41694 47684 41746
rect 47628 40404 47684 41694
rect 47740 40740 47796 42476
rect 47740 40674 47796 40684
rect 47628 40348 47796 40404
rect 47068 40178 47124 40190
rect 47068 40126 47070 40178
rect 47122 40126 47124 40178
rect 47068 39956 47124 40126
rect 47628 40180 47684 40190
rect 47068 39890 47124 39900
rect 47516 39956 47572 39966
rect 47516 39842 47572 39900
rect 47516 39790 47518 39842
rect 47570 39790 47572 39842
rect 47516 39778 47572 39790
rect 47404 39732 47460 39742
rect 47180 39618 47236 39630
rect 47180 39566 47182 39618
rect 47234 39566 47236 39618
rect 47180 39060 47236 39566
rect 47180 38994 47236 39004
rect 46956 38658 47012 38668
rect 47292 38164 47348 38174
rect 47292 38070 47348 38108
rect 47292 37938 47348 37950
rect 47292 37886 47294 37938
rect 47346 37886 47348 37938
rect 46956 37826 47012 37838
rect 46956 37774 46958 37826
rect 47010 37774 47012 37826
rect 46956 36708 47012 37774
rect 47292 37380 47348 37886
rect 47292 37314 47348 37324
rect 47068 36708 47124 36718
rect 46956 36706 47124 36708
rect 46956 36654 47070 36706
rect 47122 36654 47124 36706
rect 46956 36652 47124 36654
rect 47068 36642 47124 36652
rect 47292 36596 47348 36606
rect 47404 36596 47460 39676
rect 47628 39620 47684 40124
rect 47628 39554 47684 39564
rect 47740 39844 47796 40348
rect 47516 38836 47572 38846
rect 47516 38276 47572 38780
rect 47516 38210 47572 38220
rect 47516 37826 47572 37838
rect 47516 37774 47518 37826
rect 47570 37774 47572 37826
rect 47516 37716 47572 37774
rect 47516 37650 47572 37660
rect 47292 36594 47460 36596
rect 47292 36542 47294 36594
rect 47346 36542 47460 36594
rect 47292 36540 47460 36542
rect 47292 36530 47348 36540
rect 46956 36484 47012 36494
rect 46956 36390 47012 36428
rect 47516 36482 47572 36494
rect 47516 36430 47518 36482
rect 47570 36430 47572 36482
rect 46956 35812 47012 35822
rect 46956 35586 47012 35756
rect 47516 35812 47572 36430
rect 47516 35746 47572 35756
rect 47628 36036 47684 36046
rect 46956 35534 46958 35586
rect 47010 35534 47012 35586
rect 46956 35522 47012 35534
rect 47516 35476 47572 35486
rect 47180 35140 47236 35150
rect 47180 35046 47236 35084
rect 47404 35026 47460 35038
rect 47404 34974 47406 35026
rect 47458 34974 47460 35026
rect 46956 34914 47012 34926
rect 46956 34862 46958 34914
rect 47010 34862 47012 34914
rect 46956 34356 47012 34862
rect 47068 34804 47124 34814
rect 47068 34802 47236 34804
rect 47068 34750 47070 34802
rect 47122 34750 47236 34802
rect 47068 34748 47236 34750
rect 47068 34738 47124 34748
rect 46956 34290 47012 34300
rect 47180 34020 47236 34748
rect 47404 34692 47460 34974
rect 47404 34626 47460 34636
rect 47516 34356 47572 35420
rect 47628 34692 47684 35980
rect 47628 34626 47684 34636
rect 47516 34290 47572 34300
rect 47740 34132 47796 39788
rect 47852 35140 47908 42812
rect 47964 39620 48020 48188
rect 48076 47684 48132 47694
rect 48076 47590 48132 47628
rect 48300 47460 48356 47470
rect 48300 47366 48356 47404
rect 48188 47348 48244 47358
rect 48188 47254 48244 47292
rect 48412 46116 48468 48748
rect 48076 46060 48468 46116
rect 48524 47460 48580 47470
rect 48076 43316 48132 46060
rect 48412 45892 48468 45902
rect 48300 45780 48356 45790
rect 48188 44212 48244 44222
rect 48188 43650 48244 44156
rect 48188 43598 48190 43650
rect 48242 43598 48244 43650
rect 48188 43586 48244 43598
rect 48076 43260 48244 43316
rect 48076 41970 48132 41982
rect 48076 41918 48078 41970
rect 48130 41918 48132 41970
rect 48076 41748 48132 41918
rect 48076 41682 48132 41692
rect 48188 41410 48244 43260
rect 48188 41358 48190 41410
rect 48242 41358 48244 41410
rect 48188 41346 48244 41358
rect 48300 41410 48356 45724
rect 48412 43316 48468 45836
rect 48524 44436 48580 47404
rect 48636 47458 48692 47470
rect 48636 47406 48638 47458
rect 48690 47406 48692 47458
rect 48636 45220 48692 47406
rect 48748 46898 48804 49196
rect 48860 49028 48916 49038
rect 48860 48934 48916 48972
rect 48748 46846 48750 46898
rect 48802 46846 48804 46898
rect 48748 46834 48804 46846
rect 48860 48804 48916 48814
rect 48636 45154 48692 45164
rect 48748 45778 48804 45790
rect 48748 45726 48750 45778
rect 48802 45726 48804 45778
rect 48524 44370 48580 44380
rect 48636 44882 48692 44894
rect 48636 44830 48638 44882
rect 48690 44830 48692 44882
rect 48412 43250 48468 43260
rect 48524 44212 48580 44222
rect 48524 43204 48580 44156
rect 48636 43428 48692 44830
rect 48748 44212 48804 45726
rect 48748 44146 48804 44156
rect 48860 43540 48916 48748
rect 48972 48356 49028 49198
rect 49084 48356 49140 48366
rect 48972 48354 49140 48356
rect 48972 48302 49086 48354
rect 49138 48302 49140 48354
rect 48972 48300 49140 48302
rect 49084 48290 49140 48300
rect 49196 47796 49252 50428
rect 49308 50372 49476 50428
rect 49308 49028 49364 50372
rect 49532 49924 49588 52222
rect 49644 51604 49700 51614
rect 49644 51510 49700 51548
rect 49644 50706 49700 50718
rect 49644 50654 49646 50706
rect 49698 50654 49700 50706
rect 49644 50596 49700 50654
rect 49644 50530 49700 50540
rect 49756 50428 49812 52668
rect 49980 52500 50036 54684
rect 50092 54292 50148 54302
rect 50092 52724 50148 54236
rect 50204 53842 50260 53854
rect 50204 53790 50206 53842
rect 50258 53790 50260 53842
rect 50204 52948 50260 53790
rect 50540 53842 50596 53854
rect 50540 53790 50542 53842
rect 50594 53790 50596 53842
rect 50540 53508 50596 53790
rect 50540 53442 50596 53452
rect 50204 52892 50372 52948
rect 50204 52724 50260 52734
rect 50092 52722 50260 52724
rect 50092 52670 50206 52722
rect 50258 52670 50260 52722
rect 50092 52668 50260 52670
rect 50204 52658 50260 52668
rect 49980 52444 50260 52500
rect 50092 52276 50148 52286
rect 49980 52274 50148 52276
rect 49980 52222 50094 52274
rect 50146 52222 50148 52274
rect 49980 52220 50148 52222
rect 49868 52164 49924 52174
rect 49868 52070 49924 52108
rect 49868 51492 49924 51502
rect 49980 51492 50036 52220
rect 50092 52210 50148 52220
rect 50204 52274 50260 52444
rect 50204 52222 50206 52274
rect 50258 52222 50260 52274
rect 50204 51604 50260 52222
rect 50204 51538 50260 51548
rect 49980 51436 50148 51492
rect 49868 51398 49924 51436
rect 49868 51266 49924 51278
rect 49868 51214 49870 51266
rect 49922 51214 49924 51266
rect 49868 51156 49924 51214
rect 49868 51090 49924 51100
rect 49756 50372 50036 50428
rect 49980 50036 50036 50372
rect 49980 49970 50036 49980
rect 49532 49858 49588 49868
rect 50092 49924 50148 51436
rect 50204 51378 50260 51390
rect 50204 51326 50206 51378
rect 50258 51326 50260 51378
rect 50204 50820 50260 51326
rect 50204 50754 50260 50764
rect 50092 49858 50148 49868
rect 50204 49810 50260 49822
rect 50204 49758 50206 49810
rect 50258 49758 50260 49810
rect 49644 49698 49700 49710
rect 49644 49646 49646 49698
rect 49698 49646 49700 49698
rect 49308 48962 49364 48972
rect 49420 49586 49476 49598
rect 49420 49534 49422 49586
rect 49474 49534 49476 49586
rect 49420 48804 49476 49534
rect 49420 48738 49476 48748
rect 49532 49586 49588 49598
rect 49532 49534 49534 49586
rect 49586 49534 49588 49586
rect 49532 48468 49588 49534
rect 49532 48402 49588 48412
rect 49196 47730 49252 47740
rect 49532 47570 49588 47582
rect 49532 47518 49534 47570
rect 49586 47518 49588 47570
rect 48972 47460 49028 47470
rect 48972 46564 49028 47404
rect 49196 47348 49252 47358
rect 49196 47346 49364 47348
rect 49196 47294 49198 47346
rect 49250 47294 49364 47346
rect 49196 47292 49364 47294
rect 49196 47236 49252 47292
rect 49196 47170 49252 47180
rect 48972 46498 49028 46508
rect 49308 46452 49364 47292
rect 49532 47124 49588 47518
rect 49532 47058 49588 47068
rect 49644 46900 49700 49646
rect 49868 49476 49924 49486
rect 49868 49140 49924 49420
rect 50092 49140 50148 49150
rect 49868 49138 50148 49140
rect 49868 49086 50094 49138
rect 50146 49086 50148 49138
rect 49868 49084 50148 49086
rect 49644 46834 49700 46844
rect 49756 49028 49812 49038
rect 49756 48914 49812 48972
rect 49756 48862 49758 48914
rect 49810 48862 49812 48914
rect 49756 46786 49812 48862
rect 49868 48916 49924 49084
rect 50092 49074 50148 49084
rect 49868 48850 49924 48860
rect 49980 48468 50036 48478
rect 49756 46734 49758 46786
rect 49810 46734 49812 46786
rect 49756 46722 49812 46734
rect 49868 48242 49924 48254
rect 49868 48190 49870 48242
rect 49922 48190 49924 48242
rect 49868 47796 49924 48190
rect 49644 46674 49700 46686
rect 49644 46622 49646 46674
rect 49698 46622 49700 46674
rect 49644 46452 49700 46622
rect 49868 46676 49924 47740
rect 49980 47068 50036 48412
rect 50204 48356 50260 49758
rect 50316 49252 50372 52892
rect 50540 52722 50596 52734
rect 50540 52670 50542 52722
rect 50594 52670 50596 52722
rect 50428 52164 50484 52174
rect 50428 51602 50484 52108
rect 50428 51550 50430 51602
rect 50482 51550 50484 51602
rect 50428 51538 50484 51550
rect 50428 50482 50484 50494
rect 50428 50430 50430 50482
rect 50482 50430 50484 50482
rect 50428 50036 50484 50430
rect 50540 50372 50596 52670
rect 50652 52500 50708 54796
rect 50764 53732 50820 53742
rect 50764 53638 50820 53676
rect 51100 53060 51156 55580
rect 51212 55412 51268 55806
rect 51324 55524 51380 57344
rect 51548 55860 51604 55870
rect 51548 55766 51604 55804
rect 51324 55458 51380 55468
rect 51212 55346 51268 55356
rect 51324 54516 51380 54526
rect 51100 52994 51156 53004
rect 51212 53842 51268 53854
rect 51212 53790 51214 53842
rect 51266 53790 51268 53842
rect 51212 52948 51268 53790
rect 51212 52882 51268 52892
rect 50876 52724 50932 52734
rect 50876 52630 50932 52668
rect 51212 52722 51268 52734
rect 51212 52670 51214 52722
rect 51266 52670 51268 52722
rect 50652 52386 50708 52444
rect 50652 52334 50654 52386
rect 50706 52334 50708 52386
rect 50652 52322 50708 52334
rect 51100 52500 51156 52510
rect 50540 50306 50596 50316
rect 50652 51492 50708 51502
rect 50428 49980 50596 50036
rect 50540 49924 50596 49980
rect 50428 49812 50484 49822
rect 50428 49698 50484 49756
rect 50428 49646 50430 49698
rect 50482 49646 50484 49698
rect 50428 49634 50484 49646
rect 50316 49186 50372 49196
rect 50540 49028 50596 49868
rect 50652 49476 50708 51436
rect 50988 51378 51044 51390
rect 50988 51326 50990 51378
rect 51042 51326 51044 51378
rect 50764 50708 50820 50718
rect 50764 50614 50820 50652
rect 50988 50596 51044 51326
rect 51100 51378 51156 52444
rect 51212 52276 51268 52670
rect 51212 52210 51268 52220
rect 51324 51940 51380 54460
rect 51772 54404 51828 57344
rect 52108 57204 52164 57214
rect 51996 56868 52052 56878
rect 51884 56308 51940 56318
rect 51884 55970 51940 56252
rect 51884 55918 51886 55970
rect 51938 55918 51940 55970
rect 51884 55906 51940 55918
rect 51996 55300 52052 56812
rect 51996 55234 52052 55244
rect 51996 54404 52052 54414
rect 51772 54402 52052 54404
rect 51772 54350 51998 54402
rect 52050 54350 52052 54402
rect 51772 54348 52052 54350
rect 51996 54338 52052 54348
rect 52108 54068 52164 57148
rect 52220 56532 52276 57344
rect 52220 56466 52276 56476
rect 52668 56196 52724 57344
rect 53116 56644 53172 57344
rect 53116 56578 53172 56588
rect 53228 56756 53284 56766
rect 52668 56130 52724 56140
rect 52556 56084 52612 56094
rect 52556 55970 52612 56028
rect 52556 55918 52558 55970
rect 52610 55918 52612 55970
rect 52556 55906 52612 55918
rect 53228 55970 53284 56700
rect 53564 56308 53620 57344
rect 54012 57316 54068 57344
rect 54012 57250 54068 57260
rect 54460 56420 54516 57344
rect 54908 56980 54964 57344
rect 55356 57316 55412 57344
rect 55356 57250 55412 57260
rect 54908 56914 54964 56924
rect 54460 56354 54516 56364
rect 55020 56532 55076 56542
rect 53228 55918 53230 55970
rect 53282 55918 53284 55970
rect 53228 55906 53284 55918
rect 53452 56252 53620 56308
rect 51660 54012 52164 54068
rect 52220 55858 52276 55870
rect 52220 55806 52222 55858
rect 52274 55806 52276 55858
rect 51548 53732 51604 53742
rect 51548 53638 51604 53676
rect 51100 51326 51102 51378
rect 51154 51326 51156 51378
rect 51100 51314 51156 51326
rect 51212 51884 51380 51940
rect 51212 51268 51268 51884
rect 51436 51604 51492 51614
rect 51324 51380 51380 51390
rect 51324 51286 51380 51324
rect 51436 51378 51492 51548
rect 51436 51326 51438 51378
rect 51490 51326 51492 51378
rect 51436 51314 51492 51326
rect 51212 51202 51268 51212
rect 50988 50428 51044 50540
rect 51548 50932 51604 50942
rect 50988 50372 51156 50428
rect 50988 49810 51044 49822
rect 50988 49758 50990 49810
rect 51042 49758 51044 49810
rect 50652 49410 50708 49420
rect 50876 49698 50932 49710
rect 50876 49646 50878 49698
rect 50930 49646 50932 49698
rect 50540 48962 50596 48972
rect 50876 48580 50932 49646
rect 50876 48514 50932 48524
rect 49980 47002 50036 47012
rect 50092 48300 50260 48356
rect 50540 48468 50596 48478
rect 49868 46610 49924 46620
rect 50092 46564 50148 48300
rect 50204 48130 50260 48142
rect 50204 48078 50206 48130
rect 50258 48078 50260 48130
rect 50204 47124 50260 48078
rect 50316 48132 50372 48142
rect 50316 48038 50372 48076
rect 50204 47058 50260 47068
rect 50092 46498 50148 46508
rect 50316 47012 50372 47022
rect 49308 46396 49700 46452
rect 50204 46452 50260 46462
rect 49084 46004 49140 46014
rect 49084 45910 49140 45948
rect 49308 45218 49364 46396
rect 50204 46358 50260 46396
rect 50092 46340 50148 46350
rect 49980 46284 50092 46340
rect 49980 45892 50036 46284
rect 50092 46274 50148 46284
rect 50316 46116 50372 46956
rect 49980 45826 50036 45836
rect 50204 46060 50372 46116
rect 50092 45780 50148 45790
rect 49308 45166 49310 45218
rect 49362 45166 49364 45218
rect 49308 45154 49364 45166
rect 49532 45556 49588 45566
rect 49196 45106 49252 45118
rect 49196 45054 49198 45106
rect 49250 45054 49252 45106
rect 48972 44436 49028 44446
rect 48972 44342 49028 44380
rect 49196 44212 49252 45054
rect 49532 44578 49588 45500
rect 49196 44146 49252 44156
rect 49420 44522 49588 44578
rect 49644 45444 49700 45454
rect 49196 43540 49252 43550
rect 48860 43484 49028 43540
rect 48636 43362 48692 43372
rect 48860 43316 48916 43326
rect 48860 43222 48916 43260
rect 48524 43148 48804 43204
rect 48300 41358 48302 41410
rect 48354 41358 48356 41410
rect 48300 41346 48356 41358
rect 48524 41972 48580 41982
rect 48524 41410 48580 41916
rect 48524 41358 48526 41410
rect 48578 41358 48580 41410
rect 48524 41346 48580 41358
rect 48748 41970 48804 43148
rect 48748 41918 48750 41970
rect 48802 41918 48804 41970
rect 48076 41300 48132 41310
rect 48076 41206 48132 41244
rect 48748 41300 48804 41918
rect 48972 41412 49028 43484
rect 49196 43446 49252 43484
rect 49420 43426 49476 44522
rect 49420 43374 49422 43426
rect 49474 43374 49476 43426
rect 48972 41346 49028 41356
rect 49084 43092 49140 43102
rect 48300 41188 48356 41198
rect 48188 40178 48244 40190
rect 48188 40126 48190 40178
rect 48242 40126 48244 40178
rect 48188 39732 48244 40126
rect 48188 39638 48244 39676
rect 48076 39620 48132 39630
rect 47964 39618 48132 39620
rect 47964 39566 48078 39618
rect 48130 39566 48132 39618
rect 47964 39564 48132 39566
rect 47964 36484 48020 39564
rect 48076 39554 48132 39564
rect 48188 39060 48244 39070
rect 48300 39060 48356 41132
rect 48412 40964 48468 40974
rect 48412 39842 48468 40908
rect 48748 40852 48804 41244
rect 48972 40964 49028 41002
rect 48972 40898 49028 40908
rect 48748 40786 48804 40796
rect 48972 40740 49028 40750
rect 48412 39790 48414 39842
rect 48466 39790 48468 39842
rect 48412 39778 48468 39790
rect 48860 40402 48916 40414
rect 48860 40350 48862 40402
rect 48914 40350 48916 40402
rect 48188 39058 48356 39060
rect 48188 39006 48190 39058
rect 48242 39006 48356 39058
rect 48188 39004 48356 39006
rect 48524 39620 48580 39630
rect 48188 38994 48244 39004
rect 48300 38724 48356 38734
rect 48188 38276 48244 38286
rect 48188 38182 48244 38220
rect 48076 38164 48132 38174
rect 48076 38070 48132 38108
rect 48188 37826 48244 37838
rect 48188 37774 48190 37826
rect 48242 37774 48244 37826
rect 48188 37716 48244 37774
rect 48188 37650 48244 37660
rect 47964 36418 48020 36428
rect 48188 36036 48244 36046
rect 48188 35922 48244 35980
rect 48188 35870 48190 35922
rect 48242 35870 48244 35922
rect 48188 35858 48244 35870
rect 47852 35084 48244 35140
rect 47964 34244 48020 34254
rect 47516 34076 47796 34132
rect 47852 34132 47908 34142
rect 47068 34018 47236 34020
rect 47068 33966 47182 34018
rect 47234 33966 47236 34018
rect 47068 33964 47236 33966
rect 46956 33796 47012 33806
rect 46956 33348 47012 33740
rect 47068 33628 47124 33964
rect 47180 33954 47236 33964
rect 47292 34020 47348 34030
rect 47292 33926 47348 33964
rect 47404 33906 47460 33918
rect 47404 33854 47406 33906
rect 47458 33854 47460 33906
rect 47068 33572 47236 33628
rect 47180 33516 47348 33572
rect 47068 33348 47124 33358
rect 46956 33292 47068 33348
rect 47068 33282 47124 33292
rect 47180 33346 47236 33358
rect 47180 33294 47182 33346
rect 47234 33294 47236 33346
rect 47180 32676 47236 33294
rect 47180 32610 47236 32620
rect 46956 32452 47012 32462
rect 46956 32358 47012 32396
rect 47180 31890 47236 31902
rect 47180 31838 47182 31890
rect 47234 31838 47236 31890
rect 47068 31554 47124 31566
rect 47068 31502 47070 31554
rect 47122 31502 47124 31554
rect 47068 30996 47124 31502
rect 47180 30996 47236 31838
rect 47292 31892 47348 33516
rect 47404 32116 47460 33854
rect 47516 33628 47572 34076
rect 47852 34038 47908 34076
rect 47516 33562 47572 33572
rect 47628 33908 47684 33918
rect 47516 33460 47572 33470
rect 47516 33366 47572 33404
rect 47404 32060 47572 32116
rect 47404 31892 47460 31902
rect 47292 31890 47460 31892
rect 47292 31838 47406 31890
rect 47458 31838 47460 31890
rect 47292 31836 47460 31838
rect 47404 31826 47460 31836
rect 47516 31780 47572 32060
rect 47404 31556 47460 31566
rect 47516 31556 47572 31724
rect 47460 31500 47572 31556
rect 47180 30940 47348 30996
rect 47068 30930 47124 30940
rect 47180 30772 47236 30782
rect 46956 30770 47236 30772
rect 46956 30718 47182 30770
rect 47234 30718 47236 30770
rect 46956 30716 47236 30718
rect 46956 30436 47012 30716
rect 47180 30706 47236 30716
rect 47292 30548 47348 30940
rect 47404 30882 47460 31500
rect 47516 31220 47572 31230
rect 47516 31106 47572 31164
rect 47516 31054 47518 31106
rect 47570 31054 47572 31106
rect 47516 31042 47572 31054
rect 47628 30996 47684 33852
rect 47964 33796 48020 34188
rect 47964 33730 48020 33740
rect 48076 34132 48132 34142
rect 47852 33684 47908 33694
rect 47628 30930 47684 30940
rect 47740 33628 47852 33684
rect 47404 30830 47406 30882
rect 47458 30830 47460 30882
rect 47404 30818 47460 30830
rect 47516 30884 47572 30894
rect 47516 30790 47572 30828
rect 46956 30370 47012 30380
rect 47180 30492 47348 30548
rect 47068 30324 47124 30334
rect 46956 30212 47012 30222
rect 47068 30212 47124 30268
rect 46956 30210 47124 30212
rect 46956 30158 46958 30210
rect 47010 30158 47124 30210
rect 46956 30156 47124 30158
rect 47180 30322 47236 30492
rect 47180 30270 47182 30322
rect 47234 30270 47236 30322
rect 47180 30212 47236 30270
rect 46956 30146 47012 30156
rect 47180 30146 47236 30156
rect 47292 30324 47348 30334
rect 47292 30210 47348 30268
rect 47292 30158 47294 30210
rect 47346 30158 47348 30210
rect 47292 30146 47348 30158
rect 47404 30322 47460 30334
rect 47404 30270 47406 30322
rect 47458 30270 47460 30322
rect 47404 30212 47460 30270
rect 47404 30146 47460 30156
rect 46844 29932 47012 29988
rect 46844 29540 46900 29550
rect 46956 29540 47012 29932
rect 46956 29484 47124 29540
rect 46844 29446 46900 29484
rect 46956 29316 47012 29326
rect 46956 29222 47012 29260
rect 47068 29092 47124 29484
rect 47516 29428 47572 29438
rect 47516 29334 47572 29372
rect 46732 28814 46734 28866
rect 46786 28814 46788 28866
rect 46732 28802 46788 28814
rect 46956 29036 47124 29092
rect 46172 28588 46452 28644
rect 46396 27970 46452 28588
rect 46396 27918 46398 27970
rect 46450 27918 46452 27970
rect 46396 27906 46452 27918
rect 46060 27692 46452 27748
rect 46284 27524 46340 27534
rect 45948 26238 45950 26290
rect 46002 26238 46004 26290
rect 45948 26226 46004 26238
rect 46172 27300 46228 27310
rect 45500 26012 45780 26068
rect 45836 26012 46116 26068
rect 45388 25844 45444 25854
rect 45388 25506 45444 25788
rect 45388 25454 45390 25506
rect 45442 25454 45444 25506
rect 45388 25442 45444 25454
rect 45612 25508 45668 25518
rect 45276 25284 45332 25340
rect 45276 25228 45444 25284
rect 45388 25172 45444 25228
rect 45388 25106 45444 25116
rect 45276 24612 45332 24622
rect 45276 24050 45332 24556
rect 45388 24500 45444 24510
rect 45388 24406 45444 24444
rect 45276 23998 45278 24050
rect 45330 23998 45332 24050
rect 45276 23986 45332 23998
rect 45052 23090 45108 23100
rect 45164 23268 45220 23278
rect 45164 22484 45220 23212
rect 45164 22370 45220 22428
rect 45164 22318 45166 22370
rect 45218 22318 45220 22370
rect 45164 22306 45220 22318
rect 45500 22372 45556 22382
rect 45388 21586 45444 21598
rect 45388 21534 45390 21586
rect 45442 21534 45444 21586
rect 45388 20804 45444 21534
rect 44940 20748 45444 20804
rect 44828 18228 44884 18238
rect 44464 18060 44728 18070
rect 44520 18004 44568 18060
rect 44624 18004 44672 18060
rect 44464 17994 44728 18004
rect 43932 17838 43934 17890
rect 43986 17838 43988 17890
rect 43932 17826 43988 17838
rect 44044 17668 44100 17678
rect 44044 17574 44100 17612
rect 43804 17276 44068 17286
rect 43860 17220 43908 17276
rect 43964 17220 44012 17276
rect 43804 17210 44068 17220
rect 44156 17220 44212 17230
rect 43596 16718 43598 16770
rect 43650 16718 43652 16770
rect 43596 16706 43652 16718
rect 42700 16322 42868 16324
rect 42700 16270 42702 16322
rect 42754 16270 42868 16322
rect 42700 16268 42868 16270
rect 43372 16660 43428 16670
rect 42700 16258 42756 16268
rect 42812 16100 42868 16110
rect 42812 15426 42868 16044
rect 43260 15876 43316 15886
rect 42812 15374 42814 15426
rect 42866 15374 42868 15426
rect 42812 15362 42868 15374
rect 42924 15874 43316 15876
rect 42924 15822 43262 15874
rect 43314 15822 43316 15874
rect 42924 15820 43316 15822
rect 42924 15148 42980 15820
rect 43260 15810 43316 15820
rect 43372 15540 43428 16604
rect 43804 15708 44068 15718
rect 43860 15652 43908 15708
rect 43964 15652 44012 15708
rect 43804 15642 44068 15652
rect 43484 15540 43540 15550
rect 43372 15538 43540 15540
rect 43372 15486 43486 15538
rect 43538 15486 43540 15538
rect 43372 15484 43540 15486
rect 43484 15474 43540 15484
rect 43708 15540 43764 15550
rect 43148 15428 43204 15438
rect 42476 15092 42644 15148
rect 42476 14868 42532 14878
rect 42364 13524 42420 13534
rect 42252 12962 42308 12974
rect 42252 12910 42254 12962
rect 42306 12910 42308 12962
rect 42252 12628 42308 12910
rect 42252 12562 42308 12572
rect 42140 10098 42196 10108
rect 42252 11620 42308 11630
rect 42252 10612 42308 11564
rect 42140 8932 42196 8942
rect 42252 8932 42308 10556
rect 42140 8930 42308 8932
rect 42140 8878 42142 8930
rect 42194 8878 42308 8930
rect 42140 8876 42308 8878
rect 42140 8866 42196 8876
rect 42364 8148 42420 13468
rect 42476 11620 42532 14812
rect 42476 11554 42532 11564
rect 42476 11394 42532 11406
rect 42476 11342 42478 11394
rect 42530 11342 42532 11394
rect 42476 10052 42532 11342
rect 42588 10276 42644 15092
rect 42700 15092 42980 15148
rect 43036 15204 43092 15214
rect 42700 14530 42756 15092
rect 42700 14478 42702 14530
rect 42754 14478 42756 14530
rect 42700 14466 42756 14478
rect 43036 14532 43092 15148
rect 43036 14438 43092 14476
rect 43036 14196 43092 14206
rect 42924 13972 42980 13982
rect 42924 12180 42980 13916
rect 43036 12628 43092 14140
rect 43148 13972 43204 15372
rect 43596 15428 43652 15438
rect 43148 13906 43204 13916
rect 43372 15202 43428 15214
rect 43372 15150 43374 15202
rect 43426 15150 43428 15202
rect 43036 12562 43092 12572
rect 43148 13748 43204 13758
rect 42924 12114 42980 12124
rect 42812 11954 42868 11966
rect 42812 11902 42814 11954
rect 42866 11902 42868 11954
rect 42812 11844 42868 11902
rect 42812 11778 42868 11788
rect 43036 11620 43092 11630
rect 43036 11526 43092 11564
rect 42812 11394 42868 11406
rect 42812 11342 42814 11394
rect 42866 11342 42868 11394
rect 42812 11060 42868 11342
rect 42812 10994 42868 11004
rect 43148 10834 43204 13692
rect 43372 13636 43428 15150
rect 43484 15204 43540 15214
rect 43596 15204 43652 15372
rect 43484 15202 43652 15204
rect 43484 15150 43486 15202
rect 43538 15150 43652 15202
rect 43484 15148 43652 15150
rect 43484 15138 43540 15148
rect 43708 14980 43764 15484
rect 44156 15316 44212 17164
rect 44268 16658 44324 16670
rect 44268 16606 44270 16658
rect 44322 16606 44324 16658
rect 44268 15428 44324 16606
rect 44464 16492 44728 16502
rect 44520 16436 44568 16492
rect 44624 16436 44672 16492
rect 44464 16426 44728 16436
rect 44828 16324 44884 18172
rect 44716 16268 44884 16324
rect 44380 16210 44436 16222
rect 44380 16158 44382 16210
rect 44434 16158 44436 16210
rect 44380 15988 44436 16158
rect 44380 15922 44436 15932
rect 44716 15764 44772 16268
rect 44828 16100 44884 16110
rect 44828 16006 44884 16044
rect 44716 15708 44884 15764
rect 44268 15362 44324 15372
rect 44156 15250 44212 15260
rect 44716 15314 44772 15326
rect 44716 15262 44718 15314
rect 44770 15262 44772 15314
rect 43484 14924 43764 14980
rect 44044 15092 44100 15102
rect 43484 13970 43540 14924
rect 44044 14756 44100 15036
rect 44716 15092 44772 15262
rect 44716 15026 44772 15036
rect 44464 14924 44728 14934
rect 44520 14868 44568 14924
rect 44624 14868 44672 14924
rect 44464 14858 44728 14868
rect 43932 14532 43988 14542
rect 43932 14308 43988 14476
rect 44044 14530 44100 14700
rect 44044 14478 44046 14530
rect 44098 14478 44100 14530
rect 44044 14466 44100 14478
rect 44828 14530 44884 15708
rect 44940 15316 44996 20748
rect 45276 20578 45332 20590
rect 45276 20526 45278 20578
rect 45330 20526 45332 20578
rect 45276 20020 45332 20526
rect 45388 20020 45444 20030
rect 45276 20018 45444 20020
rect 45276 19966 45390 20018
rect 45442 19966 45444 20018
rect 45276 19964 45444 19966
rect 45388 19954 45444 19964
rect 45052 19908 45108 19918
rect 45052 19814 45108 19852
rect 45500 19572 45556 22316
rect 45612 20132 45668 25452
rect 45724 24724 45780 26012
rect 45948 25172 46004 25182
rect 45836 24724 45892 24734
rect 45724 24722 45892 24724
rect 45724 24670 45838 24722
rect 45890 24670 45892 24722
rect 45724 24668 45892 24670
rect 45724 24388 45780 24398
rect 45724 23154 45780 24332
rect 45724 23102 45726 23154
rect 45778 23102 45780 23154
rect 45724 23090 45780 23102
rect 45836 20356 45892 24668
rect 45948 22370 46004 25116
rect 46060 23156 46116 26012
rect 46172 25506 46228 27244
rect 46172 25454 46174 25506
rect 46226 25454 46228 25506
rect 46172 25442 46228 25454
rect 46060 23090 46116 23100
rect 46060 22484 46116 22494
rect 46060 22390 46116 22428
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 45948 21924 46004 22318
rect 46060 22148 46116 22158
rect 46060 22054 46116 22092
rect 45948 21858 46004 21868
rect 45948 21362 46004 21374
rect 45948 21310 45950 21362
rect 46002 21310 46004 21362
rect 45948 21252 46004 21310
rect 45948 20916 46004 21196
rect 45948 20850 46004 20860
rect 45836 20290 45892 20300
rect 45612 20066 45668 20076
rect 45836 20018 45892 20030
rect 45836 19966 45838 20018
rect 45890 19966 45892 20018
rect 45836 19796 45892 19966
rect 45836 19730 45892 19740
rect 46060 19796 46116 19806
rect 46060 19702 46116 19740
rect 45500 19506 45556 19516
rect 45164 19460 45220 19470
rect 45052 19236 45108 19246
rect 45052 17666 45108 19180
rect 45164 19234 45220 19404
rect 45276 19348 45332 19358
rect 45276 19254 45332 19292
rect 45164 19182 45166 19234
rect 45218 19182 45220 19234
rect 45164 19170 45220 19182
rect 45612 19236 45668 19246
rect 45612 18676 45668 19180
rect 45836 19236 45892 19246
rect 45836 19142 45892 19180
rect 45612 18610 45668 18620
rect 45836 18676 45892 18686
rect 45836 18562 45892 18620
rect 45836 18510 45838 18562
rect 45890 18510 45892 18562
rect 45836 18498 45892 18510
rect 45388 18452 45444 18462
rect 45388 18226 45444 18396
rect 45948 18450 46004 18462
rect 45948 18398 45950 18450
rect 46002 18398 46004 18450
rect 45388 18174 45390 18226
rect 45442 18174 45444 18226
rect 45388 18116 45444 18174
rect 45052 17614 45054 17666
rect 45106 17614 45108 17666
rect 45052 17602 45108 17614
rect 45164 18060 45444 18116
rect 45836 18228 45892 18238
rect 45052 16884 45108 16894
rect 45164 16884 45220 18060
rect 45108 16828 45220 16884
rect 45388 17780 45444 17790
rect 45052 16818 45108 16828
rect 45388 16770 45444 17724
rect 45500 17778 45556 17790
rect 45500 17726 45502 17778
rect 45554 17726 45556 17778
rect 45500 17332 45556 17726
rect 45500 17266 45556 17276
rect 45836 17220 45892 18172
rect 45836 17154 45892 17164
rect 45948 16884 46004 18398
rect 46284 17108 46340 27468
rect 46396 25060 46452 27692
rect 46620 26852 46676 26862
rect 46620 26850 46788 26852
rect 46620 26798 46622 26850
rect 46674 26798 46788 26850
rect 46620 26796 46788 26798
rect 46620 26786 46676 26796
rect 46620 26628 46676 26638
rect 46508 26516 46564 26526
rect 46508 25284 46564 26460
rect 46620 26402 46676 26572
rect 46620 26350 46622 26402
rect 46674 26350 46676 26402
rect 46620 26338 46676 26350
rect 46732 25506 46788 26796
rect 46732 25454 46734 25506
rect 46786 25454 46788 25506
rect 46732 25442 46788 25454
rect 46508 25228 46788 25284
rect 46396 24388 46452 25004
rect 46396 24322 46452 24332
rect 46508 24498 46564 24510
rect 46508 24446 46510 24498
rect 46562 24446 46564 24498
rect 46508 23940 46564 24446
rect 46508 23874 46564 23884
rect 46508 23716 46564 23726
rect 46508 23622 46564 23660
rect 46508 23156 46564 23166
rect 46508 23062 46564 23100
rect 46620 22370 46676 22382
rect 46620 22318 46622 22370
rect 46674 22318 46676 22370
rect 46396 22036 46452 22046
rect 46396 20020 46452 21980
rect 46620 21028 46676 22318
rect 46732 21588 46788 25228
rect 46956 25282 47012 29036
rect 47404 28754 47460 28766
rect 47404 28702 47406 28754
rect 47458 28702 47460 28754
rect 47292 28642 47348 28654
rect 47292 28590 47294 28642
rect 47346 28590 47348 28642
rect 47292 28196 47348 28590
rect 47404 28420 47460 28702
rect 47628 28756 47684 28766
rect 47628 28662 47684 28700
rect 47404 28354 47460 28364
rect 47180 28140 47292 28196
rect 47180 27076 47236 28140
rect 47292 28130 47348 28140
rect 47292 27524 47348 27534
rect 47292 27298 47348 27468
rect 47292 27246 47294 27298
rect 47346 27246 47348 27298
rect 47292 27234 47348 27246
rect 47404 27188 47460 27198
rect 47404 27186 47684 27188
rect 47404 27134 47406 27186
rect 47458 27134 47684 27186
rect 47404 27132 47684 27134
rect 47404 27122 47460 27132
rect 47180 27020 47348 27076
rect 47292 26908 47348 27020
rect 47180 26850 47236 26862
rect 47292 26852 47460 26908
rect 47180 26798 47182 26850
rect 47234 26798 47236 26850
rect 47180 26292 47236 26798
rect 47180 26226 47236 26236
rect 47292 25732 47348 25742
rect 47404 25732 47460 26852
rect 47628 26516 47684 27132
rect 47628 26450 47684 26460
rect 47292 25730 47460 25732
rect 47292 25678 47294 25730
rect 47346 25678 47460 25730
rect 47292 25676 47460 25678
rect 47292 25666 47348 25676
rect 46956 25230 46958 25282
rect 47010 25230 47012 25282
rect 46844 24500 46900 24510
rect 46844 24406 46900 24444
rect 46844 23604 46900 23614
rect 46844 22708 46900 23548
rect 46844 22642 46900 22652
rect 46844 22482 46900 22494
rect 46844 22430 46846 22482
rect 46898 22430 46900 22482
rect 46844 21700 46900 22430
rect 46956 21812 47012 25230
rect 47068 25284 47124 25294
rect 47068 23604 47124 25228
rect 47404 24836 47460 24846
rect 47404 24742 47460 24780
rect 47068 23538 47124 23548
rect 46956 21746 47012 21756
rect 47068 23154 47124 23166
rect 47740 23156 47796 33628
rect 47852 33618 47908 33628
rect 48076 31948 48132 34076
rect 48188 32788 48244 35084
rect 48300 34916 48356 38668
rect 48412 38276 48468 38286
rect 48412 37378 48468 38220
rect 48412 37326 48414 37378
rect 48466 37326 48468 37378
rect 48412 37314 48468 37326
rect 48300 34850 48356 34860
rect 48412 35700 48468 35710
rect 48300 34244 48356 34254
rect 48300 34150 48356 34188
rect 48188 32722 48244 32732
rect 48412 33234 48468 35644
rect 48412 33182 48414 33234
rect 48466 33182 48468 33234
rect 48188 32340 48244 32350
rect 48188 32338 48356 32340
rect 48188 32286 48190 32338
rect 48242 32286 48356 32338
rect 48188 32284 48356 32286
rect 48188 32274 48244 32284
rect 48076 31892 48244 31948
rect 48188 31890 48244 31892
rect 48188 31838 48190 31890
rect 48242 31838 48244 31890
rect 48188 31826 48244 31838
rect 48076 31778 48132 31790
rect 48076 31726 48078 31778
rect 48130 31726 48132 31778
rect 47852 31556 47908 31566
rect 47852 30994 47908 31500
rect 47852 30942 47854 30994
rect 47906 30942 47908 30994
rect 47852 30930 47908 30942
rect 48076 30212 48132 31726
rect 48300 31556 48356 32284
rect 48412 32228 48468 33182
rect 48524 33124 48580 39564
rect 48860 39620 48916 40350
rect 48972 40292 49028 40684
rect 48972 40226 49028 40236
rect 49084 40068 49140 43036
rect 49420 41972 49476 43374
rect 49420 41906 49476 41916
rect 49532 44436 49588 44446
rect 49308 41748 49364 41758
rect 49308 41746 49476 41748
rect 49308 41694 49310 41746
rect 49362 41694 49476 41746
rect 49308 41692 49476 41694
rect 49308 41682 49364 41692
rect 49420 41412 49476 41692
rect 49308 41188 49364 41198
rect 49308 41094 49364 41132
rect 48860 39526 48916 39564
rect 48972 40012 49140 40068
rect 49196 41074 49252 41086
rect 49196 41022 49198 41074
rect 49250 41022 49252 41074
rect 48748 38610 48804 38622
rect 48748 38558 48750 38610
rect 48802 38558 48804 38610
rect 48636 34020 48692 34030
rect 48636 33572 48692 33964
rect 48748 33684 48804 38558
rect 48860 37938 48916 37950
rect 48860 37886 48862 37938
rect 48914 37886 48916 37938
rect 48860 37716 48916 37886
rect 48860 36260 48916 37660
rect 48860 35810 48916 36204
rect 48860 35758 48862 35810
rect 48914 35758 48916 35810
rect 48860 34244 48916 35758
rect 48860 34178 48916 34188
rect 48748 33628 48916 33684
rect 48636 33506 48692 33516
rect 48748 33458 48804 33470
rect 48748 33406 48750 33458
rect 48802 33406 48804 33458
rect 48748 33348 48804 33406
rect 48748 33282 48804 33292
rect 48524 33068 48804 33124
rect 48636 32788 48692 32798
rect 48636 32562 48692 32732
rect 48636 32510 48638 32562
rect 48690 32510 48692 32562
rect 48636 32498 48692 32510
rect 48748 32450 48804 33068
rect 48748 32398 48750 32450
rect 48802 32398 48804 32450
rect 48748 32386 48804 32398
rect 48412 32172 48692 32228
rect 48412 31780 48468 31790
rect 48412 31686 48468 31724
rect 48524 31778 48580 31790
rect 48524 31726 48526 31778
rect 48578 31726 48580 31778
rect 48300 31490 48356 31500
rect 48524 31556 48580 31726
rect 48524 31490 48580 31500
rect 48300 31220 48356 31230
rect 48300 30996 48356 31164
rect 48524 31220 48580 31230
rect 48524 31126 48580 31164
rect 48412 30996 48468 31006
rect 48300 30994 48468 30996
rect 48300 30942 48414 30994
rect 48466 30942 48468 30994
rect 48300 30940 48468 30942
rect 48412 30930 48468 30940
rect 48524 30996 48580 31006
rect 48524 30882 48580 30940
rect 48524 30830 48526 30882
rect 48578 30830 48580 30882
rect 48524 30818 48580 30830
rect 48076 30146 48132 30156
rect 48300 30324 48356 30334
rect 48300 30210 48356 30268
rect 48300 30158 48302 30210
rect 48354 30158 48356 30210
rect 48300 30146 48356 30158
rect 48412 30212 48468 30222
rect 48636 30212 48692 32172
rect 48636 30156 48804 30212
rect 48188 29986 48244 29998
rect 48188 29934 48190 29986
rect 48242 29934 48244 29986
rect 48188 29540 48244 29934
rect 48188 29474 48244 29484
rect 48412 29428 48468 30156
rect 47964 29202 48020 29214
rect 47964 29150 47966 29202
rect 48018 29150 48020 29202
rect 47964 28532 48020 29150
rect 48412 29092 48468 29372
rect 48524 29986 48580 29998
rect 48524 29934 48526 29986
rect 48578 29934 48580 29986
rect 48524 29204 48580 29934
rect 48636 29988 48692 29998
rect 48636 29894 48692 29932
rect 48748 29764 48804 30156
rect 48524 29138 48580 29148
rect 48636 29708 48804 29764
rect 48412 29026 48468 29036
rect 48636 28868 48692 29708
rect 48412 28812 48692 28868
rect 48188 28644 48244 28654
rect 48188 28550 48244 28588
rect 47964 28466 48020 28476
rect 48076 27746 48132 27758
rect 48076 27694 48078 27746
rect 48130 27694 48132 27746
rect 47852 24612 47908 24622
rect 47852 24052 47908 24556
rect 47852 23986 47908 23996
rect 48076 23938 48132 27694
rect 48188 26964 48244 27002
rect 48188 26898 48244 26908
rect 48188 26516 48244 26526
rect 48188 25730 48244 26460
rect 48188 25678 48190 25730
rect 48242 25678 48244 25730
rect 48188 25666 48244 25678
rect 48076 23886 48078 23938
rect 48130 23886 48132 23938
rect 47068 23102 47070 23154
rect 47122 23102 47124 23154
rect 47068 21810 47124 23102
rect 47404 23100 47796 23156
rect 47852 23156 47908 23166
rect 47180 22932 47236 22942
rect 47180 22594 47236 22876
rect 47180 22542 47182 22594
rect 47234 22542 47236 22594
rect 47180 22530 47236 22542
rect 47404 22596 47460 23100
rect 47852 23062 47908 23100
rect 47740 22932 47796 22942
rect 47740 22930 48020 22932
rect 47740 22878 47742 22930
rect 47794 22878 48020 22930
rect 47740 22876 48020 22878
rect 47740 22866 47796 22876
rect 47404 22530 47460 22540
rect 47740 22596 47796 22606
rect 47516 22482 47572 22494
rect 47516 22430 47518 22482
rect 47570 22430 47572 22482
rect 47516 22372 47572 22430
rect 47068 21758 47070 21810
rect 47122 21758 47124 21810
rect 47068 21746 47124 21758
rect 47292 22316 47572 22372
rect 46844 21634 46900 21644
rect 46732 21522 46788 21532
rect 46620 20962 46676 20972
rect 46732 21364 46788 21374
rect 46508 20914 46564 20926
rect 46508 20862 46510 20914
rect 46562 20862 46564 20914
rect 46508 20580 46564 20862
rect 46508 20514 46564 20524
rect 46396 19234 46452 19964
rect 46732 20018 46788 21308
rect 47180 21028 47236 21038
rect 47180 20934 47236 20972
rect 46844 20916 46900 20926
rect 46844 20822 46900 20860
rect 47180 20468 47236 20478
rect 46732 19966 46734 20018
rect 46786 19966 46788 20018
rect 46732 19954 46788 19966
rect 46844 20356 46900 20366
rect 46396 19182 46398 19234
rect 46450 19182 46452 19234
rect 46396 19170 46452 19182
rect 46508 19908 46564 19918
rect 46508 17220 46564 19852
rect 46620 19236 46676 19246
rect 46620 17890 46676 19180
rect 46732 18564 46788 18574
rect 46732 18338 46788 18508
rect 46732 18286 46734 18338
rect 46786 18286 46788 18338
rect 46732 18274 46788 18286
rect 46620 17838 46622 17890
rect 46674 17838 46676 17890
rect 46620 17826 46676 17838
rect 46508 17154 46564 17164
rect 46844 17108 46900 20300
rect 47068 20020 47124 20030
rect 47068 19926 47124 19964
rect 47068 19796 47124 19806
rect 46956 18450 47012 18462
rect 46956 18398 46958 18450
rect 47010 18398 47012 18450
rect 46956 18340 47012 18398
rect 46956 18274 47012 18284
rect 47068 18004 47124 19740
rect 47180 18340 47236 20412
rect 47292 18788 47348 22316
rect 47404 22036 47460 22046
rect 47404 20188 47460 21980
rect 47516 21476 47572 21486
rect 47516 21026 47572 21420
rect 47740 21476 47796 22540
rect 47740 21410 47796 21420
rect 47852 22372 47908 22382
rect 47628 21364 47684 21374
rect 47628 21270 47684 21308
rect 47852 21364 47908 22316
rect 47852 21298 47908 21308
rect 47516 20974 47518 21026
rect 47570 20974 47572 21026
rect 47516 20962 47572 20974
rect 47404 20132 47684 20188
rect 47404 20020 47460 20030
rect 47404 19234 47460 19964
rect 47404 19182 47406 19234
rect 47458 19182 47460 19234
rect 47404 19170 47460 19182
rect 47292 18722 47348 18732
rect 47180 18274 47236 18284
rect 47516 18226 47572 18238
rect 47516 18174 47518 18226
rect 47570 18174 47572 18226
rect 47516 18116 47572 18174
rect 46956 17948 47124 18004
rect 47180 18060 47572 18116
rect 46956 17556 47012 17948
rect 47180 17890 47236 18060
rect 47180 17838 47182 17890
rect 47234 17838 47236 17890
rect 47180 17826 47236 17838
rect 47068 17780 47124 17790
rect 47068 17686 47124 17724
rect 47404 17666 47460 17678
rect 47404 17614 47406 17666
rect 47458 17614 47460 17666
rect 46956 17500 47236 17556
rect 46284 17052 46452 17108
rect 46844 17052 47124 17108
rect 45388 16718 45390 16770
rect 45442 16718 45444 16770
rect 45388 16706 45444 16718
rect 45836 16882 46004 16884
rect 45836 16830 45950 16882
rect 46002 16830 46004 16882
rect 45836 16828 46004 16830
rect 45500 16548 45556 16558
rect 44940 15250 44996 15260
rect 45052 16212 45108 16222
rect 44940 14980 44996 14990
rect 44940 14754 44996 14924
rect 44940 14702 44942 14754
rect 44994 14702 44996 14754
rect 44940 14690 44996 14702
rect 44828 14478 44830 14530
rect 44882 14478 44884 14530
rect 44828 14420 44884 14478
rect 44380 14364 44884 14420
rect 43932 14252 44212 14308
rect 43804 14140 44068 14150
rect 43860 14084 43908 14140
rect 43964 14084 44012 14140
rect 43804 14074 44068 14084
rect 44156 14084 44212 14252
rect 44156 14018 44212 14028
rect 43484 13918 43486 13970
rect 43538 13918 43540 13970
rect 43484 13906 43540 13918
rect 43708 13860 43764 13870
rect 43372 13570 43428 13580
rect 43596 13804 43708 13860
rect 43596 13634 43652 13804
rect 43708 13794 43764 13804
rect 44156 13860 44212 13870
rect 44380 13860 44436 14364
rect 44156 13858 44436 13860
rect 44156 13806 44158 13858
rect 44210 13806 44436 13858
rect 44156 13804 44436 13806
rect 44828 14196 44884 14206
rect 44156 13794 44212 13804
rect 44492 13748 44548 13758
rect 44492 13654 44548 13692
rect 44716 13748 44772 13758
rect 43596 13582 43598 13634
rect 43650 13582 43652 13634
rect 43596 13524 43652 13582
rect 43596 13458 43652 13468
rect 44044 13524 44100 13534
rect 44716 13524 44772 13692
rect 44100 13468 44772 13524
rect 44044 13458 44100 13468
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 43484 13188 43540 13198
rect 43372 12962 43428 12974
rect 43372 12910 43374 12962
rect 43426 12910 43428 12962
rect 43260 12740 43316 12750
rect 43260 12178 43316 12684
rect 43260 12126 43262 12178
rect 43314 12126 43316 12178
rect 43260 11844 43316 12126
rect 43260 11778 43316 11788
rect 43148 10782 43150 10834
rect 43202 10782 43204 10834
rect 43148 10770 43204 10782
rect 43372 11396 43428 12910
rect 43484 12964 43540 13132
rect 44492 13132 44660 13188
rect 44492 13074 44548 13132
rect 44492 13022 44494 13074
rect 44546 13022 44548 13074
rect 44492 13010 44548 13022
rect 44604 13076 44660 13132
rect 44604 13010 44660 13020
rect 43484 12898 43540 12908
rect 44044 12962 44100 12974
rect 44044 12910 44046 12962
rect 44098 12910 44100 12962
rect 44044 12740 44100 12910
rect 44380 12964 44436 12974
rect 44380 12740 44436 12908
rect 44604 12740 44660 12750
rect 44044 12684 44212 12740
rect 44380 12684 44604 12740
rect 43804 12572 44068 12582
rect 43484 12516 43540 12526
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 43484 11788 43540 12460
rect 43484 11732 43652 11788
rect 43372 10612 43428 11340
rect 43036 10556 43428 10612
rect 43484 11394 43540 11406
rect 43484 11342 43486 11394
rect 43538 11342 43540 11394
rect 42588 10220 42756 10276
rect 42588 10052 42644 10062
rect 42476 10050 42644 10052
rect 42476 9998 42590 10050
rect 42642 9998 42644 10050
rect 42476 9996 42644 9998
rect 42588 9986 42644 9996
rect 42700 9380 42756 10220
rect 43036 9828 43092 10556
rect 43484 10500 43540 11342
rect 43148 10444 43540 10500
rect 43148 10050 43204 10444
rect 43148 9998 43150 10050
rect 43202 9998 43204 10050
rect 43148 9986 43204 9998
rect 43596 10052 43652 11732
rect 44156 11620 44212 12684
rect 44604 12674 44660 12684
rect 44828 11956 44884 14140
rect 44940 13746 44996 13758
rect 44940 13694 44942 13746
rect 44994 13694 44996 13746
rect 44940 13636 44996 13694
rect 44940 13570 44996 13580
rect 44940 13300 44996 13310
rect 44940 13076 44996 13244
rect 44940 12628 44996 13020
rect 44940 12562 44996 12572
rect 44828 11890 44884 11900
rect 44044 11564 44212 11620
rect 44268 11844 44324 11854
rect 44268 11620 44324 11788
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44268 11564 44772 11620
rect 44044 11508 44100 11564
rect 44044 11442 44100 11452
rect 44156 11396 44212 11406
rect 44156 11302 44212 11340
rect 44044 11284 44100 11294
rect 44044 11172 44100 11228
rect 44044 11116 44212 11172
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44156 10610 44212 11116
rect 44268 11060 44324 11070
rect 44268 10722 44324 11004
rect 44268 10670 44270 10722
rect 44322 10670 44324 10722
rect 44268 10658 44324 10670
rect 44492 10948 44548 10958
rect 44492 10724 44548 10892
rect 44492 10658 44548 10668
rect 44716 10724 44772 11564
rect 45052 11394 45108 16156
rect 45388 16212 45444 16222
rect 45388 16118 45444 16156
rect 45500 16210 45556 16492
rect 45500 16158 45502 16210
rect 45554 16158 45556 16210
rect 45500 16146 45556 16158
rect 45612 16098 45668 16110
rect 45612 16046 45614 16098
rect 45666 16046 45668 16098
rect 45388 15988 45444 15998
rect 45388 15540 45444 15932
rect 45612 15988 45668 16046
rect 45612 15922 45668 15932
rect 45388 15474 45444 15484
rect 45388 15316 45444 15326
rect 45164 15204 45220 15214
rect 45388 15204 45444 15260
rect 45164 15202 45444 15204
rect 45164 15150 45166 15202
rect 45218 15150 45444 15202
rect 45164 15148 45444 15150
rect 45164 15138 45220 15148
rect 45164 14868 45220 14878
rect 45164 14754 45220 14812
rect 45164 14702 45166 14754
rect 45218 14702 45220 14754
rect 45164 14690 45220 14702
rect 45724 14532 45780 14542
rect 45836 14532 45892 16828
rect 45948 16818 46004 16828
rect 46284 16884 46340 16894
rect 46284 16790 46340 16828
rect 46396 16660 46452 17052
rect 46956 16884 47012 16894
rect 46956 16790 47012 16828
rect 45780 14476 45892 14532
rect 45948 16604 46452 16660
rect 46620 16660 46676 16670
rect 45500 13972 45556 13982
rect 45164 13524 45220 13534
rect 45164 13430 45220 13468
rect 45052 11342 45054 11394
rect 45106 11342 45108 11394
rect 45052 11330 45108 11342
rect 45164 13076 45220 13086
rect 44716 10658 44772 10668
rect 44156 10558 44158 10610
rect 44210 10558 44212 10610
rect 44156 10546 44212 10558
rect 44380 10500 44436 10510
rect 44380 10406 44436 10444
rect 44604 10388 44660 10426
rect 44604 10322 44660 10332
rect 43596 9986 43652 9996
rect 44268 10276 44324 10286
rect 44044 9940 44100 9950
rect 43932 9828 43988 9838
rect 43036 9772 43316 9828
rect 42700 9314 42756 9324
rect 42588 9044 42644 9054
rect 42588 8950 42644 8988
rect 43036 8932 43092 8942
rect 42476 8372 42532 8382
rect 42476 8278 42532 8316
rect 43036 8372 43092 8876
rect 43036 8306 43092 8316
rect 43148 8818 43204 8830
rect 43148 8766 43150 8818
rect 43202 8766 43204 8818
rect 42364 8092 42532 8148
rect 42140 7364 42196 7374
rect 42140 7270 42196 7308
rect 42252 6916 42308 6926
rect 41692 6018 41972 6020
rect 41692 5966 41918 6018
rect 41970 5966 41972 6018
rect 41692 5964 41972 5966
rect 41468 5796 41524 5806
rect 41356 5236 41412 5246
rect 41356 5142 41412 5180
rect 41132 4834 41188 4844
rect 41244 5124 41300 5134
rect 41244 4338 41300 5068
rect 41244 4286 41246 4338
rect 41298 4286 41300 4338
rect 41244 4274 41300 4286
rect 41356 4228 41412 4238
rect 41468 4228 41524 5740
rect 41356 4226 41524 4228
rect 41356 4174 41358 4226
rect 41410 4174 41524 4226
rect 41356 4172 41524 4174
rect 41356 4162 41412 4172
rect 40908 3668 40964 3678
rect 40908 3574 40964 3612
rect 41692 3444 41748 5964
rect 41916 5954 41972 5964
rect 42140 6468 42196 6478
rect 41804 5124 41860 5134
rect 42140 5124 42196 6412
rect 42252 5794 42308 6860
rect 42364 6804 42420 6814
rect 42364 6690 42420 6748
rect 42364 6638 42366 6690
rect 42418 6638 42420 6690
rect 42364 6626 42420 6638
rect 42252 5742 42254 5794
rect 42306 5742 42308 5794
rect 42252 5730 42308 5742
rect 42364 5348 42420 5358
rect 42476 5348 42532 8092
rect 42924 8146 42980 8158
rect 42924 8094 42926 8146
rect 42978 8094 42980 8146
rect 42924 7140 42980 8094
rect 43148 8148 43204 8766
rect 43148 8082 43204 8092
rect 42924 7074 42980 7084
rect 43260 6690 43316 9772
rect 43932 9604 43988 9772
rect 44044 9716 44100 9884
rect 44268 9940 44324 10220
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44492 10052 44548 10062
rect 44268 9874 44324 9884
rect 44380 9996 44492 10052
rect 44380 9938 44436 9996
rect 44492 9986 44548 9996
rect 44380 9886 44382 9938
rect 44434 9886 44436 9938
rect 44380 9874 44436 9886
rect 44828 9828 44884 9838
rect 45164 9828 45220 13020
rect 45388 12180 45444 12190
rect 44828 9826 45220 9828
rect 44828 9774 44830 9826
rect 44882 9774 45220 9826
rect 44828 9772 45220 9774
rect 45276 10612 45332 10622
rect 44828 9762 44884 9772
rect 44044 9660 44660 9716
rect 43932 9548 44212 9604
rect 43804 9436 44068 9446
rect 43484 9380 43540 9390
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 44156 9380 44212 9548
rect 43484 9154 43540 9324
rect 44156 9314 44212 9324
rect 44604 9492 44660 9660
rect 44604 9266 44660 9436
rect 44604 9214 44606 9266
rect 44658 9214 44660 9266
rect 44604 9202 44660 9214
rect 44268 9156 44324 9166
rect 43484 9102 43486 9154
rect 43538 9102 43540 9154
rect 43484 9090 43540 9102
rect 43596 9154 44324 9156
rect 43596 9102 44270 9154
rect 44322 9102 44324 9154
rect 43596 9100 44324 9102
rect 43596 9042 43652 9100
rect 44268 9090 44324 9100
rect 43596 8990 43598 9042
rect 43650 8990 43652 9042
rect 43596 8978 43652 8990
rect 44044 8932 44100 8942
rect 43372 8818 43428 8830
rect 43372 8766 43374 8818
rect 43426 8766 43428 8818
rect 43372 8260 43428 8766
rect 44044 8482 44100 8876
rect 44828 8932 44884 8942
rect 44828 8838 44884 8876
rect 44940 8708 44996 9772
rect 44464 8652 44728 8662
rect 44044 8430 44046 8482
rect 44098 8430 44100 8482
rect 43484 8260 43540 8270
rect 43372 8258 43540 8260
rect 43372 8206 43486 8258
rect 43538 8206 43540 8258
rect 43372 8204 43540 8206
rect 43372 7698 43428 8204
rect 43484 8194 43540 8204
rect 43820 8260 43876 8270
rect 43820 8166 43876 8204
rect 43932 8148 43988 8158
rect 43932 8054 43988 8092
rect 44044 8036 44100 8430
rect 44268 8596 44324 8606
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44828 8652 44940 8708
rect 44268 8484 44324 8540
rect 44828 8484 44884 8652
rect 44940 8642 44996 8652
rect 45052 9492 45108 9502
rect 44268 8428 44884 8484
rect 44044 7970 44100 7980
rect 44268 8258 44324 8270
rect 44268 8206 44270 8258
rect 44322 8206 44324 8258
rect 43372 7646 43374 7698
rect 43426 7646 43428 7698
rect 43372 7634 43428 7646
rect 43596 7924 43652 7934
rect 43596 7700 43652 7868
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 44268 7700 44324 8206
rect 44828 8258 44884 8270
rect 44828 8206 44830 8258
rect 44882 8206 44884 8258
rect 44828 7812 44884 8206
rect 44828 7746 44884 7756
rect 43596 7644 44212 7700
rect 43260 6638 43262 6690
rect 43314 6638 43316 6690
rect 43260 6626 43316 6638
rect 44156 7476 44212 7644
rect 44268 7634 44324 7644
rect 44268 7476 44324 7486
rect 44156 7474 44324 7476
rect 44156 7422 44270 7474
rect 44322 7422 44324 7474
rect 44156 7420 44324 7422
rect 44044 6580 44100 6590
rect 44156 6580 44212 7420
rect 44268 7410 44324 7420
rect 44828 7364 44884 7374
rect 44828 7270 44884 7308
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 45052 6916 45108 9436
rect 44604 6860 45108 6916
rect 45164 8930 45220 8942
rect 45164 8878 45166 8930
rect 45218 8878 45220 8930
rect 44380 6802 44436 6814
rect 44380 6750 44382 6802
rect 44434 6750 44436 6802
rect 44380 6692 44436 6750
rect 44380 6626 44436 6636
rect 44044 6578 44212 6580
rect 44044 6526 44046 6578
rect 44098 6526 44212 6578
rect 44044 6524 44212 6526
rect 44044 6514 44100 6524
rect 44492 6468 44548 6478
rect 44268 6412 44492 6468
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 44268 6130 44324 6412
rect 44492 6402 44548 6412
rect 44268 6078 44270 6130
rect 44322 6078 44324 6130
rect 44268 6066 44324 6078
rect 44604 6130 44660 6860
rect 44940 6244 44996 6254
rect 45164 6244 45220 8878
rect 45276 8370 45332 10556
rect 45388 9492 45444 12124
rect 45500 11732 45556 13916
rect 45612 13634 45668 13646
rect 45612 13582 45614 13634
rect 45666 13582 45668 13634
rect 45612 13186 45668 13582
rect 45612 13134 45614 13186
rect 45666 13134 45668 13186
rect 45612 13122 45668 13134
rect 45500 11666 45556 11676
rect 45388 9426 45444 9436
rect 45612 11508 45668 11518
rect 45612 11396 45668 11452
rect 45724 11396 45780 14476
rect 45612 11394 45780 11396
rect 45612 11342 45726 11394
rect 45778 11342 45780 11394
rect 45612 11340 45780 11342
rect 45276 8318 45278 8370
rect 45330 8318 45332 8370
rect 45276 8306 45332 8318
rect 45612 7812 45668 11340
rect 45724 11330 45780 11340
rect 45948 10724 46004 16604
rect 46620 16566 46676 16604
rect 46844 16658 46900 16670
rect 47068 16660 47124 17052
rect 46844 16606 46846 16658
rect 46898 16606 46900 16658
rect 46396 16324 46452 16334
rect 46844 16324 46900 16606
rect 46060 16322 46452 16324
rect 46060 16270 46398 16322
rect 46450 16270 46452 16322
rect 46060 16268 46452 16270
rect 46060 16098 46116 16268
rect 46396 16258 46452 16268
rect 46508 16268 46900 16324
rect 46956 16604 47124 16660
rect 46060 16046 46062 16098
rect 46114 16046 46116 16098
rect 46060 16034 46116 16046
rect 46172 16098 46228 16110
rect 46172 16046 46174 16098
rect 46226 16046 46228 16098
rect 46172 15204 46228 16046
rect 46284 15540 46340 15550
rect 46508 15540 46564 16268
rect 46284 15538 46564 15540
rect 46284 15486 46286 15538
rect 46338 15486 46564 15538
rect 46284 15484 46564 15486
rect 46620 16098 46676 16110
rect 46620 16046 46622 16098
rect 46674 16046 46676 16098
rect 46620 15988 46676 16046
rect 46732 16098 46788 16268
rect 46732 16046 46734 16098
rect 46786 16046 46788 16098
rect 46732 16034 46788 16046
rect 46284 15474 46340 15484
rect 46172 14868 46228 15148
rect 46172 14802 46228 14812
rect 46620 14980 46676 15932
rect 46844 15540 46900 15550
rect 46844 15314 46900 15484
rect 46956 15428 47012 16604
rect 47180 16436 47236 17500
rect 47404 16996 47460 17614
rect 47628 17556 47684 20132
rect 47964 20020 48020 22876
rect 48076 22260 48132 23886
rect 48188 25284 48244 25294
rect 48188 22708 48244 25228
rect 48300 23716 48356 23726
rect 48300 23154 48356 23660
rect 48300 23102 48302 23154
rect 48354 23102 48356 23154
rect 48300 23090 48356 23102
rect 48188 22652 48356 22708
rect 48188 22484 48244 22494
rect 48188 22390 48244 22428
rect 48076 22204 48244 22260
rect 48076 20020 48132 20030
rect 48020 20018 48132 20020
rect 48020 19966 48078 20018
rect 48130 19966 48132 20018
rect 48020 19964 48132 19966
rect 47964 19926 48020 19964
rect 48076 19954 48132 19964
rect 48076 19346 48132 19358
rect 48076 19294 48078 19346
rect 48130 19294 48132 19346
rect 47628 17490 47684 17500
rect 47852 19236 47908 19246
rect 47404 16930 47460 16940
rect 47516 17332 47572 17342
rect 47292 16884 47348 16894
rect 47292 16770 47348 16828
rect 47292 16718 47294 16770
rect 47346 16718 47348 16770
rect 47292 16706 47348 16718
rect 47404 16660 47460 16670
rect 47404 16566 47460 16604
rect 47180 16212 47236 16380
rect 47180 16210 47348 16212
rect 47180 16158 47182 16210
rect 47234 16158 47348 16210
rect 47180 16156 47348 16158
rect 47180 16146 47236 16156
rect 46956 15362 47012 15372
rect 46844 15262 46846 15314
rect 46898 15262 46900 15314
rect 46844 15250 46900 15262
rect 47180 15316 47236 15326
rect 47292 15316 47348 16156
rect 47404 16210 47460 16222
rect 47404 16158 47406 16210
rect 47458 16158 47460 16210
rect 47404 15540 47460 16158
rect 47516 16212 47572 17276
rect 47628 17220 47684 17230
rect 47628 16882 47684 17164
rect 47628 16830 47630 16882
rect 47682 16830 47684 16882
rect 47628 16818 47684 16830
rect 47516 16146 47572 16156
rect 47516 15876 47572 15886
rect 47516 15874 47684 15876
rect 47516 15822 47518 15874
rect 47570 15822 47684 15874
rect 47516 15820 47684 15822
rect 47516 15810 47572 15820
rect 47404 15484 47572 15540
rect 47404 15316 47460 15326
rect 47292 15314 47460 15316
rect 47292 15262 47406 15314
rect 47458 15262 47460 15314
rect 47292 15260 47460 15262
rect 46956 15204 47012 15242
rect 47180 15222 47236 15260
rect 47404 15250 47460 15260
rect 46956 15138 47012 15148
rect 47516 15202 47572 15484
rect 47516 15150 47518 15202
rect 47570 15150 47572 15202
rect 46172 14642 46228 14654
rect 46172 14590 46174 14642
rect 46226 14590 46228 14642
rect 46172 14532 46228 14590
rect 46172 14466 46228 14476
rect 46060 14420 46116 14430
rect 46060 13074 46116 14364
rect 46172 13860 46228 13870
rect 46172 13746 46228 13804
rect 46172 13694 46174 13746
rect 46226 13694 46228 13746
rect 46172 13682 46228 13694
rect 46620 13186 46676 14924
rect 47516 15092 47572 15150
rect 47180 14868 47236 14878
rect 47180 13746 47236 14812
rect 47516 14756 47572 15036
rect 47628 14868 47684 15820
rect 47740 15428 47796 15438
rect 47740 15314 47796 15372
rect 47740 15262 47742 15314
rect 47794 15262 47796 15314
rect 47740 15250 47796 15262
rect 47852 14980 47908 19180
rect 48076 19012 48132 19294
rect 48076 18946 48132 18956
rect 47852 14914 47908 14924
rect 47964 18676 48020 18686
rect 47628 14802 47684 14812
rect 47516 14690 47572 14700
rect 47404 14420 47460 14430
rect 47180 13694 47182 13746
rect 47234 13694 47236 13746
rect 47180 13682 47236 13694
rect 47292 14306 47348 14318
rect 47292 14254 47294 14306
rect 47346 14254 47348 14306
rect 47292 13636 47348 14254
rect 47404 14196 47460 14364
rect 47964 14420 48020 18620
rect 48188 17666 48244 22204
rect 48300 18676 48356 22652
rect 48412 21028 48468 28812
rect 48524 28420 48580 28430
rect 48524 26908 48580 28364
rect 48524 26852 48804 26908
rect 48748 26402 48804 26852
rect 48748 26350 48750 26402
rect 48802 26350 48804 26402
rect 48748 26338 48804 26350
rect 48860 24276 48916 33628
rect 48972 32562 49028 40012
rect 49084 38834 49140 38846
rect 49084 38782 49086 38834
rect 49138 38782 49140 38834
rect 49084 38276 49140 38782
rect 49084 38210 49140 38220
rect 49196 37940 49252 41022
rect 49420 40404 49476 41356
rect 49308 40292 49364 40302
rect 49308 40198 49364 40236
rect 49308 39844 49364 39854
rect 49420 39844 49476 40348
rect 49308 39842 49476 39844
rect 49308 39790 49310 39842
rect 49362 39790 49476 39842
rect 49308 39788 49476 39790
rect 49308 39778 49364 39788
rect 49420 38722 49476 38734
rect 49420 38670 49422 38722
rect 49474 38670 49476 38722
rect 49196 37874 49252 37884
rect 49308 38164 49364 38174
rect 49084 37716 49140 37726
rect 49084 37378 49140 37660
rect 49084 37326 49086 37378
rect 49138 37326 49140 37378
rect 49084 37314 49140 37326
rect 49084 36260 49140 36270
rect 49084 35476 49140 36204
rect 49196 36148 49252 36158
rect 49196 35586 49252 36092
rect 49308 35700 49364 38108
rect 49420 36036 49476 38670
rect 49532 38668 49588 44380
rect 49644 41186 49700 45388
rect 49756 44884 49812 44894
rect 49756 44790 49812 44828
rect 49980 44884 50036 44894
rect 49756 43428 49812 43438
rect 49756 43334 49812 43372
rect 49980 42866 50036 44828
rect 50092 44546 50148 45724
rect 50204 45668 50260 46060
rect 50316 45892 50372 45902
rect 50316 45798 50372 45836
rect 50204 45602 50260 45612
rect 50428 45668 50484 45678
rect 50428 45444 50484 45612
rect 50092 44494 50094 44546
rect 50146 44494 50148 44546
rect 50092 44482 50148 44494
rect 50204 45388 50484 45444
rect 49980 42814 49982 42866
rect 50034 42814 50036 42866
rect 49980 42802 50036 42814
rect 49644 41134 49646 41186
rect 49698 41134 49700 41186
rect 49644 41122 49700 41134
rect 49756 42420 49812 42430
rect 49756 41076 49812 42364
rect 49756 41010 49812 41020
rect 49868 41972 49924 41982
rect 49868 40628 49924 41916
rect 49980 41524 50036 41534
rect 49980 41410 50036 41468
rect 49980 41358 49982 41410
rect 50034 41358 50036 41410
rect 49980 41346 50036 41358
rect 50204 41298 50260 45388
rect 50540 44548 50596 48412
rect 50652 48242 50708 48254
rect 50652 48190 50654 48242
rect 50706 48190 50708 48242
rect 50652 47348 50708 48190
rect 50876 48244 50932 48254
rect 50876 48150 50932 48188
rect 50764 47684 50820 47694
rect 50988 47684 51044 49758
rect 51100 48468 51156 50372
rect 51436 50372 51492 50382
rect 51212 49810 51268 49822
rect 51212 49758 51214 49810
rect 51266 49758 51268 49810
rect 51212 49700 51268 49758
rect 51212 49634 51268 49644
rect 51324 49810 51380 49822
rect 51324 49758 51326 49810
rect 51378 49758 51380 49810
rect 51324 49028 51380 49758
rect 51100 48402 51156 48412
rect 51212 48972 51380 49028
rect 51100 48244 51156 48254
rect 51212 48244 51268 48972
rect 51100 48242 51268 48244
rect 51100 48190 51102 48242
rect 51154 48190 51268 48242
rect 51100 48188 51268 48190
rect 51324 48802 51380 48814
rect 51324 48750 51326 48802
rect 51378 48750 51380 48802
rect 51100 48132 51156 48188
rect 51100 48066 51156 48076
rect 50764 47682 51044 47684
rect 50764 47630 50766 47682
rect 50818 47630 51044 47682
rect 50764 47628 51044 47630
rect 50764 47618 50820 47628
rect 51212 47572 51268 47582
rect 51324 47572 51380 48750
rect 51212 47570 51380 47572
rect 51212 47518 51214 47570
rect 51266 47518 51380 47570
rect 51212 47516 51380 47518
rect 51212 47506 51268 47516
rect 51436 47460 51492 50316
rect 51548 49364 51604 50876
rect 51548 49298 51604 49308
rect 51660 48804 51716 54012
rect 51884 53842 51940 53854
rect 51884 53790 51886 53842
rect 51938 53790 51940 53842
rect 51884 53620 51940 53790
rect 51884 53554 51940 53564
rect 52108 53730 52164 53742
rect 52108 53678 52110 53730
rect 52162 53678 52164 53730
rect 51996 52724 52052 52734
rect 51772 52722 52052 52724
rect 51772 52670 51998 52722
rect 52050 52670 52052 52722
rect 51772 52668 52052 52670
rect 51772 51492 51828 52668
rect 51996 52658 52052 52668
rect 51996 52500 52052 52510
rect 51884 52276 51940 52286
rect 51884 52182 51940 52220
rect 51772 51426 51828 51436
rect 51996 50818 52052 52444
rect 52108 51604 52164 53678
rect 52220 53172 52276 55806
rect 52892 55860 52948 55870
rect 52892 55766 52948 55804
rect 52668 55524 52724 55534
rect 52668 54402 52724 55468
rect 53452 55076 53508 56252
rect 54572 56084 54628 56094
rect 54124 56082 54628 56084
rect 54124 56030 54574 56082
rect 54626 56030 54628 56082
rect 54124 56028 54628 56030
rect 53564 55972 53620 55982
rect 53564 55878 53620 55916
rect 53676 55412 53732 55422
rect 53452 55010 53508 55020
rect 53564 55410 53732 55412
rect 53564 55358 53678 55410
rect 53730 55358 53732 55410
rect 53564 55356 53732 55358
rect 53004 54516 53060 54526
rect 53004 54514 53508 54516
rect 53004 54462 53006 54514
rect 53058 54462 53508 54514
rect 53004 54460 53508 54462
rect 53004 54450 53060 54460
rect 52668 54350 52670 54402
rect 52722 54350 52724 54402
rect 52668 54338 52724 54350
rect 52332 54292 52388 54302
rect 52332 54290 52612 54292
rect 52332 54238 52334 54290
rect 52386 54238 52612 54290
rect 52332 54236 52612 54238
rect 52332 54226 52388 54236
rect 52556 54068 52612 54236
rect 53340 54290 53396 54302
rect 53340 54238 53342 54290
rect 53394 54238 53396 54290
rect 52556 54012 53284 54068
rect 53228 53954 53284 54012
rect 53228 53902 53230 53954
rect 53282 53902 53284 53954
rect 53228 53890 53284 53902
rect 52892 53842 52948 53854
rect 52892 53790 52894 53842
rect 52946 53790 52948 53842
rect 52556 53732 52612 53742
rect 52556 53638 52612 53676
rect 52556 53508 52612 53518
rect 52220 53116 52500 53172
rect 52332 52948 52388 52958
rect 52332 52834 52388 52892
rect 52332 52782 52334 52834
rect 52386 52782 52388 52834
rect 52332 52770 52388 52782
rect 52220 52724 52276 52734
rect 52220 52388 52276 52668
rect 52220 52332 52388 52388
rect 52220 52052 52276 52062
rect 52220 51958 52276 51996
rect 52108 51548 52276 51604
rect 52108 51380 52164 51390
rect 52108 51286 52164 51324
rect 51996 50766 51998 50818
rect 52050 50766 52052 50818
rect 51996 50754 52052 50766
rect 52108 51156 52164 51166
rect 52108 50698 52164 51100
rect 52220 50932 52276 51548
rect 52332 51266 52388 52332
rect 52332 51214 52334 51266
rect 52386 51214 52388 51266
rect 52332 51202 52388 51214
rect 52220 50876 52388 50932
rect 51884 50642 52164 50698
rect 52220 50708 52276 50718
rect 51884 49700 51940 50642
rect 51884 49634 51940 49644
rect 52108 49924 52164 49934
rect 51996 49586 52052 49598
rect 51996 49534 51998 49586
rect 52050 49534 52052 49586
rect 51996 49140 52052 49534
rect 51996 49074 52052 49084
rect 51660 48738 51716 48748
rect 51884 48802 51940 48814
rect 51884 48750 51886 48802
rect 51938 48750 51940 48802
rect 51772 48580 51828 48590
rect 51660 48244 51716 48254
rect 51548 48018 51604 48030
rect 51548 47966 51550 48018
rect 51602 47966 51604 48018
rect 51548 47684 51604 47966
rect 51548 47618 51604 47628
rect 51436 47394 51492 47404
rect 51548 47460 51604 47470
rect 51660 47460 51716 48188
rect 51548 47458 51716 47460
rect 51548 47406 51550 47458
rect 51602 47406 51716 47458
rect 51548 47404 51716 47406
rect 50652 47292 51380 47348
rect 50764 46900 50820 46910
rect 50652 46676 50708 46686
rect 50652 44884 50708 46620
rect 50764 46340 50820 46844
rect 51324 46898 51380 47292
rect 51324 46846 51326 46898
rect 51378 46846 51380 46898
rect 51324 46834 51380 46846
rect 51436 47236 51492 47246
rect 51436 46676 51492 47180
rect 50764 46274 50820 46284
rect 50876 46620 51492 46676
rect 50764 45892 50820 45902
rect 50764 45798 50820 45836
rect 50876 45556 50932 46620
rect 51436 46452 51492 46462
rect 51436 46228 51492 46396
rect 51436 46114 51492 46172
rect 51436 46062 51438 46114
rect 51490 46062 51492 46114
rect 51436 46050 51492 46062
rect 50988 45892 51044 45902
rect 51212 45892 51268 45902
rect 50988 45798 51044 45836
rect 51100 45890 51268 45892
rect 51100 45838 51214 45890
rect 51266 45838 51268 45890
rect 51100 45836 51268 45838
rect 50652 44818 50708 44828
rect 50764 45500 50932 45556
rect 50764 44660 50820 45500
rect 51100 45444 51156 45836
rect 51212 45826 51268 45836
rect 50876 45388 51156 45444
rect 51324 45778 51380 45790
rect 51324 45726 51326 45778
rect 51378 45726 51380 45778
rect 51324 45444 51380 45726
rect 50876 45330 50932 45388
rect 51324 45378 51380 45388
rect 50876 45278 50878 45330
rect 50930 45278 50932 45330
rect 50876 45266 50932 45278
rect 50764 44594 50820 44604
rect 50876 44996 50932 45006
rect 51324 44996 51380 45006
rect 50652 44548 50708 44558
rect 50540 44546 50708 44548
rect 50540 44494 50654 44546
rect 50706 44494 50708 44546
rect 50540 44492 50708 44494
rect 50652 44482 50708 44492
rect 50204 41246 50206 41298
rect 50258 41246 50260 41298
rect 50204 41234 50260 41246
rect 50316 44436 50372 44446
rect 49980 41076 50036 41086
rect 49980 40982 50036 41020
rect 49756 40572 49924 40628
rect 49756 40068 49812 40572
rect 49868 40404 49924 40414
rect 49868 40292 49924 40348
rect 50092 40404 50148 40414
rect 49868 40236 50036 40292
rect 49756 40002 49812 40012
rect 49868 38722 49924 38734
rect 49868 38670 49870 38722
rect 49922 38670 49924 38722
rect 49532 38612 49700 38668
rect 49532 37044 49588 37054
rect 49532 36950 49588 36988
rect 49420 35970 49476 35980
rect 49532 36482 49588 36494
rect 49532 36430 49534 36482
rect 49586 36430 49588 36482
rect 49308 35644 49476 35700
rect 49196 35534 49198 35586
rect 49250 35534 49252 35586
rect 49196 35522 49252 35534
rect 49084 35410 49140 35420
rect 49420 33572 49476 35644
rect 49532 35364 49588 36430
rect 49532 35298 49588 35308
rect 49420 33506 49476 33516
rect 49532 34244 49588 34254
rect 48972 32510 48974 32562
rect 49026 32510 49028 32562
rect 48972 32498 49028 32510
rect 49308 32450 49364 32462
rect 49308 32398 49310 32450
rect 49362 32398 49364 32450
rect 49084 31778 49140 31790
rect 49084 31726 49086 31778
rect 49138 31726 49140 31778
rect 49084 31668 49140 31726
rect 49084 31602 49140 31612
rect 49308 31220 49364 32398
rect 49420 31890 49476 31902
rect 49420 31838 49422 31890
rect 49474 31838 49476 31890
rect 49420 31444 49476 31838
rect 49420 31378 49476 31388
rect 49308 31154 49364 31164
rect 49084 31108 49140 31118
rect 49532 31108 49588 34188
rect 49644 31668 49700 38612
rect 49756 37380 49812 37390
rect 49756 31948 49812 37324
rect 49868 35812 49924 38670
rect 49980 36932 50036 40236
rect 50092 38948 50148 40348
rect 50316 39732 50372 44380
rect 50428 44212 50484 44222
rect 50428 43314 50484 44156
rect 50876 44100 50932 44940
rect 51100 44994 51380 44996
rect 51100 44942 51326 44994
rect 51378 44942 51380 44994
rect 51100 44940 51380 44942
rect 50988 44884 51044 44894
rect 50988 44322 51044 44828
rect 50988 44270 50990 44322
rect 51042 44270 51044 44322
rect 50988 44258 51044 44270
rect 50876 44034 50932 44044
rect 51100 43876 51156 44940
rect 51324 44930 51380 44940
rect 51436 44882 51492 44894
rect 51436 44830 51438 44882
rect 51490 44830 51492 44882
rect 51212 44660 51268 44670
rect 51212 44100 51268 44604
rect 51436 44548 51492 44830
rect 51212 44034 51268 44044
rect 51324 44492 51492 44548
rect 50764 43820 51156 43876
rect 50764 43678 50820 43820
rect 51324 43708 51380 44492
rect 51548 44436 51604 47404
rect 51548 44370 51604 44380
rect 51660 46676 51716 46686
rect 51660 45892 51716 46620
rect 51436 44324 51492 44334
rect 51436 44230 51492 44268
rect 50652 43622 50820 43678
rect 50876 43652 50932 43662
rect 50428 43262 50430 43314
rect 50482 43262 50484 43314
rect 50428 43250 50484 43262
rect 50540 43538 50596 43550
rect 50540 43486 50542 43538
rect 50594 43486 50596 43538
rect 50540 43316 50596 43486
rect 50540 43250 50596 43260
rect 50652 43138 50708 43622
rect 50764 43540 50820 43550
rect 50764 43446 50820 43484
rect 50428 43082 50708 43138
rect 50764 43316 50820 43326
rect 50428 42194 50484 43082
rect 50764 42980 50820 43260
rect 50428 42142 50430 42194
rect 50482 42142 50484 42194
rect 50428 42130 50484 42142
rect 50652 42924 50820 42980
rect 50428 41186 50484 41198
rect 50428 41134 50430 41186
rect 50482 41134 50484 41186
rect 50428 41076 50484 41134
rect 50428 41010 50484 41020
rect 50428 40180 50484 40190
rect 50428 40086 50484 40124
rect 50316 39666 50372 39676
rect 50428 39394 50484 39406
rect 50428 39342 50430 39394
rect 50482 39342 50484 39394
rect 50092 38882 50148 38892
rect 50204 39172 50260 39182
rect 49980 36866 50036 36876
rect 50092 37940 50148 37950
rect 50092 36708 50148 37884
rect 50092 36642 50148 36652
rect 49868 35746 49924 35756
rect 50092 35476 50148 35486
rect 49980 35026 50036 35038
rect 49980 34974 49982 35026
rect 50034 34974 50036 35026
rect 49868 33908 49924 33918
rect 49868 33814 49924 33852
rect 49980 33684 50036 34974
rect 49980 33618 50036 33628
rect 49868 33572 49924 33582
rect 49868 32676 49924 33516
rect 49868 32610 49924 32620
rect 49980 33122 50036 33134
rect 49980 33070 49982 33122
rect 50034 33070 50036 33122
rect 49868 32452 49924 32462
rect 49980 32452 50036 33070
rect 50092 32786 50148 35420
rect 50204 33460 50260 39116
rect 50428 38836 50484 39342
rect 50428 38770 50484 38780
rect 50540 38834 50596 38846
rect 50540 38782 50542 38834
rect 50594 38782 50596 38834
rect 50428 38276 50484 38286
rect 50540 38276 50596 38782
rect 50428 38274 50596 38276
rect 50428 38222 50430 38274
rect 50482 38222 50596 38274
rect 50428 38220 50596 38222
rect 50428 38210 50484 38220
rect 50652 38164 50708 42924
rect 50876 41748 50932 43596
rect 50876 41682 50932 41692
rect 51100 43652 51380 43708
rect 51436 44100 51492 44110
rect 51100 43426 51156 43652
rect 51100 43374 51102 43426
rect 51154 43374 51156 43426
rect 50764 41412 50820 41422
rect 50764 39284 50820 41356
rect 50876 41188 50932 41198
rect 50876 40740 50932 41132
rect 51100 41188 51156 43374
rect 51212 43540 51268 43550
rect 51212 42082 51268 43484
rect 51324 43428 51380 43438
rect 51324 43334 51380 43372
rect 51436 42196 51492 44044
rect 51660 44100 51716 45836
rect 51772 44660 51828 48524
rect 51884 47460 51940 48750
rect 52108 48242 52164 49868
rect 52220 49812 52276 50652
rect 52332 49924 52388 50876
rect 52332 49858 52388 49868
rect 52220 49746 52276 49756
rect 52332 49588 52388 49598
rect 52332 49494 52388 49532
rect 52332 49140 52388 49150
rect 52108 48190 52110 48242
rect 52162 48190 52164 48242
rect 52108 48178 52164 48190
rect 52220 48804 52276 48814
rect 52220 47796 52276 48748
rect 52332 48468 52388 49084
rect 52332 48402 52388 48412
rect 52108 47740 52276 47796
rect 51996 47460 52052 47470
rect 51884 47458 52052 47460
rect 51884 47406 51998 47458
rect 52050 47406 52052 47458
rect 51884 47404 52052 47406
rect 51996 47394 52052 47404
rect 51884 47012 51940 47022
rect 51884 45892 51940 46956
rect 51884 45826 51940 45836
rect 51996 45780 52052 45790
rect 51996 45686 52052 45724
rect 51884 45668 51940 45678
rect 51884 45574 51940 45612
rect 52108 45108 52164 47740
rect 52220 47570 52276 47582
rect 52220 47518 52222 47570
rect 52274 47518 52276 47570
rect 52220 46004 52276 47518
rect 52444 47012 52500 53116
rect 52556 51604 52612 53452
rect 52668 53284 52724 53294
rect 52668 53170 52724 53228
rect 52668 53118 52670 53170
rect 52722 53118 52724 53170
rect 52668 53106 52724 53118
rect 52892 52948 52948 53790
rect 52668 52892 52948 52948
rect 53340 52948 53396 54238
rect 52668 52052 52724 52892
rect 53340 52882 53396 52892
rect 52780 52722 52836 52734
rect 52780 52670 52782 52722
rect 52834 52670 52836 52722
rect 52780 52164 52836 52670
rect 52892 52722 52948 52734
rect 53340 52724 53396 52734
rect 52892 52670 52894 52722
rect 52946 52670 52948 52722
rect 52892 52500 52948 52670
rect 52892 52434 52948 52444
rect 53004 52722 53396 52724
rect 53004 52670 53342 52722
rect 53394 52670 53396 52722
rect 53004 52668 53396 52670
rect 52780 52098 52836 52108
rect 52892 52164 52948 52174
rect 53004 52164 53060 52668
rect 53340 52658 53396 52668
rect 52892 52162 53060 52164
rect 52892 52110 52894 52162
rect 52946 52110 53060 52162
rect 52892 52108 53060 52110
rect 53116 52274 53172 52286
rect 53116 52222 53118 52274
rect 53170 52222 53172 52274
rect 52892 52098 52948 52108
rect 52668 51986 52724 51996
rect 53116 52052 53172 52222
rect 53116 51986 53172 51996
rect 52556 51538 52612 51548
rect 52780 51436 53172 51492
rect 52668 51380 52724 51390
rect 52444 46946 52500 46956
rect 52556 51378 52724 51380
rect 52556 51326 52670 51378
rect 52722 51326 52724 51378
rect 52556 51324 52724 51326
rect 52332 46674 52388 46686
rect 52332 46622 52334 46674
rect 52386 46622 52388 46674
rect 52332 46116 52388 46622
rect 52444 46676 52500 46686
rect 52444 46582 52500 46620
rect 52444 46116 52500 46126
rect 52332 46114 52500 46116
rect 52332 46062 52446 46114
rect 52498 46062 52500 46114
rect 52332 46060 52500 46062
rect 52444 46050 52500 46060
rect 52220 45948 52388 46004
rect 52332 45332 52388 45948
rect 52444 45332 52500 45342
rect 52332 45330 52500 45332
rect 52332 45278 52446 45330
rect 52498 45278 52500 45330
rect 52332 45276 52500 45278
rect 52444 45266 52500 45276
rect 51996 45052 52164 45108
rect 51772 44604 51940 44660
rect 51660 43204 51716 44044
rect 51772 44434 51828 44446
rect 51772 44382 51774 44434
rect 51826 44382 51828 44434
rect 51772 43764 51828 44382
rect 51772 43698 51828 43708
rect 51660 43138 51716 43148
rect 51436 42130 51492 42140
rect 51212 42030 51214 42082
rect 51266 42030 51268 42082
rect 51212 42018 51268 42030
rect 51884 41972 51940 44604
rect 51996 43652 52052 45052
rect 52108 44884 52164 44894
rect 52108 44790 52164 44828
rect 52332 44098 52388 44110
rect 52332 44046 52334 44098
rect 52386 44046 52388 44098
rect 52332 43764 52388 44046
rect 52332 43698 52388 43708
rect 52556 43678 52612 51324
rect 52668 51314 52724 51324
rect 52780 50820 52836 51436
rect 53116 51380 53172 51436
rect 53340 51380 53396 51390
rect 53116 51378 53396 51380
rect 53116 51326 53342 51378
rect 53394 51326 53396 51378
rect 53116 51324 53396 51326
rect 53340 51314 53396 51324
rect 53004 51266 53060 51278
rect 53004 51214 53006 51266
rect 53058 51214 53060 51266
rect 52892 51154 52948 51166
rect 52892 51102 52894 51154
rect 52946 51102 52948 51154
rect 52892 50878 52948 51102
rect 53004 51156 53060 51214
rect 53452 51268 53508 54460
rect 53564 53956 53620 55356
rect 53676 55346 53732 55356
rect 54012 55300 54068 55310
rect 54012 55206 54068 55244
rect 53676 54740 53732 54750
rect 54124 54740 54180 56028
rect 54572 56018 54628 56028
rect 55020 56082 55076 56476
rect 55020 56030 55022 56082
rect 55074 56030 55076 56082
rect 55020 56018 55076 56030
rect 54348 55860 54404 55870
rect 54348 55766 54404 55804
rect 55356 55858 55412 55870
rect 55356 55806 55358 55858
rect 55410 55806 55412 55858
rect 53732 54684 54180 54740
rect 54236 55748 54292 55758
rect 53676 54674 53732 54684
rect 54012 54402 54068 54414
rect 54012 54350 54014 54402
rect 54066 54350 54068 54402
rect 53564 53890 53620 53900
rect 53676 54290 53732 54302
rect 53676 54238 53678 54290
rect 53730 54238 53732 54290
rect 53564 53730 53620 53742
rect 53564 53678 53566 53730
rect 53618 53678 53620 53730
rect 53564 53508 53620 53678
rect 53564 53442 53620 53452
rect 53676 52948 53732 54238
rect 53900 54292 53956 54302
rect 54012 54292 54068 54350
rect 53956 54236 54068 54292
rect 53900 54226 53956 54236
rect 54236 54180 54292 55692
rect 54684 55412 54740 55422
rect 54684 55318 54740 55356
rect 54908 55300 54964 55310
rect 54796 55298 54964 55300
rect 54796 55246 54910 55298
rect 54962 55246 54964 55298
rect 54796 55244 54964 55246
rect 54348 54292 54404 54302
rect 54348 54198 54404 54236
rect 54012 54124 54292 54180
rect 53900 53732 53956 53742
rect 53900 53638 53956 53676
rect 54012 53284 54068 54124
rect 54796 54068 54852 55244
rect 54908 55234 54964 55244
rect 55356 54516 55412 55806
rect 55692 55860 55748 55870
rect 55692 55766 55748 55804
rect 55804 55524 55860 57344
rect 56252 56868 56308 57344
rect 56252 56802 56308 56812
rect 55804 55458 55860 55468
rect 56028 55858 56084 55870
rect 56028 55806 56030 55858
rect 56082 55806 56084 55858
rect 55244 54460 55412 54516
rect 55916 55410 55972 55422
rect 55916 55358 55918 55410
rect 55970 55358 55972 55410
rect 55020 54292 55076 54302
rect 53900 53228 54068 53284
rect 54124 54012 54852 54068
rect 54908 54290 55076 54292
rect 54908 54238 55022 54290
rect 55074 54238 55076 54290
rect 54908 54236 55076 54238
rect 53564 52892 53732 52948
rect 53788 53060 53844 53070
rect 53564 51604 53620 52892
rect 53788 52836 53844 53004
rect 53676 52780 53844 52836
rect 53676 52722 53732 52780
rect 53676 52670 53678 52722
rect 53730 52670 53732 52722
rect 53676 52658 53732 52670
rect 53676 52274 53732 52286
rect 53676 52222 53678 52274
rect 53730 52222 53732 52274
rect 53676 51716 53732 52222
rect 53676 51650 53732 51660
rect 53564 51538 53620 51548
rect 53452 51212 53620 51268
rect 53004 51090 53060 51100
rect 53452 51044 53508 51054
rect 52892 50822 53396 50878
rect 52668 50764 52836 50820
rect 52668 48244 52724 50764
rect 52892 50706 52948 50718
rect 52892 50654 52894 50706
rect 52946 50654 52948 50706
rect 52780 50484 52836 50522
rect 52780 50418 52836 50428
rect 52668 48178 52724 48188
rect 52668 48020 52724 48030
rect 52668 48018 52836 48020
rect 52668 47966 52670 48018
rect 52722 47966 52836 48018
rect 52668 47964 52836 47966
rect 52668 47954 52724 47964
rect 52668 47684 52724 47694
rect 52668 46562 52724 47628
rect 52668 46510 52670 46562
rect 52722 46510 52724 46562
rect 52668 46498 52724 46510
rect 52780 45444 52836 47964
rect 52892 47908 52948 50654
rect 53116 50372 53172 50382
rect 53116 50370 53284 50372
rect 53116 50318 53118 50370
rect 53170 50318 53284 50370
rect 53116 50316 53284 50318
rect 53116 50306 53172 50316
rect 53004 49924 53060 49934
rect 53004 49810 53060 49868
rect 53004 49758 53006 49810
rect 53058 49758 53060 49810
rect 53004 49746 53060 49758
rect 53116 49812 53172 49822
rect 53004 49140 53060 49150
rect 53116 49140 53172 49756
rect 53060 49084 53172 49140
rect 53004 49046 53060 49084
rect 52892 47852 53172 47908
rect 52892 47684 52948 47694
rect 52892 47458 52948 47628
rect 52892 47406 52894 47458
rect 52946 47406 52948 47458
rect 52892 47394 52948 47406
rect 52892 47012 52948 47022
rect 52892 46228 52948 46956
rect 53116 46676 53172 47852
rect 53116 46610 53172 46620
rect 53004 46562 53060 46574
rect 53004 46510 53006 46562
rect 53058 46510 53060 46562
rect 53004 46452 53060 46510
rect 53004 46386 53060 46396
rect 53116 46450 53172 46462
rect 53116 46398 53118 46450
rect 53170 46398 53172 46450
rect 52892 46172 53060 46228
rect 52780 45378 52836 45388
rect 52892 45106 52948 45118
rect 52892 45054 52894 45106
rect 52946 45054 52948 45106
rect 52892 44434 52948 45054
rect 52892 44382 52894 44434
rect 52946 44382 52948 44434
rect 52892 44212 52948 44382
rect 52892 44146 52948 44156
rect 52668 44100 52724 44110
rect 52668 44098 52836 44100
rect 52668 44046 52670 44098
rect 52722 44046 52836 44098
rect 52668 44044 52836 44046
rect 52668 44034 52724 44044
rect 52780 43764 52836 44044
rect 52780 43708 52948 43764
rect 52556 43622 52724 43678
rect 51996 43586 52052 43596
rect 52108 43540 52164 43550
rect 52108 43446 52164 43484
rect 52556 43538 52612 43550
rect 52556 43486 52558 43538
rect 52610 43486 52612 43538
rect 51996 43426 52052 43438
rect 51996 43374 51998 43426
rect 52050 43374 52052 43426
rect 51996 43204 52052 43374
rect 51996 43138 52052 43148
rect 52220 43428 52276 43438
rect 52108 42754 52164 42766
rect 52108 42702 52110 42754
rect 52162 42702 52164 42754
rect 51884 41916 52052 41972
rect 51436 41860 51492 41870
rect 51436 41858 51940 41860
rect 51436 41806 51438 41858
rect 51490 41806 51940 41858
rect 51436 41804 51940 41806
rect 51436 41794 51492 41804
rect 51212 41748 51268 41758
rect 51212 41654 51268 41692
rect 51324 41300 51380 41310
rect 51324 41206 51380 41244
rect 51100 41122 51156 41132
rect 51772 41188 51828 41198
rect 50988 40740 51044 40750
rect 50876 40684 50988 40740
rect 50988 40674 51044 40684
rect 51212 40516 51268 40526
rect 51212 40514 51492 40516
rect 51212 40462 51214 40514
rect 51266 40462 51492 40514
rect 51212 40460 51492 40462
rect 51212 40450 51268 40460
rect 51324 40290 51380 40302
rect 51324 40238 51326 40290
rect 51378 40238 51380 40290
rect 50764 39218 50820 39228
rect 50876 40178 50932 40190
rect 50876 40126 50878 40178
rect 50930 40126 50932 40178
rect 50876 39060 50932 40126
rect 51100 40178 51156 40190
rect 51100 40126 51102 40178
rect 51154 40126 51156 40178
rect 50988 39620 51044 39630
rect 50988 39526 51044 39564
rect 51100 39396 51156 40126
rect 51100 39330 51156 39340
rect 50876 38994 50932 39004
rect 51212 39172 51268 39182
rect 50764 38948 50820 38958
rect 50764 38854 50820 38892
rect 51212 38834 51268 39116
rect 51212 38782 51214 38834
rect 51266 38782 51268 38834
rect 51212 38770 51268 38782
rect 50988 38612 51044 38622
rect 50540 38108 50708 38164
rect 50876 38610 51044 38612
rect 50876 38558 50990 38610
rect 51042 38558 51044 38610
rect 50876 38556 51044 38558
rect 50428 35474 50484 35486
rect 50428 35422 50430 35474
rect 50482 35422 50484 35474
rect 50428 34804 50484 35422
rect 50316 34748 50484 34804
rect 50316 34354 50372 34748
rect 50540 34692 50596 38108
rect 50652 37492 50708 37502
rect 50876 37492 50932 38556
rect 50988 38546 51044 38556
rect 51100 38610 51156 38622
rect 51100 38558 51102 38610
rect 51154 38558 51156 38610
rect 51100 38052 51156 38558
rect 51324 38500 51380 40238
rect 51324 38434 51380 38444
rect 51436 38164 51492 40460
rect 51548 39730 51604 39742
rect 51548 39678 51550 39730
rect 51602 39678 51604 39730
rect 51548 38388 51604 39678
rect 51772 38836 51828 41132
rect 51884 39060 51940 41804
rect 51996 40516 52052 41916
rect 51996 40450 52052 40460
rect 51884 38994 51940 39004
rect 51996 40180 52052 40190
rect 51996 39058 52052 40124
rect 51996 39006 51998 39058
rect 52050 39006 52052 39058
rect 51996 38994 52052 39006
rect 51772 38780 51940 38836
rect 51548 38322 51604 38332
rect 51436 38108 51604 38164
rect 51100 37986 51156 37996
rect 51436 37938 51492 37950
rect 51436 37886 51438 37938
rect 51490 37886 51492 37938
rect 50652 37490 50932 37492
rect 50652 37438 50654 37490
rect 50706 37438 50932 37490
rect 50652 37436 50932 37438
rect 51100 37828 51156 37838
rect 50652 37426 50708 37436
rect 51100 37266 51156 37772
rect 51436 37716 51492 37886
rect 51436 37650 51492 37660
rect 51100 37214 51102 37266
rect 51154 37214 51156 37266
rect 51100 37202 51156 37214
rect 51436 37042 51492 37054
rect 51436 36990 51438 37042
rect 51490 36990 51492 37042
rect 51324 36484 51380 36494
rect 50876 35586 50932 35598
rect 50876 35534 50878 35586
rect 50930 35534 50932 35586
rect 50876 35252 50932 35534
rect 51212 35586 51268 35598
rect 51212 35534 51214 35586
rect 51266 35534 51268 35586
rect 50988 35476 51044 35486
rect 50988 35382 51044 35420
rect 50876 35186 50932 35196
rect 51212 35140 51268 35534
rect 51212 35074 51268 35084
rect 51324 35026 51380 36428
rect 51436 36148 51492 36990
rect 51436 36082 51492 36092
rect 51548 35924 51604 38108
rect 51772 38162 51828 38174
rect 51772 38110 51774 38162
rect 51826 38110 51828 38162
rect 51548 35858 51604 35868
rect 51660 38052 51716 38062
rect 51324 34974 51326 35026
rect 51378 34974 51380 35026
rect 51324 34962 51380 34974
rect 51436 35586 51492 35598
rect 51436 35534 51438 35586
rect 51490 35534 51492 35586
rect 50316 34302 50318 34354
rect 50370 34302 50372 34354
rect 50316 34290 50372 34302
rect 50428 34636 50596 34692
rect 50876 34916 50932 34926
rect 50428 33460 50484 34636
rect 50764 34580 50820 34590
rect 50764 34356 50820 34524
rect 50540 34300 50820 34356
rect 50540 34130 50596 34300
rect 50876 34242 50932 34860
rect 50876 34190 50878 34242
rect 50930 34190 50932 34242
rect 50876 34178 50932 34190
rect 50540 34078 50542 34130
rect 50594 34078 50596 34130
rect 50540 34066 50596 34078
rect 50764 34020 50820 34030
rect 50764 33926 50820 33964
rect 50988 34020 51044 34058
rect 50988 33954 51044 33964
rect 51100 33796 51156 33806
rect 50540 33684 50596 33694
rect 50540 33572 50596 33628
rect 50540 33506 50596 33516
rect 50876 33628 50932 33638
rect 50204 33394 50260 33404
rect 50316 33404 50484 33460
rect 50652 33460 50708 33470
rect 50092 32734 50094 32786
rect 50146 32734 50148 32786
rect 50092 32722 50148 32734
rect 49868 32450 50036 32452
rect 49868 32398 49870 32450
rect 49922 32398 50036 32450
rect 49868 32396 50036 32398
rect 49868 32386 49924 32396
rect 50092 32228 50148 32238
rect 49756 31892 50036 31948
rect 49644 31602 49700 31612
rect 49756 31778 49812 31790
rect 49756 31726 49758 31778
rect 49810 31726 49812 31778
rect 49084 30772 49140 31052
rect 49420 31052 49588 31108
rect 49196 30996 49252 31006
rect 49420 30996 49476 31052
rect 49196 30994 49476 30996
rect 49196 30942 49198 30994
rect 49250 30942 49476 30994
rect 49196 30940 49476 30942
rect 49196 30930 49252 30940
rect 49084 30716 49476 30772
rect 48972 30324 49028 30334
rect 48972 30230 49028 30268
rect 49084 29986 49140 29998
rect 49084 29934 49086 29986
rect 49138 29934 49140 29986
rect 49084 29764 49140 29934
rect 49084 29698 49140 29708
rect 49084 29204 49140 29214
rect 49140 29148 49252 29204
rect 49084 29110 49140 29148
rect 48972 28642 49028 28654
rect 48972 28590 48974 28642
rect 49026 28590 49028 28642
rect 48972 24946 49028 28590
rect 48972 24894 48974 24946
rect 49026 24894 49028 24946
rect 48972 24882 49028 24894
rect 49084 27412 49140 27422
rect 48748 24220 48916 24276
rect 48748 23268 48804 24220
rect 48860 24052 48916 24062
rect 48860 23958 48916 23996
rect 48748 23202 48804 23212
rect 48972 23156 49028 23166
rect 48748 23044 48804 23054
rect 48748 22950 48804 22988
rect 48860 21812 48916 21822
rect 48748 21476 48804 21486
rect 48748 21382 48804 21420
rect 48748 21028 48804 21038
rect 48412 20972 48580 21028
rect 48412 20020 48468 20030
rect 48412 19458 48468 19964
rect 48412 19406 48414 19458
rect 48466 19406 48468 19458
rect 48412 19394 48468 19406
rect 48300 18610 48356 18620
rect 48188 17614 48190 17666
rect 48242 17614 48244 17666
rect 48188 17602 48244 17614
rect 48076 17556 48132 17566
rect 48076 14756 48132 17500
rect 48300 17556 48356 17566
rect 48188 17332 48244 17342
rect 48188 16994 48244 17276
rect 48188 16942 48190 16994
rect 48242 16942 48244 16994
rect 48188 16930 48244 16942
rect 48300 16772 48356 17500
rect 48300 16706 48356 16716
rect 48188 16098 48244 16110
rect 48188 16046 48190 16098
rect 48242 16046 48244 16098
rect 48188 15316 48244 16046
rect 48300 15540 48356 15550
rect 48300 15446 48356 15484
rect 48188 15250 48244 15260
rect 48076 14690 48132 14700
rect 48524 14756 48580 20972
rect 48636 20692 48692 20702
rect 48636 20598 48692 20636
rect 48748 20018 48804 20972
rect 48860 20802 48916 21756
rect 48860 20750 48862 20802
rect 48914 20750 48916 20802
rect 48860 20738 48916 20750
rect 48748 19966 48750 20018
rect 48802 19966 48804 20018
rect 48748 19954 48804 19966
rect 48972 19906 49028 23100
rect 49084 23044 49140 27356
rect 49196 26402 49252 29148
rect 49308 28980 49364 28990
rect 49308 28754 49364 28924
rect 49308 28702 49310 28754
rect 49362 28702 49364 28754
rect 49308 28690 49364 28702
rect 49420 27412 49476 30716
rect 49532 30212 49588 31052
rect 49756 31332 49812 31726
rect 49644 30770 49700 30782
rect 49644 30718 49646 30770
rect 49698 30718 49700 30770
rect 49644 30660 49700 30718
rect 49644 30594 49700 30604
rect 49532 30146 49588 30156
rect 49532 29988 49588 29998
rect 49532 29428 49588 29932
rect 49756 29876 49812 31276
rect 49868 31220 49924 31230
rect 49868 30660 49924 31164
rect 49868 30594 49924 30604
rect 49532 29334 49588 29372
rect 49644 29820 49812 29876
rect 49644 29204 49700 29820
rect 49868 29316 49924 29326
rect 49420 27346 49476 27356
rect 49532 29148 49700 29204
rect 49756 29204 49812 29214
rect 49420 27186 49476 27198
rect 49420 27134 49422 27186
rect 49474 27134 49476 27186
rect 49420 27076 49476 27134
rect 49420 27010 49476 27020
rect 49532 26908 49588 29148
rect 49756 29110 49812 29148
rect 49420 26852 49588 26908
rect 49644 28980 49700 28990
rect 49196 26350 49198 26402
rect 49250 26350 49252 26402
rect 49196 26338 49252 26350
rect 49308 26516 49364 26526
rect 49308 25956 49364 26460
rect 49420 26402 49476 26852
rect 49420 26350 49422 26402
rect 49474 26350 49476 26402
rect 49420 26292 49476 26350
rect 49420 26236 49588 26292
rect 49532 25956 49588 26236
rect 49084 22978 49140 22988
rect 49196 25900 49364 25956
rect 49420 25900 49588 25956
rect 49084 22372 49140 22382
rect 49196 22372 49252 25900
rect 49308 25732 49364 25742
rect 49308 25638 49364 25676
rect 49308 22596 49364 22606
rect 49308 22502 49364 22540
rect 49196 22316 49364 22372
rect 49084 21868 49140 22316
rect 49084 21812 49252 21868
rect 49196 21588 49252 21812
rect 48972 19854 48974 19906
rect 49026 19854 49028 19906
rect 48972 19842 49028 19854
rect 49084 21586 49252 21588
rect 49084 21534 49198 21586
rect 49250 21534 49252 21586
rect 49084 21532 49252 21534
rect 48860 19572 48916 19582
rect 48748 18338 48804 18350
rect 48748 18286 48750 18338
rect 48802 18286 48804 18338
rect 48748 17892 48804 18286
rect 48860 18116 48916 19516
rect 48972 19236 49028 19246
rect 48972 19142 49028 19180
rect 49084 18564 49140 21532
rect 49196 21522 49252 21532
rect 49196 21252 49252 21262
rect 49196 21026 49252 21196
rect 49196 20974 49198 21026
rect 49250 20974 49252 21026
rect 49196 20962 49252 20974
rect 49196 19460 49252 19470
rect 49196 19366 49252 19404
rect 49084 18470 49140 18508
rect 49308 18452 49364 22316
rect 49420 20580 49476 25900
rect 49644 25508 49700 28924
rect 49756 28644 49812 28654
rect 49756 28550 49812 28588
rect 49868 28420 49924 29260
rect 49756 28364 49924 28420
rect 49756 26908 49812 28364
rect 49868 27300 49924 27310
rect 49868 27074 49924 27244
rect 49868 27022 49870 27074
rect 49922 27022 49924 27074
rect 49868 27010 49924 27022
rect 49756 26852 49924 26908
rect 49756 26516 49812 26526
rect 49868 26516 49924 26852
rect 49756 26514 49924 26516
rect 49756 26462 49758 26514
rect 49810 26462 49924 26514
rect 49756 26460 49924 26462
rect 49756 26450 49812 26460
rect 49868 25732 49924 25742
rect 49756 25508 49812 25518
rect 49644 25452 49756 25508
rect 49756 25394 49812 25452
rect 49756 25342 49758 25394
rect 49810 25342 49812 25394
rect 49756 24836 49812 25342
rect 49756 24770 49812 24780
rect 49532 24498 49588 24510
rect 49532 24446 49534 24498
rect 49586 24446 49588 24498
rect 49532 20804 49588 24446
rect 49868 24052 49924 25676
rect 49756 23996 49924 24052
rect 49644 23268 49700 23278
rect 49644 23174 49700 23212
rect 49756 22484 49812 23996
rect 49868 23828 49924 23838
rect 49868 22596 49924 23772
rect 49980 22932 50036 31892
rect 50092 31778 50148 32172
rect 50204 32004 50260 32014
rect 50316 32004 50372 33404
rect 50652 33346 50708 33404
rect 50652 33294 50654 33346
rect 50706 33294 50708 33346
rect 50652 33282 50708 33294
rect 50428 33234 50484 33246
rect 50428 33182 50430 33234
rect 50482 33182 50484 33234
rect 50428 33124 50484 33182
rect 50876 33236 50932 33572
rect 50876 33170 50932 33180
rect 50428 33068 50820 33124
rect 50428 32564 50484 32574
rect 50764 32564 50820 33068
rect 50988 33122 51044 33134
rect 50988 33070 50990 33122
rect 51042 33070 51044 33122
rect 50988 33012 51044 33070
rect 50988 32946 51044 32956
rect 51100 32788 51156 33740
rect 51436 33572 51492 35534
rect 51660 34692 51716 37996
rect 51772 37380 51828 38110
rect 51772 37314 51828 37324
rect 51660 34626 51716 34636
rect 51772 36148 51828 36158
rect 51772 34356 51828 36092
rect 51772 34290 51828 34300
rect 51884 34132 51940 38780
rect 52108 36484 52164 42702
rect 52220 41076 52276 43372
rect 52332 43426 52388 43438
rect 52332 43374 52334 43426
rect 52386 43374 52388 43426
rect 52332 42084 52388 43374
rect 52556 43316 52612 43486
rect 52556 43250 52612 43260
rect 52444 43092 52500 43102
rect 52444 42196 52500 43036
rect 52444 42130 52500 42140
rect 52556 42308 52612 42318
rect 52332 42018 52388 42028
rect 52444 41972 52500 41982
rect 52556 41972 52612 42252
rect 52668 42196 52724 43622
rect 52780 43538 52836 43550
rect 52780 43486 52782 43538
rect 52834 43486 52836 43538
rect 52780 43428 52836 43486
rect 52780 43092 52836 43372
rect 52780 43026 52836 43036
rect 52668 42130 52724 42140
rect 52892 41972 52948 43708
rect 52444 41970 52612 41972
rect 52444 41918 52446 41970
rect 52498 41918 52612 41970
rect 52444 41916 52612 41918
rect 52780 41916 52948 41972
rect 52332 41748 52388 41758
rect 52332 41188 52388 41692
rect 52332 41122 52388 41132
rect 52220 41010 52276 41020
rect 52220 40740 52276 40750
rect 52220 40514 52276 40684
rect 52444 40740 52500 41916
rect 52780 41636 52836 41916
rect 52892 41748 52948 41758
rect 52892 41654 52948 41692
rect 52780 41570 52836 41580
rect 52892 41524 52948 41534
rect 52892 41412 52948 41468
rect 52780 41356 52948 41412
rect 52556 41076 52612 41086
rect 52556 40982 52612 41020
rect 52444 40674 52500 40684
rect 52780 40516 52836 41356
rect 52220 40462 52222 40514
rect 52274 40462 52276 40514
rect 52220 40450 52276 40462
rect 52444 40460 52836 40516
rect 52892 41188 52948 41198
rect 52444 39284 52500 40460
rect 52668 40178 52724 40190
rect 52668 40126 52670 40178
rect 52722 40126 52724 40178
rect 52668 39844 52724 40126
rect 52668 39778 52724 39788
rect 52444 39218 52500 39228
rect 52556 39732 52612 39742
rect 52556 39172 52612 39676
rect 52668 39396 52724 39406
rect 52668 39302 52724 39340
rect 52220 38948 52276 38958
rect 52220 38854 52276 38892
rect 52444 38836 52500 38874
rect 52556 38836 52612 39116
rect 52780 39172 52836 39182
rect 52668 38836 52724 38846
rect 52556 38834 52724 38836
rect 52556 38782 52670 38834
rect 52722 38782 52724 38834
rect 52556 38780 52724 38782
rect 52444 38770 52500 38780
rect 52556 38610 52612 38622
rect 52556 38558 52558 38610
rect 52610 38558 52612 38610
rect 52444 38052 52500 38062
rect 52444 37716 52500 37996
rect 52444 37378 52500 37660
rect 52444 37326 52446 37378
rect 52498 37326 52500 37378
rect 52444 37314 52500 37326
rect 52556 36932 52612 38558
rect 52556 36866 52612 36876
rect 52108 36418 52164 36428
rect 52444 36820 52500 36830
rect 52220 36370 52276 36382
rect 52220 36318 52222 36370
rect 52274 36318 52276 36370
rect 51996 35924 52052 35934
rect 51996 35476 52052 35868
rect 52108 35700 52164 35710
rect 52108 35606 52164 35644
rect 51996 35410 52052 35420
rect 52220 34914 52276 36318
rect 52332 35700 52388 35710
rect 52332 35606 52388 35644
rect 52220 34862 52222 34914
rect 52274 34862 52276 34914
rect 52220 34850 52276 34862
rect 52444 34692 52500 36764
rect 52668 36708 52724 38780
rect 52668 36642 52724 36652
rect 52780 36484 52836 39116
rect 52892 38612 52948 41132
rect 53004 38668 53060 46172
rect 53116 46004 53172 46398
rect 53228 46004 53284 50316
rect 53340 46900 53396 50822
rect 53452 50818 53508 50988
rect 53452 50766 53454 50818
rect 53506 50766 53508 50818
rect 53452 50754 53508 50766
rect 53564 50708 53620 51212
rect 53676 51156 53732 51166
rect 53676 51154 53844 51156
rect 53676 51102 53678 51154
rect 53730 51102 53844 51154
rect 53676 51100 53844 51102
rect 53676 51090 53732 51100
rect 53564 50642 53620 50652
rect 53676 50594 53732 50606
rect 53676 50542 53678 50594
rect 53730 50542 53732 50594
rect 53676 50372 53732 50542
rect 53676 50306 53732 50316
rect 53452 49924 53508 49934
rect 53452 49026 53508 49868
rect 53564 49588 53620 49598
rect 53564 49494 53620 49532
rect 53452 48974 53454 49026
rect 53506 48974 53508 49026
rect 53452 48962 53508 48974
rect 53788 48244 53844 51100
rect 53900 50148 53956 53228
rect 54012 52164 54068 52174
rect 54012 52070 54068 52108
rect 54124 51492 54180 54012
rect 54236 53842 54292 53854
rect 54236 53790 54238 53842
rect 54290 53790 54292 53842
rect 54236 53060 54292 53790
rect 54236 52994 54292 53004
rect 54684 53732 54740 53742
rect 54684 52946 54740 53676
rect 54684 52894 54686 52946
rect 54738 52894 54740 52946
rect 54684 52882 54740 52894
rect 54572 52836 54628 52846
rect 54348 52722 54404 52734
rect 54348 52670 54350 52722
rect 54402 52670 54404 52722
rect 54348 52500 54404 52670
rect 54348 52434 54404 52444
rect 54124 51426 54180 51436
rect 54236 52388 54292 52398
rect 54236 51380 54292 52332
rect 54348 52274 54404 52286
rect 54348 52222 54350 52274
rect 54402 52222 54404 52274
rect 54348 51940 54404 52222
rect 54348 51874 54404 51884
rect 54572 51492 54628 52780
rect 54908 52388 54964 54236
rect 55020 54226 55076 54236
rect 55132 54180 55188 54190
rect 55132 53956 55188 54124
rect 55132 53890 55188 53900
rect 55020 53730 55076 53742
rect 55020 53678 55022 53730
rect 55074 53678 55076 53730
rect 55020 52948 55076 53678
rect 55244 53284 55300 54460
rect 55916 54404 55972 55358
rect 56028 54516 56084 55806
rect 56252 55858 56308 55870
rect 56252 55806 56254 55858
rect 56306 55806 56308 55858
rect 56252 55636 56308 55806
rect 56252 55570 56308 55580
rect 56028 54450 56084 54460
rect 56252 55298 56308 55310
rect 56252 55246 56254 55298
rect 56306 55246 56308 55298
rect 55916 54338 55972 54348
rect 55356 54290 55412 54302
rect 55356 54238 55358 54290
rect 55410 54238 55412 54290
rect 55356 54180 55412 54238
rect 56028 54292 56084 54302
rect 56028 54198 56084 54236
rect 55356 54114 55412 54124
rect 55244 53218 55300 53228
rect 55356 53842 55412 53854
rect 55356 53790 55358 53842
rect 55410 53790 55412 53842
rect 55020 52882 55076 52892
rect 55356 52948 55412 53790
rect 56028 53732 56084 53742
rect 55356 52882 55412 52892
rect 55804 53730 56084 53732
rect 55804 53678 56030 53730
rect 56082 53678 56084 53730
rect 55804 53676 56084 53678
rect 55020 52724 55076 52734
rect 55356 52724 55412 52734
rect 55020 52722 55300 52724
rect 55020 52670 55022 52722
rect 55074 52670 55300 52722
rect 55020 52668 55300 52670
rect 55020 52658 55076 52668
rect 54908 52332 55076 52388
rect 54684 52162 54740 52174
rect 54684 52110 54686 52162
rect 54738 52110 54740 52162
rect 54684 51716 54740 52110
rect 54684 51650 54740 51660
rect 54796 52052 54852 52062
rect 54572 51426 54628 51436
rect 54236 51324 54404 51380
rect 54124 51268 54180 51278
rect 54124 51044 54180 51212
rect 54236 51156 54292 51166
rect 54236 51062 54292 51100
rect 54124 50978 54180 50988
rect 54236 50484 54292 50522
rect 54236 50418 54292 50428
rect 54348 50260 54404 51324
rect 54572 51268 54628 51306
rect 54572 51202 54628 51212
rect 54460 51044 54516 51054
rect 54460 50818 54516 50988
rect 54460 50766 54462 50818
rect 54514 50766 54516 50818
rect 54460 50754 54516 50766
rect 54684 50820 54740 50830
rect 54572 50484 54628 50494
rect 54684 50484 54740 50764
rect 54572 50482 54740 50484
rect 54572 50430 54574 50482
rect 54626 50430 54740 50482
rect 54572 50428 54740 50430
rect 54572 50418 54628 50428
rect 54348 50194 54404 50204
rect 53900 50082 53956 50092
rect 54684 49586 54740 49598
rect 54684 49534 54686 49586
rect 54738 49534 54740 49586
rect 54348 49140 54404 49150
rect 54124 49138 54404 49140
rect 54124 49086 54350 49138
rect 54402 49086 54404 49138
rect 54124 49084 54404 49086
rect 53788 48178 53844 48188
rect 54012 49026 54068 49038
rect 54012 48974 54014 49026
rect 54066 48974 54068 49026
rect 53900 48132 53956 48142
rect 53788 48020 53844 48030
rect 53452 48018 53844 48020
rect 53452 47966 53790 48018
rect 53842 47966 53844 48018
rect 53452 47964 53844 47966
rect 53452 47458 53508 47964
rect 53788 47954 53844 47964
rect 53452 47406 53454 47458
rect 53506 47406 53508 47458
rect 53452 47394 53508 47406
rect 53788 47796 53844 47806
rect 53788 47348 53844 47740
rect 53788 47282 53844 47292
rect 53340 46844 53508 46900
rect 53340 46676 53396 46686
rect 53340 46582 53396 46620
rect 53228 45948 53396 46004
rect 53116 45938 53172 45948
rect 53228 45780 53284 45790
rect 53116 45668 53172 45678
rect 53116 40292 53172 45612
rect 53228 44994 53284 45724
rect 53228 44942 53230 44994
rect 53282 44942 53284 44994
rect 53228 44930 53284 44942
rect 53228 43314 53284 43326
rect 53228 43262 53230 43314
rect 53282 43262 53284 43314
rect 53228 42532 53284 43262
rect 53228 42466 53284 42476
rect 53228 41074 53284 41086
rect 53228 41022 53230 41074
rect 53282 41022 53284 41074
rect 53228 40516 53284 41022
rect 53228 40450 53284 40460
rect 53116 40226 53172 40236
rect 53340 39732 53396 45948
rect 53452 45780 53508 46844
rect 53788 46676 53844 46686
rect 53788 46582 53844 46620
rect 53676 46452 53732 46462
rect 53564 46228 53620 46238
rect 53564 46114 53620 46172
rect 53564 46062 53566 46114
rect 53618 46062 53620 46114
rect 53564 46050 53620 46062
rect 53452 45724 53620 45780
rect 53452 44434 53508 44446
rect 53452 44382 53454 44434
rect 53506 44382 53508 44434
rect 53452 42644 53508 44382
rect 53564 43652 53620 45724
rect 53676 43764 53732 46396
rect 53788 46228 53844 46238
rect 53788 45668 53844 46172
rect 53788 45602 53844 45612
rect 53788 45332 53844 45342
rect 53900 45332 53956 48076
rect 54012 46004 54068 48974
rect 54124 46116 54180 49084
rect 54348 49074 54404 49084
rect 54684 48916 54740 49534
rect 54460 48860 54740 48916
rect 54236 48132 54292 48142
rect 54236 48038 54292 48076
rect 54348 48018 54404 48030
rect 54348 47966 54350 48018
rect 54402 47966 54404 48018
rect 54348 47684 54404 47966
rect 54236 47628 54404 47684
rect 54236 46676 54292 47628
rect 54348 47460 54404 47470
rect 54460 47460 54516 48860
rect 54796 48804 54852 51996
rect 54908 51380 54964 51390
rect 54908 51266 54964 51324
rect 54908 51214 54910 51266
rect 54962 51214 54964 51266
rect 54908 51202 54964 51214
rect 54908 50932 54964 50942
rect 54908 49476 54964 50876
rect 55020 50820 55076 52332
rect 55132 52162 55188 52174
rect 55132 52110 55134 52162
rect 55186 52110 55188 52162
rect 55132 50820 55188 52110
rect 55244 51492 55300 52668
rect 55356 52722 55748 52724
rect 55356 52670 55358 52722
rect 55410 52670 55748 52722
rect 55356 52668 55748 52670
rect 55356 52658 55412 52668
rect 55356 52274 55412 52286
rect 55356 52222 55358 52274
rect 55410 52222 55412 52274
rect 55356 51716 55412 52222
rect 55356 51650 55412 51660
rect 55244 51436 55412 51492
rect 55244 51154 55300 51166
rect 55244 51102 55246 51154
rect 55298 51102 55300 51154
rect 55244 51044 55300 51102
rect 55356 51044 55412 51436
rect 55580 51154 55636 51166
rect 55580 51102 55582 51154
rect 55634 51102 55636 51154
rect 55356 50988 55524 51044
rect 55244 50978 55300 50988
rect 55356 50820 55412 50830
rect 55132 50818 55412 50820
rect 55132 50766 55358 50818
rect 55410 50766 55412 50818
rect 55132 50764 55412 50766
rect 55020 50754 55076 50764
rect 55356 50754 55412 50764
rect 55020 50596 55076 50606
rect 55468 50596 55524 50988
rect 55020 50502 55076 50540
rect 55132 50540 55524 50596
rect 54908 49410 54964 49420
rect 54684 48748 54852 48804
rect 55020 49026 55076 49038
rect 55020 48974 55022 49026
rect 55074 48974 55076 49026
rect 55020 48804 55076 48974
rect 54684 48580 54740 48748
rect 55020 48738 55076 48748
rect 54348 47458 54516 47460
rect 54348 47406 54350 47458
rect 54402 47406 54516 47458
rect 54348 47404 54516 47406
rect 54572 48524 54740 48580
rect 54348 47394 54404 47404
rect 54236 46610 54292 46620
rect 54572 46228 54628 48524
rect 54460 46172 54628 46228
rect 54684 48356 54740 48366
rect 54124 46060 54292 46116
rect 54012 45948 54180 46004
rect 53788 45330 53956 45332
rect 53788 45278 53790 45330
rect 53842 45278 53956 45330
rect 53788 45276 53956 45278
rect 54012 45778 54068 45790
rect 54012 45726 54014 45778
rect 54066 45726 54068 45778
rect 54012 45668 54068 45726
rect 53788 45266 53844 45276
rect 54012 44772 54068 45612
rect 54124 45332 54180 45948
rect 54236 45444 54292 46060
rect 54460 45556 54516 46172
rect 54684 46004 54740 48300
rect 54796 48244 54852 48254
rect 54796 48242 54964 48244
rect 54796 48190 54798 48242
rect 54850 48190 54964 48242
rect 54796 48188 54964 48190
rect 54796 48178 54852 48188
rect 54796 47460 54852 47470
rect 54796 47366 54852 47404
rect 54236 45378 54292 45388
rect 54348 45500 54516 45556
rect 54572 45948 54740 46004
rect 54796 46676 54852 46686
rect 54908 46676 54964 48188
rect 55020 48132 55076 48142
rect 55020 48038 55076 48076
rect 55132 47908 55188 50540
rect 55580 49812 55636 51102
rect 55692 50148 55748 52668
rect 55692 50082 55748 50092
rect 55580 49756 55748 49812
rect 55020 47852 55188 47908
rect 55244 49586 55300 49598
rect 55580 49588 55636 49598
rect 55244 49534 55246 49586
rect 55298 49534 55300 49586
rect 55020 47012 55076 47852
rect 55132 47684 55188 47694
rect 55244 47684 55300 49534
rect 55468 49586 55636 49588
rect 55468 49534 55582 49586
rect 55634 49534 55636 49586
rect 55468 49532 55636 49534
rect 55356 49252 55412 49262
rect 55356 49158 55412 49196
rect 55132 47682 55300 47684
rect 55132 47630 55134 47682
rect 55186 47630 55300 47682
rect 55132 47628 55300 47630
rect 55356 48018 55412 48030
rect 55356 47966 55358 48018
rect 55410 47966 55412 48018
rect 55132 47618 55188 47628
rect 55356 47068 55412 47966
rect 55020 46946 55076 46956
rect 55244 47012 55412 47068
rect 55244 46676 55300 47012
rect 54908 46620 55076 46676
rect 54572 45890 54628 45948
rect 54572 45838 54574 45890
rect 54626 45838 54628 45890
rect 54124 45266 54180 45276
rect 54012 44706 54068 44716
rect 54348 44548 54404 45500
rect 54572 44548 54628 45838
rect 54796 45890 54852 46620
rect 54908 46452 54964 46462
rect 54908 46358 54964 46396
rect 55020 46228 55076 46620
rect 55244 46610 55300 46620
rect 55356 46674 55412 46686
rect 55356 46622 55358 46674
rect 55410 46622 55412 46674
rect 54796 45838 54798 45890
rect 54850 45838 54852 45890
rect 54796 45826 54852 45838
rect 54908 46172 55076 46228
rect 55244 46452 55300 46462
rect 54684 45780 54740 45790
rect 54684 45686 54740 45724
rect 54796 45332 54852 45342
rect 54796 44578 54852 45276
rect 54908 45108 54964 46172
rect 55132 45890 55188 45902
rect 55132 45838 55134 45890
rect 55186 45838 55188 45890
rect 55132 45780 55188 45838
rect 55132 45714 55188 45724
rect 54908 45052 55188 45108
rect 54908 44884 54964 44894
rect 54908 44790 54964 44828
rect 54348 44492 54516 44548
rect 54572 44492 54740 44548
rect 54796 44522 54964 44578
rect 54460 44436 54516 44492
rect 53676 43698 53732 43708
rect 53788 44342 54292 44398
rect 54460 44370 54516 44380
rect 53564 43586 53620 43596
rect 53564 43316 53620 43326
rect 53564 43222 53620 43260
rect 53676 42868 53732 42878
rect 53676 42774 53732 42812
rect 53452 42578 53508 42588
rect 53452 42196 53508 42206
rect 53452 41076 53508 42140
rect 53788 42196 53844 44342
rect 54236 44324 54292 44342
rect 54348 44324 54404 44334
rect 54236 44322 54404 44324
rect 54236 44270 54350 44322
rect 54402 44270 54404 44322
rect 54236 44268 54404 44270
rect 54348 44258 54404 44268
rect 54572 44322 54628 44334
rect 54572 44270 54574 44322
rect 54626 44270 54628 44322
rect 54124 44212 54180 44222
rect 54012 44210 54180 44212
rect 54012 44158 54126 44210
rect 54178 44158 54180 44210
rect 54012 44156 54180 44158
rect 53900 44098 53956 44110
rect 53900 44046 53902 44098
rect 53954 44046 53956 44098
rect 53900 43876 53956 44046
rect 54012 44100 54068 44156
rect 54124 44146 54180 44156
rect 54460 44210 54516 44222
rect 54460 44158 54462 44210
rect 54514 44158 54516 44210
rect 54012 44034 54068 44044
rect 54460 43988 54516 44158
rect 54124 43932 54516 43988
rect 53900 43820 54068 43876
rect 53900 43652 53956 43662
rect 53900 42866 53956 43596
rect 53900 42814 53902 42866
rect 53954 42814 53956 42866
rect 53900 42802 53956 42814
rect 53788 42130 53844 42140
rect 54012 42194 54068 43820
rect 54124 43678 54180 43932
rect 54572 43764 54628 44270
rect 54684 43764 54740 44492
rect 54796 43764 54852 43774
rect 54684 43708 54796 43764
rect 54572 43698 54628 43708
rect 54796 43698 54852 43708
rect 54124 43622 54292 43678
rect 54124 43540 54180 43550
rect 54124 43446 54180 43484
rect 54124 42756 54180 42766
rect 54236 42756 54292 43622
rect 54460 43652 54516 43662
rect 54460 43428 54516 43596
rect 54572 43428 54628 43438
rect 54460 43426 54628 43428
rect 54460 43374 54574 43426
rect 54626 43374 54628 43426
rect 54460 43372 54628 43374
rect 54572 43362 54628 43372
rect 54124 42754 54292 42756
rect 54124 42702 54126 42754
rect 54178 42702 54292 42754
rect 54124 42700 54292 42702
rect 54348 43092 54404 43102
rect 54348 42754 54404 43036
rect 54908 42958 54964 44522
rect 54348 42702 54350 42754
rect 54402 42702 54404 42754
rect 54796 42902 54964 42958
rect 55020 44322 55076 44334
rect 55020 44270 55022 44322
rect 55074 44270 55076 44322
rect 54124 42690 54180 42700
rect 54348 42690 54404 42702
rect 54572 42698 54628 42710
rect 54460 42644 54516 42654
rect 54460 42550 54516 42588
rect 54572 42646 54574 42698
rect 54626 42646 54628 42698
rect 54572 42532 54628 42646
rect 54572 42466 54628 42476
rect 54012 42142 54014 42194
rect 54066 42142 54068 42194
rect 54012 42130 54068 42142
rect 54572 42196 54628 42206
rect 54572 42102 54628 42140
rect 53564 41300 53620 41310
rect 53564 41206 53620 41244
rect 54012 41300 54068 41310
rect 53452 41010 53508 41020
rect 53788 40180 53844 40190
rect 53564 40178 53844 40180
rect 53564 40126 53790 40178
rect 53842 40126 53844 40178
rect 53564 40124 53844 40126
rect 53564 39842 53620 40124
rect 53788 40114 53844 40124
rect 53564 39790 53566 39842
rect 53618 39790 53620 39842
rect 53564 39778 53620 39790
rect 53340 39676 53508 39732
rect 53452 39620 53508 39676
rect 53676 39620 53732 39630
rect 53452 39618 53732 39620
rect 53452 39566 53678 39618
rect 53730 39566 53732 39618
rect 53452 39564 53732 39566
rect 53676 39554 53732 39564
rect 53788 39620 53844 39630
rect 53900 39620 53956 39630
rect 53788 39618 53900 39620
rect 53788 39566 53790 39618
rect 53842 39566 53900 39618
rect 53788 39564 53900 39566
rect 53788 39554 53844 39564
rect 53340 39508 53396 39518
rect 53340 39506 53508 39508
rect 53340 39454 53342 39506
rect 53394 39454 53508 39506
rect 53340 39452 53508 39454
rect 53340 39442 53396 39452
rect 53116 39396 53172 39434
rect 53116 39330 53172 39340
rect 53116 39172 53172 39182
rect 53116 38946 53172 39116
rect 53116 38894 53118 38946
rect 53170 38894 53172 38946
rect 53116 38882 53172 38894
rect 53340 39060 53396 39070
rect 53340 38668 53396 39004
rect 53452 38948 53508 39452
rect 53788 39396 53844 39406
rect 53452 38882 53508 38892
rect 53564 39284 53620 39294
rect 53564 38724 53620 39228
rect 53004 38612 53172 38668
rect 52892 38546 52948 38556
rect 53116 38052 53172 38612
rect 52892 37996 53172 38052
rect 53228 38612 53284 38622
rect 53340 38612 53508 38668
rect 53564 38658 53620 38668
rect 53676 38948 53732 38958
rect 52892 37604 52948 37996
rect 53004 37828 53060 37838
rect 53004 37826 53172 37828
rect 53004 37774 53006 37826
rect 53058 37774 53172 37826
rect 53004 37772 53172 37774
rect 53004 37762 53060 37772
rect 52892 37548 53060 37604
rect 52892 37044 52948 37054
rect 52892 36950 52948 36988
rect 52668 36428 52836 36484
rect 52668 36036 52724 36428
rect 52668 35970 52724 35980
rect 52780 36260 52836 36270
rect 52556 35812 52612 35822
rect 52556 35718 52612 35756
rect 52668 35700 52724 35710
rect 52780 35700 52836 36204
rect 52668 35698 52836 35700
rect 52668 35646 52670 35698
rect 52722 35646 52836 35698
rect 52668 35644 52836 35646
rect 52668 35634 52724 35644
rect 52892 35586 52948 35598
rect 52892 35534 52894 35586
rect 52946 35534 52948 35586
rect 52892 35476 52948 35534
rect 52892 35410 52948 35420
rect 51772 34076 51940 34132
rect 52108 34636 52500 34692
rect 52780 35140 52836 35150
rect 51436 33506 51492 33516
rect 51660 33572 51716 33582
rect 50988 32732 51156 32788
rect 51212 33460 51268 33470
rect 50876 32564 50932 32574
rect 50484 32562 50932 32564
rect 50484 32510 50878 32562
rect 50930 32510 50932 32562
rect 50484 32508 50932 32510
rect 50428 32498 50484 32508
rect 50876 32498 50932 32508
rect 50204 32002 50372 32004
rect 50204 31950 50206 32002
rect 50258 31950 50372 32002
rect 50204 31948 50372 31950
rect 50428 32338 50484 32350
rect 50428 32286 50430 32338
rect 50482 32286 50484 32338
rect 50428 32004 50484 32286
rect 50204 31938 50260 31948
rect 50428 31938 50484 31948
rect 50652 32116 50708 32126
rect 50652 31890 50708 32060
rect 50652 31838 50654 31890
rect 50706 31838 50708 31890
rect 50652 31826 50708 31838
rect 50092 31726 50094 31778
rect 50146 31726 50148 31778
rect 50092 31714 50148 31726
rect 50428 31780 50484 31790
rect 50428 31686 50484 31724
rect 50316 31668 50372 31678
rect 50204 31556 50260 31566
rect 50092 30436 50148 30446
rect 50092 29652 50148 30380
rect 50204 30324 50260 31500
rect 50204 30258 50260 30268
rect 50316 30100 50372 31612
rect 50764 31332 50820 31342
rect 50988 31332 51044 32732
rect 51100 32564 51156 32574
rect 51212 32564 51268 33404
rect 51100 32562 51268 32564
rect 51100 32510 51102 32562
rect 51154 32510 51268 32562
rect 51100 32508 51268 32510
rect 51100 32498 51156 32508
rect 50820 31276 51044 31332
rect 50764 31266 50820 31276
rect 51212 30996 51268 32508
rect 51324 33346 51380 33358
rect 51324 33294 51326 33346
rect 51378 33294 51380 33346
rect 51324 31892 51380 33294
rect 51548 33346 51604 33358
rect 51548 33294 51550 33346
rect 51602 33294 51604 33346
rect 51436 33234 51492 33246
rect 51436 33182 51438 33234
rect 51490 33182 51492 33234
rect 51436 32788 51492 33182
rect 51436 32722 51492 32732
rect 51548 32676 51604 33294
rect 51548 32610 51604 32620
rect 51436 32338 51492 32350
rect 51436 32286 51438 32338
rect 51490 32286 51492 32338
rect 51436 32228 51492 32286
rect 51436 32162 51492 32172
rect 51548 32340 51604 32350
rect 51548 32004 51604 32284
rect 51548 31938 51604 31948
rect 51324 31836 51492 31892
rect 51324 31668 51380 31678
rect 51324 31574 51380 31612
rect 51324 31220 51380 31230
rect 51324 31126 51380 31164
rect 51212 30902 51268 30940
rect 50764 30770 50820 30782
rect 50764 30718 50766 30770
rect 50818 30718 50820 30770
rect 50764 30212 50820 30718
rect 51324 30772 51380 30782
rect 51324 30678 51380 30716
rect 51436 30436 51492 31836
rect 51660 30884 51716 33516
rect 51772 32116 51828 34076
rect 51996 34020 52052 34030
rect 51884 34018 52052 34020
rect 51884 33966 51998 34018
rect 52050 33966 52052 34018
rect 51884 33964 52052 33966
rect 51884 33572 51940 33964
rect 51996 33954 52052 33964
rect 51884 33506 51940 33516
rect 52108 33460 52164 34636
rect 52556 34244 52612 34254
rect 52556 34150 52612 34188
rect 52220 34130 52276 34142
rect 52220 34078 52222 34130
rect 52274 34078 52276 34130
rect 52220 33572 52276 34078
rect 52220 33506 52276 33516
rect 51996 33404 52164 33460
rect 52668 33460 52724 33470
rect 51884 33346 51940 33358
rect 51884 33294 51886 33346
rect 51938 33294 51940 33346
rect 51884 32564 51940 33294
rect 51884 32498 51940 32508
rect 51996 32562 52052 33404
rect 52668 33366 52724 33404
rect 52220 33348 52276 33358
rect 51996 32510 51998 32562
rect 52050 32510 52052 32562
rect 51996 32498 52052 32510
rect 52108 33346 52276 33348
rect 52108 33294 52222 33346
rect 52274 33294 52276 33346
rect 52108 33292 52276 33294
rect 51772 32060 52052 32116
rect 51660 30818 51716 30828
rect 51772 31892 51828 31902
rect 51324 30380 51492 30436
rect 51548 30772 51604 30782
rect 51212 30324 51268 30334
rect 51212 30230 51268 30268
rect 50764 30146 50820 30156
rect 50092 29586 50148 29596
rect 50204 30044 50372 30100
rect 50204 29540 50260 30044
rect 50204 29474 50260 29484
rect 50316 29428 50372 29438
rect 50316 29334 50372 29372
rect 50764 29426 50820 29438
rect 50764 29374 50766 29426
rect 50818 29374 50820 29426
rect 50204 29314 50260 29326
rect 50204 29262 50206 29314
rect 50258 29262 50260 29314
rect 50092 28754 50148 28766
rect 50092 28702 50094 28754
rect 50146 28702 50148 28754
rect 50092 24836 50148 28702
rect 50204 28084 50260 29262
rect 50764 29316 50820 29374
rect 50764 29250 50820 29260
rect 50988 29426 51044 29438
rect 50988 29374 50990 29426
rect 51042 29374 51044 29426
rect 50204 28018 50260 28028
rect 50316 29092 50372 29102
rect 50316 27858 50372 29036
rect 50988 28644 51044 29374
rect 51100 29204 51156 29214
rect 51324 29204 51380 30380
rect 51548 30100 51604 30716
rect 51660 30212 51716 30222
rect 51660 30118 51716 30156
rect 51100 29202 51380 29204
rect 51100 29150 51102 29202
rect 51154 29150 51380 29202
rect 51100 29148 51380 29150
rect 51436 30044 51604 30100
rect 51100 29138 51156 29148
rect 50988 28578 51044 28588
rect 51100 28980 51156 28990
rect 51100 28866 51156 28924
rect 51100 28814 51102 28866
rect 51154 28814 51156 28866
rect 50316 27806 50318 27858
rect 50370 27806 50372 27858
rect 50316 27794 50372 27806
rect 50652 28530 50708 28542
rect 50652 28478 50654 28530
rect 50706 28478 50708 28530
rect 50428 27074 50484 27086
rect 50428 27022 50430 27074
rect 50482 27022 50484 27074
rect 50428 26852 50484 27022
rect 50652 26908 50708 28478
rect 50876 27412 50932 27422
rect 50876 27186 50932 27356
rect 50876 27134 50878 27186
rect 50930 27134 50932 27186
rect 50876 27122 50932 27134
rect 51100 27076 51156 28814
rect 51100 27010 51156 27020
rect 51436 26908 51492 30044
rect 51772 29988 51828 31836
rect 50316 26796 50484 26852
rect 50540 26852 50708 26908
rect 50988 26852 51492 26908
rect 51548 29932 51828 29988
rect 51884 31220 51940 31230
rect 51884 30210 51940 31164
rect 51884 30158 51886 30210
rect 51938 30158 51940 30210
rect 50204 26066 50260 26078
rect 50204 26014 50206 26066
rect 50258 26014 50260 26066
rect 50204 25284 50260 26014
rect 50316 25732 50372 26796
rect 50540 26516 50596 26852
rect 50316 25666 50372 25676
rect 50428 26460 50596 26516
rect 50204 25218 50260 25228
rect 50316 24948 50372 24958
rect 50092 24780 50260 24836
rect 50092 22932 50148 22942
rect 49980 22876 50092 22932
rect 50092 22838 50148 22876
rect 50204 22820 50260 24780
rect 50204 22754 50260 22764
rect 49868 22540 50036 22596
rect 49756 22428 49924 22484
rect 49644 22372 49700 22382
rect 49700 22316 49812 22372
rect 49644 22306 49700 22316
rect 49756 22258 49812 22316
rect 49756 22206 49758 22258
rect 49810 22206 49812 22258
rect 49756 22194 49812 22206
rect 49532 20738 49588 20748
rect 49644 22148 49700 22158
rect 49420 20524 49588 20580
rect 49420 18452 49476 18462
rect 49308 18396 49420 18452
rect 48860 18050 48916 18060
rect 48748 17826 48804 17836
rect 48860 17554 48916 17566
rect 48860 17502 48862 17554
rect 48914 17502 48916 17554
rect 48860 17218 48916 17502
rect 48860 17162 49364 17218
rect 49196 16996 49252 17006
rect 48636 16772 48692 16782
rect 48636 16678 48692 16716
rect 48860 16436 48916 16446
rect 48860 16322 48916 16380
rect 48860 16270 48862 16322
rect 48914 16270 48916 16322
rect 48636 16098 48692 16110
rect 48636 16046 48638 16098
rect 48690 16046 48692 16098
rect 48636 15540 48692 16046
rect 48748 15988 48804 15998
rect 48748 15894 48804 15932
rect 48636 15474 48692 15484
rect 48524 14690 48580 14700
rect 48636 14980 48692 14990
rect 48636 14642 48692 14924
rect 48636 14590 48638 14642
rect 48690 14590 48692 14642
rect 48636 14578 48692 14590
rect 48748 14868 48804 14878
rect 48748 14642 48804 14812
rect 48748 14590 48750 14642
rect 48802 14590 48804 14642
rect 48748 14578 48804 14590
rect 47964 14354 48020 14364
rect 48412 14420 48468 14430
rect 48412 14326 48468 14364
rect 48188 14306 48244 14318
rect 48188 14254 48190 14306
rect 48242 14254 48244 14306
rect 48188 14196 48244 14254
rect 47404 14130 47460 14140
rect 47628 14140 48244 14196
rect 46956 13188 47012 13198
rect 46620 13134 46622 13186
rect 46674 13134 46676 13186
rect 46620 13122 46676 13134
rect 46844 13186 47012 13188
rect 46844 13134 46958 13186
rect 47010 13134 47012 13186
rect 46844 13132 47012 13134
rect 46060 13022 46062 13074
rect 46114 13022 46116 13074
rect 46060 12292 46116 13022
rect 46172 13076 46228 13086
rect 46172 12982 46228 13020
rect 46844 13076 46900 13132
rect 46956 13122 47012 13132
rect 47180 13186 47236 13198
rect 47180 13134 47182 13186
rect 47234 13134 47236 13186
rect 47180 13076 47236 13134
rect 47292 13188 47348 13580
rect 47404 13188 47460 13198
rect 47292 13186 47460 13188
rect 47292 13134 47406 13186
rect 47458 13134 47460 13186
rect 47292 13132 47460 13134
rect 47404 13122 47460 13132
rect 47180 13020 47348 13076
rect 46844 13010 46900 13020
rect 46508 12962 46564 12974
rect 46508 12910 46510 12962
rect 46562 12910 46564 12962
rect 46508 12628 46564 12910
rect 47292 12964 47348 13020
rect 47292 12908 47460 12964
rect 47068 12852 47124 12862
rect 47068 12850 47348 12852
rect 47068 12798 47070 12850
rect 47122 12798 47348 12850
rect 47068 12796 47348 12798
rect 47068 12786 47124 12796
rect 46508 12562 46564 12572
rect 46844 12516 46900 12526
rect 46060 12236 46228 12292
rect 45836 10668 46004 10724
rect 45836 7924 45892 10668
rect 45836 7858 45892 7868
rect 45948 10500 46004 10510
rect 45612 7746 45668 7756
rect 45836 7700 45892 7710
rect 44996 6188 45220 6244
rect 44940 6178 44996 6188
rect 44604 6078 44606 6130
rect 44658 6078 44660 6130
rect 44156 5796 44212 5806
rect 44604 5796 44660 6078
rect 44212 5740 44660 5796
rect 45052 5906 45108 5918
rect 45052 5854 45054 5906
rect 45106 5854 45108 5906
rect 44156 5730 44212 5740
rect 43484 5684 43540 5694
rect 42364 5346 42532 5348
rect 42364 5294 42366 5346
rect 42418 5294 42532 5346
rect 42364 5292 42532 5294
rect 43036 5682 43540 5684
rect 43036 5630 43486 5682
rect 43538 5630 43540 5682
rect 43036 5628 43540 5630
rect 42364 5282 42420 5292
rect 41804 5122 41972 5124
rect 41804 5070 41806 5122
rect 41858 5070 41972 5122
rect 41804 5068 41972 5070
rect 41804 5058 41860 5068
rect 40796 3332 40964 3388
rect 40684 2930 40740 2940
rect 40572 2716 40740 2772
rect 40572 2436 40628 2446
rect 40460 2098 40516 2110
rect 40460 2046 40462 2098
rect 40514 2046 40516 2098
rect 40012 1652 40068 1662
rect 40012 1202 40068 1596
rect 40012 1150 40014 1202
rect 40066 1150 40068 1202
rect 40012 1138 40068 1150
rect 39788 980 39844 990
rect 39788 886 39844 924
rect 40236 980 40292 990
rect 40236 532 40292 924
rect 40460 756 40516 2046
rect 40460 690 40516 700
rect 40124 476 40292 532
rect 40124 112 40180 476
rect 40572 112 40628 2380
rect 40684 1314 40740 2716
rect 40796 2212 40852 2222
rect 40796 2118 40852 2156
rect 40684 1262 40686 1314
rect 40738 1262 40740 1314
rect 40684 1250 40740 1262
rect 40908 1092 40964 3332
rect 41692 2770 41748 3388
rect 41804 4226 41860 4238
rect 41804 4174 41806 4226
rect 41858 4174 41860 4226
rect 41804 2996 41860 4174
rect 41916 4228 41972 5068
rect 42140 5030 42196 5068
rect 42588 5236 42644 5246
rect 42588 4338 42644 5180
rect 43036 5122 43092 5628
rect 43484 5618 43540 5628
rect 43596 5572 43652 5582
rect 43596 5460 43652 5516
rect 43036 5070 43038 5122
rect 43090 5070 43092 5122
rect 43036 5058 43092 5070
rect 43372 5404 43652 5460
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 44828 5460 44884 5470
rect 42588 4286 42590 4338
rect 42642 4286 42644 4338
rect 42588 4274 42644 4286
rect 42812 5012 42868 5022
rect 41916 4172 42196 4228
rect 42140 3778 42196 4172
rect 42140 3726 42142 3778
rect 42194 3726 42196 3778
rect 42140 3714 42196 3726
rect 42812 3778 42868 4956
rect 43372 4338 43428 5404
rect 44828 5346 44884 5404
rect 44828 5294 44830 5346
rect 44882 5294 44884 5346
rect 44828 5282 44884 5294
rect 43484 5124 43540 5134
rect 43484 5030 43540 5068
rect 44380 5124 44436 5162
rect 44380 5058 44436 5068
rect 44604 5124 44660 5134
rect 45052 5124 45108 5854
rect 45164 5794 45220 6188
rect 45612 6804 45668 6814
rect 45612 6466 45668 6748
rect 45836 6692 45892 7644
rect 45948 7698 46004 10444
rect 45948 7646 45950 7698
rect 46002 7646 46004 7698
rect 45948 6916 46004 7646
rect 46060 10388 46116 10398
rect 46060 6916 46116 10332
rect 46172 9154 46228 12236
rect 46396 12180 46452 12190
rect 46284 11506 46340 11518
rect 46284 11454 46286 11506
rect 46338 11454 46340 11506
rect 46284 11284 46340 11454
rect 46284 11218 46340 11228
rect 46396 10164 46452 12124
rect 46732 11844 46788 11854
rect 46732 11396 46788 11788
rect 46396 10098 46452 10108
rect 46620 11340 46788 11396
rect 46172 9102 46174 9154
rect 46226 9102 46228 9154
rect 46172 9090 46228 9102
rect 46508 9042 46564 9054
rect 46508 8990 46510 9042
rect 46562 8990 46564 9042
rect 46508 8482 46564 8990
rect 46508 8430 46510 8482
rect 46562 8430 46564 8482
rect 46508 8418 46564 8430
rect 46508 7812 46564 7822
rect 46508 7474 46564 7756
rect 46508 7422 46510 7474
rect 46562 7422 46564 7474
rect 46508 7410 46564 7422
rect 46620 7140 46676 11340
rect 46732 11172 46788 11182
rect 46732 10500 46788 11116
rect 46732 10434 46788 10444
rect 46844 9044 46900 12460
rect 46956 12180 47012 12190
rect 46956 11060 47012 12124
rect 47292 12178 47348 12796
rect 47292 12126 47294 12178
rect 47346 12126 47348 12178
rect 47292 12114 47348 12126
rect 47404 12068 47460 12908
rect 47628 12852 47684 14140
rect 47964 13972 48020 13982
rect 47964 13746 48020 13916
rect 48524 13972 48580 13982
rect 48524 13878 48580 13916
rect 48860 13972 48916 16270
rect 49196 16322 49252 16940
rect 49196 16270 49198 16322
rect 49250 16270 49252 16322
rect 49196 16258 49252 16270
rect 49308 16322 49364 17162
rect 49420 16772 49476 18396
rect 49420 16706 49476 16716
rect 49308 16270 49310 16322
rect 49362 16270 49364 16322
rect 49308 16258 49364 16270
rect 49420 16210 49476 16222
rect 49420 16158 49422 16210
rect 49474 16158 49476 16210
rect 49420 15988 49476 16158
rect 49420 15922 49476 15932
rect 48972 15764 49028 15774
rect 48972 15316 49028 15708
rect 48972 14642 49028 15260
rect 49420 15316 49476 15326
rect 49420 15202 49476 15260
rect 49420 15150 49422 15202
rect 49474 15150 49476 15202
rect 49420 15138 49476 15150
rect 49532 14980 49588 20524
rect 49644 18452 49700 22092
rect 49756 21362 49812 21374
rect 49756 21310 49758 21362
rect 49810 21310 49812 21362
rect 49756 21028 49812 21310
rect 49756 20962 49812 20972
rect 49756 20690 49812 20702
rect 49756 20638 49758 20690
rect 49810 20638 49812 20690
rect 49756 20018 49812 20638
rect 49756 19966 49758 20018
rect 49810 19966 49812 20018
rect 49756 19122 49812 19966
rect 49756 19070 49758 19122
rect 49810 19070 49812 19122
rect 49756 18900 49812 19070
rect 49756 18834 49812 18844
rect 49868 18564 49924 22428
rect 49980 21586 50036 22540
rect 49980 21534 49982 21586
rect 50034 21534 50036 21586
rect 49980 21522 50036 21534
rect 50204 21028 50260 21038
rect 50204 20934 50260 20972
rect 50092 20132 50148 20142
rect 50092 19906 50148 20076
rect 50092 19854 50094 19906
rect 50146 19854 50148 19906
rect 50092 19842 50148 19854
rect 50204 19346 50260 19358
rect 50204 19294 50206 19346
rect 50258 19294 50260 19346
rect 50204 19012 50260 19294
rect 50204 18946 50260 18956
rect 50316 18788 50372 24892
rect 50428 23268 50484 26460
rect 50540 26292 50596 26302
rect 50540 26290 50708 26292
rect 50540 26238 50542 26290
rect 50594 26238 50708 26290
rect 50540 26236 50708 26238
rect 50540 26226 50596 26236
rect 50540 25732 50596 25742
rect 50540 25508 50596 25676
rect 50540 25414 50596 25452
rect 50652 24948 50708 26236
rect 50988 26180 51044 26852
rect 50652 24882 50708 24892
rect 50764 26124 51044 26180
rect 51212 26290 51268 26302
rect 51212 26238 51214 26290
rect 51266 26238 51268 26290
rect 50652 24724 50708 24734
rect 50652 24610 50708 24668
rect 50652 24558 50654 24610
rect 50706 24558 50708 24610
rect 50652 24546 50708 24558
rect 50764 24276 50820 26124
rect 50988 25618 51044 25630
rect 50988 25566 50990 25618
rect 51042 25566 51044 25618
rect 50988 25508 51044 25566
rect 50988 25442 51044 25452
rect 50428 23202 50484 23212
rect 50652 24220 50820 24276
rect 50988 24948 51044 24958
rect 50540 22260 50596 22270
rect 50428 21362 50484 21374
rect 50428 21310 50430 21362
rect 50482 21310 50484 21362
rect 50428 20244 50484 21310
rect 50428 20178 50484 20188
rect 50316 18722 50372 18732
rect 50428 19572 50484 19582
rect 50428 18900 50484 19516
rect 50540 19460 50596 22204
rect 50540 19394 50596 19404
rect 49868 18508 50148 18564
rect 49644 18358 49700 18396
rect 49980 18338 50036 18350
rect 49980 18286 49982 18338
rect 50034 18286 50036 18338
rect 49756 18226 49812 18238
rect 49756 18174 49758 18226
rect 49810 18174 49812 18226
rect 49756 16996 49812 18174
rect 49644 16940 49812 16996
rect 49868 18226 49924 18238
rect 49868 18174 49870 18226
rect 49922 18174 49924 18226
rect 49644 16322 49700 16940
rect 49868 16884 49924 18174
rect 49980 16996 50036 18286
rect 50092 18228 50148 18508
rect 50092 17780 50148 18172
rect 50092 17714 50148 17724
rect 50204 18452 50260 18462
rect 49980 16930 50036 16940
rect 50092 17332 50148 17342
rect 49756 16828 49924 16884
rect 49756 16770 49812 16828
rect 49756 16718 49758 16770
rect 49810 16718 49812 16770
rect 49756 16706 49812 16718
rect 50092 16324 50148 17276
rect 50204 16882 50260 18396
rect 50316 18450 50372 18462
rect 50316 18398 50318 18450
rect 50370 18398 50372 18450
rect 50316 17106 50372 18398
rect 50428 17332 50484 18844
rect 50652 17892 50708 24220
rect 50988 23826 51044 24892
rect 50988 23774 50990 23826
rect 51042 23774 51044 23826
rect 50988 23762 51044 23774
rect 51100 24836 51156 24846
rect 50764 23268 50820 23278
rect 50764 22370 50820 23212
rect 51100 23156 51156 24780
rect 51212 23378 51268 26238
rect 51324 26178 51380 26190
rect 51324 26126 51326 26178
rect 51378 26126 51380 26178
rect 51324 25284 51380 26126
rect 51324 25218 51380 25228
rect 51548 25172 51604 29932
rect 51548 25106 51604 25116
rect 51660 29540 51716 29550
rect 51660 24612 51716 29484
rect 51884 29092 51940 30158
rect 51772 29036 51940 29092
rect 51772 26908 51828 29036
rect 51996 28980 52052 32060
rect 52108 30772 52164 33292
rect 52220 33282 52276 33292
rect 52444 33348 52500 33358
rect 52780 33348 52836 35084
rect 52444 33346 52612 33348
rect 52444 33294 52446 33346
rect 52498 33294 52612 33346
rect 52444 33292 52612 33294
rect 52444 33282 52500 33292
rect 52332 33234 52388 33246
rect 52332 33182 52334 33234
rect 52386 33182 52388 33234
rect 52220 33012 52276 33022
rect 52220 32340 52276 32956
rect 52332 32564 52388 33182
rect 52332 32508 52500 32564
rect 52332 32340 52388 32350
rect 52220 32338 52388 32340
rect 52220 32286 52334 32338
rect 52386 32286 52388 32338
rect 52220 32284 52388 32286
rect 52332 32274 52388 32284
rect 52332 31892 52388 31902
rect 52220 31668 52276 31678
rect 52220 30996 52276 31612
rect 52220 30902 52276 30940
rect 52108 30716 52276 30772
rect 52220 30434 52276 30716
rect 52220 30382 52222 30434
rect 52274 30382 52276 30434
rect 52220 30370 52276 30382
rect 52332 30434 52388 31836
rect 52332 30382 52334 30434
rect 52386 30382 52388 30434
rect 52108 30324 52164 30334
rect 52108 30230 52164 30268
rect 52332 29764 52388 30382
rect 51884 28924 52052 28980
rect 52108 29426 52164 29438
rect 52108 29374 52110 29426
rect 52162 29374 52164 29426
rect 51884 27748 51940 28924
rect 52108 28868 52164 29374
rect 52332 29092 52388 29708
rect 52444 29314 52500 32508
rect 52556 32228 52612 33292
rect 52780 33282 52836 33292
rect 52892 34244 52948 34254
rect 52892 32676 52948 34188
rect 53004 34020 53060 37548
rect 53116 37044 53172 37772
rect 53116 36978 53172 36988
rect 53116 36708 53172 36718
rect 53116 35588 53172 36652
rect 53116 35522 53172 35532
rect 53228 35810 53284 38556
rect 53228 35758 53230 35810
rect 53282 35758 53284 35810
rect 53004 33954 53060 33964
rect 53116 34130 53172 34142
rect 53116 34078 53118 34130
rect 53170 34078 53172 34130
rect 53116 33908 53172 34078
rect 53228 34132 53284 35758
rect 53340 37268 53396 37278
rect 53340 35140 53396 37212
rect 53452 35698 53508 38612
rect 53564 38052 53620 38062
rect 53564 37958 53620 37996
rect 53564 37044 53620 37054
rect 53564 36484 53620 36988
rect 53676 36708 53732 38892
rect 53788 37268 53844 39340
rect 53788 37202 53844 37212
rect 53900 37044 53956 39564
rect 54012 38834 54068 41244
rect 54796 41188 54852 42902
rect 54908 42754 54964 42766
rect 54908 42702 54910 42754
rect 54962 42702 54964 42754
rect 54908 41412 54964 42702
rect 55020 42084 55076 44270
rect 55020 42018 55076 42028
rect 54908 41346 54964 41356
rect 54684 41132 54852 41188
rect 54348 40180 54404 40190
rect 54348 40178 54628 40180
rect 54348 40126 54350 40178
rect 54402 40126 54628 40178
rect 54348 40124 54628 40126
rect 54348 40114 54404 40124
rect 54572 39842 54628 40124
rect 54572 39790 54574 39842
rect 54626 39790 54628 39842
rect 54572 39778 54628 39790
rect 54348 39620 54404 39630
rect 54348 39526 54404 39564
rect 54460 39506 54516 39518
rect 54460 39454 54462 39506
rect 54514 39454 54516 39506
rect 54012 38782 54014 38834
rect 54066 38782 54068 38834
rect 54012 38770 54068 38782
rect 54236 39060 54292 39070
rect 54124 38162 54180 38174
rect 54124 38110 54126 38162
rect 54178 38110 54180 38162
rect 53676 36642 53732 36652
rect 53788 36988 53956 37044
rect 54012 37042 54068 37054
rect 54012 36990 54014 37042
rect 54066 36990 54068 37042
rect 53676 36484 53732 36494
rect 53564 36482 53732 36484
rect 53564 36430 53678 36482
rect 53730 36430 53732 36482
rect 53564 36428 53732 36430
rect 53676 36418 53732 36428
rect 53788 36260 53844 36988
rect 53900 36708 53956 36718
rect 54012 36708 54068 36990
rect 54124 37044 54180 38110
rect 54124 36978 54180 36988
rect 54124 36708 54180 36718
rect 54012 36706 54180 36708
rect 54012 36654 54126 36706
rect 54178 36654 54180 36706
rect 54012 36652 54180 36654
rect 53900 36482 53956 36652
rect 54124 36642 54180 36652
rect 54236 36706 54292 39004
rect 54460 38836 54516 39454
rect 54460 38770 54516 38780
rect 54572 38948 54628 38958
rect 54348 38724 54404 38762
rect 54572 38668 54628 38892
rect 54684 38836 54740 41132
rect 54796 40964 54852 40974
rect 54796 40962 55076 40964
rect 54796 40910 54798 40962
rect 54850 40910 55076 40962
rect 54796 40908 55076 40910
rect 54796 40898 54852 40908
rect 54796 39732 54852 39742
rect 54796 39618 54852 39676
rect 54796 39566 54798 39618
rect 54850 39566 54852 39618
rect 54796 39554 54852 39566
rect 55020 39618 55076 40908
rect 55020 39566 55022 39618
rect 55074 39566 55076 39618
rect 55020 39554 55076 39566
rect 54684 38780 54964 38836
rect 54348 38658 54404 38668
rect 54236 36654 54238 36706
rect 54290 36654 54292 36706
rect 54236 36642 54292 36654
rect 54460 38612 54628 38668
rect 54908 38722 54964 38780
rect 54908 38670 54910 38722
rect 54962 38670 54964 38722
rect 54908 38658 54964 38670
rect 54684 38612 54740 38622
rect 53900 36430 53902 36482
rect 53954 36430 53956 36482
rect 53900 36418 53956 36430
rect 54348 36484 54404 36494
rect 54348 36390 54404 36428
rect 54460 36260 54516 38612
rect 54684 38518 54740 38556
rect 54796 38500 54852 38510
rect 54572 38052 54628 38062
rect 54572 37266 54628 37996
rect 54572 37214 54574 37266
rect 54626 37214 54628 37266
rect 54572 37202 54628 37214
rect 54796 36706 54852 38444
rect 55132 37604 55188 45052
rect 55244 44436 55300 46396
rect 55356 45668 55412 46622
rect 55356 45218 55412 45612
rect 55356 45166 55358 45218
rect 55410 45166 55412 45218
rect 55356 45154 55412 45166
rect 55468 45220 55524 49532
rect 55580 49522 55636 49532
rect 55580 48242 55636 48254
rect 55580 48190 55582 48242
rect 55634 48190 55636 48242
rect 55580 47572 55636 48190
rect 55692 47684 55748 49756
rect 55804 48132 55860 53676
rect 56028 53666 56084 53676
rect 56028 52724 56084 52734
rect 55916 52722 56084 52724
rect 55916 52670 56030 52722
rect 56082 52670 56084 52722
rect 55916 52668 56084 52670
rect 55916 51380 55972 52668
rect 56028 52658 56084 52668
rect 56028 52388 56084 52398
rect 56028 52294 56084 52332
rect 55916 51314 55972 51324
rect 56028 51156 56084 51166
rect 55916 51154 56084 51156
rect 55916 51102 56030 51154
rect 56082 51102 56084 51154
rect 55916 51100 56084 51102
rect 55916 50428 55972 51100
rect 56028 51090 56084 51100
rect 56140 50594 56196 50606
rect 56140 50542 56142 50594
rect 56194 50542 56196 50594
rect 55916 50372 56084 50428
rect 55804 48066 55860 48076
rect 55916 49586 55972 49598
rect 55916 49534 55918 49586
rect 55970 49534 55972 49586
rect 55916 47908 55972 49534
rect 56028 49252 56084 50372
rect 56140 49252 56196 50542
rect 56252 49812 56308 55246
rect 56364 54292 56420 54302
rect 56364 54290 56532 54292
rect 56364 54238 56366 54290
rect 56418 54238 56532 54290
rect 56364 54236 56532 54238
rect 56364 54226 56420 54236
rect 56364 53842 56420 53854
rect 56364 53790 56366 53842
rect 56418 53790 56420 53842
rect 56364 52948 56420 53790
rect 56364 52882 56420 52892
rect 56364 52724 56420 52734
rect 56364 52630 56420 52668
rect 56364 52274 56420 52286
rect 56364 52222 56366 52274
rect 56418 52222 56420 52274
rect 56364 51604 56420 52222
rect 56364 51538 56420 51548
rect 56364 51156 56420 51166
rect 56364 51062 56420 51100
rect 56364 50708 56420 50718
rect 56364 50614 56420 50652
rect 56252 49746 56308 49756
rect 56252 49588 56308 49598
rect 56252 49494 56308 49532
rect 56364 49252 56420 49262
rect 56140 49250 56420 49252
rect 56140 49198 56366 49250
rect 56418 49198 56420 49250
rect 56140 49196 56420 49198
rect 56028 49186 56084 49196
rect 56364 49186 56420 49196
rect 55916 47842 55972 47852
rect 56028 49028 56084 49038
rect 56028 47796 56084 48972
rect 56028 47730 56084 47740
rect 56140 48242 56196 48254
rect 56140 48190 56142 48242
rect 56194 48190 56196 48242
rect 55692 47618 55748 47628
rect 55580 47506 55636 47516
rect 56028 47460 56084 47470
rect 55692 47458 56084 47460
rect 55692 47406 56030 47458
rect 56082 47406 56084 47458
rect 55692 47404 56084 47406
rect 55468 45164 55636 45220
rect 55356 44436 55412 44446
rect 55244 44434 55412 44436
rect 55244 44382 55358 44434
rect 55410 44382 55412 44434
rect 55244 44380 55412 44382
rect 55356 44370 55412 44380
rect 55468 43316 55524 43326
rect 55244 42980 55300 42990
rect 55244 42886 55300 42924
rect 55244 42756 55300 42766
rect 55244 42532 55300 42700
rect 55244 42466 55300 42476
rect 55468 41860 55524 43260
rect 55468 41794 55524 41804
rect 55356 41188 55412 41198
rect 55356 41094 55412 41132
rect 55244 40962 55300 40974
rect 55244 40910 55246 40962
rect 55298 40910 55300 40962
rect 55244 39172 55300 40910
rect 55244 39106 55300 39116
rect 55356 40292 55412 40302
rect 55244 38722 55300 38734
rect 55244 38670 55246 38722
rect 55298 38670 55300 38722
rect 55244 38612 55300 38670
rect 55244 38546 55300 38556
rect 55132 37538 55188 37548
rect 55244 37826 55300 37838
rect 55244 37774 55246 37826
rect 55298 37774 55300 37826
rect 55132 37044 55188 37054
rect 55132 36950 55188 36988
rect 54796 36654 54798 36706
rect 54850 36654 54852 36706
rect 54796 36642 54852 36654
rect 53788 36204 53956 36260
rect 53452 35646 53454 35698
rect 53506 35646 53508 35698
rect 53452 35252 53508 35646
rect 53788 35474 53844 35486
rect 53788 35422 53790 35474
rect 53842 35422 53844 35474
rect 53452 35186 53508 35196
rect 53676 35364 53732 35374
rect 53340 35074 53396 35084
rect 53228 34066 53284 34076
rect 53564 35028 53620 35038
rect 53564 34132 53620 34972
rect 53564 34018 53620 34076
rect 53564 33966 53566 34018
rect 53618 33966 53620 34018
rect 53564 33954 53620 33966
rect 53116 33852 53284 33908
rect 53228 33796 53284 33852
rect 53228 33740 53620 33796
rect 53116 33684 53172 33694
rect 53116 33348 53172 33628
rect 53564 33572 53620 33740
rect 53676 33684 53732 35308
rect 53788 35252 53844 35422
rect 53788 33908 53844 35196
rect 53900 34804 53956 36204
rect 54236 36204 54516 36260
rect 54684 36484 54740 36494
rect 54236 35810 54292 36204
rect 54236 35758 54238 35810
rect 54290 35758 54292 35810
rect 54236 35746 54292 35758
rect 54124 35700 54180 35710
rect 54124 35606 54180 35644
rect 54124 35476 54180 35486
rect 54124 35364 54180 35420
rect 53900 34738 53956 34748
rect 54012 35308 54180 35364
rect 54684 35474 54740 36428
rect 54908 36484 54964 36494
rect 54796 36036 54852 36046
rect 54796 35810 54852 35980
rect 54796 35758 54798 35810
rect 54850 35758 54852 35810
rect 54796 35746 54852 35758
rect 54908 35698 54964 36428
rect 55132 36260 55188 36270
rect 54908 35646 54910 35698
rect 54962 35646 54964 35698
rect 54908 35634 54964 35646
rect 55020 36258 55188 36260
rect 55020 36206 55134 36258
rect 55186 36206 55188 36258
rect 55020 36204 55188 36206
rect 54684 35422 54686 35474
rect 54738 35422 54740 35474
rect 54012 34356 54068 35308
rect 54684 35252 54740 35422
rect 54740 35196 54852 35252
rect 54684 35186 54740 35196
rect 54796 35138 54852 35196
rect 54796 35086 54798 35138
rect 54850 35086 54852 35138
rect 54796 35074 54852 35086
rect 54684 35028 54740 35038
rect 54684 34934 54740 34972
rect 54572 34914 54628 34926
rect 54572 34862 54574 34914
rect 54626 34862 54628 34914
rect 54348 34804 54404 34814
rect 54348 34710 54404 34748
rect 54124 34692 54180 34702
rect 54124 34690 54292 34692
rect 54124 34638 54126 34690
rect 54178 34638 54292 34690
rect 54124 34636 54292 34638
rect 54124 34626 54180 34636
rect 54236 34580 54292 34636
rect 54572 34580 54628 34862
rect 55020 34804 55076 36204
rect 55132 36194 55188 36204
rect 55244 35924 55300 37774
rect 55356 36596 55412 40236
rect 55468 40178 55524 40190
rect 55468 40126 55470 40178
rect 55522 40126 55524 40178
rect 55468 37156 55524 40126
rect 55580 39508 55636 45164
rect 55692 42980 55748 47404
rect 56028 47394 56084 47404
rect 56028 46452 56084 46462
rect 56028 46358 56084 46396
rect 55916 46002 55972 46014
rect 55916 45950 55918 46002
rect 55970 45950 55972 46002
rect 55804 45332 55860 45342
rect 55804 45218 55860 45276
rect 55804 45166 55806 45218
rect 55858 45166 55860 45218
rect 55804 45154 55860 45166
rect 55804 43428 55860 43438
rect 55804 43334 55860 43372
rect 55692 42914 55748 42924
rect 55804 42420 55860 42430
rect 55692 41748 55748 41758
rect 55692 41654 55748 41692
rect 55804 40964 55860 42364
rect 55916 41412 55972 45950
rect 56028 45220 56084 45230
rect 56028 45106 56084 45164
rect 56028 45054 56030 45106
rect 56082 45054 56084 45106
rect 56028 45042 56084 45054
rect 56140 44548 56196 48190
rect 56252 48244 56308 48254
rect 56252 46788 56308 48188
rect 56476 48132 56532 54236
rect 56700 50428 56756 57344
rect 56588 50372 56756 50428
rect 56812 55636 56868 55646
rect 56588 48692 56644 50372
rect 56812 49028 56868 55580
rect 56812 48962 56868 48972
rect 57036 53060 57092 53070
rect 56588 48626 56644 48636
rect 56476 48076 56868 48132
rect 56364 48020 56420 48030
rect 56364 48018 56644 48020
rect 56364 47966 56366 48018
rect 56418 47966 56644 48018
rect 56364 47964 56644 47966
rect 56364 47954 56420 47964
rect 56476 47796 56532 47806
rect 56364 47572 56420 47582
rect 56364 47478 56420 47516
rect 56252 46722 56308 46732
rect 56364 46450 56420 46462
rect 56364 46398 56366 46450
rect 56418 46398 56420 46450
rect 56252 45890 56308 45902
rect 56252 45838 56254 45890
rect 56306 45838 56308 45890
rect 56252 45444 56308 45838
rect 56252 45378 56308 45388
rect 56364 45332 56420 46398
rect 56364 45266 56420 45276
rect 56476 45220 56532 47740
rect 56588 47068 56644 47964
rect 56588 47012 56756 47068
rect 56476 45154 56532 45164
rect 56364 44996 56420 45006
rect 56364 44994 56532 44996
rect 56364 44942 56366 44994
rect 56418 44942 56532 44994
rect 56364 44940 56532 44942
rect 56364 44930 56420 44940
rect 56252 44882 56308 44894
rect 56252 44830 56254 44882
rect 56306 44830 56308 44882
rect 56252 44772 56308 44830
rect 56252 44706 56308 44716
rect 56028 44492 56196 44548
rect 56028 42980 56084 44492
rect 56364 44436 56420 44446
rect 56364 44342 56420 44380
rect 56140 44324 56196 44334
rect 56140 44322 56308 44324
rect 56140 44270 56142 44322
rect 56194 44270 56308 44322
rect 56140 44268 56308 44270
rect 56140 44258 56196 44268
rect 56252 43652 56308 44268
rect 56476 43988 56532 44940
rect 56476 43922 56532 43932
rect 56252 43596 56532 43652
rect 56364 43428 56420 43438
rect 56364 43334 56420 43372
rect 56252 43314 56308 43326
rect 56252 43262 56254 43314
rect 56306 43262 56308 43314
rect 56028 42924 56196 42980
rect 55916 41346 55972 41356
rect 56028 42754 56084 42766
rect 56028 42702 56030 42754
rect 56082 42702 56084 42754
rect 55916 41188 55972 41198
rect 55916 41094 55972 41132
rect 55804 40898 55860 40908
rect 55916 40516 55972 40526
rect 55916 40422 55972 40460
rect 56028 39844 56084 42702
rect 56140 42532 56196 42924
rect 56252 42756 56308 43262
rect 56252 42690 56308 42700
rect 56364 42866 56420 42878
rect 56364 42814 56366 42866
rect 56418 42814 56420 42866
rect 56140 42476 56308 42532
rect 56140 42084 56196 42094
rect 56140 41990 56196 42028
rect 56252 41410 56308 42476
rect 56252 41358 56254 41410
rect 56306 41358 56308 41410
rect 56252 41346 56308 41358
rect 56364 41412 56420 42814
rect 56364 41346 56420 41356
rect 56476 41188 56532 43596
rect 56252 41132 56532 41188
rect 56028 39788 56196 39844
rect 56028 39620 56084 39630
rect 56028 39526 56084 39564
rect 55580 39442 55636 39452
rect 55804 39060 55860 39070
rect 55692 38948 55748 38958
rect 55692 38854 55748 38892
rect 55580 38836 55636 38846
rect 55580 38742 55636 38780
rect 55804 38834 55860 39004
rect 55804 38782 55806 38834
rect 55858 38782 55860 38834
rect 55804 38770 55860 38782
rect 55468 37090 55524 37100
rect 55580 38612 55636 38622
rect 55356 36540 55524 36596
rect 55356 36372 55412 36382
rect 55356 36278 55412 36316
rect 55468 36036 55524 36540
rect 55468 35970 55524 35980
rect 55356 35924 55412 35934
rect 55244 35922 55412 35924
rect 55244 35870 55358 35922
rect 55410 35870 55412 35922
rect 55244 35868 55412 35870
rect 55356 35858 55412 35868
rect 55132 35698 55188 35710
rect 55132 35646 55134 35698
rect 55186 35646 55188 35698
rect 55132 35588 55188 35646
rect 55132 35522 55188 35532
rect 55244 35700 55300 35710
rect 55244 35138 55300 35644
rect 55244 35086 55246 35138
rect 55298 35086 55300 35138
rect 55244 35074 55300 35086
rect 55356 34804 55412 34814
rect 55020 34738 55076 34748
rect 55132 34802 55412 34804
rect 55132 34750 55358 34802
rect 55410 34750 55412 34802
rect 55132 34748 55412 34750
rect 54236 34524 54404 34580
rect 54572 34524 55076 34580
rect 54348 34356 54404 34524
rect 54684 34356 54740 34366
rect 54012 34300 54292 34356
rect 54348 34354 54740 34356
rect 54348 34302 54686 34354
rect 54738 34302 54740 34354
rect 54348 34300 54740 34302
rect 53788 33842 53844 33852
rect 54012 34020 54068 34030
rect 53676 33628 53956 33684
rect 53564 33516 53732 33572
rect 53116 33282 53172 33292
rect 53452 33236 53508 33246
rect 53676 33236 53732 33516
rect 53900 33570 53956 33628
rect 53900 33518 53902 33570
rect 53954 33518 53956 33570
rect 53452 33234 53732 33236
rect 53452 33182 53454 33234
rect 53506 33182 53732 33234
rect 53452 33180 53732 33182
rect 53452 33170 53508 33180
rect 52668 32564 52724 32574
rect 52668 32562 52836 32564
rect 52668 32510 52670 32562
rect 52722 32510 52836 32562
rect 52668 32508 52836 32510
rect 52668 32498 52724 32508
rect 52556 32172 52724 32228
rect 52556 32004 52612 32014
rect 52556 29538 52612 31948
rect 52668 31780 52724 32172
rect 52780 32004 52836 32508
rect 52892 32562 52948 32620
rect 52892 32510 52894 32562
rect 52946 32510 52948 32562
rect 52892 32498 52948 32510
rect 53564 32564 53620 32574
rect 53340 32452 53396 32462
rect 53340 32450 53508 32452
rect 53340 32398 53342 32450
rect 53394 32398 53508 32450
rect 53340 32396 53508 32398
rect 53340 32386 53396 32396
rect 53116 32338 53172 32350
rect 53116 32286 53118 32338
rect 53170 32286 53172 32338
rect 52892 32004 52948 32014
rect 52780 32002 52948 32004
rect 52780 31950 52894 32002
rect 52946 31950 52948 32002
rect 52780 31948 52948 31950
rect 52892 31938 52948 31948
rect 53116 32004 53172 32286
rect 53116 31938 53172 31948
rect 53228 32338 53284 32350
rect 53228 32286 53230 32338
rect 53282 32286 53284 32338
rect 53228 31780 53284 32286
rect 53340 32228 53396 32238
rect 53452 32228 53508 32396
rect 53396 32172 53508 32228
rect 53340 32162 53396 32172
rect 52668 31724 53284 31780
rect 53004 31332 53060 31342
rect 52668 30884 52724 30894
rect 52668 30790 52724 30828
rect 52556 29486 52558 29538
rect 52610 29486 52612 29538
rect 52556 29474 52612 29486
rect 52668 30100 52724 30110
rect 52444 29262 52446 29314
rect 52498 29262 52500 29314
rect 52444 29250 52500 29262
rect 52332 29026 52388 29036
rect 52556 29204 52612 29214
rect 52668 29204 52724 30044
rect 52780 29428 52836 29438
rect 52780 29334 52836 29372
rect 53004 29316 53060 31276
rect 53228 30100 53284 30110
rect 53228 29650 53284 30044
rect 53340 30098 53396 30110
rect 53340 30046 53342 30098
rect 53394 30046 53396 30098
rect 53340 29876 53396 30046
rect 53340 29810 53396 29820
rect 53228 29598 53230 29650
rect 53282 29598 53284 29650
rect 53228 29586 53284 29598
rect 53340 29540 53396 29550
rect 53340 29426 53396 29484
rect 53340 29374 53342 29426
rect 53394 29374 53396 29426
rect 53340 29362 53396 29374
rect 53004 29260 53284 29316
rect 52668 29148 52836 29204
rect 52108 28802 52164 28812
rect 52556 28868 52612 29148
rect 52556 28802 52612 28812
rect 51996 28756 52052 28766
rect 51996 28082 52052 28700
rect 52220 28420 52276 28430
rect 52668 28420 52724 28430
rect 52220 28326 52276 28364
rect 52332 28418 52724 28420
rect 52332 28366 52670 28418
rect 52722 28366 52724 28418
rect 52332 28364 52724 28366
rect 51996 28030 51998 28082
rect 52050 28030 52052 28082
rect 51996 28018 52052 28030
rect 52108 28196 52164 28206
rect 52108 27858 52164 28140
rect 52108 27806 52110 27858
rect 52162 27806 52164 27858
rect 52108 27794 52164 27806
rect 52220 27970 52276 27982
rect 52220 27918 52222 27970
rect 52274 27918 52276 27970
rect 51884 27682 51940 27692
rect 51772 26852 51940 26908
rect 51884 26292 51940 26852
rect 52108 26850 52164 26862
rect 52108 26798 52110 26850
rect 52162 26798 52164 26850
rect 51996 26516 52052 26526
rect 52108 26516 52164 26798
rect 52220 26628 52276 27918
rect 52220 26562 52276 26572
rect 51996 26514 52164 26516
rect 51996 26462 51998 26514
rect 52050 26462 52164 26514
rect 51996 26460 52164 26462
rect 51996 26450 52052 26460
rect 52220 26292 52276 26302
rect 51884 26290 52276 26292
rect 51884 26238 52222 26290
rect 52274 26238 52276 26290
rect 51884 26236 52276 26238
rect 52220 26068 52276 26236
rect 52220 26002 52276 26012
rect 52332 25844 52388 28364
rect 52668 28354 52724 28364
rect 52780 28196 52836 29148
rect 53228 29202 53284 29260
rect 53228 29150 53230 29202
rect 53282 29150 53284 29202
rect 53228 29138 53284 29150
rect 53340 29092 53396 29102
rect 53340 28866 53396 29036
rect 53340 28814 53342 28866
rect 53394 28814 53396 28866
rect 53340 28802 53396 28814
rect 52892 28756 52948 28766
rect 52892 28642 52948 28700
rect 52892 28590 52894 28642
rect 52946 28590 52948 28642
rect 52892 28578 52948 28590
rect 53116 28642 53172 28654
rect 53116 28590 53118 28642
rect 53170 28590 53172 28642
rect 52780 28140 52948 28196
rect 52556 27860 52612 27870
rect 52556 27766 52612 27804
rect 52780 27858 52836 27870
rect 52780 27806 52782 27858
rect 52834 27806 52836 27858
rect 52780 27524 52836 27806
rect 52780 27458 52836 27468
rect 52668 27188 52724 27198
rect 52668 27094 52724 27132
rect 52892 26908 52948 28140
rect 53116 27188 53172 28590
rect 53228 28530 53284 28542
rect 53228 28478 53230 28530
rect 53282 28478 53284 28530
rect 53228 27300 53284 28478
rect 53564 28308 53620 32508
rect 53676 31666 53732 33180
rect 53788 33460 53844 33470
rect 53788 32450 53844 33404
rect 53900 32900 53956 33518
rect 54012 33124 54068 33964
rect 54012 33058 54068 33068
rect 53900 32834 53956 32844
rect 53788 32398 53790 32450
rect 53842 32398 53844 32450
rect 53788 32386 53844 32398
rect 54124 32338 54180 32350
rect 54124 32286 54126 32338
rect 54178 32286 54180 32338
rect 54012 32228 54068 32238
rect 53676 31614 53678 31666
rect 53730 31614 53732 31666
rect 53676 30996 53732 31614
rect 53788 32004 53844 32014
rect 53788 31218 53844 31948
rect 53788 31166 53790 31218
rect 53842 31166 53844 31218
rect 53788 31154 53844 31166
rect 53676 30930 53732 30940
rect 53676 30772 53732 30782
rect 53676 30322 53732 30716
rect 53676 30270 53678 30322
rect 53730 30270 53732 30322
rect 53676 30258 53732 30270
rect 53900 29876 53956 29886
rect 53900 29426 53956 29820
rect 53900 29374 53902 29426
rect 53954 29374 53956 29426
rect 53900 29316 53956 29374
rect 53900 29250 53956 29260
rect 53564 28242 53620 28252
rect 53676 29204 53732 29214
rect 53340 28084 53396 28094
rect 53340 27990 53396 28028
rect 53340 27748 53396 27758
rect 53340 27654 53396 27692
rect 53452 27746 53508 27758
rect 53452 27694 53454 27746
rect 53506 27694 53508 27746
rect 53228 27234 53284 27244
rect 53116 27122 53172 27132
rect 52780 26852 52948 26908
rect 53452 26964 53508 27694
rect 53452 26898 53508 26908
rect 53564 27188 53620 27198
rect 52444 26628 52500 26638
rect 52444 26290 52500 26572
rect 52556 26404 52612 26414
rect 52556 26310 52612 26348
rect 52444 26238 52446 26290
rect 52498 26238 52500 26290
rect 52444 26226 52500 26238
rect 52668 26292 52724 26302
rect 52668 26198 52724 26236
rect 52108 25788 52388 25844
rect 52556 26180 52612 26190
rect 52108 25730 52164 25788
rect 52108 25678 52110 25730
rect 52162 25678 52164 25730
rect 52108 25666 52164 25678
rect 52556 25732 52612 26124
rect 52668 25732 52724 25742
rect 52556 25730 52724 25732
rect 52556 25678 52670 25730
rect 52722 25678 52724 25730
rect 52556 25676 52724 25678
rect 52668 25666 52724 25676
rect 52780 25508 52836 26852
rect 52668 25452 52836 25508
rect 52892 26628 52948 26638
rect 51212 23326 51214 23378
rect 51266 23326 51268 23378
rect 51212 23314 51268 23326
rect 51324 24388 51380 24398
rect 50988 23100 51156 23156
rect 50764 22318 50766 22370
rect 50818 22318 50820 22370
rect 50764 22306 50820 22318
rect 50876 23044 50932 23054
rect 50876 22596 50932 22988
rect 50764 21476 50820 21486
rect 50764 21382 50820 21420
rect 50876 20132 50932 22540
rect 50988 22372 51044 23100
rect 50988 22306 51044 22316
rect 51100 22932 51156 22942
rect 50652 17826 50708 17836
rect 50764 20076 50932 20132
rect 50428 17266 50484 17276
rect 50764 17108 50820 20076
rect 50876 19908 50932 19918
rect 50876 18564 50932 19852
rect 51100 19236 51156 22876
rect 51324 22594 51380 24332
rect 51548 23828 51604 23838
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 22530 51380 22542
rect 51436 23714 51492 23726
rect 51436 23662 51438 23714
rect 51490 23662 51492 23714
rect 51212 21924 51268 21934
rect 51212 21586 51268 21868
rect 51212 21534 51214 21586
rect 51266 21534 51268 21586
rect 51212 21522 51268 21534
rect 51324 21476 51380 21486
rect 51436 21476 51492 23662
rect 51548 21586 51604 23772
rect 51548 21534 51550 21586
rect 51602 21534 51604 21586
rect 51548 21522 51604 21534
rect 51324 21474 51492 21476
rect 51324 21422 51326 21474
rect 51378 21422 51492 21474
rect 51324 21420 51492 21422
rect 51324 21410 51380 21420
rect 51660 20804 51716 24556
rect 51772 25396 51828 25406
rect 51772 22596 51828 25340
rect 52108 25396 52164 25406
rect 52108 25060 52164 25340
rect 52108 24994 52164 25004
rect 52444 24948 52500 24958
rect 52444 24854 52500 24892
rect 52108 24498 52164 24510
rect 52108 24446 52110 24498
rect 52162 24446 52164 24498
rect 52108 24052 52164 24446
rect 52556 24388 52612 24398
rect 52556 24162 52612 24332
rect 52556 24110 52558 24162
rect 52610 24110 52612 24162
rect 52556 24098 52612 24110
rect 52108 23986 52164 23996
rect 52668 23828 52724 25452
rect 51772 22530 51828 22540
rect 52108 23772 52724 23828
rect 52780 24610 52836 24622
rect 52780 24558 52782 24610
rect 52834 24558 52836 24610
rect 51660 20738 51716 20748
rect 51324 20580 51380 20590
rect 51212 20578 51380 20580
rect 51212 20526 51326 20578
rect 51378 20526 51380 20578
rect 51212 20524 51380 20526
rect 51212 19348 51268 20524
rect 51324 20514 51380 20524
rect 51884 20578 51940 20590
rect 51884 20526 51886 20578
rect 51938 20526 51940 20578
rect 51324 20244 51380 20254
rect 51324 20150 51380 20188
rect 51884 20244 51940 20526
rect 51996 20580 52052 20590
rect 51996 20486 52052 20524
rect 51884 20178 51940 20188
rect 52108 20188 52164 23772
rect 52220 23268 52276 23278
rect 52220 23174 52276 23212
rect 52668 23044 52724 23054
rect 52668 22950 52724 22988
rect 52444 22148 52500 22158
rect 52444 22146 52724 22148
rect 52444 22094 52446 22146
rect 52498 22094 52724 22146
rect 52444 22092 52724 22094
rect 52444 22082 52500 22092
rect 52332 21362 52388 21374
rect 52332 21310 52334 21362
rect 52386 21310 52388 21362
rect 52332 21140 52388 21310
rect 52332 21074 52388 21084
rect 52444 21362 52500 21374
rect 52444 21310 52446 21362
rect 52498 21310 52500 21362
rect 52332 20914 52388 20926
rect 52332 20862 52334 20914
rect 52386 20862 52388 20914
rect 52108 20132 52276 20188
rect 52108 19908 52164 19918
rect 52108 19814 52164 19852
rect 51884 19572 51940 19582
rect 51884 19348 51940 19516
rect 51212 19292 51828 19348
rect 51100 19180 51492 19236
rect 51324 19010 51380 19022
rect 51324 18958 51326 19010
rect 51378 18958 51380 19010
rect 51324 18676 51380 18958
rect 51324 18610 51380 18620
rect 50876 18498 50932 18508
rect 51212 18564 51268 18574
rect 51212 18470 51268 18508
rect 51324 18452 51380 18462
rect 51324 18358 51380 18396
rect 50876 18340 50932 18350
rect 50876 18246 50932 18284
rect 51100 18228 51156 18238
rect 51100 18226 51268 18228
rect 51100 18174 51102 18226
rect 51154 18174 51268 18226
rect 51100 18172 51268 18174
rect 51100 18162 51156 18172
rect 51100 17668 51156 17678
rect 50988 17556 51044 17566
rect 50316 17054 50318 17106
rect 50370 17054 50372 17106
rect 50316 17042 50372 17054
rect 50652 17052 50820 17108
rect 50876 17554 51044 17556
rect 50876 17502 50990 17554
rect 51042 17502 51044 17554
rect 50876 17500 51044 17502
rect 50204 16830 50206 16882
rect 50258 16830 50260 16882
rect 50204 16818 50260 16830
rect 50316 16658 50372 16670
rect 50316 16606 50318 16658
rect 50370 16606 50372 16658
rect 50316 16436 50372 16606
rect 50316 16370 50372 16380
rect 49644 16270 49646 16322
rect 49698 16270 49700 16322
rect 49644 16258 49700 16270
rect 49980 16268 50148 16324
rect 49644 15540 49700 15550
rect 49644 15316 49700 15484
rect 49644 15250 49700 15260
rect 49980 15314 50036 16268
rect 50204 16212 50260 16222
rect 50652 16212 50708 17052
rect 50764 16882 50820 16894
rect 50764 16830 50766 16882
rect 50818 16830 50820 16882
rect 50764 16660 50820 16830
rect 50764 16594 50820 16604
rect 50092 15988 50148 15998
rect 50092 15894 50148 15932
rect 50204 15986 50260 16156
rect 50204 15934 50206 15986
rect 50258 15934 50260 15986
rect 49980 15262 49982 15314
rect 50034 15262 50036 15314
rect 49980 15148 50036 15262
rect 50204 15204 50260 15934
rect 49532 14914 49588 14924
rect 49868 15092 49924 15102
rect 49980 15092 50148 15148
rect 50204 15138 50260 15148
rect 50316 16156 50708 16212
rect 50876 16212 50932 17500
rect 50988 17490 51044 17500
rect 50988 16884 51044 16894
rect 50988 16790 51044 16828
rect 49868 14754 49924 15036
rect 49868 14702 49870 14754
rect 49922 14702 49924 14754
rect 49868 14690 49924 14702
rect 48972 14590 48974 14642
rect 49026 14590 49028 14642
rect 48972 14578 49028 14590
rect 49532 14644 49588 14654
rect 49532 14550 49588 14588
rect 48860 13906 48916 13916
rect 48972 14420 49028 14430
rect 47964 13694 47966 13746
rect 48018 13694 48020 13746
rect 47964 13682 48020 13694
rect 48076 13522 48132 13534
rect 48076 13470 48078 13522
rect 48130 13470 48132 13522
rect 48076 13188 48132 13470
rect 48972 13300 49028 14364
rect 50092 14420 50148 15092
rect 50316 14980 50372 16156
rect 50876 16146 50932 16156
rect 50540 15986 50596 15998
rect 50540 15934 50542 15986
rect 50594 15934 50596 15986
rect 50428 15876 50484 15886
rect 50428 15202 50484 15820
rect 50540 15540 50596 15934
rect 50540 15474 50596 15484
rect 50652 15988 50708 15998
rect 50652 15314 50708 15932
rect 50764 15874 50820 15886
rect 50764 15822 50766 15874
rect 50818 15822 50820 15874
rect 50764 15764 50820 15822
rect 50876 15876 50932 15886
rect 50876 15782 50932 15820
rect 50764 15698 50820 15708
rect 50652 15262 50654 15314
rect 50706 15262 50708 15314
rect 50652 15250 50708 15262
rect 50428 15150 50430 15202
rect 50482 15150 50484 15202
rect 50428 15138 50484 15150
rect 51100 15202 51156 17612
rect 51212 16212 51268 18172
rect 51324 17108 51380 17118
rect 51324 17014 51380 17052
rect 51436 16884 51492 19180
rect 51772 19018 51828 19292
rect 51884 19234 51940 19292
rect 51884 19182 51886 19234
rect 51938 19182 51940 19234
rect 51884 19170 51940 19182
rect 51772 18962 52052 19018
rect 51660 18788 51716 18798
rect 51548 17554 51604 17566
rect 51548 17502 51550 17554
rect 51602 17502 51604 17554
rect 51548 17332 51604 17502
rect 51548 17266 51604 17276
rect 51212 16146 51268 16156
rect 51324 16828 51492 16884
rect 51100 15150 51102 15202
rect 51154 15150 51156 15202
rect 51100 15138 51156 15150
rect 50316 14924 50596 14980
rect 48972 13234 49028 13244
rect 49196 14196 49252 14206
rect 48076 13122 48132 13132
rect 48636 13188 48692 13198
rect 48636 12962 48692 13132
rect 48860 13188 48916 13198
rect 48860 13094 48916 13132
rect 48636 12910 48638 12962
rect 48690 12910 48692 12962
rect 47628 12796 48132 12852
rect 48076 12738 48132 12796
rect 48076 12686 48078 12738
rect 48130 12686 48132 12738
rect 47852 12516 47908 12526
rect 47908 12460 48020 12516
rect 47852 12450 47908 12460
rect 47964 12178 48020 12460
rect 47964 12126 47966 12178
rect 48018 12126 48020 12178
rect 47964 12114 48020 12126
rect 47516 12068 47572 12078
rect 47404 12066 47572 12068
rect 47404 12014 47518 12066
rect 47570 12014 47572 12066
rect 47404 12012 47572 12014
rect 46956 10994 47012 11004
rect 47068 11956 47124 11966
rect 46956 9044 47012 9054
rect 46844 9042 47012 9044
rect 46844 8990 46958 9042
rect 47010 8990 47012 9042
rect 46844 8988 47012 8990
rect 46956 8978 47012 8988
rect 46844 8820 46900 8830
rect 46844 7140 46900 8764
rect 46956 7924 47012 7934
rect 47068 7924 47124 11900
rect 47292 11844 47348 11854
rect 47292 10050 47348 11788
rect 47404 11508 47460 12012
rect 47516 12002 47572 12012
rect 47740 12068 47796 12078
rect 47740 12066 47908 12068
rect 47740 12014 47742 12066
rect 47794 12014 47908 12066
rect 47740 12012 47908 12014
rect 47740 12002 47796 12012
rect 47852 11956 47908 12012
rect 47852 11890 47908 11900
rect 47404 11414 47460 11452
rect 47852 11396 47908 11406
rect 48076 11396 48132 12686
rect 48300 12740 48356 12750
rect 48300 12738 48468 12740
rect 48300 12686 48302 12738
rect 48354 12686 48468 12738
rect 48300 12684 48468 12686
rect 48300 12674 48356 12684
rect 48412 12628 48468 12684
rect 48412 12572 48580 12628
rect 48300 12516 48356 12526
rect 48300 12290 48356 12460
rect 48300 12238 48302 12290
rect 48354 12238 48356 12290
rect 48300 12226 48356 12238
rect 48300 12068 48356 12078
rect 48524 12068 48580 12572
rect 48356 12012 48468 12068
rect 48300 12002 48356 12012
rect 48188 11954 48244 11966
rect 48188 11902 48190 11954
rect 48242 11902 48244 11954
rect 48188 11618 48244 11902
rect 48412 11954 48468 12012
rect 48412 11902 48414 11954
rect 48466 11902 48468 11954
rect 48412 11890 48468 11902
rect 48300 11844 48356 11854
rect 48300 11732 48356 11788
rect 48524 11732 48580 12012
rect 48636 12066 48692 12910
rect 48636 12014 48638 12066
rect 48690 12014 48692 12066
rect 48636 12002 48692 12014
rect 48748 12962 48804 12974
rect 48748 12910 48750 12962
rect 48802 12910 48804 12962
rect 48748 11956 48804 12910
rect 48972 12962 49028 12974
rect 48972 12910 48974 12962
rect 49026 12910 49028 12962
rect 48972 12516 49028 12910
rect 48972 12450 49028 12460
rect 48748 11890 48804 11900
rect 48300 11676 48580 11732
rect 48636 11844 48692 11854
rect 48188 11566 48190 11618
rect 48242 11566 48244 11618
rect 48188 11554 48244 11566
rect 48524 11396 48580 11406
rect 48076 11340 48244 11396
rect 47628 11060 47684 11070
rect 47292 9998 47294 10050
rect 47346 9998 47348 10050
rect 47292 9986 47348 9998
rect 47404 10164 47460 10174
rect 47404 10050 47460 10108
rect 47404 9998 47406 10050
rect 47458 9998 47460 10050
rect 47404 9716 47460 9998
rect 47404 9650 47460 9660
rect 47180 9604 47236 9614
rect 47180 9510 47236 9548
rect 47628 9492 47684 11004
rect 47740 10612 47796 10622
rect 47740 10518 47796 10556
rect 47852 9828 47908 11340
rect 47964 10500 48020 10510
rect 47964 10406 48020 10444
rect 48076 10498 48132 10510
rect 48076 10446 48078 10498
rect 48130 10446 48132 10498
rect 48076 10164 48132 10446
rect 48076 10098 48132 10108
rect 48188 10108 48244 11340
rect 48524 11302 48580 11340
rect 48524 11060 48580 11070
rect 48412 10612 48468 10622
rect 48412 10518 48468 10556
rect 48524 10498 48580 11004
rect 48524 10446 48526 10498
rect 48578 10446 48580 10498
rect 48524 10164 48580 10446
rect 48188 10052 48356 10108
rect 48524 10098 48580 10108
rect 48188 9940 48244 9950
rect 47852 9762 47908 9772
rect 48076 9938 48244 9940
rect 48076 9886 48190 9938
rect 48242 9886 48244 9938
rect 48076 9884 48244 9886
rect 47628 9436 47908 9492
rect 47740 9042 47796 9054
rect 47740 8990 47742 9042
rect 47794 8990 47796 9042
rect 47180 8932 47236 8942
rect 47180 8838 47236 8876
rect 47516 8372 47572 8382
rect 47180 7924 47236 7934
rect 47068 7868 47180 7924
rect 46956 7362 47012 7868
rect 47180 7858 47236 7868
rect 46956 7310 46958 7362
rect 47010 7310 47012 7362
rect 46956 7298 47012 7310
rect 47180 7476 47236 7486
rect 46844 7084 47012 7140
rect 46620 7074 46676 7084
rect 46172 6916 46228 6926
rect 46060 6914 46228 6916
rect 46060 6862 46174 6914
rect 46226 6862 46228 6914
rect 46060 6860 46228 6862
rect 45948 6850 46004 6860
rect 46172 6850 46228 6860
rect 46620 6916 46676 6926
rect 46284 6804 46340 6814
rect 46284 6710 46340 6748
rect 46620 6802 46676 6860
rect 46620 6750 46622 6802
rect 46674 6750 46676 6802
rect 46620 6738 46676 6750
rect 46060 6692 46116 6702
rect 45836 6690 46116 6692
rect 45836 6638 46062 6690
rect 46114 6638 46116 6690
rect 45836 6636 46116 6638
rect 46060 6626 46116 6636
rect 46508 6690 46564 6702
rect 46508 6638 46510 6690
rect 46562 6638 46564 6690
rect 45612 6414 45614 6466
rect 45666 6414 45668 6466
rect 45388 5908 45444 5918
rect 45612 5908 45668 6414
rect 45388 5906 45668 5908
rect 45388 5854 45390 5906
rect 45442 5854 45668 5906
rect 45388 5852 45668 5854
rect 45836 6356 45892 6366
rect 45388 5842 45444 5852
rect 45164 5742 45166 5794
rect 45218 5742 45220 5794
rect 45164 5730 45220 5742
rect 45836 5236 45892 6300
rect 44156 4900 44212 4910
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 43372 4286 43374 4338
rect 43426 4286 43428 4338
rect 43372 4274 43428 4286
rect 44156 4338 44212 4844
rect 44604 4452 44660 5068
rect 44604 4386 44660 4396
rect 44716 5068 45108 5124
rect 45724 5180 45892 5236
rect 44156 4286 44158 4338
rect 44210 4286 44212 4338
rect 44156 4274 44212 4286
rect 44492 4340 44548 4350
rect 44492 4246 44548 4284
rect 42812 3726 42814 3778
rect 42866 3726 42868 3778
rect 41804 2940 42308 2996
rect 41692 2718 41694 2770
rect 41746 2718 41748 2770
rect 41692 2706 41748 2718
rect 42140 2772 42196 2782
rect 41132 2660 41188 2670
rect 41132 2566 41188 2604
rect 41468 2548 41524 2558
rect 41468 2210 41524 2492
rect 41468 2158 41470 2210
rect 41522 2158 41524 2210
rect 41468 2146 41524 2158
rect 42140 2210 42196 2716
rect 42140 2158 42142 2210
rect 42194 2158 42196 2210
rect 42140 2146 42196 2158
rect 41132 2098 41188 2110
rect 41132 2046 41134 2098
rect 41186 2046 41188 2098
rect 41132 1428 41188 2046
rect 41132 1362 41188 1372
rect 41916 1764 41972 1774
rect 41020 1092 41076 1102
rect 40908 1090 41076 1092
rect 40908 1038 41022 1090
rect 41074 1038 41076 1090
rect 40908 1036 41076 1038
rect 41020 1026 41076 1036
rect 41468 1092 41524 1102
rect 41020 532 41076 542
rect 41020 112 41076 476
rect 41468 112 41524 1036
rect 41916 112 41972 1708
rect 42252 1426 42308 2940
rect 42812 2770 42868 3726
rect 44044 4228 44100 4238
rect 42812 2718 42814 2770
rect 42866 2718 42868 2770
rect 42812 2706 42868 2718
rect 43036 3666 43092 3678
rect 43036 3614 43038 3666
rect 43090 3614 43092 3666
rect 42476 2546 42532 2558
rect 42476 2494 42478 2546
rect 42530 2494 42532 2546
rect 42476 1988 42532 2494
rect 43036 2436 43092 3614
rect 43372 3554 43428 3566
rect 43372 3502 43374 3554
rect 43426 3502 43428 3554
rect 43372 2660 43428 3502
rect 44044 3444 44100 4172
rect 44268 4116 44324 4126
rect 44716 4116 44772 5068
rect 44940 4900 44996 4910
rect 44268 4114 44772 4116
rect 44268 4062 44270 4114
rect 44322 4062 44772 4114
rect 44268 4060 44772 4062
rect 44828 4564 44884 4574
rect 44828 4450 44884 4508
rect 44828 4398 44830 4450
rect 44882 4398 44884 4450
rect 44268 4050 44324 4060
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 44828 3778 44884 4398
rect 44828 3726 44830 3778
rect 44882 3726 44884 3778
rect 44828 3714 44884 3726
rect 44156 3668 44212 3678
rect 44156 3574 44212 3612
rect 44492 3668 44548 3678
rect 44044 3378 44100 3388
rect 43804 3164 44068 3174
rect 43484 3108 43540 3118
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 43484 2882 43540 3052
rect 43484 2830 43486 2882
rect 43538 2830 43540 2882
rect 43484 2818 43540 2830
rect 43596 2772 43652 2782
rect 43596 2678 43652 2716
rect 44492 2770 44548 3612
rect 44492 2718 44494 2770
rect 44546 2718 44548 2770
rect 44492 2706 44548 2718
rect 44828 3332 44884 3342
rect 44828 2770 44884 3276
rect 44828 2718 44830 2770
rect 44882 2718 44884 2770
rect 43372 2594 43428 2604
rect 44156 2660 44212 2670
rect 44156 2566 44212 2604
rect 43148 2548 43204 2558
rect 43148 2454 43204 2492
rect 43932 2548 43988 2558
rect 42476 1922 42532 1932
rect 42812 2380 43092 2436
rect 42252 1374 42254 1426
rect 42306 1374 42308 1426
rect 42252 1362 42308 1374
rect 42364 868 42420 878
rect 42364 112 42420 812
rect 42812 112 42868 2380
rect 42924 2212 42980 2222
rect 42924 1314 42980 2156
rect 43932 2210 43988 2492
rect 43932 2158 43934 2210
rect 43986 2158 43988 2210
rect 43932 2146 43988 2158
rect 44268 2548 44324 2558
rect 44268 2210 44324 2492
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 44268 2158 44270 2210
rect 44322 2158 44324 2210
rect 42924 1262 42926 1314
rect 42978 1262 42980 1314
rect 42924 1250 42980 1262
rect 43260 2098 43316 2110
rect 43260 2046 43262 2098
rect 43314 2046 43316 2098
rect 43260 1204 43316 2046
rect 43484 2100 43540 2110
rect 43260 1138 43316 1148
rect 43372 1876 43428 1886
rect 43148 978 43204 990
rect 43372 980 43428 1820
rect 43484 1202 43540 2044
rect 43484 1150 43486 1202
rect 43538 1150 43540 1202
rect 43484 1138 43540 1150
rect 43596 2098 43652 2110
rect 43596 2046 43598 2098
rect 43650 2046 43652 2098
rect 43596 1092 43652 2046
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 44268 1314 44324 2158
rect 44604 2098 44660 2110
rect 44604 2046 44606 2098
rect 44658 2046 44660 2098
rect 44604 1652 44660 2046
rect 44604 1586 44660 1596
rect 44268 1262 44270 1314
rect 44322 1262 44324 1314
rect 44268 1250 44324 1262
rect 44828 1314 44884 2718
rect 44940 2210 44996 4844
rect 45164 3666 45220 3678
rect 45164 3614 45166 3666
rect 45218 3614 45220 3666
rect 45164 3556 45220 3614
rect 45164 3490 45220 3500
rect 45500 3666 45556 3678
rect 45500 3614 45502 3666
rect 45554 3614 45556 3666
rect 45500 3388 45556 3614
rect 45276 3332 45556 3388
rect 45276 2772 45332 3332
rect 45724 2996 45780 5180
rect 46284 4338 46340 4350
rect 46284 4286 46286 4338
rect 46338 4286 46340 4338
rect 46172 3892 46228 3902
rect 46172 3778 46228 3836
rect 46172 3726 46174 3778
rect 46226 3726 46228 3778
rect 46172 3714 46228 3726
rect 45836 3554 45892 3566
rect 45836 3502 45838 3554
rect 45890 3502 45892 3554
rect 45836 3388 45892 3502
rect 45836 3332 46116 3388
rect 45724 2930 45780 2940
rect 44940 2158 44942 2210
rect 44994 2158 44996 2210
rect 44940 2146 44996 2158
rect 45052 2716 45332 2772
rect 45500 2772 45556 2782
rect 44828 1262 44830 1314
rect 44882 1262 44884 1314
rect 44828 1250 44884 1262
rect 45052 1204 45108 2716
rect 45500 2678 45556 2716
rect 45724 2772 45780 2782
rect 45388 2660 45444 2670
rect 45164 2546 45220 2558
rect 45164 2494 45166 2546
rect 45218 2494 45220 2546
rect 45164 2324 45220 2494
rect 45164 2258 45220 2268
rect 45276 2100 45332 2110
rect 45164 2098 45332 2100
rect 45164 2046 45278 2098
rect 45330 2046 45332 2098
rect 45164 2044 45332 2046
rect 45164 1540 45220 2044
rect 45276 2034 45332 2044
rect 45164 1474 45220 1484
rect 44940 1148 45108 1204
rect 45276 1428 45332 1438
rect 45276 1202 45332 1372
rect 45276 1150 45278 1202
rect 45330 1150 45332 1202
rect 43596 1026 43652 1036
rect 44044 1092 44100 1102
rect 43148 926 43150 978
rect 43202 926 43204 978
rect 43148 420 43204 926
rect 43148 354 43204 364
rect 43260 924 43428 980
rect 43260 112 43316 924
rect 44044 644 44100 1036
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 44940 644 44996 1148
rect 45276 1138 45332 1150
rect 45052 980 45108 990
rect 45388 980 45444 2604
rect 45612 2212 45668 2222
rect 45612 2118 45668 2156
rect 45724 1316 45780 2716
rect 46060 2660 46116 3332
rect 46284 2884 46340 4286
rect 46508 4340 46564 6638
rect 46508 4274 46564 4284
rect 46620 5124 46676 5134
rect 46508 4116 46564 4126
rect 46620 4116 46676 5068
rect 46508 4114 46676 4116
rect 46508 4062 46510 4114
rect 46562 4062 46676 4114
rect 46508 4060 46676 4062
rect 46844 5012 46900 5022
rect 46508 4050 46564 4060
rect 46508 3892 46564 3902
rect 46284 2818 46340 2828
rect 46396 3668 46452 3678
rect 46172 2660 46228 2670
rect 46060 2658 46228 2660
rect 46060 2606 46174 2658
rect 46226 2606 46228 2658
rect 46060 2604 46228 2606
rect 46172 2594 46228 2604
rect 45836 2548 45892 2558
rect 45836 2454 45892 2492
rect 45948 2436 46004 2446
rect 45836 1988 45892 1998
rect 45836 1894 45892 1932
rect 45052 886 45108 924
rect 45164 924 45444 980
rect 45500 1260 45780 1316
rect 45164 756 45220 924
rect 44044 578 44100 588
rect 44604 588 44996 644
rect 45052 700 45220 756
rect 44156 420 44212 430
rect 43820 308 43876 318
rect 43708 252 43820 308
rect 43708 112 43764 252
rect 43820 242 43876 252
rect 44156 112 44212 364
rect 44604 112 44660 588
rect 45052 112 45108 700
rect 45500 112 45556 1260
rect 45948 112 46004 2380
rect 46284 2212 46340 2222
rect 46284 1314 46340 2156
rect 46284 1262 46286 1314
rect 46338 1262 46340 1314
rect 46284 1250 46340 1262
rect 46396 112 46452 3612
rect 46508 2770 46564 3836
rect 46844 3778 46900 4956
rect 46844 3726 46846 3778
rect 46898 3726 46900 3778
rect 46508 2718 46510 2770
rect 46562 2718 46564 2770
rect 46508 2706 46564 2718
rect 46732 3556 46788 3566
rect 46620 2098 46676 2110
rect 46620 2046 46622 2098
rect 46674 2046 46676 2098
rect 46620 1988 46676 2046
rect 46620 1922 46676 1932
rect 46732 1428 46788 3500
rect 46844 2770 46900 3726
rect 46956 3108 47012 7084
rect 47180 6580 47236 7420
rect 47180 6514 47236 6524
rect 47068 6132 47124 6142
rect 47068 3892 47124 6076
rect 47068 3826 47124 3836
rect 47068 3668 47124 3678
rect 47068 3574 47124 3612
rect 47404 3556 47460 3566
rect 47404 3462 47460 3500
rect 47516 3220 47572 8316
rect 47740 8036 47796 8990
rect 47740 7970 47796 7980
rect 47852 3668 47908 9436
rect 48076 8932 48132 9884
rect 48188 9874 48244 9884
rect 48076 8866 48132 8876
rect 48188 9716 48244 9726
rect 48188 9044 48244 9660
rect 47964 8260 48020 8298
rect 48188 8260 48244 8988
rect 48300 8482 48356 10052
rect 48412 9828 48468 9838
rect 48412 9042 48468 9772
rect 48636 9380 48692 11788
rect 49084 11620 49140 11630
rect 48748 11508 48804 11518
rect 48748 11414 48804 11452
rect 49084 11506 49140 11564
rect 49084 11454 49086 11506
rect 49138 11454 49140 11506
rect 48748 10612 48804 10622
rect 48972 10612 49028 10622
rect 48748 10610 49028 10612
rect 48748 10558 48750 10610
rect 48802 10558 48974 10610
rect 49026 10558 49028 10610
rect 48748 10556 49028 10558
rect 48748 10546 48804 10556
rect 48972 10546 49028 10556
rect 48860 10276 48916 10286
rect 48412 8990 48414 9042
rect 48466 8990 48468 9042
rect 48412 8978 48468 8990
rect 48524 9324 48692 9380
rect 48748 9938 48804 9950
rect 48748 9886 48750 9938
rect 48802 9886 48804 9938
rect 48300 8430 48302 8482
rect 48354 8430 48356 8482
rect 48300 8418 48356 8430
rect 48300 8260 48356 8270
rect 48188 8258 48356 8260
rect 48188 8206 48302 8258
rect 48354 8206 48356 8258
rect 48188 8204 48356 8206
rect 47964 8194 48020 8204
rect 48300 8194 48356 8204
rect 48188 8036 48244 8046
rect 48188 7698 48244 7980
rect 48188 7646 48190 7698
rect 48242 7646 48244 7698
rect 48188 7634 48244 7646
rect 48300 7812 48356 7822
rect 48300 7476 48356 7756
rect 48300 7410 48356 7420
rect 47852 3602 47908 3612
rect 48412 6244 48468 6254
rect 47516 3154 47572 3164
rect 46956 3042 47012 3052
rect 48412 2996 48468 6188
rect 48412 2930 48468 2940
rect 46844 2718 46846 2770
rect 46898 2718 46900 2770
rect 46844 2706 46900 2718
rect 48412 2770 48468 2782
rect 48412 2718 48414 2770
rect 48466 2718 48468 2770
rect 47180 2546 47236 2558
rect 47180 2494 47182 2546
rect 47234 2494 47236 2546
rect 47180 2212 47236 2494
rect 47516 2546 47572 2558
rect 47516 2494 47518 2546
rect 47570 2494 47572 2546
rect 47516 2436 47572 2494
rect 47852 2548 47908 2558
rect 47852 2454 47908 2492
rect 48188 2548 48244 2558
rect 48188 2454 48244 2492
rect 47516 2370 47572 2380
rect 48412 2436 48468 2718
rect 48412 2370 48468 2380
rect 47180 2146 47236 2156
rect 47292 2324 47348 2334
rect 47292 2210 47348 2268
rect 47292 2158 47294 2210
rect 47346 2158 47348 2210
rect 47292 2146 47348 2158
rect 48076 2212 48132 2222
rect 46956 2098 47012 2110
rect 46956 2046 46958 2098
rect 47010 2046 47012 2098
rect 46956 1876 47012 2046
rect 46956 1810 47012 1820
rect 46732 1362 46788 1372
rect 47404 1764 47460 1774
rect 46956 1204 47012 1214
rect 46956 1110 47012 1148
rect 47292 1092 47348 1102
rect 46732 978 46788 990
rect 46732 926 46734 978
rect 46786 926 46788 978
rect 46732 532 46788 926
rect 46732 466 46788 476
rect 46844 980 46900 990
rect 46844 112 46900 924
rect 47292 112 47348 1036
rect 47404 1090 47460 1708
rect 47628 1652 47684 1662
rect 47628 1202 47684 1596
rect 48076 1314 48132 2156
rect 48412 2212 48468 2222
rect 48412 2118 48468 2156
rect 48076 1262 48078 1314
rect 48130 1262 48132 1314
rect 48076 1250 48132 1262
rect 48188 1876 48244 1886
rect 47628 1150 47630 1202
rect 47682 1150 47684 1202
rect 47628 1138 47684 1150
rect 47404 1038 47406 1090
rect 47458 1038 47460 1090
rect 47404 1026 47460 1038
rect 47740 756 47796 766
rect 47740 112 47796 700
rect 48188 112 48244 1820
rect 48300 978 48356 990
rect 48300 926 48302 978
rect 48354 926 48356 978
rect 48300 644 48356 926
rect 48524 756 48580 9324
rect 48636 8596 48692 8606
rect 48636 8370 48692 8540
rect 48636 8318 48638 8370
rect 48690 8318 48692 8370
rect 48636 8306 48692 8318
rect 48748 7698 48804 9886
rect 48748 7646 48750 7698
rect 48802 7646 48804 7698
rect 48748 7634 48804 7646
rect 48860 7364 48916 10220
rect 48972 9940 49028 9950
rect 48972 9826 49028 9884
rect 48972 9774 48974 9826
rect 49026 9774 49028 9826
rect 48972 8596 49028 9774
rect 49084 9044 49140 11454
rect 49196 9716 49252 14140
rect 49532 13972 49588 13982
rect 49308 13748 49364 13758
rect 49308 11844 49364 13692
rect 49420 12404 49476 12414
rect 49420 12066 49476 12348
rect 49420 12014 49422 12066
rect 49474 12014 49476 12066
rect 49420 12002 49476 12014
rect 49308 11788 49476 11844
rect 49420 10724 49476 11788
rect 49420 10658 49476 10668
rect 49532 10722 49588 13916
rect 49756 13748 49812 13758
rect 49644 13524 49700 13534
rect 49644 11956 49700 13468
rect 49756 12178 49812 13692
rect 50092 13746 50148 14364
rect 50092 13694 50094 13746
rect 50146 13694 50148 13746
rect 49756 12126 49758 12178
rect 49810 12126 49812 12178
rect 49756 12114 49812 12126
rect 49868 12852 49924 12862
rect 50092 12852 50148 13694
rect 50204 14868 50260 14878
rect 50204 13074 50260 14812
rect 50428 14420 50484 14430
rect 50428 14326 50484 14364
rect 50204 13022 50206 13074
rect 50258 13022 50260 13074
rect 50204 13010 50260 13022
rect 49868 12850 50148 12852
rect 49868 12798 49870 12850
rect 49922 12798 50148 12850
rect 49868 12796 50148 12798
rect 50428 12964 50484 12974
rect 49644 11900 49812 11956
rect 49532 10670 49534 10722
rect 49586 10670 49588 10722
rect 49532 10658 49588 10670
rect 49308 10612 49364 10622
rect 49308 10518 49364 10556
rect 49420 10388 49476 10398
rect 49308 10386 49476 10388
rect 49308 10334 49422 10386
rect 49474 10334 49476 10386
rect 49308 10332 49476 10334
rect 49308 10164 49364 10332
rect 49420 10322 49476 10332
rect 49644 10386 49700 10398
rect 49644 10334 49646 10386
rect 49698 10334 49700 10386
rect 49308 10098 49364 10108
rect 49644 10164 49700 10334
rect 49644 10098 49700 10108
rect 49420 9940 49476 9950
rect 49308 9828 49364 9838
rect 49308 9734 49364 9772
rect 49196 9650 49252 9660
rect 49308 9268 49364 9278
rect 49196 9044 49252 9054
rect 49084 9042 49252 9044
rect 49084 8990 49198 9042
rect 49250 8990 49252 9042
rect 49084 8988 49252 8990
rect 49196 8978 49252 8988
rect 48972 8530 49028 8540
rect 48860 7298 48916 7308
rect 48748 5908 48804 5918
rect 48636 5684 48692 5694
rect 48636 2884 48692 5628
rect 48748 4564 48804 5852
rect 48748 4498 48804 4508
rect 48972 5796 49028 5806
rect 48636 2818 48692 2828
rect 48748 3556 48804 3566
rect 48748 2210 48804 3500
rect 48860 2772 48916 2782
rect 48860 2658 48916 2716
rect 48860 2606 48862 2658
rect 48914 2606 48916 2658
rect 48860 2594 48916 2606
rect 48748 2158 48750 2210
rect 48802 2158 48804 2210
rect 48748 2146 48804 2158
rect 48972 1988 49028 5740
rect 49084 3444 49140 3454
rect 49084 2210 49140 3388
rect 49308 2660 49364 9212
rect 49420 8260 49476 9884
rect 49756 9940 49812 11900
rect 49756 9874 49812 9884
rect 49868 10276 49924 12796
rect 50316 12068 50372 12078
rect 50316 11974 50372 12012
rect 50204 11844 50260 11854
rect 50204 10498 50260 11788
rect 50204 10446 50206 10498
rect 50258 10446 50260 10498
rect 50204 10434 50260 10446
rect 50316 11282 50372 11294
rect 50316 11230 50318 11282
rect 50370 11230 50372 11282
rect 50316 10276 50372 11230
rect 50428 10610 50484 12908
rect 50428 10558 50430 10610
rect 50482 10558 50484 10610
rect 50428 10546 50484 10558
rect 49868 10220 50372 10276
rect 49532 8820 49588 8830
rect 49532 8482 49588 8764
rect 49532 8430 49534 8482
rect 49586 8430 49588 8482
rect 49532 8418 49588 8430
rect 49420 8204 49588 8260
rect 49420 5236 49476 5246
rect 49420 3108 49476 5180
rect 49532 3332 49588 8204
rect 49868 8036 49924 10220
rect 50204 10052 50260 10062
rect 49980 9602 50036 9614
rect 49980 9550 49982 9602
rect 50034 9550 50036 9602
rect 49980 9268 50036 9550
rect 49980 9202 50036 9212
rect 50204 9266 50260 9996
rect 50204 9214 50206 9266
rect 50258 9214 50260 9266
rect 50204 9202 50260 9214
rect 50316 9602 50372 9614
rect 50316 9550 50318 9602
rect 50370 9550 50372 9602
rect 50316 8820 50372 9550
rect 50540 9492 50596 14924
rect 50876 14756 50932 14766
rect 50876 14662 50932 14700
rect 51100 13746 51156 13758
rect 51100 13694 51102 13746
rect 51154 13694 51156 13746
rect 50764 13636 50820 13646
rect 50652 12404 50708 12414
rect 50652 12066 50708 12348
rect 50764 12292 50820 13580
rect 50876 13636 50932 13646
rect 50876 13634 51044 13636
rect 50876 13582 50878 13634
rect 50930 13582 51044 13634
rect 50876 13580 51044 13582
rect 50876 13570 50932 13580
rect 50876 13412 50932 13422
rect 50876 12404 50932 13356
rect 50988 12740 51044 13580
rect 50988 12674 51044 12684
rect 50988 12404 51044 12414
rect 50876 12402 51044 12404
rect 50876 12350 50990 12402
rect 51042 12350 51044 12402
rect 50876 12348 51044 12350
rect 50988 12338 51044 12348
rect 51100 12404 51156 13694
rect 51100 12338 51156 12348
rect 50764 12236 50932 12292
rect 50652 12014 50654 12066
rect 50706 12014 50708 12066
rect 50652 10724 50708 12014
rect 50764 11620 50820 11630
rect 50764 11526 50820 11564
rect 50652 10668 50820 10724
rect 50316 8754 50372 8764
rect 50428 9436 50596 9492
rect 50652 10498 50708 10510
rect 50652 10446 50654 10498
rect 50706 10446 50708 10498
rect 49868 7970 49924 7980
rect 49980 8708 50036 8718
rect 49868 7700 49924 7710
rect 49868 7362 49924 7644
rect 49868 7310 49870 7362
rect 49922 7310 49924 7362
rect 49868 7298 49924 7310
rect 49532 3266 49588 3276
rect 49756 5124 49812 5134
rect 49420 3052 49588 3108
rect 49308 2594 49364 2604
rect 49084 2158 49086 2210
rect 49138 2158 49140 2210
rect 49084 2146 49140 2158
rect 49196 2546 49252 2558
rect 49196 2494 49198 2546
rect 49250 2494 49252 2546
rect 49196 2212 49252 2494
rect 49196 2146 49252 2156
rect 49420 2098 49476 2110
rect 49420 2046 49422 2098
rect 49474 2046 49476 2098
rect 49196 1988 49252 1998
rect 48972 1932 49140 1988
rect 48636 1540 48692 1550
rect 48636 1202 48692 1484
rect 48636 1150 48638 1202
rect 48690 1150 48692 1202
rect 48636 1138 48692 1150
rect 48972 978 49028 990
rect 48972 926 48974 978
rect 49026 926 49028 978
rect 48524 700 48692 756
rect 48300 578 48356 588
rect 48636 112 48692 700
rect 48972 308 49028 926
rect 48972 242 49028 252
rect 49084 112 49140 1932
rect 49196 1202 49252 1932
rect 49196 1150 49198 1202
rect 49250 1150 49252 1202
rect 49196 1138 49252 1150
rect 49420 1092 49476 2046
rect 49420 1026 49476 1036
rect 49532 112 49588 3052
rect 49756 2210 49812 5068
rect 49756 2158 49758 2210
rect 49810 2158 49812 2210
rect 49756 2146 49812 2158
rect 49868 1428 49924 1438
rect 49868 1202 49924 1372
rect 49868 1150 49870 1202
rect 49922 1150 49924 1202
rect 49868 1138 49924 1150
rect 49644 978 49700 990
rect 49644 926 49646 978
rect 49698 926 49700 978
rect 49644 420 49700 926
rect 49980 868 50036 8652
rect 50316 8036 50372 8046
rect 50316 7476 50372 7980
rect 50204 7474 50372 7476
rect 50204 7422 50318 7474
rect 50370 7422 50372 7474
rect 50204 7420 50372 7422
rect 50204 6690 50260 7420
rect 50316 7410 50372 7420
rect 50204 6638 50206 6690
rect 50258 6638 50260 6690
rect 50204 6626 50260 6638
rect 50204 4004 50260 4014
rect 50204 3388 50260 3948
rect 50204 3332 50372 3388
rect 49980 812 50148 868
rect 50092 756 50148 812
rect 50092 690 50148 700
rect 49644 354 49700 364
rect 49980 644 50036 654
rect 49980 196 50036 588
rect 50316 308 50372 3332
rect 50316 242 50372 252
rect 49980 112 50036 140
rect 50428 112 50484 9436
rect 50540 9268 50596 9278
rect 50540 9174 50596 9212
rect 50652 9044 50708 10446
rect 50764 9828 50820 10668
rect 50764 9734 50820 9772
rect 50764 9044 50820 9054
rect 50652 8988 50764 9044
rect 50764 8930 50820 8988
rect 50764 8878 50766 8930
rect 50818 8878 50820 8930
rect 50652 8370 50708 8382
rect 50652 8318 50654 8370
rect 50706 8318 50708 8370
rect 50652 8148 50708 8318
rect 50652 8082 50708 8092
rect 50540 6802 50596 6814
rect 50540 6750 50542 6802
rect 50594 6750 50596 6802
rect 50540 6692 50596 6750
rect 50540 6626 50596 6636
rect 50764 6356 50820 8878
rect 50764 6290 50820 6300
rect 50764 3780 50820 3790
rect 50764 1202 50820 3724
rect 50876 1316 50932 12236
rect 51324 12180 51380 16828
rect 51548 16436 51604 16446
rect 51548 16210 51604 16380
rect 51548 16158 51550 16210
rect 51602 16158 51604 16210
rect 51548 16146 51604 16158
rect 51436 16100 51492 16110
rect 51436 16006 51492 16044
rect 51660 15876 51716 18732
rect 51996 18450 52052 18962
rect 52108 18564 52164 18574
rect 52108 18470 52164 18508
rect 51996 18398 51998 18450
rect 52050 18398 52052 18450
rect 51996 18386 52052 18398
rect 52108 18340 52164 18350
rect 51996 17892 52052 17902
rect 51996 17798 52052 17836
rect 52108 17668 52164 18284
rect 52108 16436 52164 17612
rect 52108 16370 52164 16380
rect 51996 16098 52052 16110
rect 51996 16046 51998 16098
rect 52050 16046 52052 16098
rect 51436 15820 51716 15876
rect 51884 15874 51940 15886
rect 51884 15822 51886 15874
rect 51938 15822 51940 15874
rect 51436 15314 51492 15820
rect 51436 15262 51438 15314
rect 51490 15262 51492 15314
rect 51436 15250 51492 15262
rect 51884 13972 51940 15822
rect 51996 14756 52052 16046
rect 52108 15540 52164 15550
rect 52108 15446 52164 15484
rect 51996 14690 52052 14700
rect 51884 13906 51940 13916
rect 51996 14306 52052 14318
rect 51996 14254 51998 14306
rect 52050 14254 52052 14306
rect 51996 13860 52052 14254
rect 51996 13794 52052 13804
rect 51996 13634 52052 13646
rect 51996 13582 51998 13634
rect 52050 13582 52052 13634
rect 51436 13524 51492 13534
rect 51436 13522 51940 13524
rect 51436 13470 51438 13522
rect 51490 13470 51940 13522
rect 51436 13468 51940 13470
rect 51436 13458 51492 13468
rect 51884 13074 51940 13468
rect 51884 13022 51886 13074
rect 51938 13022 51940 13074
rect 51884 13010 51940 13022
rect 51772 12852 51828 12862
rect 51436 12740 51492 12750
rect 51436 12646 51492 12684
rect 51212 12124 51380 12180
rect 50988 10610 51044 10622
rect 50988 10558 50990 10610
rect 51042 10558 51044 10610
rect 50988 8372 51044 10558
rect 51212 10164 51268 12124
rect 51324 11954 51380 11966
rect 51324 11902 51326 11954
rect 51378 11902 51380 11954
rect 51324 11844 51380 11902
rect 51324 11778 51380 11788
rect 51324 10388 51380 10398
rect 51324 10386 51492 10388
rect 51324 10334 51326 10386
rect 51378 10334 51492 10386
rect 51324 10332 51492 10334
rect 51324 10322 51380 10332
rect 51212 10108 51380 10164
rect 51100 9940 51156 9950
rect 51100 9938 51268 9940
rect 51100 9886 51102 9938
rect 51154 9886 51268 9938
rect 51100 9884 51268 9886
rect 51100 9874 51156 9884
rect 51100 8930 51156 8942
rect 51100 8878 51102 8930
rect 51154 8878 51156 8930
rect 51100 8372 51156 8878
rect 51212 8484 51268 9884
rect 51324 9268 51380 10108
rect 51436 10052 51492 10332
rect 51436 9986 51492 9996
rect 51660 10164 51716 10174
rect 51660 10050 51716 10108
rect 51660 9998 51662 10050
rect 51714 9998 51716 10050
rect 51660 9986 51716 9998
rect 51772 9604 51828 12796
rect 51996 12404 52052 13582
rect 52108 13522 52164 13534
rect 52108 13470 52110 13522
rect 52162 13470 52164 13522
rect 52108 13186 52164 13470
rect 52220 13412 52276 20132
rect 52332 18564 52388 20862
rect 52444 20580 52500 21310
rect 52556 21364 52612 21374
rect 52556 21270 52612 21308
rect 52668 20916 52724 22092
rect 52780 21252 52836 24558
rect 52892 23268 52948 26572
rect 53564 26290 53620 27132
rect 53676 26740 53732 29148
rect 54012 29092 54068 32172
rect 54124 32116 54180 32286
rect 54236 32340 54292 34300
rect 54684 34290 54740 34300
rect 54236 32274 54292 32284
rect 54348 34132 54404 34142
rect 54124 32060 54292 32116
rect 54124 31892 54180 31902
rect 54124 31798 54180 31836
rect 54236 31332 54292 32060
rect 54348 31668 54404 34076
rect 54348 31602 54404 31612
rect 54460 34020 54516 34030
rect 54460 31444 54516 33964
rect 55020 33570 55076 34524
rect 55020 33518 55022 33570
rect 55074 33518 55076 33570
rect 55020 33506 55076 33518
rect 54572 32564 54628 32574
rect 54572 32562 54740 32564
rect 54572 32510 54574 32562
rect 54626 32510 54740 32562
rect 54572 32508 54740 32510
rect 54572 32498 54628 32508
rect 54460 31378 54516 31388
rect 54236 31266 54292 31276
rect 54348 30996 54404 31006
rect 54236 29988 54292 29998
rect 54236 29314 54292 29932
rect 54236 29262 54238 29314
rect 54290 29262 54292 29314
rect 54236 29250 54292 29262
rect 54348 29316 54404 30940
rect 54684 30772 54740 32508
rect 54796 32562 54852 32574
rect 55132 32564 55188 34748
rect 55356 34738 55412 34748
rect 55580 34692 55636 38556
rect 56028 38610 56084 38622
rect 56028 38558 56030 38610
rect 56082 38558 56084 38610
rect 56028 38276 56084 38558
rect 55804 38220 56084 38276
rect 55692 36932 55748 36942
rect 55692 35698 55748 36876
rect 55804 36372 55860 38220
rect 56028 38052 56084 38062
rect 56028 37958 56084 37996
rect 56140 36820 56196 39788
rect 56252 39842 56308 41132
rect 56252 39790 56254 39842
rect 56306 39790 56308 39842
rect 56252 39778 56308 39790
rect 56588 41076 56644 41086
rect 56476 39508 56532 39518
rect 56476 38668 56532 39452
rect 56252 38612 56532 38668
rect 56588 38612 56644 41020
rect 56252 37268 56308 38612
rect 56588 38546 56644 38556
rect 56700 38500 56756 47012
rect 56812 42084 56868 48076
rect 57036 47796 57092 53004
rect 57260 52948 57316 52958
rect 57260 50428 57316 52892
rect 57260 50372 57428 50428
rect 57036 47730 57092 47740
rect 57148 47908 57204 47918
rect 57036 47572 57092 47582
rect 56812 42018 56868 42028
rect 56924 44436 56980 44446
rect 56812 41636 56868 41646
rect 56812 38724 56868 41580
rect 56812 38658 56868 38668
rect 56700 38434 56756 38444
rect 56588 38388 56644 38398
rect 56364 38164 56420 38174
rect 56364 38070 56420 38108
rect 56476 37380 56532 37390
rect 56252 37212 56420 37268
rect 56028 36764 56196 36820
rect 56252 37042 56308 37054
rect 56252 36990 56254 37042
rect 56306 36990 56308 37042
rect 55916 36596 55972 36606
rect 55916 36502 55972 36540
rect 55804 36306 55860 36316
rect 55804 35924 55860 35934
rect 55804 35810 55860 35868
rect 55804 35758 55806 35810
rect 55858 35758 55860 35810
rect 55804 35746 55860 35758
rect 55692 35646 55694 35698
rect 55746 35646 55748 35698
rect 55692 35634 55748 35646
rect 55916 35474 55972 35486
rect 55916 35422 55918 35474
rect 55970 35422 55972 35474
rect 55916 34916 55972 35422
rect 55916 34850 55972 34860
rect 55468 34636 55636 34692
rect 55916 34692 55972 34702
rect 55468 34580 55524 34636
rect 55916 34598 55972 34636
rect 55244 34524 55524 34580
rect 55244 34132 55300 34524
rect 56028 34356 56084 36764
rect 56140 36594 56196 36606
rect 56140 36542 56142 36594
rect 56194 36542 56196 36594
rect 56140 36372 56196 36542
rect 56252 36484 56308 36990
rect 56252 36418 56308 36428
rect 56140 35476 56196 36316
rect 56252 36260 56308 36270
rect 56252 36166 56308 36204
rect 56140 35382 56196 35420
rect 56140 35028 56196 35038
rect 56140 34934 56196 34972
rect 56140 34804 56196 34814
rect 56140 34710 56196 34748
rect 55804 34300 56084 34356
rect 55692 34244 55748 34254
rect 55692 34150 55748 34188
rect 55244 34066 55300 34076
rect 55356 34132 55412 34142
rect 55356 34130 55636 34132
rect 55356 34078 55358 34130
rect 55410 34078 55636 34130
rect 55356 34076 55636 34078
rect 55356 34066 55412 34076
rect 55244 33908 55300 33918
rect 55244 33906 55412 33908
rect 55244 33854 55246 33906
rect 55298 33854 55412 33906
rect 55244 33852 55412 33854
rect 55244 33842 55300 33852
rect 54796 32510 54798 32562
rect 54850 32510 54852 32562
rect 54796 31220 54852 32510
rect 54796 31154 54852 31164
rect 54908 32508 55188 32564
rect 54908 30996 54964 32508
rect 55020 32338 55076 32350
rect 55020 32286 55022 32338
rect 55074 32286 55076 32338
rect 55020 32004 55076 32286
rect 55132 32340 55188 32350
rect 55132 32246 55188 32284
rect 55244 32338 55300 32350
rect 55244 32286 55246 32338
rect 55298 32286 55300 32338
rect 55244 32228 55300 32286
rect 55244 32162 55300 32172
rect 55356 32116 55412 33852
rect 55356 32050 55412 32060
rect 55468 33906 55524 33918
rect 55468 33854 55470 33906
rect 55522 33854 55524 33906
rect 55020 31948 55188 32004
rect 55132 31668 55188 31948
rect 55244 31892 55300 31902
rect 55468 31892 55524 33854
rect 55244 31890 55524 31892
rect 55244 31838 55246 31890
rect 55298 31838 55524 31890
rect 55244 31836 55524 31838
rect 55244 31826 55300 31836
rect 55132 31612 55524 31668
rect 54908 30940 55076 30996
rect 54684 30716 54852 30772
rect 54796 30212 54852 30716
rect 54908 30770 54964 30782
rect 54908 30718 54910 30770
rect 54962 30718 54964 30770
rect 54908 30548 54964 30718
rect 54908 30482 54964 30492
rect 54908 30212 54964 30222
rect 54796 30210 54964 30212
rect 54796 30158 54910 30210
rect 54962 30158 54964 30210
rect 54796 30156 54964 30158
rect 54908 30146 54964 30156
rect 55020 29764 55076 30940
rect 55020 29698 55076 29708
rect 55468 29650 55524 31612
rect 55580 31108 55636 34076
rect 55804 33124 55860 34300
rect 55916 34130 55972 34142
rect 55916 34078 55918 34130
rect 55970 34078 55972 34130
rect 55916 33236 55972 34078
rect 56364 33908 56420 37212
rect 56476 36148 56532 37324
rect 56476 36082 56532 36092
rect 56364 33842 56420 33852
rect 56588 33684 56644 38332
rect 56812 38164 56868 38174
rect 56588 33618 56644 33628
rect 56700 38052 56756 38062
rect 56028 33460 56084 33470
rect 56364 33460 56420 33470
rect 56028 33458 56308 33460
rect 56028 33406 56030 33458
rect 56082 33406 56308 33458
rect 56028 33404 56308 33406
rect 56028 33394 56084 33404
rect 55916 33180 56196 33236
rect 55804 33068 56084 33124
rect 55692 32452 55748 32462
rect 55692 32358 55748 32396
rect 56028 32450 56084 33068
rect 56028 32398 56030 32450
rect 56082 32398 56084 32450
rect 56028 32386 56084 32398
rect 56028 31778 56084 31790
rect 56028 31726 56030 31778
rect 56082 31726 56084 31778
rect 56028 31556 56084 31726
rect 56028 31490 56084 31500
rect 56028 31220 56084 31230
rect 56140 31220 56196 33180
rect 56028 31218 56196 31220
rect 56028 31166 56030 31218
rect 56082 31166 56196 31218
rect 56028 31164 56196 31166
rect 56028 31154 56084 31164
rect 55580 31052 55972 31108
rect 55468 29598 55470 29650
rect 55522 29598 55524 29650
rect 55468 29586 55524 29598
rect 55580 30660 55636 30670
rect 54348 29092 54404 29260
rect 53900 29036 54068 29092
rect 54236 29036 54404 29092
rect 55132 29092 55188 29102
rect 53900 28644 53956 29036
rect 53788 28642 53956 28644
rect 53788 28590 53902 28642
rect 53954 28590 53956 28642
rect 53788 28588 53956 28590
rect 53788 27860 53844 28588
rect 53900 28578 53956 28588
rect 54124 28642 54180 28654
rect 54124 28590 54126 28642
rect 54178 28590 54180 28642
rect 54012 28532 54068 28542
rect 54012 28438 54068 28476
rect 54124 28196 54180 28590
rect 54124 28130 54180 28140
rect 53900 28084 53956 28094
rect 53900 27990 53956 28028
rect 53788 27804 53956 27860
rect 53676 26674 53732 26684
rect 53788 27412 53844 27422
rect 53788 27298 53844 27356
rect 53788 27246 53790 27298
rect 53842 27246 53844 27298
rect 53788 26516 53844 27246
rect 53788 26450 53844 26460
rect 53564 26238 53566 26290
rect 53618 26238 53620 26290
rect 53564 26180 53620 26238
rect 53900 26292 53956 27804
rect 54236 27188 54292 29036
rect 55020 28868 55076 28878
rect 55020 28774 55076 28812
rect 54348 28756 54404 28766
rect 54348 28642 54404 28700
rect 54348 28590 54350 28642
rect 54402 28590 54404 28642
rect 54348 28578 54404 28590
rect 54796 28644 54852 28654
rect 54572 28418 54628 28430
rect 54572 28366 54574 28418
rect 54626 28366 54628 28418
rect 54572 27636 54628 28366
rect 54236 27122 54292 27132
rect 54460 27580 54628 27636
rect 54236 26962 54292 26974
rect 54236 26910 54238 26962
rect 54290 26910 54292 26962
rect 53900 26226 53956 26236
rect 54012 26852 54068 26862
rect 53564 25732 53620 26124
rect 54012 26178 54068 26796
rect 54012 26126 54014 26178
rect 54066 26126 54068 26178
rect 54012 26114 54068 26126
rect 54236 26180 54292 26910
rect 54460 26740 54516 27580
rect 54796 27300 54852 28588
rect 54908 28418 54964 28430
rect 54908 28366 54910 28418
rect 54962 28366 54964 28418
rect 54908 28308 54964 28366
rect 54908 28242 54964 28252
rect 55020 27748 55076 27758
rect 55020 27654 55076 27692
rect 54908 27300 54964 27310
rect 54796 27298 54964 27300
rect 54796 27246 54910 27298
rect 54962 27246 54964 27298
rect 54796 27244 54964 27246
rect 54908 27234 54964 27244
rect 55020 27300 55076 27310
rect 55020 27206 55076 27244
rect 55132 27076 55188 29036
rect 55580 28644 55636 30604
rect 55916 30322 55972 31052
rect 56140 30436 56196 30446
rect 56140 30342 56196 30380
rect 55916 30270 55918 30322
rect 55970 30270 55972 30322
rect 55916 30258 55972 30270
rect 55580 28578 55636 28588
rect 55804 30212 55860 30222
rect 54460 26674 54516 26684
rect 54572 27020 55188 27076
rect 55244 28418 55300 28430
rect 55244 28366 55246 28418
rect 55298 28366 55300 28418
rect 55244 27076 55300 28366
rect 54236 26114 54292 26124
rect 53004 25620 53060 25630
rect 53004 25618 53172 25620
rect 53004 25566 53006 25618
rect 53058 25566 53172 25618
rect 53004 25564 53172 25566
rect 53004 25554 53060 25564
rect 53004 24052 53060 24062
rect 53004 23938 53060 23996
rect 53004 23886 53006 23938
rect 53058 23886 53060 23938
rect 53004 23874 53060 23886
rect 52892 23202 52948 23212
rect 53116 22932 53172 25564
rect 53564 25396 53620 25676
rect 54348 26068 54404 26078
rect 53900 25620 53956 25630
rect 53900 25526 53956 25564
rect 53564 25394 53844 25396
rect 53564 25342 53566 25394
rect 53618 25342 53844 25394
rect 53564 25340 53844 25342
rect 53564 25330 53620 25340
rect 53788 24724 53844 25340
rect 54012 25172 54068 25182
rect 53900 24724 53956 24734
rect 53788 24722 53956 24724
rect 53788 24670 53902 24722
rect 53954 24670 53956 24722
rect 53788 24668 53956 24670
rect 53228 24612 53284 24622
rect 53228 24610 53732 24612
rect 53228 24558 53230 24610
rect 53282 24558 53732 24610
rect 53228 24556 53732 24558
rect 53228 24546 53284 24556
rect 53340 24388 53396 24398
rect 53116 22866 53172 22876
rect 53228 23940 53284 23950
rect 53004 22484 53060 22494
rect 52892 22482 53060 22484
rect 52892 22430 53006 22482
rect 53058 22430 53060 22482
rect 52892 22428 53060 22430
rect 52892 21812 52948 22428
rect 53004 22418 53060 22428
rect 53116 22370 53172 22382
rect 53116 22318 53118 22370
rect 53170 22318 53172 22370
rect 53004 22148 53060 22158
rect 53004 22054 53060 22092
rect 52892 21746 52948 21756
rect 52780 21186 52836 21196
rect 53004 21586 53060 21598
rect 53004 21534 53006 21586
rect 53058 21534 53060 21586
rect 52892 21140 52948 21150
rect 52780 20916 52836 20926
rect 52668 20914 52836 20916
rect 52668 20862 52782 20914
rect 52834 20862 52836 20914
rect 52668 20860 52836 20862
rect 52780 20850 52836 20860
rect 52556 20804 52612 20814
rect 52556 20710 52612 20748
rect 52892 20690 52948 21084
rect 52892 20638 52894 20690
rect 52946 20638 52948 20690
rect 52892 20626 52948 20638
rect 53004 20692 53060 21534
rect 53004 20626 53060 20636
rect 52444 20524 52836 20580
rect 52444 20356 52500 20366
rect 52444 19458 52500 20300
rect 52780 20244 52836 20524
rect 52892 20244 52948 20254
rect 52780 20242 52948 20244
rect 52780 20190 52894 20242
rect 52946 20190 52948 20242
rect 52780 20188 52948 20190
rect 52892 20178 52948 20188
rect 52668 19908 52724 19918
rect 52668 19814 52724 19852
rect 52444 19406 52446 19458
rect 52498 19406 52500 19458
rect 52444 19394 52500 19406
rect 52780 19572 52836 19582
rect 52332 18508 52500 18564
rect 52444 18452 52500 18508
rect 52332 18340 52388 18350
rect 52444 18340 52500 18396
rect 52668 18452 52724 18462
rect 52556 18340 52612 18350
rect 52444 18338 52612 18340
rect 52444 18286 52558 18338
rect 52610 18286 52612 18338
rect 52444 18284 52612 18286
rect 52332 18246 52388 18284
rect 52556 18274 52612 18284
rect 52444 18004 52500 18014
rect 52332 17780 52388 17790
rect 52332 16994 52388 17724
rect 52332 16942 52334 16994
rect 52386 16942 52388 16994
rect 52332 16930 52388 16942
rect 52444 17220 52500 17948
rect 52668 18004 52724 18396
rect 52668 17938 52724 17948
rect 52780 17780 52836 19516
rect 53116 19124 53172 22318
rect 53228 20130 53284 23884
rect 53228 20078 53230 20130
rect 53282 20078 53284 20130
rect 53228 20066 53284 20078
rect 53228 19908 53284 19918
rect 53228 19348 53284 19852
rect 53228 19282 53284 19292
rect 53004 18676 53060 18686
rect 53004 18582 53060 18620
rect 53116 18564 53172 19068
rect 53116 18498 53172 18508
rect 52892 18450 52948 18462
rect 53340 18452 53396 24332
rect 53676 24162 53732 24556
rect 53676 24110 53678 24162
rect 53730 24110 53732 24162
rect 53676 24098 53732 24110
rect 53564 23268 53620 23278
rect 53564 22370 53620 23212
rect 53788 23268 53844 23278
rect 53788 23174 53844 23212
rect 53564 22318 53566 22370
rect 53618 22318 53620 22370
rect 53564 22306 53620 22318
rect 53676 22258 53732 22270
rect 53676 22206 53678 22258
rect 53730 22206 53732 22258
rect 53564 21812 53620 21822
rect 53452 21586 53508 21598
rect 53452 21534 53454 21586
rect 53506 21534 53508 21586
rect 53452 19908 53508 21534
rect 53452 19842 53508 19852
rect 53564 19572 53620 21756
rect 53676 20802 53732 22206
rect 53788 21588 53844 21598
rect 53788 21474 53844 21532
rect 53788 21422 53790 21474
rect 53842 21422 53844 21474
rect 53788 21410 53844 21422
rect 53900 21252 53956 24668
rect 54012 23940 54068 25116
rect 54236 24612 54292 24622
rect 54236 24518 54292 24556
rect 54012 23846 54068 23884
rect 54236 24050 54292 24062
rect 54236 23998 54238 24050
rect 54290 23998 54292 24050
rect 54236 23828 54292 23998
rect 54236 23762 54292 23772
rect 54348 23044 54404 26012
rect 54572 24836 54628 27020
rect 55244 27010 55300 27020
rect 55468 28084 55524 28094
rect 55356 26964 55412 26974
rect 54796 26850 54852 26862
rect 54796 26798 54798 26850
rect 54850 26798 54852 26850
rect 54796 26404 54852 26798
rect 55244 26740 55300 26750
rect 55244 26514 55300 26684
rect 55244 26462 55246 26514
rect 55298 26462 55300 26514
rect 55244 26450 55300 26462
rect 54796 26338 54852 26348
rect 55132 25284 55188 25294
rect 54572 24770 54628 24780
rect 54684 25282 55188 25284
rect 54684 25230 55134 25282
rect 55186 25230 55188 25282
rect 54684 25228 55188 25230
rect 54572 24052 54628 24062
rect 54460 24050 54628 24052
rect 54460 23998 54574 24050
rect 54626 23998 54628 24050
rect 54460 23996 54628 23998
rect 54460 23268 54516 23996
rect 54572 23986 54628 23996
rect 54572 23380 54628 23390
rect 54684 23380 54740 25228
rect 55132 25218 55188 25228
rect 55356 25060 55412 26908
rect 55468 25508 55524 28028
rect 55580 27858 55636 27870
rect 55580 27806 55582 27858
rect 55634 27806 55636 27858
rect 55580 26628 55636 27806
rect 55580 26292 55636 26572
rect 55580 26226 55636 26236
rect 55804 26180 55860 30156
rect 56028 30098 56084 30110
rect 56028 30046 56030 30098
rect 56082 30046 56084 30098
rect 56028 29428 56084 30046
rect 56252 29428 56308 33404
rect 56364 33458 56644 33460
rect 56364 33406 56366 33458
rect 56418 33406 56644 33458
rect 56364 33404 56644 33406
rect 56364 33394 56420 33404
rect 56476 32340 56532 32350
rect 56028 29362 56084 29372
rect 56140 29372 56308 29428
rect 56364 31890 56420 31902
rect 56364 31838 56366 31890
rect 56418 31838 56420 31890
rect 56364 29428 56420 31838
rect 56476 30436 56532 32284
rect 56476 30370 56532 30380
rect 56588 29876 56644 33404
rect 56588 29810 56644 29820
rect 56700 29428 56756 37996
rect 56812 30324 56868 38108
rect 56924 31220 56980 44380
rect 57036 41188 57092 47516
rect 57148 41636 57204 47852
rect 57148 41570 57204 41580
rect 57260 45332 57316 45342
rect 57260 41412 57316 45276
rect 57036 41122 57092 41132
rect 57148 41356 57316 41412
rect 57036 38500 57092 38510
rect 57036 32564 57092 38444
rect 57036 32498 57092 32508
rect 57148 31668 57204 41356
rect 57260 39732 57316 39742
rect 57260 37268 57316 39676
rect 57260 37202 57316 37212
rect 57260 37044 57316 37054
rect 57372 37044 57428 50372
rect 57316 36988 57428 37044
rect 57260 36978 57316 36988
rect 57260 36820 57316 36830
rect 57260 32116 57316 36764
rect 57260 32050 57316 32060
rect 57372 33684 57428 33694
rect 57148 31602 57204 31612
rect 56924 31154 56980 31164
rect 57260 30772 57316 30782
rect 57372 30772 57428 33628
rect 57316 30716 57428 30772
rect 57260 30706 57316 30716
rect 56812 30258 56868 30268
rect 55916 29204 55972 29214
rect 55916 29110 55972 29148
rect 55916 28868 55972 28906
rect 56140 28868 56196 29372
rect 56364 29362 56420 29372
rect 56476 29372 56756 29428
rect 56252 29204 56308 29214
rect 56476 29204 56532 29372
rect 56252 29202 56532 29204
rect 56252 29150 56254 29202
rect 56306 29150 56532 29202
rect 56252 29148 56532 29150
rect 56252 29138 56308 29148
rect 56364 28980 56420 28990
rect 56252 28868 56308 28878
rect 56140 28866 56308 28868
rect 56140 28814 56254 28866
rect 56306 28814 56308 28866
rect 56140 28812 56308 28814
rect 55916 28802 55972 28812
rect 56252 28802 56308 28812
rect 55916 28644 55972 28654
rect 55916 27188 55972 28588
rect 56140 28532 56196 28542
rect 56028 27636 56084 27646
rect 56028 27542 56084 27580
rect 56140 27298 56196 28476
rect 56364 27746 56420 28924
rect 56364 27694 56366 27746
rect 56418 27694 56420 27746
rect 56364 27682 56420 27694
rect 56476 28532 56532 28542
rect 56140 27246 56142 27298
rect 56194 27246 56196 27298
rect 56140 27234 56196 27246
rect 55916 27132 56084 27188
rect 55916 26964 55972 27002
rect 55916 26898 55972 26908
rect 55916 26180 55972 26190
rect 55804 26178 55972 26180
rect 55804 26126 55918 26178
rect 55970 26126 55972 26178
rect 55804 26124 55972 26126
rect 55916 26114 55972 26124
rect 56028 25956 56084 27132
rect 56140 27076 56196 27086
rect 56140 26962 56196 27020
rect 56140 26910 56142 26962
rect 56194 26910 56196 26962
rect 56140 26898 56196 26910
rect 56140 26292 56196 26302
rect 56140 26198 56196 26236
rect 55804 25900 56084 25956
rect 55692 25844 55748 25854
rect 55468 25452 55636 25508
rect 55132 25004 55412 25060
rect 55468 25284 55524 25294
rect 54572 23378 54740 23380
rect 54572 23326 54574 23378
rect 54626 23326 54740 23378
rect 54572 23324 54740 23326
rect 55020 24500 55076 24510
rect 54572 23314 54628 23324
rect 54460 23202 54516 23212
rect 54796 23156 54852 23166
rect 54572 23154 54852 23156
rect 54572 23102 54798 23154
rect 54850 23102 54852 23154
rect 54572 23100 54852 23102
rect 54572 23044 54628 23100
rect 54796 23090 54852 23100
rect 55020 23154 55076 24444
rect 55132 23266 55188 25004
rect 55468 24948 55524 25228
rect 55356 24892 55524 24948
rect 55132 23214 55134 23266
rect 55186 23214 55188 23266
rect 55132 23202 55188 23214
rect 55244 24836 55300 24846
rect 55020 23102 55022 23154
rect 55074 23102 55076 23154
rect 55020 23090 55076 23102
rect 55244 23154 55300 24780
rect 55244 23102 55246 23154
rect 55298 23102 55300 23154
rect 55244 23090 55300 23102
rect 54348 22988 54628 23044
rect 54908 22932 54964 22942
rect 54684 22820 54740 22830
rect 54124 22596 54180 22606
rect 54124 22502 54180 22540
rect 53676 20750 53678 20802
rect 53730 20750 53732 20802
rect 53676 19908 53732 20750
rect 53676 19842 53732 19852
rect 53788 21196 53956 21252
rect 54012 22148 54068 22158
rect 54012 21588 54068 22092
rect 53564 19516 53732 19572
rect 53564 19348 53620 19358
rect 53564 19254 53620 19292
rect 52892 18398 52894 18450
rect 52946 18398 52948 18450
rect 52892 18228 52948 18398
rect 52892 18162 52948 18172
rect 53228 18396 53396 18452
rect 53452 19236 53508 19246
rect 52444 16882 52500 17164
rect 52444 16830 52446 16882
rect 52498 16830 52500 16882
rect 52444 16818 52500 16830
rect 52668 17724 52836 17780
rect 52332 16100 52388 16110
rect 52332 16006 52388 16044
rect 52556 14868 52612 14878
rect 52556 14754 52612 14812
rect 52556 14702 52558 14754
rect 52610 14702 52612 14754
rect 52556 14690 52612 14702
rect 52668 14532 52724 17724
rect 53116 17444 53172 17454
rect 52892 17442 53172 17444
rect 52892 17390 53118 17442
rect 53170 17390 53172 17442
rect 52892 17388 53172 17390
rect 52780 16770 52836 16782
rect 52780 16718 52782 16770
rect 52834 16718 52836 16770
rect 52780 14980 52836 16718
rect 52892 16770 52948 17388
rect 53116 17378 53172 17388
rect 52892 16718 52894 16770
rect 52946 16718 52948 16770
rect 52892 16706 52948 16718
rect 53004 17220 53060 17230
rect 52780 14914 52836 14924
rect 52892 16548 52948 16558
rect 52892 14756 52948 16492
rect 53004 15540 53060 17164
rect 53116 16772 53172 16782
rect 53116 16678 53172 16716
rect 53004 15474 53060 15484
rect 53228 15204 53284 18396
rect 53340 18228 53396 18238
rect 53452 18228 53508 19180
rect 53676 18676 53732 19516
rect 53676 18610 53732 18620
rect 53340 18226 53508 18228
rect 53340 18174 53342 18226
rect 53394 18174 53508 18226
rect 53340 18172 53508 18174
rect 53564 18564 53620 18574
rect 53340 18162 53396 18172
rect 53452 18004 53508 18014
rect 53452 16548 53508 17948
rect 53564 17892 53620 18508
rect 53676 18226 53732 18238
rect 53676 18174 53678 18226
rect 53730 18174 53732 18226
rect 53676 18116 53732 18174
rect 53676 18050 53732 18060
rect 53676 17892 53732 17902
rect 53564 17890 53732 17892
rect 53564 17838 53678 17890
rect 53730 17838 53732 17890
rect 53564 17836 53732 17838
rect 53676 17826 53732 17836
rect 53564 17556 53620 17566
rect 53564 17554 53732 17556
rect 53564 17502 53566 17554
rect 53618 17502 53732 17554
rect 53564 17500 53732 17502
rect 53564 17490 53620 17500
rect 53564 17108 53620 17118
rect 53564 17014 53620 17052
rect 53676 16548 53732 17500
rect 53452 16492 53620 16548
rect 53340 16436 53396 16446
rect 53340 15988 53396 16380
rect 53452 16324 53508 16334
rect 53452 16230 53508 16268
rect 53340 15932 53508 15988
rect 53116 15148 53284 15204
rect 53340 15316 53396 15326
rect 53340 15202 53396 15260
rect 53340 15150 53342 15202
rect 53394 15150 53396 15202
rect 52668 14466 52724 14476
rect 52780 14700 52948 14756
rect 53004 14980 53060 14990
rect 52332 13804 52724 13860
rect 52332 13746 52388 13804
rect 52332 13694 52334 13746
rect 52386 13694 52388 13746
rect 52332 13682 52388 13694
rect 52556 13636 52612 13646
rect 52556 13542 52612 13580
rect 52220 13346 52276 13356
rect 52444 13188 52500 13198
rect 52108 13134 52110 13186
rect 52162 13134 52164 13186
rect 52108 13122 52164 13134
rect 52220 13186 52500 13188
rect 52220 13134 52446 13186
rect 52498 13134 52500 13186
rect 52220 13132 52500 13134
rect 52220 12964 52276 13132
rect 52444 13122 52500 13132
rect 51996 12338 52052 12348
rect 52108 12908 52276 12964
rect 52332 12964 52388 12974
rect 52108 12402 52164 12908
rect 52332 12870 52388 12908
rect 52444 12850 52500 12862
rect 52444 12798 52446 12850
rect 52498 12798 52500 12850
rect 52444 12404 52500 12798
rect 52108 12350 52110 12402
rect 52162 12350 52164 12402
rect 52108 12338 52164 12350
rect 52220 12348 52500 12404
rect 52556 12404 52612 12414
rect 52108 11844 52164 11854
rect 51884 11620 51940 11630
rect 51884 11526 51940 11564
rect 51996 10612 52052 10622
rect 51996 10518 52052 10556
rect 51884 10164 51940 10174
rect 51884 9604 51940 10108
rect 51996 10052 52052 10062
rect 51996 9826 52052 9996
rect 51996 9774 51998 9826
rect 52050 9774 52052 9826
rect 51996 9762 52052 9774
rect 51884 9548 52052 9604
rect 51772 9538 51828 9548
rect 51324 9212 51940 9268
rect 51772 8484 51828 8494
rect 51212 8482 51828 8484
rect 51212 8430 51774 8482
rect 51826 8430 51828 8482
rect 51212 8428 51828 8430
rect 51772 8418 51828 8428
rect 51100 8316 51268 8372
rect 50988 8306 51044 8316
rect 51100 8146 51156 8158
rect 51100 8094 51102 8146
rect 51154 8094 51156 8146
rect 51100 7924 51156 8094
rect 51100 7858 51156 7868
rect 51100 7250 51156 7262
rect 51100 7198 51102 7250
rect 51154 7198 51156 7250
rect 51100 3444 51156 7198
rect 51212 6244 51268 8316
rect 51436 7700 51492 7710
rect 51436 7474 51492 7644
rect 51436 7422 51438 7474
rect 51490 7422 51492 7474
rect 51436 7410 51492 7422
rect 51548 7476 51604 7486
rect 51212 6178 51268 6188
rect 51324 7140 51380 7150
rect 51100 3378 51156 3388
rect 50876 1250 50932 1260
rect 50764 1150 50766 1202
rect 50818 1150 50820 1202
rect 50764 1138 50820 1150
rect 50876 1092 50932 1102
rect 50540 980 50596 990
rect 50540 886 50596 924
rect 50876 112 50932 1036
rect 51324 112 51380 7084
rect 51548 4788 51604 7420
rect 51772 6466 51828 6478
rect 51772 6414 51774 6466
rect 51826 6414 51828 6466
rect 51772 6132 51828 6414
rect 51772 6066 51828 6076
rect 51548 4722 51604 4732
rect 51884 1428 51940 9212
rect 51996 8148 52052 9548
rect 51996 8082 52052 8092
rect 52108 7364 52164 11788
rect 52220 10836 52276 12348
rect 52444 12180 52500 12190
rect 52332 12178 52500 12180
rect 52332 12126 52446 12178
rect 52498 12126 52500 12178
rect 52332 12124 52500 12126
rect 52332 11620 52388 12124
rect 52444 12114 52500 12124
rect 52556 12068 52612 12348
rect 52668 12292 52724 13804
rect 52780 13076 52836 14700
rect 52892 14532 52948 14542
rect 52892 14438 52948 14476
rect 52892 13860 52948 13870
rect 53004 13860 53060 14924
rect 53116 14084 53172 15148
rect 53340 15138 53396 15150
rect 53340 14756 53396 14766
rect 53340 14662 53396 14700
rect 53116 14018 53172 14028
rect 53452 13972 53508 15932
rect 53564 15204 53620 16492
rect 53676 16482 53732 16492
rect 53788 16212 53844 21196
rect 53900 20018 53956 20030
rect 53900 19966 53902 20018
rect 53954 19966 53956 20018
rect 53900 19908 53956 19966
rect 53900 19842 53956 19852
rect 54012 19460 54068 21532
rect 54124 21812 54180 21822
rect 54124 21026 54180 21756
rect 54124 20974 54126 21026
rect 54178 20974 54180 21026
rect 54124 20962 54180 20974
rect 54460 20804 54516 20814
rect 53900 19404 54068 19460
rect 54124 20692 54180 20702
rect 54124 19458 54180 20636
rect 54460 20244 54516 20748
rect 54348 19796 54404 19806
rect 54348 19702 54404 19740
rect 54460 19460 54516 20188
rect 54124 19406 54126 19458
rect 54178 19406 54180 19458
rect 53900 16548 53956 19404
rect 54124 19394 54180 19406
rect 54348 19404 54516 19460
rect 54572 19796 54628 19806
rect 54236 19348 54292 19358
rect 54236 19254 54292 19292
rect 54012 19234 54068 19246
rect 54012 19182 54014 19234
rect 54066 19182 54068 19234
rect 54012 18228 54068 19182
rect 54012 18162 54068 18172
rect 54124 18450 54180 18462
rect 54124 18398 54126 18450
rect 54178 18398 54180 18450
rect 54012 17554 54068 17566
rect 54012 17502 54014 17554
rect 54066 17502 54068 17554
rect 54012 17108 54068 17502
rect 54124 17332 54180 18398
rect 54124 17266 54180 17276
rect 54236 17668 54292 17678
rect 54348 17668 54404 19404
rect 54460 19236 54516 19246
rect 54460 19142 54516 19180
rect 54236 17666 54404 17668
rect 54236 17614 54238 17666
rect 54290 17614 54404 17666
rect 54236 17612 54404 17614
rect 54460 18228 54516 18238
rect 54012 17042 54068 17052
rect 54236 16772 54292 17612
rect 54236 16706 54292 16716
rect 54348 17442 54404 17454
rect 54348 17390 54350 17442
rect 54402 17390 54404 17442
rect 54348 16548 54404 17390
rect 53900 16492 54404 16548
rect 53788 16156 54068 16212
rect 53900 15986 53956 15998
rect 53900 15934 53902 15986
rect 53954 15934 53956 15986
rect 53676 15540 53732 15550
rect 53900 15540 53956 15934
rect 54012 15652 54068 16156
rect 54348 15876 54404 16492
rect 54348 15810 54404 15820
rect 54012 15596 54404 15652
rect 53732 15484 53956 15540
rect 53676 15426 53732 15484
rect 53676 15374 53678 15426
rect 53730 15374 53732 15426
rect 53676 15362 53732 15374
rect 53564 15138 53620 15148
rect 53788 14420 53844 14430
rect 53228 13916 53508 13972
rect 53676 14084 53732 14094
rect 52892 13858 53060 13860
rect 52892 13806 52894 13858
rect 52946 13806 53060 13858
rect 52892 13804 53060 13806
rect 53116 13860 53172 13870
rect 52892 13794 52948 13804
rect 53004 13636 53060 13646
rect 53004 13186 53060 13580
rect 53004 13134 53006 13186
rect 53058 13134 53060 13186
rect 53004 13122 53060 13134
rect 52892 13076 52948 13086
rect 52780 13074 52948 13076
rect 52780 13022 52894 13074
rect 52946 13022 52948 13074
rect 52780 13020 52948 13022
rect 52892 13010 52948 13020
rect 53116 12404 53172 13804
rect 53228 13186 53284 13916
rect 53452 13524 53508 13534
rect 53452 13430 53508 13468
rect 53228 13134 53230 13186
rect 53282 13134 53284 13186
rect 53228 13122 53284 13134
rect 53340 12852 53396 12862
rect 53116 12348 53284 12404
rect 52668 12236 53172 12292
rect 52668 12068 52724 12078
rect 52556 12066 52724 12068
rect 52556 12014 52670 12066
rect 52722 12014 52724 12066
rect 52556 12012 52724 12014
rect 52668 12002 52724 12012
rect 53004 12066 53060 12078
rect 53004 12014 53006 12066
rect 53058 12014 53060 12066
rect 52332 11554 52388 11564
rect 52444 11844 52500 11854
rect 52444 11618 52500 11788
rect 53004 11844 53060 12014
rect 53004 11778 53060 11788
rect 52444 11566 52446 11618
rect 52498 11566 52500 11618
rect 52444 11554 52500 11566
rect 52556 11620 52612 11630
rect 53116 11620 53172 12236
rect 52332 10836 52388 10846
rect 52220 10834 52388 10836
rect 52220 10782 52334 10834
rect 52386 10782 52388 10834
rect 52220 10780 52388 10782
rect 52332 10770 52388 10780
rect 52220 10388 52276 10398
rect 52220 10294 52276 10332
rect 52220 9828 52276 9838
rect 52556 9828 52612 11564
rect 52668 11564 53172 11620
rect 52668 10834 52724 11564
rect 53228 11508 53284 12348
rect 52668 10782 52670 10834
rect 52722 10782 52724 10834
rect 52668 10770 52724 10782
rect 52780 11452 53284 11508
rect 52780 10722 52836 11452
rect 53116 11284 53172 11294
rect 52780 10670 52782 10722
rect 52834 10670 52836 10722
rect 52780 10658 52836 10670
rect 53004 11060 53060 11070
rect 52892 10612 52948 10622
rect 52220 8820 52276 9772
rect 52444 9772 52612 9828
rect 52668 10500 52724 10510
rect 52668 9826 52724 10444
rect 52668 9774 52670 9826
rect 52722 9774 52724 9826
rect 52332 9156 52388 9166
rect 52332 8930 52388 9100
rect 52332 8878 52334 8930
rect 52386 8878 52388 8930
rect 52332 8866 52388 8878
rect 52220 8754 52276 8764
rect 52332 8148 52388 8158
rect 52220 7924 52276 7934
rect 52220 7586 52276 7868
rect 52220 7534 52222 7586
rect 52274 7534 52276 7586
rect 52220 7522 52276 7534
rect 52108 7308 52276 7364
rect 52108 6244 52164 6254
rect 52108 6130 52164 6188
rect 52108 6078 52110 6130
rect 52162 6078 52164 6130
rect 52108 6066 52164 6078
rect 51884 1362 51940 1372
rect 52108 2996 52164 3006
rect 51772 756 51828 766
rect 51772 112 51828 700
rect 52108 756 52164 2940
rect 52108 690 52164 700
rect 52220 112 52276 7308
rect 52332 4116 52388 8092
rect 52444 6356 52500 9772
rect 52668 9762 52724 9774
rect 52780 9938 52836 9950
rect 52780 9886 52782 9938
rect 52834 9886 52836 9938
rect 52556 9604 52612 9614
rect 52556 7588 52612 9548
rect 52668 9044 52724 9054
rect 52668 8950 52724 8988
rect 52668 8820 52724 8830
rect 52668 8036 52724 8764
rect 52780 8484 52836 9886
rect 52892 9380 52948 10556
rect 52892 9314 52948 9324
rect 52780 8418 52836 8428
rect 52892 8370 52948 8382
rect 52892 8318 52894 8370
rect 52946 8318 52948 8370
rect 52892 8260 52948 8318
rect 52892 8194 52948 8204
rect 52668 7980 52948 8036
rect 52556 7532 52724 7588
rect 52556 7364 52612 7374
rect 52556 7270 52612 7308
rect 52444 6300 52612 6356
rect 52444 6132 52500 6142
rect 52444 6038 52500 6076
rect 52556 5236 52612 6300
rect 52668 6132 52724 7532
rect 52668 6066 52724 6076
rect 52780 6802 52836 6814
rect 52780 6750 52782 6802
rect 52834 6750 52836 6802
rect 52556 5170 52612 5180
rect 52332 4050 52388 4060
rect 52556 4788 52612 4798
rect 52556 868 52612 4732
rect 52668 4564 52724 4574
rect 52668 1092 52724 4508
rect 52668 1026 52724 1036
rect 52780 868 52836 6750
rect 52892 5906 52948 7980
rect 53004 7700 53060 11004
rect 53004 7634 53060 7644
rect 53116 6914 53172 11228
rect 53228 9042 53284 9054
rect 53228 8990 53230 9042
rect 53282 8990 53284 9042
rect 53228 8820 53284 8990
rect 53340 9044 53396 12796
rect 53564 12738 53620 12750
rect 53564 12686 53566 12738
rect 53618 12686 53620 12738
rect 53452 12180 53508 12190
rect 53452 10610 53508 12124
rect 53564 12068 53620 12686
rect 53564 12002 53620 12012
rect 53676 11732 53732 14028
rect 53564 11676 53732 11732
rect 53564 11620 53620 11676
rect 53564 11554 53620 11564
rect 53676 11506 53732 11518
rect 53676 11454 53678 11506
rect 53730 11454 53732 11506
rect 53452 10558 53454 10610
rect 53506 10558 53508 10610
rect 53452 10052 53508 10558
rect 53452 9986 53508 9996
rect 53564 10948 53620 10958
rect 53340 8978 53396 8988
rect 53452 9156 53508 9166
rect 53564 9156 53620 10892
rect 53676 10612 53732 11454
rect 53788 10948 53844 14364
rect 53900 11396 53956 15484
rect 54348 15148 54404 15596
rect 54236 15092 54404 15148
rect 54124 13300 54180 13310
rect 54012 12180 54068 12190
rect 54012 12086 54068 12124
rect 54012 11396 54068 11406
rect 53900 11394 54068 11396
rect 53900 11342 54014 11394
rect 54066 11342 54068 11394
rect 53900 11340 54068 11342
rect 54012 11330 54068 11340
rect 53788 10882 53844 10892
rect 53676 10546 53732 10556
rect 53788 10724 53844 10734
rect 53788 10498 53844 10668
rect 53788 10446 53790 10498
rect 53842 10446 53844 10498
rect 53788 10434 53844 10446
rect 53676 10052 53732 10062
rect 53676 9716 53732 9996
rect 54012 9940 54068 9950
rect 54012 9846 54068 9884
rect 53676 9714 53844 9716
rect 53676 9662 53678 9714
rect 53730 9662 53844 9714
rect 53676 9660 53844 9662
rect 53676 9650 53732 9660
rect 53564 9100 53732 9156
rect 53228 8754 53284 8764
rect 53340 8146 53396 8158
rect 53340 8094 53342 8146
rect 53394 8094 53396 8146
rect 53340 7924 53396 8094
rect 53340 7700 53396 7868
rect 53340 7634 53396 7644
rect 53116 6862 53118 6914
rect 53170 6862 53172 6914
rect 53116 6850 53172 6862
rect 53228 7252 53284 7262
rect 52892 5854 52894 5906
rect 52946 5854 52948 5906
rect 52892 5842 52948 5854
rect 53116 5906 53172 5918
rect 53116 5854 53118 5906
rect 53170 5854 53172 5906
rect 53116 5124 53172 5854
rect 53228 5794 53284 7196
rect 53228 5742 53230 5794
rect 53282 5742 53284 5794
rect 53228 5730 53284 5742
rect 53340 6580 53396 6590
rect 53340 5346 53396 6524
rect 53452 6356 53508 9100
rect 53564 8932 53620 8942
rect 53564 8838 53620 8876
rect 53676 7924 53732 9100
rect 53788 8820 53844 9660
rect 54124 9268 54180 13244
rect 54124 9202 54180 9212
rect 53788 8754 53844 8764
rect 53676 7858 53732 7868
rect 53900 8484 53956 8494
rect 53564 7588 53620 7598
rect 53564 6692 53620 7532
rect 53788 7252 53844 7262
rect 53788 7158 53844 7196
rect 53564 6626 53620 6636
rect 53676 6580 53732 6590
rect 53676 6486 53732 6524
rect 53452 6300 53732 6356
rect 53340 5294 53342 5346
rect 53394 5294 53396 5346
rect 53340 5282 53396 5294
rect 53564 6020 53620 6030
rect 53116 5058 53172 5068
rect 53564 4340 53620 5964
rect 53676 5346 53732 6300
rect 53788 6132 53844 6142
rect 53900 6132 53956 8428
rect 54124 8372 54180 8382
rect 54124 8278 54180 8316
rect 54124 6916 54180 6926
rect 54124 6822 54180 6860
rect 53788 6130 53956 6132
rect 53788 6078 53790 6130
rect 53842 6078 53956 6130
rect 53788 6076 53956 6078
rect 53788 6066 53844 6076
rect 53676 5294 53678 5346
rect 53730 5294 53732 5346
rect 53676 5282 53732 5294
rect 54124 5906 54180 5918
rect 54124 5854 54126 5906
rect 54178 5854 54180 5906
rect 54124 5346 54180 5854
rect 54236 5572 54292 15092
rect 54460 14868 54516 18172
rect 54572 16324 54628 19740
rect 54684 19460 54740 22764
rect 54684 19394 54740 19404
rect 54684 19234 54740 19246
rect 54684 19182 54686 19234
rect 54738 19182 54740 19234
rect 54684 18452 54740 19182
rect 54684 18386 54740 18396
rect 54796 18340 54852 18350
rect 54684 18226 54740 18238
rect 54684 18174 54686 18226
rect 54738 18174 54740 18226
rect 54684 17556 54740 18174
rect 54684 17490 54740 17500
rect 54796 17442 54852 18284
rect 54908 18228 54964 22876
rect 55244 22148 55300 22158
rect 55244 22054 55300 22092
rect 55356 22036 55412 24892
rect 55468 24500 55524 24510
rect 55468 24406 55524 24444
rect 55356 21970 55412 21980
rect 55468 21588 55524 21598
rect 55244 21586 55524 21588
rect 55244 21534 55470 21586
rect 55522 21534 55524 21586
rect 55244 21532 55524 21534
rect 55020 21364 55076 21374
rect 55020 21362 55188 21364
rect 55020 21310 55022 21362
rect 55074 21310 55188 21362
rect 55020 21308 55188 21310
rect 55020 21298 55076 21308
rect 55020 20244 55076 20254
rect 55020 19458 55076 20188
rect 55020 19406 55022 19458
rect 55074 19406 55076 19458
rect 55020 19394 55076 19406
rect 54908 18172 55076 18228
rect 55020 17892 55076 18172
rect 55132 18004 55188 21308
rect 55244 21026 55300 21532
rect 55468 21522 55524 21532
rect 55244 20974 55246 21026
rect 55298 20974 55300 21026
rect 55244 20962 55300 20974
rect 55580 21028 55636 25452
rect 55692 21924 55748 25788
rect 55804 24164 55860 25900
rect 56252 25620 56308 25630
rect 56028 25618 56308 25620
rect 56028 25566 56254 25618
rect 56306 25566 56308 25618
rect 56028 25564 56308 25566
rect 55916 25506 55972 25518
rect 55916 25454 55918 25506
rect 55970 25454 55972 25506
rect 55916 25396 55972 25454
rect 55916 25330 55972 25340
rect 55916 24164 55972 24174
rect 55804 24162 55972 24164
rect 55804 24110 55918 24162
rect 55970 24110 55972 24162
rect 55804 24108 55972 24110
rect 55916 24098 55972 24108
rect 55916 23492 55972 23502
rect 55916 23154 55972 23436
rect 55916 23102 55918 23154
rect 55970 23102 55972 23154
rect 55916 23090 55972 23102
rect 56028 22596 56084 25564
rect 56252 25554 56308 25564
rect 56140 24722 56196 24734
rect 56140 24670 56142 24722
rect 56194 24670 56196 24722
rect 56140 23044 56196 24670
rect 56364 24612 56420 24622
rect 56476 24612 56532 28476
rect 57148 27636 57204 27646
rect 57036 27188 57092 27198
rect 56364 24610 56532 24612
rect 56364 24558 56366 24610
rect 56418 24558 56532 24610
rect 56364 24556 56532 24558
rect 56588 26740 56644 26750
rect 56364 24546 56420 24556
rect 56588 24388 56644 26684
rect 56924 26292 56980 26302
rect 56364 24332 56644 24388
rect 56812 24948 56868 24958
rect 56252 24050 56308 24062
rect 56252 23998 56254 24050
rect 56306 23998 56308 24050
rect 56252 23268 56308 23998
rect 56252 23202 56308 23212
rect 56252 23044 56308 23054
rect 56140 23042 56308 23044
rect 56140 22990 56254 23042
rect 56306 22990 56308 23042
rect 56140 22988 56308 22990
rect 56252 22978 56308 22988
rect 56364 22820 56420 24332
rect 55692 21858 55748 21868
rect 55804 22540 56084 22596
rect 56252 22764 56420 22820
rect 56588 23940 56644 23950
rect 56252 22594 56308 22764
rect 56252 22542 56254 22594
rect 56306 22542 56308 22594
rect 55692 21700 55748 21738
rect 55692 21634 55748 21644
rect 55580 20962 55636 20972
rect 55692 21252 55748 21262
rect 55356 20244 55412 20254
rect 55356 19460 55412 20188
rect 55468 19796 55524 19806
rect 55468 19702 55524 19740
rect 55356 19404 55524 19460
rect 55244 19346 55300 19358
rect 55244 19294 55246 19346
rect 55298 19294 55300 19346
rect 55244 18228 55300 19294
rect 55356 19234 55412 19246
rect 55356 19182 55358 19234
rect 55410 19182 55412 19234
rect 55356 19124 55412 19182
rect 55356 19058 55412 19068
rect 55468 18900 55524 19404
rect 55244 18162 55300 18172
rect 55356 18844 55524 18900
rect 55132 17948 55300 18004
rect 55020 17836 55188 17892
rect 54908 17780 54964 17790
rect 54908 17686 54964 17724
rect 55020 17668 55076 17678
rect 55020 17574 55076 17612
rect 55132 17444 55188 17836
rect 54796 17390 54798 17442
rect 54850 17390 54852 17442
rect 54796 17378 54852 17390
rect 55020 17388 55188 17444
rect 54684 16996 54740 17006
rect 54684 16770 54740 16940
rect 54684 16718 54686 16770
rect 54738 16718 54740 16770
rect 54684 16706 54740 16718
rect 54908 16772 54964 16782
rect 54796 16324 54852 16334
rect 54572 16322 54852 16324
rect 54572 16270 54798 16322
rect 54850 16270 54852 16322
rect 54572 16268 54852 16270
rect 54796 16258 54852 16268
rect 54572 16098 54628 16110
rect 54572 16046 54574 16098
rect 54626 16046 54628 16098
rect 54572 15876 54628 16046
rect 54684 16100 54740 16110
rect 54684 16006 54740 16044
rect 54908 16098 54964 16716
rect 55020 16324 55076 17388
rect 55132 17220 55188 17230
rect 55132 16994 55188 17164
rect 55132 16942 55134 16994
rect 55186 16942 55188 16994
rect 55132 16930 55188 16942
rect 55020 16258 55076 16268
rect 55132 16660 55188 16670
rect 54908 16046 54910 16098
rect 54962 16046 54964 16098
rect 54908 16034 54964 16046
rect 54572 15810 54628 15820
rect 54572 15540 54628 15550
rect 54572 15428 54628 15484
rect 54572 15426 54852 15428
rect 54572 15374 54574 15426
rect 54626 15374 54852 15426
rect 54572 15372 54852 15374
rect 54572 15362 54628 15372
rect 54348 14812 54516 14868
rect 54348 13636 54404 14812
rect 54460 14644 54516 14654
rect 54460 14550 54516 14588
rect 54796 14532 54852 15372
rect 54908 15204 54964 15214
rect 54908 15110 54964 15148
rect 54908 14532 54964 14542
rect 54796 14530 54964 14532
rect 54796 14478 54910 14530
rect 54962 14478 54964 14530
rect 54796 14476 54964 14478
rect 54908 14466 54964 14476
rect 54348 13570 54404 13580
rect 54572 14196 54628 14206
rect 54572 13634 54628 14140
rect 54572 13582 54574 13634
rect 54626 13582 54628 13634
rect 54572 13570 54628 13582
rect 55020 13746 55076 13758
rect 55020 13694 55022 13746
rect 55074 13694 55076 13746
rect 54908 13300 54964 13310
rect 54684 13188 54740 13198
rect 54684 13094 54740 13132
rect 54460 12068 54516 12078
rect 54460 11974 54516 12012
rect 54460 10388 54516 10398
rect 54348 8820 54404 8830
rect 54348 7476 54404 8764
rect 54460 8258 54516 10332
rect 54796 8820 54852 8830
rect 54460 8206 54462 8258
rect 54514 8206 54516 8258
rect 54460 8194 54516 8206
rect 54572 8818 54852 8820
rect 54572 8766 54798 8818
rect 54850 8766 54852 8818
rect 54572 8764 54852 8766
rect 54460 7476 54516 7486
rect 54348 7474 54516 7476
rect 54348 7422 54462 7474
rect 54514 7422 54516 7474
rect 54348 7420 54516 7422
rect 54460 6468 54516 7420
rect 54460 6402 54516 6412
rect 54348 6356 54404 6366
rect 54348 5794 54404 6300
rect 54348 5742 54350 5794
rect 54402 5742 54404 5794
rect 54348 5730 54404 5742
rect 54236 5516 54404 5572
rect 54124 5294 54126 5346
rect 54178 5294 54180 5346
rect 54124 5282 54180 5294
rect 53564 4274 53620 4284
rect 53564 4116 53620 4126
rect 52556 812 52724 868
rect 52668 112 52724 812
rect 52780 802 52836 812
rect 53116 3108 53172 3118
rect 53116 112 53172 3052
rect 53564 112 53620 4060
rect 54124 4116 54180 4126
rect 54124 4114 54292 4116
rect 54124 4062 54126 4114
rect 54178 4062 54292 4114
rect 54124 4060 54292 4062
rect 54124 4050 54180 4060
rect 54012 3780 54068 3790
rect 54012 112 54068 3724
rect 54236 196 54292 4060
rect 54348 1540 54404 5516
rect 54460 5012 54516 5022
rect 54572 5012 54628 8764
rect 54796 8754 54852 8764
rect 54908 8484 54964 13244
rect 55020 12852 55076 13694
rect 55132 13524 55188 16604
rect 55244 16098 55300 17948
rect 55356 17892 55412 18844
rect 55692 18452 55748 21196
rect 55804 21028 55860 22540
rect 56252 22530 56308 22542
rect 56588 22484 56644 23884
rect 56812 23940 56868 24892
rect 56812 23874 56868 23884
rect 56476 22428 56644 22484
rect 56700 23828 56756 23838
rect 56028 22372 56084 22382
rect 56028 22370 56196 22372
rect 56028 22318 56030 22370
rect 56082 22318 56196 22370
rect 56028 22316 56196 22318
rect 56028 22306 56084 22316
rect 56028 22148 56084 22158
rect 55916 21588 55972 21598
rect 56028 21588 56084 22092
rect 55916 21586 56084 21588
rect 55916 21534 55918 21586
rect 55970 21534 56084 21586
rect 55916 21532 56084 21534
rect 56140 21588 56196 22316
rect 56140 21532 56308 21588
rect 55916 21522 55972 21532
rect 56028 21364 56084 21374
rect 56028 21270 56084 21308
rect 56140 21362 56196 21374
rect 56140 21310 56142 21362
rect 56194 21310 56196 21362
rect 56028 21028 56084 21038
rect 55804 21026 56084 21028
rect 55804 20974 56030 21026
rect 56082 20974 56084 21026
rect 55804 20972 56084 20974
rect 56028 20962 56084 20972
rect 56140 20244 56196 21310
rect 56140 20178 56196 20188
rect 56252 19906 56308 21532
rect 56364 21028 56420 21038
rect 56364 20934 56420 20972
rect 56252 19854 56254 19906
rect 56306 19854 56308 19906
rect 56252 19842 56308 19854
rect 55916 19794 55972 19806
rect 55916 19742 55918 19794
rect 55970 19742 55972 19794
rect 55916 19684 55972 19742
rect 55916 19618 55972 19628
rect 56028 19460 56084 19470
rect 56028 19366 56084 19404
rect 56364 19460 56420 19470
rect 56364 19366 56420 19404
rect 56252 19236 56308 19246
rect 55692 18396 56084 18452
rect 55356 17826 55412 17836
rect 55468 18228 55524 18238
rect 55244 16046 55246 16098
rect 55298 16046 55300 16098
rect 55244 16034 55300 16046
rect 55356 17666 55412 17678
rect 55356 17614 55358 17666
rect 55410 17614 55412 17666
rect 55132 13458 55188 13468
rect 55244 15764 55300 15774
rect 55132 12852 55188 12862
rect 55020 12850 55188 12852
rect 55020 12798 55134 12850
rect 55186 12798 55188 12850
rect 55020 12796 55188 12798
rect 55132 12180 55188 12796
rect 55132 12114 55188 12124
rect 55132 11956 55188 11966
rect 55020 11732 55076 11742
rect 55020 11618 55076 11676
rect 55020 11566 55022 11618
rect 55074 11566 55076 11618
rect 55020 11554 55076 11566
rect 55020 10388 55076 10398
rect 55020 10294 55076 10332
rect 55132 10164 55188 11900
rect 54460 5010 54628 5012
rect 54460 4958 54462 5010
rect 54514 4958 54628 5010
rect 54460 4956 54628 4958
rect 54684 8428 54964 8484
rect 55020 10108 55188 10164
rect 54460 4946 54516 4956
rect 54684 4788 54740 8428
rect 55020 8370 55076 10108
rect 55244 9828 55300 15708
rect 55356 15540 55412 17614
rect 55356 15474 55412 15484
rect 55356 11506 55412 11518
rect 55356 11454 55358 11506
rect 55410 11454 55412 11506
rect 55356 10612 55412 11454
rect 55356 10546 55412 10556
rect 55132 9772 55300 9828
rect 55132 8932 55188 9772
rect 55244 9604 55300 9614
rect 55244 9602 55412 9604
rect 55244 9550 55246 9602
rect 55298 9550 55412 9602
rect 55244 9548 55412 9550
rect 55244 9538 55300 9548
rect 55244 8932 55300 8942
rect 55132 8930 55300 8932
rect 55132 8878 55246 8930
rect 55298 8878 55300 8930
rect 55132 8876 55300 8878
rect 55244 8866 55300 8876
rect 55020 8318 55022 8370
rect 55074 8318 55076 8370
rect 55020 8306 55076 8318
rect 54908 8258 54964 8270
rect 54908 8206 54910 8258
rect 54962 8206 54964 8258
rect 54908 8148 54964 8206
rect 54908 8092 55076 8148
rect 54796 8036 54852 8046
rect 54796 7362 54852 7980
rect 54796 7310 54798 7362
rect 54850 7310 54852 7362
rect 54796 7298 54852 7310
rect 54908 5796 54964 5806
rect 54908 5702 54964 5740
rect 54460 4732 54740 4788
rect 54908 5124 54964 5134
rect 55020 5124 55076 8092
rect 55356 6692 55412 9548
rect 55468 9042 55524 18172
rect 55804 18226 55860 18238
rect 55804 18174 55806 18226
rect 55858 18174 55860 18226
rect 55692 18004 55748 18014
rect 55692 16882 55748 17948
rect 55804 17780 55860 18174
rect 55804 17714 55860 17724
rect 55692 16830 55694 16882
rect 55746 16830 55748 16882
rect 55692 16818 55748 16830
rect 55804 17332 55860 17342
rect 55580 14868 55636 14878
rect 55580 13970 55636 14812
rect 55580 13918 55582 13970
rect 55634 13918 55636 13970
rect 55580 13906 55636 13918
rect 55692 13972 55748 13982
rect 55692 13858 55748 13916
rect 55692 13806 55694 13858
rect 55746 13806 55748 13858
rect 55692 13794 55748 13806
rect 55692 12404 55748 12414
rect 55580 11956 55636 11966
rect 55580 11862 55636 11900
rect 55692 11732 55748 12348
rect 55468 8990 55470 9042
rect 55522 8990 55524 9042
rect 55468 8978 55524 8990
rect 55580 11676 55748 11732
rect 54964 5068 55076 5124
rect 55132 6636 55412 6692
rect 55468 8596 55524 8606
rect 54460 4338 54516 4732
rect 54460 4286 54462 4338
rect 54514 4286 54516 4338
rect 54460 4274 54516 4286
rect 54908 4338 54964 5068
rect 54908 4286 54910 4338
rect 54962 4286 54964 4338
rect 54908 4274 54964 4286
rect 55020 4676 55076 4686
rect 55020 3778 55076 4620
rect 55132 4226 55188 6636
rect 55468 6580 55524 8540
rect 55468 6514 55524 6524
rect 55244 6466 55300 6478
rect 55244 6414 55246 6466
rect 55298 6414 55300 6466
rect 55244 5234 55300 6414
rect 55468 5682 55524 5694
rect 55468 5630 55470 5682
rect 55522 5630 55524 5682
rect 55468 5348 55524 5630
rect 55468 5282 55524 5292
rect 55244 5182 55246 5234
rect 55298 5182 55300 5234
rect 55244 5170 55300 5182
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 4162 55188 4174
rect 55020 3726 55022 3778
rect 55074 3726 55076 3778
rect 55020 3714 55076 3726
rect 55356 3780 55412 3790
rect 55356 3686 55412 3724
rect 54348 1474 54404 1484
rect 54908 3668 54964 3678
rect 54236 130 54292 140
rect 54460 1428 54516 1438
rect 54460 112 54516 1372
rect 54908 112 54964 3612
rect 55580 2770 55636 11676
rect 55804 5906 55860 17276
rect 56028 16884 56084 18396
rect 56252 18450 56308 19180
rect 56252 18398 56254 18450
rect 56306 18398 56308 18450
rect 56252 18386 56308 18398
rect 56364 18340 56420 18350
rect 56364 18246 56420 18284
rect 56364 17892 56420 17902
rect 56364 17798 56420 17836
rect 56140 17668 56196 17678
rect 56140 17666 56308 17668
rect 56140 17614 56142 17666
rect 56194 17614 56308 17666
rect 56140 17612 56308 17614
rect 56140 17602 56196 17612
rect 56028 16828 56196 16884
rect 56028 16660 56084 16670
rect 55916 16658 56084 16660
rect 55916 16606 56030 16658
rect 56082 16606 56084 16658
rect 55916 16604 56084 16606
rect 55916 13300 55972 16604
rect 56028 16594 56084 16604
rect 56028 16324 56084 16334
rect 56028 16230 56084 16268
rect 56028 16100 56084 16110
rect 56028 15316 56084 16044
rect 56140 15876 56196 16828
rect 56252 16212 56308 17612
rect 56364 16324 56420 16334
rect 56364 16230 56420 16268
rect 56252 16146 56308 16156
rect 56140 15820 56420 15876
rect 56140 15540 56196 15550
rect 56140 15446 56196 15484
rect 56028 15260 56308 15316
rect 56028 14756 56084 14766
rect 56028 14662 56084 14700
rect 56140 14308 56196 14318
rect 56140 13746 56196 14252
rect 56140 13694 56142 13746
rect 56194 13694 56196 13746
rect 56140 13682 56196 13694
rect 56140 13524 56196 13534
rect 55916 13244 56084 13300
rect 55916 12962 55972 12974
rect 55916 12910 55918 12962
rect 55970 12910 55972 12962
rect 55916 12292 55972 12910
rect 55916 12226 55972 12236
rect 56028 12178 56084 13244
rect 56028 12126 56030 12178
rect 56082 12126 56084 12178
rect 56028 12114 56084 12126
rect 56028 11394 56084 11406
rect 56028 11342 56030 11394
rect 56082 11342 56084 11394
rect 56028 11172 56084 11342
rect 56028 11106 56084 11116
rect 56028 10612 56084 10622
rect 56028 10518 56084 10556
rect 56140 10388 56196 13468
rect 56252 13186 56308 15260
rect 56364 14754 56420 15820
rect 56364 14702 56366 14754
rect 56418 14702 56420 14754
rect 56364 14690 56420 14702
rect 56364 14420 56420 14430
rect 56364 13634 56420 14364
rect 56364 13582 56366 13634
rect 56418 13582 56420 13634
rect 56364 13570 56420 13582
rect 56252 13134 56254 13186
rect 56306 13134 56308 13186
rect 56252 13122 56308 13134
rect 56364 12068 56420 12078
rect 56476 12068 56532 22428
rect 56700 21868 56756 23772
rect 56588 21812 56756 21868
rect 56812 23268 56868 23278
rect 56588 14532 56644 21812
rect 56700 19236 56756 19246
rect 56700 16324 56756 19180
rect 56700 16258 56756 16268
rect 56588 14466 56644 14476
rect 56812 14308 56868 23212
rect 56924 19348 56980 26236
rect 56924 19282 56980 19292
rect 56812 14242 56868 14252
rect 56924 19124 56980 19134
rect 56364 12066 56532 12068
rect 56364 12014 56366 12066
rect 56418 12014 56532 12066
rect 56364 12012 56532 12014
rect 56588 13076 56644 13086
rect 56364 12002 56420 12012
rect 56140 10322 56196 10332
rect 56252 11956 56308 11966
rect 56140 9828 56196 9838
rect 56028 9826 56196 9828
rect 56028 9774 56142 9826
rect 56194 9774 56196 9826
rect 56028 9772 56196 9774
rect 55916 9716 55972 9726
rect 55916 8932 55972 9660
rect 56028 9156 56084 9772
rect 56140 9762 56196 9772
rect 56028 9090 56084 9100
rect 56028 8932 56084 8942
rect 55916 8930 56084 8932
rect 55916 8878 56030 8930
rect 56082 8878 56084 8930
rect 55916 8876 56084 8878
rect 56028 8866 56084 8876
rect 56252 8820 56308 11900
rect 56364 11620 56420 11630
rect 56364 11526 56420 11564
rect 56364 10500 56420 10510
rect 56364 10406 56420 10444
rect 56364 10052 56420 10062
rect 56364 9958 56420 9996
rect 56364 9044 56420 9054
rect 56364 8930 56420 8988
rect 56364 8878 56366 8930
rect 56418 8878 56420 8930
rect 56364 8866 56420 8878
rect 56140 8764 56308 8820
rect 56028 8370 56084 8382
rect 56028 8318 56030 8370
rect 56082 8318 56084 8370
rect 56028 7812 56084 8318
rect 56028 7746 56084 7756
rect 56028 7250 56084 7262
rect 56028 7198 56030 7250
rect 56082 7198 56084 7250
rect 55916 6802 55972 6814
rect 55916 6750 55918 6802
rect 55970 6750 55972 6802
rect 55916 6692 55972 6750
rect 55916 6626 55972 6636
rect 55804 5854 55806 5906
rect 55858 5854 55860 5906
rect 55804 5842 55860 5854
rect 55916 5234 55972 5246
rect 55916 5182 55918 5234
rect 55970 5182 55972 5234
rect 55916 5012 55972 5182
rect 55916 4946 55972 4956
rect 55692 4564 55748 4574
rect 56028 4564 56084 7198
rect 56140 6692 56196 8764
rect 56588 8708 56644 13020
rect 56252 8652 56644 8708
rect 56252 7140 56308 8652
rect 56364 8484 56420 8494
rect 56924 8484 56980 19068
rect 57036 17892 57092 27132
rect 57148 19460 57204 27580
rect 57260 25396 57316 25406
rect 57260 23828 57316 25340
rect 57260 23762 57316 23772
rect 57260 22708 57316 22718
rect 57316 22652 57428 22708
rect 57260 22642 57316 22652
rect 57148 19394 57204 19404
rect 57036 17826 57092 17836
rect 57148 17780 57204 17790
rect 56364 8482 56980 8484
rect 56364 8430 56366 8482
rect 56418 8430 56980 8482
rect 56364 8428 56980 8430
rect 57036 14644 57092 14654
rect 56364 8418 56420 8428
rect 56252 7074 56308 7084
rect 56364 8260 56420 8270
rect 57036 8260 57092 14588
rect 56252 6916 56308 6926
rect 56364 6916 56420 8204
rect 56252 6914 56420 6916
rect 56252 6862 56254 6914
rect 56306 6862 56420 6914
rect 56252 6860 56420 6862
rect 56476 8204 57092 8260
rect 57148 8260 57204 17724
rect 56252 6850 56308 6860
rect 56140 6636 56420 6692
rect 56252 6468 56308 6478
rect 55692 4562 56084 4564
rect 55692 4510 55694 4562
rect 55746 4510 56084 4562
rect 55692 4508 56084 4510
rect 56140 5796 56196 5806
rect 55692 4498 55748 4508
rect 56028 4340 56084 4350
rect 56140 4340 56196 5740
rect 56252 5124 56308 6412
rect 56252 5030 56308 5068
rect 56364 4900 56420 6636
rect 56028 4338 56196 4340
rect 56028 4286 56030 4338
rect 56082 4286 56196 4338
rect 56028 4284 56196 4286
rect 56252 4844 56420 4900
rect 56028 4274 56084 4284
rect 55916 4228 55972 4238
rect 55916 3780 55972 4172
rect 56028 3780 56084 3790
rect 55916 3778 56084 3780
rect 55916 3726 56030 3778
rect 56082 3726 56084 3778
rect 55916 3724 56084 3726
rect 56028 3714 56084 3724
rect 56252 3388 56308 4844
rect 56364 3780 56420 3790
rect 56476 3780 56532 8204
rect 57148 8194 57204 8204
rect 57260 14196 57316 14206
rect 56364 3778 56532 3780
rect 56364 3726 56366 3778
rect 56418 3726 56532 3778
rect 56364 3724 56532 3726
rect 56588 7700 56644 7710
rect 56364 3714 56420 3724
rect 56140 3332 56308 3388
rect 56588 3388 56644 7644
rect 57260 6804 57316 14140
rect 57372 9044 57428 22652
rect 57372 8978 57428 8988
rect 56924 6748 57316 6804
rect 56588 3332 56756 3388
rect 55580 2718 55582 2770
rect 55634 2718 55636 2770
rect 55580 2706 55636 2718
rect 55804 3220 55860 3230
rect 55244 2660 55300 2670
rect 55244 2566 55300 2604
rect 55804 2212 55860 3164
rect 55916 2884 55972 2894
rect 55916 2658 55972 2828
rect 55916 2606 55918 2658
rect 55970 2606 55972 2658
rect 55916 2594 55972 2606
rect 55916 2212 55972 2222
rect 55804 2210 55972 2212
rect 55804 2158 55918 2210
rect 55970 2158 55972 2210
rect 55804 2156 55972 2158
rect 55916 2146 55972 2156
rect 56140 1986 56196 3332
rect 56252 3108 56308 3118
rect 56252 2770 56308 3052
rect 56252 2718 56254 2770
rect 56306 2718 56308 2770
rect 56252 2706 56308 2718
rect 56700 2548 56756 3332
rect 56924 3108 56980 6748
rect 56924 3042 56980 3052
rect 57036 5124 57092 5134
rect 56140 1934 56142 1986
rect 56194 1934 56196 1986
rect 56140 1922 56196 1934
rect 56252 2492 56756 2548
rect 55804 1540 55860 1550
rect 55356 1316 55412 1326
rect 55356 112 55412 1260
rect 55804 112 55860 1484
rect 56252 112 56308 2492
rect 57036 2436 57092 5068
rect 56700 2380 57092 2436
rect 56700 112 56756 2380
rect 24220 84 24332 94
rect 24220 28 24276 84
rect 24276 18 24332 28
rect 24416 0 24528 112
rect 24864 0 24976 112
rect 25312 0 25424 112
rect 25760 0 25872 112
rect 26208 0 26320 112
rect 26656 0 26768 112
rect 27104 0 27216 112
rect 27552 0 27664 112
rect 28000 0 28112 112
rect 28448 0 28560 112
rect 28896 0 29008 112
rect 29344 0 29456 112
rect 29792 0 29904 112
rect 30240 0 30352 112
rect 30688 0 30800 112
rect 31136 0 31248 112
rect 31584 0 31696 112
rect 32032 0 32144 112
rect 32480 0 32592 112
rect 32928 0 33040 112
rect 33376 0 33488 112
rect 33824 0 33936 112
rect 34272 0 34384 112
rect 34720 0 34832 112
rect 35168 0 35280 112
rect 35616 0 35728 112
rect 36064 0 36176 112
rect 36512 0 36624 112
rect 36960 0 37072 112
rect 37408 0 37520 112
rect 37856 0 37968 112
rect 38304 0 38416 112
rect 38752 0 38864 112
rect 39200 0 39312 112
rect 39648 0 39760 112
rect 40096 0 40208 112
rect 40544 0 40656 112
rect 40992 0 41104 112
rect 41440 0 41552 112
rect 41888 0 42000 112
rect 42336 0 42448 112
rect 42784 0 42896 112
rect 43232 0 43344 112
rect 43680 0 43792 112
rect 44128 0 44240 112
rect 44576 0 44688 112
rect 45024 0 45136 112
rect 45472 0 45584 112
rect 45920 0 46032 112
rect 46368 0 46480 112
rect 46816 0 46928 112
rect 47264 0 47376 112
rect 47712 0 47824 112
rect 48160 0 48272 112
rect 48608 0 48720 112
rect 49056 0 49168 112
rect 49504 0 49616 112
rect 49952 0 50064 112
rect 50400 0 50512 112
rect 50848 0 50960 112
rect 51296 0 51408 112
rect 51744 0 51856 112
rect 52192 0 52304 112
rect 52640 0 52752 112
rect 53088 0 53200 112
rect 53536 0 53648 112
rect 53984 0 54096 112
rect 54432 0 54544 112
rect 54880 0 54992 112
rect 55328 0 55440 112
rect 55776 0 55888 112
rect 56224 0 56336 112
rect 56672 0 56784 112
<< via2 >>
rect 588 56812 644 56868
rect 476 52668 532 52724
rect 140 51324 196 51380
rect 140 43932 196 43988
rect 252 49532 308 49588
rect 140 43708 196 43764
rect 364 48188 420 48244
rect 364 46508 420 46564
rect 364 43372 420 43428
rect 140 43036 196 43092
rect 252 39116 308 39172
rect 700 56700 756 56756
rect 924 57148 980 57204
rect 700 55692 756 55748
rect 1596 57036 1652 57092
rect 1708 56924 1764 56980
rect 1148 55692 1204 55748
rect 1260 55356 1316 55412
rect 924 54348 980 54404
rect 700 54124 756 54180
rect 1148 53900 1204 53956
rect 924 53564 980 53620
rect 812 53116 868 53172
rect 588 50540 644 50596
rect 700 50876 756 50932
rect 588 48748 644 48804
rect 700 43596 756 43652
rect 588 43484 644 43540
rect 476 38892 532 38948
rect 140 29372 196 29428
rect 252 38332 308 38388
rect 252 18956 308 19012
rect 364 31836 420 31892
rect 252 18620 308 18676
rect 140 12796 196 12852
rect 28 12124 84 12180
rect 700 38668 756 38724
rect 700 34076 756 34132
rect 588 32956 644 33012
rect 588 30380 644 30436
rect 1036 52780 1092 52836
rect 1148 52332 1204 52388
rect 1260 53564 1316 53620
rect 1596 52834 1652 52836
rect 1596 52782 1598 52834
rect 1598 52782 1650 52834
rect 1650 52782 1652 52834
rect 1596 52780 1652 52782
rect 1484 52556 1540 52612
rect 1260 51100 1316 51156
rect 1148 49250 1204 49252
rect 1148 49198 1150 49250
rect 1150 49198 1202 49250
rect 1202 49198 1204 49250
rect 1148 49196 1204 49198
rect 1036 48636 1092 48692
rect 1148 48354 1204 48356
rect 1148 48302 1150 48354
rect 1150 48302 1202 48354
rect 1202 48302 1204 48354
rect 1148 48300 1204 48302
rect 1148 46732 1204 46788
rect 1484 50764 1540 50820
rect 1932 54684 1988 54740
rect 1820 54290 1876 54292
rect 1820 54238 1822 54290
rect 1822 54238 1874 54290
rect 1874 54238 1876 54290
rect 1820 54236 1876 54238
rect 1932 53730 1988 53732
rect 1932 53678 1934 53730
rect 1934 53678 1986 53730
rect 1986 53678 1988 53730
rect 1932 53676 1988 53678
rect 2156 57148 2212 57204
rect 2380 57148 2436 57204
rect 2380 56812 2436 56868
rect 2380 56252 2436 56308
rect 2268 56140 2324 56196
rect 2268 55468 2324 55524
rect 2044 52220 2100 52276
rect 1708 51548 1764 51604
rect 1932 51884 1988 51940
rect 1484 50540 1540 50596
rect 1596 49868 1652 49924
rect 1820 51266 1876 51268
rect 1820 51214 1822 51266
rect 1822 51214 1874 51266
rect 1874 51214 1876 51266
rect 1820 51212 1876 51214
rect 1596 49698 1652 49700
rect 1596 49646 1598 49698
rect 1598 49646 1650 49698
rect 1650 49646 1652 49698
rect 1596 49644 1652 49646
rect 1596 49308 1652 49364
rect 1484 48636 1540 48692
rect 1596 47964 1652 48020
rect 1820 50764 1876 50820
rect 1932 49756 1988 49812
rect 1820 48636 1876 48692
rect 1372 46114 1428 46116
rect 1372 46062 1374 46114
rect 1374 46062 1426 46114
rect 1426 46062 1428 46114
rect 1372 46060 1428 46062
rect 1260 44940 1316 44996
rect 1036 42812 1092 42868
rect 1596 46562 1652 46564
rect 1596 46510 1598 46562
rect 1598 46510 1650 46562
rect 1650 46510 1652 46562
rect 1596 46508 1652 46510
rect 1260 42252 1316 42308
rect 1596 43372 1652 43428
rect 1484 42252 1540 42308
rect 1036 41468 1092 41524
rect 1148 40460 1204 40516
rect 1148 40290 1204 40292
rect 1148 40238 1150 40290
rect 1150 40238 1202 40290
rect 1202 40238 1204 40290
rect 1148 40236 1204 40238
rect 1372 40012 1428 40068
rect 924 32732 980 32788
rect 1036 34300 1092 34356
rect 1260 38946 1316 38948
rect 1260 38894 1262 38946
rect 1262 38894 1314 38946
rect 1314 38894 1316 38946
rect 1260 38892 1316 38894
rect 1820 44940 1876 44996
rect 1932 47068 1988 47124
rect 2940 56028 2996 56084
rect 3052 56812 3108 56868
rect 3388 56364 3444 56420
rect 3612 56700 3668 56756
rect 4284 57148 4340 57204
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4284 56476 4340 56532
rect 4012 56420 4068 56422
rect 4172 56364 4228 56420
rect 3948 55970 4004 55972
rect 3948 55918 3950 55970
rect 3950 55918 4002 55970
rect 4002 55918 4004 55970
rect 3948 55916 4004 55918
rect 3500 55804 3556 55860
rect 2604 54572 2660 54628
rect 2716 54514 2772 54516
rect 2716 54462 2718 54514
rect 2718 54462 2770 54514
rect 2770 54462 2772 54514
rect 2716 54460 2772 54462
rect 2156 51772 2212 51828
rect 2828 53116 2884 53172
rect 2940 54348 2996 54404
rect 2940 52892 2996 52948
rect 2716 52220 2772 52276
rect 2940 52668 2996 52724
rect 2940 52220 2996 52276
rect 2828 52108 2884 52164
rect 2604 51996 2660 52052
rect 2940 51154 2996 51156
rect 2940 51102 2942 51154
rect 2942 51102 2994 51154
rect 2994 51102 2996 51154
rect 2940 51100 2996 51102
rect 2828 50876 2884 50932
rect 3276 55132 3332 55188
rect 3500 55410 3556 55412
rect 3500 55358 3502 55410
rect 3502 55358 3554 55410
rect 3554 55358 3556 55410
rect 3500 55356 3556 55358
rect 4060 55186 4116 55188
rect 4060 55134 4062 55186
rect 4062 55134 4114 55186
rect 4114 55134 4116 55186
rect 4060 55132 4116 55134
rect 3388 55020 3444 55076
rect 3804 54906 3860 54908
rect 3276 54460 3332 54516
rect 3164 54402 3220 54404
rect 3164 54350 3166 54402
rect 3166 54350 3218 54402
rect 3218 54350 3220 54402
rect 3164 54348 3220 54350
rect 3388 54796 3444 54852
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 4732 56252 4788 56308
rect 5068 56476 5124 56532
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 4508 55468 4564 55524
rect 4508 55244 4564 55300
rect 4956 55580 5012 55636
rect 4844 55020 4900 55076
rect 4956 55356 5012 55412
rect 4284 54796 4340 54852
rect 4284 54514 4340 54516
rect 4284 54462 4286 54514
rect 4286 54462 4338 54514
rect 4338 54462 4340 54514
rect 4284 54460 4340 54462
rect 3164 53788 3220 53844
rect 3388 53452 3444 53508
rect 3276 53116 3332 53172
rect 4464 54122 4520 54124
rect 3724 54012 3780 54068
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3612 53788 3668 53844
rect 4060 53900 4116 53956
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 5068 55132 5124 55188
rect 5068 53900 5124 53956
rect 5628 56028 5684 56084
rect 5740 57036 5796 57092
rect 6076 56252 6132 56308
rect 6300 56028 6356 56084
rect 5292 55020 5348 55076
rect 5180 53788 5236 53844
rect 5292 54124 5348 54180
rect 5404 54012 5460 54068
rect 3388 52722 3444 52724
rect 3388 52670 3390 52722
rect 3390 52670 3442 52722
rect 3442 52670 3444 52722
rect 3388 52668 3444 52670
rect 3276 52444 3332 52500
rect 3500 52556 3556 52612
rect 3612 52444 3668 52500
rect 3164 51884 3220 51940
rect 4956 52892 5012 52948
rect 4172 52780 4228 52836
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 4396 52722 4452 52724
rect 4396 52670 4398 52722
rect 4398 52670 4450 52722
rect 4450 52670 4452 52722
rect 4396 52668 4452 52670
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 4732 52274 4788 52276
rect 4732 52222 4734 52274
rect 4734 52222 4786 52274
rect 4786 52222 4788 52274
rect 4732 52220 4788 52222
rect 4284 51884 4340 51940
rect 4396 51996 4452 52052
rect 3388 51100 3444 51156
rect 3500 50876 3556 50932
rect 2492 49196 2548 49252
rect 2268 48972 2324 49028
rect 2156 48524 2212 48580
rect 2044 46284 2100 46340
rect 2044 46002 2100 46004
rect 2044 45950 2046 46002
rect 2046 45950 2098 46002
rect 2098 45950 2100 46002
rect 2044 45948 2100 45950
rect 2492 48914 2548 48916
rect 2492 48862 2494 48914
rect 2494 48862 2546 48914
rect 2546 48862 2548 48914
rect 2492 48860 2548 48862
rect 2492 46620 2548 46676
rect 2268 45388 2324 45444
rect 1932 44492 1988 44548
rect 1820 44434 1876 44436
rect 1820 44382 1822 44434
rect 1822 44382 1874 44434
rect 1874 44382 1876 44434
rect 1820 44380 1876 44382
rect 2268 45052 2324 45108
rect 2044 44268 2100 44324
rect 2156 44492 2212 44548
rect 1820 44156 1876 44212
rect 1820 43372 1876 43428
rect 1820 42978 1876 42980
rect 1820 42926 1822 42978
rect 1822 42926 1874 42978
rect 1874 42926 1876 42978
rect 1820 42924 1876 42926
rect 1932 42588 1988 42644
rect 2044 43596 2100 43652
rect 1708 41916 1764 41972
rect 1596 41858 1652 41860
rect 1596 41806 1598 41858
rect 1598 41806 1650 41858
rect 1650 41806 1652 41858
rect 1596 41804 1652 41806
rect 1708 41020 1764 41076
rect 1596 40402 1652 40404
rect 1596 40350 1598 40402
rect 1598 40350 1650 40402
rect 1650 40350 1652 40402
rect 1596 40348 1652 40350
rect 1932 40684 1988 40740
rect 1708 38722 1764 38724
rect 1708 38670 1710 38722
rect 1710 38670 1762 38722
rect 1762 38670 1764 38722
rect 1708 38668 1764 38670
rect 2268 42924 2324 42980
rect 2380 42364 2436 42420
rect 2828 50482 2884 50484
rect 2828 50430 2830 50482
rect 2830 50430 2882 50482
rect 2882 50430 2884 50482
rect 2828 50428 2884 50430
rect 3052 49980 3108 50036
rect 4172 51378 4228 51380
rect 4172 51326 4174 51378
rect 4174 51326 4226 51378
rect 4226 51326 4228 51378
rect 4172 51324 4228 51326
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 4508 50428 4564 50484
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 3500 49698 3556 49700
rect 3500 49646 3502 49698
rect 3502 49646 3554 49698
rect 3554 49646 3556 49698
rect 3500 49644 3556 49646
rect 3164 49532 3220 49588
rect 2828 49196 2884 49252
rect 2940 49308 2996 49364
rect 2940 48748 2996 48804
rect 2940 48300 2996 48356
rect 2716 48242 2772 48244
rect 2716 48190 2718 48242
rect 2718 48190 2770 48242
rect 2770 48190 2772 48242
rect 2716 48188 2772 48190
rect 2828 47682 2884 47684
rect 2828 47630 2830 47682
rect 2830 47630 2882 47682
rect 2882 47630 2884 47682
rect 2828 47628 2884 47630
rect 2716 45724 2772 45780
rect 2828 45836 2884 45892
rect 2604 45276 2660 45332
rect 2716 45388 2772 45444
rect 2604 44940 2660 44996
rect 2604 43036 2660 43092
rect 3388 49586 3444 49588
rect 3388 49534 3390 49586
rect 3390 49534 3442 49586
rect 3442 49534 3444 49586
rect 3388 49532 3444 49534
rect 3388 48636 3444 48692
rect 3052 48188 3108 48244
rect 3052 47404 3108 47460
rect 3164 47964 3220 48020
rect 3052 47068 3108 47124
rect 3164 46620 3220 46676
rect 3388 48300 3444 48356
rect 3500 48972 3556 49028
rect 3388 47852 3444 47908
rect 3052 46172 3108 46228
rect 3164 46396 3220 46452
rect 3164 45388 3220 45444
rect 3164 44940 3220 44996
rect 3052 44828 3108 44884
rect 2940 43148 2996 43204
rect 3388 46562 3444 46564
rect 3388 46510 3390 46562
rect 3390 46510 3442 46562
rect 3442 46510 3444 46562
rect 3388 46508 3444 46510
rect 5292 52834 5348 52836
rect 5292 52782 5294 52834
rect 5294 52782 5346 52834
rect 5346 52782 5348 52834
rect 5292 52780 5348 52782
rect 5964 55468 6020 55524
rect 5628 53618 5684 53620
rect 5628 53566 5630 53618
rect 5630 53566 5682 53618
rect 5682 53566 5684 53618
rect 5628 53564 5684 53566
rect 7420 56364 7476 56420
rect 7868 56364 7924 56420
rect 6748 55580 6804 55636
rect 6524 55468 6580 55524
rect 6076 55298 6132 55300
rect 6076 55246 6078 55298
rect 6078 55246 6130 55298
rect 6130 55246 6132 55298
rect 6076 55244 6132 55246
rect 5740 53340 5796 53396
rect 5964 54402 6020 54404
rect 5964 54350 5966 54402
rect 5966 54350 6018 54402
rect 6018 54350 6020 54402
rect 5964 54348 6020 54350
rect 5516 52556 5572 52612
rect 5404 52444 5460 52500
rect 5628 51154 5684 51156
rect 5628 51102 5630 51154
rect 5630 51102 5682 51154
rect 5682 51102 5684 51154
rect 5628 51100 5684 51102
rect 5628 50652 5684 50708
rect 4732 50204 4788 50260
rect 5068 49980 5124 50036
rect 4396 49810 4452 49812
rect 4396 49758 4398 49810
rect 4398 49758 4450 49810
rect 4450 49758 4452 49810
rect 4396 49756 4452 49758
rect 3948 49420 4004 49476
rect 4172 49532 4228 49588
rect 4060 49308 4116 49364
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 3948 48972 4004 49028
rect 3836 48748 3892 48804
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 4172 48524 4228 48580
rect 4508 48412 4564 48468
rect 4956 48412 5012 48468
rect 4172 47852 4228 47908
rect 5068 47964 5124 48020
rect 4464 47850 4520 47852
rect 4284 47740 4340 47796
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4956 47852 5012 47908
rect 4672 47796 4728 47798
rect 3724 47180 3780 47236
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4172 47068 4228 47124
rect 4012 47012 4068 47014
rect 4620 47628 4676 47684
rect 4396 47458 4452 47460
rect 4396 47406 4398 47458
rect 4398 47406 4450 47458
rect 4450 47406 4452 47458
rect 4396 47404 4452 47406
rect 5068 47570 5124 47572
rect 5068 47518 5070 47570
rect 5070 47518 5122 47570
rect 5122 47518 5124 47570
rect 5068 47516 5124 47518
rect 6188 53058 6244 53060
rect 6188 53006 6190 53058
rect 6190 53006 6242 53058
rect 6242 53006 6244 53058
rect 6188 53004 6244 53006
rect 6412 54908 6468 54964
rect 6524 55244 6580 55300
rect 6300 51772 6356 51828
rect 5404 49420 5460 49476
rect 5404 49196 5460 49252
rect 5516 48860 5572 48916
rect 5628 48972 5684 49028
rect 5292 48242 5348 48244
rect 5292 48190 5294 48242
rect 5294 48190 5346 48242
rect 5346 48190 5348 48242
rect 5292 48188 5348 48190
rect 5180 47404 5236 47460
rect 4956 47068 5012 47124
rect 5180 47068 5236 47124
rect 3948 46562 4004 46564
rect 3948 46510 3950 46562
rect 3950 46510 4002 46562
rect 4002 46510 4004 46562
rect 3948 46508 4004 46510
rect 4060 46284 4116 46340
rect 3836 46172 3892 46228
rect 3388 45612 3444 45668
rect 4060 46002 4116 46004
rect 4060 45950 4062 46002
rect 4062 45950 4114 46002
rect 4114 45950 4116 46002
rect 4060 45948 4116 45950
rect 3948 45612 4004 45668
rect 3500 45276 3556 45332
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 4284 46396 4340 46452
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 4172 45388 4228 45444
rect 3388 44994 3444 44996
rect 3388 44942 3390 44994
rect 3390 44942 3442 44994
rect 3442 44942 3444 44994
rect 3388 44940 3444 44942
rect 3500 44828 3556 44884
rect 2716 42812 2772 42868
rect 2492 41804 2548 41860
rect 2268 41468 2324 41524
rect 3164 43650 3220 43652
rect 3164 43598 3166 43650
rect 3166 43598 3218 43650
rect 3218 43598 3220 43650
rect 3164 43596 3220 43598
rect 2604 41132 2660 41188
rect 2156 40684 2212 40740
rect 2380 40908 2436 40964
rect 1596 38162 1652 38164
rect 1596 38110 1598 38162
rect 1598 38110 1650 38162
rect 1650 38110 1652 38162
rect 1596 38108 1652 38110
rect 2044 39842 2100 39844
rect 2044 39790 2046 39842
rect 2046 39790 2098 39842
rect 2098 39790 2100 39842
rect 2044 39788 2100 39790
rect 2716 41692 2772 41748
rect 2828 41020 2884 41076
rect 2828 40348 2884 40404
rect 2604 39900 2660 39956
rect 3388 43148 3444 43204
rect 3164 42028 3220 42084
rect 3276 42700 3332 42756
rect 3388 42476 3444 42532
rect 3948 45106 4004 45108
rect 3948 45054 3950 45106
rect 3950 45054 4002 45106
rect 4002 45054 4004 45106
rect 3948 45052 4004 45054
rect 4396 45276 4452 45332
rect 4620 45276 4676 45332
rect 4172 44716 4228 44772
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4172 43932 4228 43988
rect 4012 43876 4068 43878
rect 4060 43538 4116 43540
rect 4060 43486 4062 43538
rect 4062 43486 4114 43538
rect 4114 43486 4116 43538
rect 4060 43484 4116 43486
rect 4284 43538 4340 43540
rect 4284 43486 4286 43538
rect 4286 43486 4338 43538
rect 4338 43486 4340 43538
rect 4284 43484 4340 43486
rect 3500 41916 3556 41972
rect 3164 41804 3220 41860
rect 2716 40124 2772 40180
rect 3052 41692 3108 41748
rect 2156 38780 2212 38836
rect 2380 39452 2436 39508
rect 1596 36764 1652 36820
rect 1484 36204 1540 36260
rect 1260 34130 1316 34132
rect 1260 34078 1262 34130
rect 1262 34078 1314 34130
rect 1314 34078 1316 34130
rect 1260 34076 1316 34078
rect 1036 32620 1092 32676
rect 812 32284 868 32340
rect 924 32508 980 32564
rect 812 32060 868 32116
rect 1148 32508 1204 32564
rect 1372 33570 1428 33572
rect 1372 33518 1374 33570
rect 1374 33518 1426 33570
rect 1426 33518 1428 33570
rect 1372 33516 1428 33518
rect 1708 35308 1764 35364
rect 1708 33906 1764 33908
rect 1708 33854 1710 33906
rect 1710 33854 1762 33906
rect 1762 33854 1764 33906
rect 1708 33852 1764 33854
rect 1820 33628 1876 33684
rect 1820 33068 1876 33124
rect 1484 32956 1540 33012
rect 924 31164 980 31220
rect 1484 32732 1540 32788
rect 1372 32284 1428 32340
rect 1708 32450 1764 32452
rect 1708 32398 1710 32450
rect 1710 32398 1762 32450
rect 1762 32398 1764 32450
rect 1708 32396 1764 32398
rect 1596 32284 1652 32340
rect 476 28364 532 28420
rect 700 29708 756 29764
rect 588 22876 644 22932
rect 364 18508 420 18564
rect 476 21532 532 21588
rect 812 25676 868 25732
rect 700 22204 756 22260
rect 812 25452 868 25508
rect 924 23212 980 23268
rect 1036 28364 1092 28420
rect 1036 27020 1092 27076
rect 1372 27858 1428 27860
rect 1372 27806 1374 27858
rect 1374 27806 1426 27858
rect 1426 27806 1428 27858
rect 1372 27804 1428 27806
rect 2156 36764 2212 36820
rect 2044 33458 2100 33460
rect 2044 33406 2046 33458
rect 2046 33406 2098 33458
rect 2098 33406 2100 33458
rect 2044 33404 2100 33406
rect 1596 29314 1652 29316
rect 1596 29262 1598 29314
rect 1598 29262 1650 29314
rect 1650 29262 1652 29314
rect 1596 29260 1652 29262
rect 1596 27468 1652 27524
rect 1932 29484 1988 29540
rect 2044 32956 2100 33012
rect 1708 27132 1764 27188
rect 1372 26012 1428 26068
rect 1708 26066 1764 26068
rect 1708 26014 1710 26066
rect 1710 26014 1762 26066
rect 1762 26014 1764 26066
rect 1708 26012 1764 26014
rect 1260 25506 1316 25508
rect 1260 25454 1262 25506
rect 1262 25454 1314 25506
rect 1314 25454 1316 25506
rect 1260 25452 1316 25454
rect 1148 24610 1204 24612
rect 1148 24558 1150 24610
rect 1150 24558 1202 24610
rect 1202 24558 1204 24610
rect 1148 24556 1204 24558
rect 1036 21362 1092 21364
rect 1036 21310 1038 21362
rect 1038 21310 1090 21362
rect 1090 21310 1092 21362
rect 1036 21308 1092 21310
rect 812 20860 868 20916
rect 1372 21644 1428 21700
rect 1372 21474 1428 21476
rect 1372 21422 1374 21474
rect 1374 21422 1426 21474
rect 1426 21422 1428 21474
rect 1372 21420 1428 21422
rect 1260 20188 1316 20244
rect 1372 21084 1428 21140
rect 1148 19794 1204 19796
rect 1148 19742 1150 19794
rect 1150 19742 1202 19794
rect 1202 19742 1204 19794
rect 1148 19740 1204 19742
rect 700 18844 756 18900
rect 812 19068 868 19124
rect 588 16828 644 16884
rect 476 16716 532 16772
rect 588 16380 644 16436
rect 252 10220 308 10276
rect 364 14364 420 14420
rect 252 7308 308 7364
rect 476 9212 532 9268
rect 700 14588 756 14644
rect 700 11116 756 11172
rect 924 18172 980 18228
rect 1820 25730 1876 25732
rect 1820 25678 1822 25730
rect 1822 25678 1874 25730
rect 1874 25678 1876 25730
rect 1820 25676 1876 25678
rect 1820 24332 1876 24388
rect 1708 23772 1764 23828
rect 1484 19740 1540 19796
rect 1596 23660 1652 23716
rect 1484 19346 1540 19348
rect 1484 19294 1486 19346
rect 1486 19294 1538 19346
rect 1538 19294 1540 19346
rect 1484 19292 1540 19294
rect 1372 18226 1428 18228
rect 1372 18174 1374 18226
rect 1374 18174 1426 18226
rect 1426 18174 1428 18226
rect 1372 18172 1428 18174
rect 1372 17500 1428 17556
rect 1260 16716 1316 16772
rect 1372 16268 1428 16324
rect 1260 16098 1316 16100
rect 1260 16046 1262 16098
rect 1262 16046 1314 16098
rect 1314 16046 1316 16098
rect 1260 16044 1316 16046
rect 1260 15708 1316 15764
rect 1148 14530 1204 14532
rect 1148 14478 1150 14530
rect 1150 14478 1202 14530
rect 1202 14478 1204 14530
rect 1148 14476 1204 14478
rect 1036 14418 1092 14420
rect 1036 14366 1038 14418
rect 1038 14366 1090 14418
rect 1090 14366 1092 14418
rect 1036 14364 1092 14366
rect 1708 21474 1764 21476
rect 1708 21422 1710 21474
rect 1710 21422 1762 21474
rect 1762 21422 1764 21474
rect 1708 21420 1764 21422
rect 1932 22370 1988 22372
rect 1932 22318 1934 22370
rect 1934 22318 1986 22370
rect 1986 22318 1988 22370
rect 1932 22316 1988 22318
rect 2156 27804 2212 27860
rect 2380 38444 2436 38500
rect 2492 37996 2548 38052
rect 2716 37772 2772 37828
rect 3388 41858 3444 41860
rect 3388 41806 3390 41858
rect 3390 41806 3442 41858
rect 3442 41806 3444 41858
rect 3388 41804 3444 41806
rect 3724 43036 3780 43092
rect 5068 46620 5124 46676
rect 4956 45500 5012 45556
rect 5292 45500 5348 45556
rect 5180 45388 5236 45444
rect 4956 44994 5012 44996
rect 4956 44942 4958 44994
rect 4958 44942 5010 44994
rect 5010 44942 5012 44994
rect 4956 44940 5012 44942
rect 5068 44882 5124 44884
rect 5068 44830 5070 44882
rect 5070 44830 5122 44882
rect 5122 44830 5124 44882
rect 5068 44828 5124 44830
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 4956 44716 5012 44772
rect 3948 42476 4004 42532
rect 4284 42754 4340 42756
rect 4284 42702 4286 42754
rect 4286 42702 4338 42754
rect 4338 42702 4340 42754
rect 4284 42700 4340 42702
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 3276 39900 3332 39956
rect 3388 41020 3444 41076
rect 4060 41970 4116 41972
rect 4060 41918 4062 41970
rect 4062 41918 4114 41970
rect 4114 41918 4116 41970
rect 4060 41916 4116 41918
rect 3836 41020 3892 41076
rect 4284 42028 4340 42084
rect 4284 41580 4340 41636
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 4508 41298 4564 41300
rect 4508 41246 4510 41298
rect 4510 41246 4562 41298
rect 4562 41246 4564 41298
rect 4508 41244 4564 41246
rect 4844 41244 4900 41300
rect 5292 45164 5348 45220
rect 5292 44604 5348 44660
rect 5180 44268 5236 44324
rect 5628 48412 5684 48468
rect 5740 47740 5796 47796
rect 5628 47180 5684 47236
rect 5404 44156 5460 44212
rect 5292 43820 5348 43876
rect 5068 41468 5124 41524
rect 3500 40796 3556 40852
rect 4284 41020 4340 41076
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4172 40796 4228 40852
rect 4732 40796 4788 40852
rect 4012 40740 4068 40742
rect 3500 40460 3556 40516
rect 3276 39618 3332 39620
rect 3276 39566 3278 39618
rect 3278 39566 3330 39618
rect 3330 39566 3332 39618
rect 3276 39564 3332 39566
rect 3164 39452 3220 39508
rect 3388 39452 3444 39508
rect 3276 38892 3332 38948
rect 4284 40348 4340 40404
rect 4956 40796 5012 40852
rect 5068 41186 5124 41188
rect 5068 41134 5070 41186
rect 5070 41134 5122 41186
rect 5122 41134 5124 41186
rect 5068 41132 5124 41134
rect 4172 39900 4228 39956
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 3612 38332 3668 38388
rect 3612 38050 3668 38052
rect 3612 37998 3614 38050
rect 3614 37998 3666 38050
rect 3666 37998 3668 38050
rect 3612 37996 3668 37998
rect 3836 38834 3892 38836
rect 3836 38782 3838 38834
rect 3838 38782 3890 38834
rect 3890 38782 3892 38834
rect 3836 38780 3892 38782
rect 4060 38780 4116 38836
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 5292 41858 5348 41860
rect 5292 41806 5294 41858
rect 5294 41806 5346 41858
rect 5346 41806 5348 41858
rect 5292 41804 5348 41806
rect 5516 42140 5572 42196
rect 5740 46450 5796 46452
rect 5740 46398 5742 46450
rect 5742 46398 5794 46450
rect 5794 46398 5796 46450
rect 5740 46396 5796 46398
rect 5964 48748 6020 48804
rect 6076 49644 6132 49700
rect 5964 48130 6020 48132
rect 5964 48078 5966 48130
rect 5966 48078 6018 48130
rect 6018 48078 6020 48130
rect 5964 48076 6020 48078
rect 5964 47740 6020 47796
rect 5964 47180 6020 47236
rect 5964 46956 6020 47012
rect 5964 46732 6020 46788
rect 6636 54124 6692 54180
rect 6972 55858 7028 55860
rect 6972 55806 6974 55858
rect 6974 55806 7026 55858
rect 7026 55806 7028 55858
rect 6972 55804 7028 55806
rect 7308 55580 7364 55636
rect 6972 55410 7028 55412
rect 6972 55358 6974 55410
rect 6974 55358 7026 55410
rect 7026 55358 7028 55410
rect 6972 55356 7028 55358
rect 6860 53228 6916 53284
rect 6972 55132 7028 55188
rect 6524 52946 6580 52948
rect 6524 52894 6526 52946
rect 6526 52894 6578 52946
rect 6578 52894 6580 52946
rect 6524 52892 6580 52894
rect 6412 51212 6468 51268
rect 6748 52892 6804 52948
rect 6300 50764 6356 50820
rect 6300 50092 6356 50148
rect 6188 47740 6244 47796
rect 6076 45948 6132 46004
rect 6188 46956 6244 47012
rect 5740 42364 5796 42420
rect 5852 44604 5908 44660
rect 5628 41916 5684 41972
rect 5628 41468 5684 41524
rect 5516 41186 5572 41188
rect 5516 41134 5518 41186
rect 5518 41134 5570 41186
rect 5570 41134 5572 41186
rect 5516 41132 5572 41134
rect 5404 40684 5460 40740
rect 5516 40402 5572 40404
rect 5516 40350 5518 40402
rect 5518 40350 5570 40402
rect 5570 40350 5572 40402
rect 5516 40348 5572 40350
rect 5404 40178 5460 40180
rect 5404 40126 5406 40178
rect 5406 40126 5458 40178
rect 5458 40126 5460 40178
rect 5404 40124 5460 40126
rect 5628 40124 5684 40180
rect 5964 43708 6020 43764
rect 5964 42700 6020 42756
rect 4284 38780 4340 38836
rect 4396 39116 4452 39172
rect 5180 39564 5236 39620
rect 5068 38780 5124 38836
rect 4732 38668 4788 38724
rect 4956 38722 5012 38724
rect 4956 38670 4958 38722
rect 4958 38670 5010 38722
rect 5010 38670 5012 38722
rect 4956 38668 5012 38670
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4844 38444 4900 38500
rect 4672 38388 4728 38390
rect 3948 38220 4004 38276
rect 5068 37996 5124 38052
rect 3388 37548 3444 37604
rect 2828 37100 2884 37156
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 3668 36988 3724 37044
rect 2716 36764 2772 36820
rect 4396 37772 4452 37828
rect 4396 37154 4452 37156
rect 4396 37102 4398 37154
rect 4398 37102 4450 37154
rect 4450 37102 4452 37154
rect 4396 37100 4452 37102
rect 4956 37660 5012 37716
rect 5404 39116 5460 39172
rect 5180 37548 5236 37604
rect 5068 37324 5124 37380
rect 4620 37100 4676 37156
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 5068 36988 5124 37044
rect 2492 36204 2548 36260
rect 2828 36482 2884 36484
rect 2828 36430 2830 36482
rect 2830 36430 2882 36482
rect 2882 36430 2884 36482
rect 2828 36428 2884 36430
rect 2940 36316 2996 36372
rect 2380 35420 2436 35476
rect 2604 35196 2660 35252
rect 2828 35026 2884 35028
rect 2828 34974 2830 35026
rect 2830 34974 2882 35026
rect 2882 34974 2884 35026
rect 2828 34972 2884 34974
rect 2604 34188 2660 34244
rect 2716 34860 2772 34916
rect 2492 33404 2548 33460
rect 2828 33404 2884 33460
rect 3276 36370 3332 36372
rect 3276 36318 3278 36370
rect 3278 36318 3330 36370
rect 3330 36318 3332 36370
rect 3276 36316 3332 36318
rect 3500 35868 3556 35924
rect 4060 36316 4116 36372
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 3948 35868 4004 35924
rect 3836 35532 3892 35588
rect 3836 35308 3892 35364
rect 3724 35196 3780 35252
rect 3500 35084 3556 35140
rect 3500 34914 3556 34916
rect 3500 34862 3502 34914
rect 3502 34862 3554 34914
rect 3554 34862 3556 34914
rect 3500 34860 3556 34862
rect 3724 34914 3780 34916
rect 3724 34862 3726 34914
rect 3726 34862 3778 34914
rect 3778 34862 3780 34914
rect 3724 34860 3780 34862
rect 3052 34076 3108 34132
rect 3724 34636 3780 34692
rect 3948 34636 4004 34692
rect 3804 34522 3860 34524
rect 3612 34412 3668 34468
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 4732 36482 4788 36484
rect 4732 36430 4734 36482
rect 4734 36430 4786 36482
rect 4786 36430 4788 36482
rect 4732 36428 4788 36430
rect 4508 36316 4564 36372
rect 4396 36092 4452 36148
rect 4284 35868 4340 35924
rect 4508 35980 4564 36036
rect 4508 35532 4564 35588
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 5068 36092 5124 36148
rect 4956 35810 5012 35812
rect 4956 35758 4958 35810
rect 4958 35758 5010 35810
rect 5010 35758 5012 35810
rect 4956 35756 5012 35758
rect 4844 35084 4900 35140
rect 3500 33740 3556 33796
rect 3164 33516 3220 33572
rect 2604 32732 2660 32788
rect 3388 32450 3444 32452
rect 3388 32398 3390 32450
rect 3390 32398 3442 32450
rect 3442 32398 3444 32450
rect 3388 32396 3444 32398
rect 2828 32060 2884 32116
rect 4284 34524 4340 34580
rect 3948 34130 4004 34132
rect 3948 34078 3950 34130
rect 3950 34078 4002 34130
rect 4002 34078 4004 34130
rect 3948 34076 4004 34078
rect 4396 34412 4452 34468
rect 5068 35196 5124 35252
rect 4956 34412 5012 34468
rect 5068 34636 5124 34692
rect 4396 34018 4452 34020
rect 4396 33966 4398 34018
rect 4398 33966 4450 34018
rect 4450 33966 4452 34018
rect 4396 33964 4452 33966
rect 3836 33852 3892 33908
rect 3948 33570 4004 33572
rect 3948 33518 3950 33570
rect 3950 33518 4002 33570
rect 4002 33518 4004 33570
rect 3948 33516 4004 33518
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4060 33068 4116 33124
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4284 32956 4340 33012
rect 4012 32900 4068 32902
rect 4732 33292 4788 33348
rect 4620 32956 4676 33012
rect 5068 33068 5124 33124
rect 4844 32956 4900 33012
rect 4396 32844 4452 32900
rect 3948 32620 4004 32676
rect 3612 32284 3668 32340
rect 4172 32674 4228 32676
rect 4172 32622 4174 32674
rect 4174 32622 4226 32674
rect 4226 32622 4228 32674
rect 4172 32620 4228 32622
rect 4620 32508 4676 32564
rect 4060 32396 4116 32452
rect 3836 32172 3892 32228
rect 3500 32060 3556 32116
rect 3388 31836 3444 31892
rect 3164 31500 3220 31556
rect 3276 31724 3332 31780
rect 3052 31276 3108 31332
rect 2716 30268 2772 30324
rect 2940 30156 2996 30212
rect 2828 29426 2884 29428
rect 2828 29374 2830 29426
rect 2830 29374 2882 29426
rect 2882 29374 2884 29426
rect 2828 29372 2884 29374
rect 2604 29260 2660 29316
rect 2380 28028 2436 28084
rect 2604 28924 2660 28980
rect 2492 27916 2548 27972
rect 2268 25116 2324 25172
rect 2156 24668 2212 24724
rect 1820 21308 1876 21364
rect 1708 21026 1764 21028
rect 1708 20974 1710 21026
rect 1710 20974 1762 21026
rect 1762 20974 1764 21026
rect 1708 20972 1764 20974
rect 1820 20300 1876 20356
rect 1708 18226 1764 18228
rect 1708 18174 1710 18226
rect 1710 18174 1762 18226
rect 1762 18174 1764 18226
rect 1708 18172 1764 18174
rect 2044 20524 2100 20580
rect 1932 20076 1988 20132
rect 1820 16994 1876 16996
rect 1820 16942 1822 16994
rect 1822 16942 1874 16994
rect 1874 16942 1876 16994
rect 1820 16940 1876 16942
rect 1820 16044 1876 16100
rect 2156 19068 2212 19124
rect 2268 21308 2324 21364
rect 2828 28866 2884 28868
rect 2828 28814 2830 28866
rect 2830 28814 2882 28866
rect 2882 28814 2884 28866
rect 2828 28812 2884 28814
rect 2716 27804 2772 27860
rect 2940 27746 2996 27748
rect 2940 27694 2942 27746
rect 2942 27694 2994 27746
rect 2994 27694 2996 27746
rect 2940 27692 2996 27694
rect 3276 30940 3332 30996
rect 3388 30604 3444 30660
rect 4172 32338 4228 32340
rect 4172 32286 4174 32338
rect 4174 32286 4226 32338
rect 4226 32286 4228 32338
rect 4172 32284 4228 32286
rect 3948 32060 4004 32116
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 3612 31724 3668 31780
rect 4284 31778 4340 31780
rect 4284 31726 4286 31778
rect 4286 31726 4338 31778
rect 4338 31726 4340 31778
rect 4284 31724 4340 31726
rect 3612 31276 3668 31332
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4284 31388 4340 31444
rect 4012 31332 4068 31334
rect 4508 31276 4564 31332
rect 4508 31052 4564 31108
rect 3612 30716 3668 30772
rect 3948 30994 4004 30996
rect 3948 30942 3950 30994
rect 3950 30942 4002 30994
rect 4002 30942 4004 30994
rect 3948 30940 4004 30942
rect 4060 30604 4116 30660
rect 4172 30492 4228 30548
rect 4060 30210 4116 30212
rect 4060 30158 4062 30210
rect 4062 30158 4114 30210
rect 4114 30158 4116 30210
rect 4060 30156 4116 30158
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 3276 29484 3332 29540
rect 3164 29260 3220 29316
rect 3836 29426 3892 29428
rect 3836 29374 3838 29426
rect 3838 29374 3890 29426
rect 3890 29374 3892 29426
rect 3836 29372 3892 29374
rect 3388 28924 3444 28980
rect 3276 28812 3332 28868
rect 3276 28364 3332 28420
rect 3612 28642 3668 28644
rect 3612 28590 3614 28642
rect 3614 28590 3666 28642
rect 3666 28590 3668 28642
rect 3612 28588 3668 28590
rect 4060 29596 4116 29652
rect 5292 37324 5348 37380
rect 5292 35868 5348 35924
rect 5292 35026 5348 35028
rect 5292 34974 5294 35026
rect 5294 34974 5346 35026
rect 5346 34974 5348 35026
rect 5292 34972 5348 34974
rect 5292 34524 5348 34580
rect 5292 33628 5348 33684
rect 5628 38050 5684 38052
rect 5628 37998 5630 38050
rect 5630 37998 5682 38050
rect 5682 37998 5684 38050
rect 5628 37996 5684 37998
rect 6188 45276 6244 45332
rect 6188 45052 6244 45108
rect 6412 48412 6468 48468
rect 6636 52220 6692 52276
rect 6636 51884 6692 51940
rect 6748 52108 6804 52164
rect 6636 51548 6692 51604
rect 6636 50092 6692 50148
rect 6860 51548 6916 51604
rect 7084 54514 7140 54516
rect 7084 54462 7086 54514
rect 7086 54462 7138 54514
rect 7138 54462 7140 54514
rect 7084 54460 7140 54462
rect 7308 53788 7364 53844
rect 7644 55580 7700 55636
rect 7420 53564 7476 53620
rect 7532 54348 7588 54404
rect 7196 53506 7252 53508
rect 7196 53454 7198 53506
rect 7198 53454 7250 53506
rect 7250 53454 7252 53506
rect 7196 53452 7252 53454
rect 7644 54290 7700 54292
rect 7644 54238 7646 54290
rect 7646 54238 7698 54290
rect 7698 54238 7700 54290
rect 7644 54236 7700 54238
rect 8092 55298 8148 55300
rect 8092 55246 8094 55298
rect 8094 55246 8146 55298
rect 8146 55246 8148 55298
rect 8092 55244 8148 55246
rect 9212 56924 9268 56980
rect 9324 56364 9380 56420
rect 8764 55468 8820 55524
rect 9100 55298 9156 55300
rect 9100 55246 9102 55298
rect 9102 55246 9154 55298
rect 9154 55246 9156 55298
rect 9100 55244 9156 55246
rect 8316 55132 8372 55188
rect 7980 53900 8036 53956
rect 7644 53340 7700 53396
rect 7084 52668 7140 52724
rect 7196 51436 7252 51492
rect 7308 51266 7364 51268
rect 7308 51214 7310 51266
rect 7310 51214 7362 51266
rect 7362 51214 7364 51266
rect 7308 51212 7364 51214
rect 7084 50988 7140 51044
rect 6972 50764 7028 50820
rect 6860 50706 6916 50708
rect 6860 50654 6862 50706
rect 6862 50654 6914 50706
rect 6914 50654 6916 50706
rect 6860 50652 6916 50654
rect 7196 50652 7252 50708
rect 6860 50204 6916 50260
rect 6748 49084 6804 49140
rect 6524 48188 6580 48244
rect 6300 43820 6356 43876
rect 6412 47404 6468 47460
rect 6188 43596 6244 43652
rect 6300 43036 6356 43092
rect 6748 48524 6804 48580
rect 6748 46956 6804 47012
rect 6972 49868 7028 49924
rect 7196 49868 7252 49924
rect 7196 48636 7252 48692
rect 6524 45500 6580 45556
rect 6636 44380 6692 44436
rect 6412 42754 6468 42756
rect 6412 42702 6414 42754
rect 6414 42702 6466 42754
rect 6466 42702 6468 42754
rect 6412 42700 6468 42702
rect 6300 42252 6356 42308
rect 6188 42194 6244 42196
rect 6188 42142 6190 42194
rect 6190 42142 6242 42194
rect 6242 42142 6244 42194
rect 6188 42140 6244 42142
rect 6188 40796 6244 40852
rect 6300 40514 6356 40516
rect 6300 40462 6302 40514
rect 6302 40462 6354 40514
rect 6354 40462 6356 40514
rect 6300 40460 6356 40462
rect 5964 37548 6020 37604
rect 6188 38108 6244 38164
rect 6188 37772 6244 37828
rect 6188 37154 6244 37156
rect 6188 37102 6190 37154
rect 6190 37102 6242 37154
rect 6242 37102 6244 37154
rect 6188 37100 6244 37102
rect 5516 35308 5572 35364
rect 5404 33516 5460 33572
rect 5292 32060 5348 32116
rect 5516 35084 5572 35140
rect 5516 32508 5572 32564
rect 5516 32338 5572 32340
rect 5516 32286 5518 32338
rect 5518 32286 5570 32338
rect 5570 32286 5572 32338
rect 5516 32284 5572 32286
rect 4844 31778 4900 31780
rect 4844 31726 4846 31778
rect 4846 31726 4898 31778
rect 4898 31726 4900 31778
rect 4844 31724 4900 31726
rect 4732 31052 4788 31108
rect 5068 31388 5124 31444
rect 5180 31500 5236 31556
rect 5068 31106 5124 31108
rect 5068 31054 5070 31106
rect 5070 31054 5122 31106
rect 5122 31054 5124 31106
rect 5068 31052 5124 31054
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4956 30604 5012 30660
rect 4672 30548 4728 30550
rect 4844 30492 4900 30548
rect 4508 30210 4564 30212
rect 4508 30158 4510 30210
rect 4510 30158 4562 30210
rect 4562 30158 4564 30210
rect 4508 30156 4564 30158
rect 4396 30044 4452 30100
rect 4396 29820 4452 29876
rect 4284 29708 4340 29764
rect 4844 30156 4900 30212
rect 4172 29036 4228 29092
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 3948 28642 4004 28644
rect 3948 28590 3950 28642
rect 3950 28590 4002 28642
rect 4002 28590 4004 28642
rect 3948 28588 4004 28590
rect 6636 42028 6692 42084
rect 6524 40796 6580 40852
rect 6860 46562 6916 46564
rect 6860 46510 6862 46562
rect 6862 46510 6914 46562
rect 6914 46510 6916 46562
rect 6860 46508 6916 46510
rect 7196 47516 7252 47572
rect 7084 47458 7140 47460
rect 7084 47406 7086 47458
rect 7086 47406 7138 47458
rect 7138 47406 7140 47458
rect 7084 47404 7140 47406
rect 7084 44604 7140 44660
rect 6972 44380 7028 44436
rect 6860 44044 6916 44100
rect 6972 43932 7028 43988
rect 6860 42252 6916 42308
rect 7644 52556 7700 52612
rect 7532 50594 7588 50596
rect 7532 50542 7534 50594
rect 7534 50542 7586 50594
rect 7586 50542 7588 50594
rect 7532 50540 7588 50542
rect 7420 48412 7476 48468
rect 7532 50204 7588 50260
rect 7532 49868 7588 49924
rect 7420 47740 7476 47796
rect 7756 51548 7812 51604
rect 7980 53116 8036 53172
rect 7980 52108 8036 52164
rect 8988 54572 9044 54628
rect 8204 52162 8260 52164
rect 8204 52110 8206 52162
rect 8206 52110 8258 52162
rect 8258 52110 8260 52162
rect 8204 52108 8260 52110
rect 8092 50988 8148 51044
rect 8428 52444 8484 52500
rect 8428 51660 8484 51716
rect 8092 50764 8148 50820
rect 7868 49756 7924 49812
rect 7756 47570 7812 47572
rect 7756 47518 7758 47570
rect 7758 47518 7810 47570
rect 7810 47518 7812 47570
rect 7756 47516 7812 47518
rect 7532 46956 7588 47012
rect 7756 46732 7812 46788
rect 7980 48300 8036 48356
rect 7980 47458 8036 47460
rect 7980 47406 7982 47458
rect 7982 47406 8034 47458
rect 8034 47406 8036 47458
rect 7980 47404 8036 47406
rect 7868 46620 7924 46676
rect 7980 47180 8036 47236
rect 7980 46732 8036 46788
rect 7532 45500 7588 45556
rect 7420 45388 7476 45444
rect 7756 45052 7812 45108
rect 7532 44044 7588 44100
rect 7196 43148 7252 43204
rect 7084 42252 7140 42308
rect 7420 43426 7476 43428
rect 7420 43374 7422 43426
rect 7422 43374 7474 43426
rect 7474 43374 7476 43426
rect 7420 43372 7476 43374
rect 6972 42028 7028 42084
rect 6748 41132 6804 41188
rect 6860 41580 6916 41636
rect 6636 39564 6692 39620
rect 6860 40012 6916 40068
rect 6748 39116 6804 39172
rect 7084 41468 7140 41524
rect 7532 42476 7588 42532
rect 7420 42028 7476 42084
rect 7420 41804 7476 41860
rect 7308 41186 7364 41188
rect 7308 41134 7310 41186
rect 7310 41134 7362 41186
rect 7362 41134 7364 41186
rect 7308 41132 7364 41134
rect 7420 40124 7476 40180
rect 7308 39900 7364 39956
rect 7868 43484 7924 43540
rect 7756 41468 7812 41524
rect 7756 40908 7812 40964
rect 8428 51378 8484 51380
rect 8428 51326 8430 51378
rect 8430 51326 8482 51378
rect 8482 51326 8484 51378
rect 8428 51324 8484 51326
rect 8316 50594 8372 50596
rect 8316 50542 8318 50594
rect 8318 50542 8370 50594
rect 8370 50542 8372 50594
rect 8316 50540 8372 50542
rect 8652 52444 8708 52500
rect 8876 53452 8932 53508
rect 9436 56140 9492 56196
rect 10108 57260 10164 57316
rect 10108 56364 10164 56420
rect 9660 55468 9716 55524
rect 9548 55356 9604 55412
rect 10444 55468 10500 55524
rect 9884 55356 9940 55412
rect 9772 54460 9828 54516
rect 10444 55298 10500 55300
rect 10444 55246 10446 55298
rect 10446 55246 10498 55298
rect 10498 55246 10500 55298
rect 10444 55244 10500 55246
rect 9772 54290 9828 54292
rect 9772 54238 9774 54290
rect 9774 54238 9826 54290
rect 9826 54238 9828 54290
rect 9772 54236 9828 54238
rect 10220 54908 10276 54964
rect 9884 53900 9940 53956
rect 9660 53564 9716 53620
rect 9772 53452 9828 53508
rect 9324 53228 9380 53284
rect 9324 52780 9380 52836
rect 8988 52386 9044 52388
rect 8988 52334 8990 52386
rect 8990 52334 9042 52386
rect 9042 52334 9044 52386
rect 8988 52332 9044 52334
rect 9100 52220 9156 52276
rect 8876 51772 8932 51828
rect 8764 51548 8820 51604
rect 8764 50428 8820 50484
rect 8204 49980 8260 50036
rect 8316 49868 8372 49924
rect 8428 49532 8484 49588
rect 8316 49084 8372 49140
rect 8204 49026 8260 49028
rect 8204 48974 8206 49026
rect 8206 48974 8258 49026
rect 8258 48974 8260 49026
rect 8204 48972 8260 48974
rect 8204 47068 8260 47124
rect 8204 45500 8260 45556
rect 8092 45052 8148 45108
rect 8092 44716 8148 44772
rect 8204 44434 8260 44436
rect 8204 44382 8206 44434
rect 8206 44382 8258 44434
rect 8258 44382 8260 44434
rect 8204 44380 8260 44382
rect 8092 44322 8148 44324
rect 8092 44270 8094 44322
rect 8094 44270 8146 44322
rect 8146 44270 8148 44322
rect 8092 44268 8148 44270
rect 8204 44098 8260 44100
rect 8204 44046 8206 44098
rect 8206 44046 8258 44098
rect 8258 44046 8260 44098
rect 8204 44044 8260 44046
rect 8652 48300 8708 48356
rect 8764 49532 8820 49588
rect 8540 47516 8596 47572
rect 8652 46508 8708 46564
rect 9324 52332 9380 52388
rect 9548 51884 9604 51940
rect 9548 51548 9604 51604
rect 9548 51212 9604 51268
rect 9324 50204 9380 50260
rect 9324 49980 9380 50036
rect 9212 49420 9268 49476
rect 8876 48802 8932 48804
rect 8876 48750 8878 48802
rect 8878 48750 8930 48802
rect 8930 48750 8932 48802
rect 8876 48748 8932 48750
rect 9100 48860 9156 48916
rect 8988 47628 9044 47684
rect 9436 48972 9492 49028
rect 8988 47404 9044 47460
rect 9212 47180 9268 47236
rect 8764 46284 8820 46340
rect 8988 45666 9044 45668
rect 8988 45614 8990 45666
rect 8990 45614 9042 45666
rect 9042 45614 9044 45666
rect 8988 45612 9044 45614
rect 8652 45052 8708 45108
rect 9324 46956 9380 47012
rect 9212 46060 9268 46116
rect 9212 45836 9268 45892
rect 9212 45388 9268 45444
rect 8764 45276 8820 45332
rect 8540 44604 8596 44660
rect 8428 43932 8484 43988
rect 8764 43372 8820 43428
rect 8428 43148 8484 43204
rect 8204 43036 8260 43092
rect 8092 42588 8148 42644
rect 8428 42252 8484 42308
rect 8092 41410 8148 41412
rect 8092 41358 8094 41410
rect 8094 41358 8146 41410
rect 8146 41358 8148 41410
rect 8092 41356 8148 41358
rect 8316 40796 8372 40852
rect 8204 40348 8260 40404
rect 8988 43260 9044 43316
rect 8764 41916 8820 41972
rect 8876 42252 8932 42308
rect 9212 43036 9268 43092
rect 9324 43596 9380 43652
rect 9100 42252 9156 42308
rect 8988 42194 9044 42196
rect 8988 42142 8990 42194
rect 8990 42142 9042 42194
rect 9042 42142 9044 42194
rect 8988 42140 9044 42142
rect 9324 42140 9380 42196
rect 9436 44716 9492 44772
rect 8540 41244 8596 41300
rect 8764 41132 8820 41188
rect 6412 38220 6468 38276
rect 5852 36428 5908 36484
rect 5740 35756 5796 35812
rect 5852 35532 5908 35588
rect 5740 35196 5796 35252
rect 5964 35474 6020 35476
rect 5964 35422 5966 35474
rect 5966 35422 6018 35474
rect 6018 35422 6020 35474
rect 5964 35420 6020 35422
rect 5740 33740 5796 33796
rect 5852 34524 5908 34580
rect 6524 37548 6580 37604
rect 6076 34524 6132 34580
rect 6188 36092 6244 36148
rect 6076 34130 6132 34132
rect 6076 34078 6078 34130
rect 6078 34078 6130 34130
rect 6130 34078 6132 34130
rect 6076 34076 6132 34078
rect 5740 31948 5796 32004
rect 5628 31836 5684 31892
rect 5516 31500 5572 31556
rect 5292 30940 5348 30996
rect 5964 32396 6020 32452
rect 6412 35586 6468 35588
rect 6412 35534 6414 35586
rect 6414 35534 6466 35586
rect 6466 35534 6468 35586
rect 6412 35532 6468 35534
rect 6300 34076 6356 34132
rect 6188 31948 6244 32004
rect 6188 31388 6244 31444
rect 6412 33964 6468 34020
rect 6636 34748 6692 34804
rect 6524 33628 6580 33684
rect 6636 33458 6692 33460
rect 6636 33406 6638 33458
rect 6638 33406 6690 33458
rect 6690 33406 6692 33458
rect 6636 33404 6692 33406
rect 6636 32956 6692 33012
rect 6188 31106 6244 31108
rect 6188 31054 6190 31106
rect 6190 31054 6242 31106
rect 6242 31054 6244 31106
rect 6188 31052 6244 31054
rect 6412 31052 6468 31108
rect 5628 30210 5684 30212
rect 5628 30158 5630 30210
rect 5630 30158 5682 30210
rect 5682 30158 5684 30210
rect 5628 30156 5684 30158
rect 5180 29596 5236 29652
rect 5964 30604 6020 30660
rect 6076 30156 6132 30212
rect 5404 29484 5460 29540
rect 4956 29314 5012 29316
rect 4956 29262 4958 29314
rect 4958 29262 5010 29314
rect 5010 29262 5012 29314
rect 4956 29260 5012 29262
rect 4956 28754 5012 28756
rect 4956 28702 4958 28754
rect 4958 28702 5010 28754
rect 5010 28702 5012 28754
rect 4956 28700 5012 28702
rect 4396 28364 4452 28420
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 4172 28140 4228 28196
rect 3500 27858 3556 27860
rect 3500 27806 3502 27858
rect 3502 27806 3554 27858
rect 3554 27806 3556 27858
rect 3500 27804 3556 27806
rect 3724 27804 3780 27860
rect 3724 27356 3780 27412
rect 3948 27858 4004 27860
rect 3948 27806 3950 27858
rect 3950 27806 4002 27858
rect 4002 27806 4004 27858
rect 3948 27804 4004 27806
rect 3052 27244 3108 27300
rect 3164 27132 3220 27188
rect 2828 26796 2884 26852
rect 2492 26124 2548 26180
rect 3052 25900 3108 25956
rect 2492 24556 2548 24612
rect 2492 22540 2548 22596
rect 3612 27186 3668 27188
rect 3612 27134 3614 27186
rect 3614 27134 3666 27186
rect 3666 27134 3668 27186
rect 3612 27132 3668 27134
rect 3948 27244 4004 27300
rect 3948 26908 4004 26964
rect 3500 26572 3556 26628
rect 3276 25900 3332 25956
rect 3836 26796 3892 26852
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 4396 28028 4452 28084
rect 4396 27692 4452 27748
rect 4732 28140 4788 28196
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 4956 27468 5012 27524
rect 4620 27020 4676 27076
rect 4956 27186 5012 27188
rect 4956 27134 4958 27186
rect 4958 27134 5010 27186
rect 5010 27134 5012 27186
rect 4956 27132 5012 27134
rect 4956 26908 5012 26964
rect 4396 26572 4452 26628
rect 4956 26348 5012 26404
rect 4396 26290 4452 26292
rect 4396 26238 4398 26290
rect 4398 26238 4450 26290
rect 4450 26238 4452 26290
rect 4396 26236 4452 26238
rect 5068 26236 5124 26292
rect 4464 25898 4520 25900
rect 3836 25788 3892 25844
rect 4284 25788 4340 25844
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 4844 25788 4900 25844
rect 4620 25564 4676 25620
rect 3388 25452 3444 25508
rect 4172 25452 4228 25508
rect 3612 25340 3668 25396
rect 3388 25116 3444 25172
rect 3276 24722 3332 24724
rect 3276 24670 3278 24722
rect 3278 24670 3330 24722
rect 3330 24670 3332 24722
rect 3276 24668 3332 24670
rect 3164 24556 3220 24612
rect 2716 22652 2772 22708
rect 2828 23100 2884 23156
rect 2716 22258 2772 22260
rect 2716 22206 2718 22258
rect 2718 22206 2770 22258
rect 2770 22206 2772 22258
rect 2716 22204 2772 22206
rect 2828 22092 2884 22148
rect 2716 21698 2772 21700
rect 2716 21646 2718 21698
rect 2718 21646 2770 21698
rect 2770 21646 2772 21698
rect 2716 21644 2772 21646
rect 2380 20636 2436 20692
rect 2380 19234 2436 19236
rect 2380 19182 2382 19234
rect 2382 19182 2434 19234
rect 2434 19182 2436 19234
rect 2380 19180 2436 19182
rect 2044 18844 2100 18900
rect 2156 17666 2212 17668
rect 2156 17614 2158 17666
rect 2158 17614 2210 17666
rect 2210 17614 2212 17666
rect 2156 17612 2212 17614
rect 2268 16770 2324 16772
rect 2268 16718 2270 16770
rect 2270 16718 2322 16770
rect 2322 16718 2324 16770
rect 2268 16716 2324 16718
rect 1932 15708 1988 15764
rect 2156 16604 2212 16660
rect 1932 15260 1988 15316
rect 1484 15148 1540 15204
rect 1820 14642 1876 14644
rect 1820 14590 1822 14642
rect 1822 14590 1874 14642
rect 1874 14590 1876 14642
rect 1820 14588 1876 14590
rect 1596 14476 1652 14532
rect 1708 13858 1764 13860
rect 1708 13806 1710 13858
rect 1710 13806 1762 13858
rect 1762 13806 1764 13858
rect 1708 13804 1764 13806
rect 1148 12290 1204 12292
rect 1148 12238 1150 12290
rect 1150 12238 1202 12290
rect 1202 12238 1204 12290
rect 1148 12236 1204 12238
rect 1148 11900 1204 11956
rect 812 8316 868 8372
rect 364 7196 420 7252
rect 476 7532 532 7588
rect 252 6188 308 6244
rect 700 6972 756 7028
rect 476 3388 532 3444
rect 476 2604 532 2660
rect 812 3612 868 3668
rect 1260 11788 1316 11844
rect 1260 11564 1316 11620
rect 1372 10892 1428 10948
rect 1260 9042 1316 9044
rect 1260 8990 1262 9042
rect 1262 8990 1314 9042
rect 1314 8990 1316 9042
rect 1260 8988 1316 8990
rect 1260 7196 1316 7252
rect 1148 6860 1204 6916
rect 700 2828 756 2884
rect 1932 12178 1988 12180
rect 1932 12126 1934 12178
rect 1934 12126 1986 12178
rect 1986 12126 1988 12178
rect 1932 12124 1988 12126
rect 1820 11564 1876 11620
rect 1596 11506 1652 11508
rect 1596 11454 1598 11506
rect 1598 11454 1650 11506
rect 1650 11454 1652 11506
rect 1596 11452 1652 11454
rect 1596 11116 1652 11172
rect 2268 15708 2324 15764
rect 2492 18844 2548 18900
rect 2492 18620 2548 18676
rect 2492 15260 2548 15316
rect 2380 14754 2436 14756
rect 2380 14702 2382 14754
rect 2382 14702 2434 14754
rect 2434 14702 2436 14754
rect 2380 14700 2436 14702
rect 2268 14588 2324 14644
rect 2492 14642 2548 14644
rect 2492 14590 2494 14642
rect 2494 14590 2546 14642
rect 2546 14590 2548 14642
rect 2492 14588 2548 14590
rect 2156 14364 2212 14420
rect 3052 20860 3108 20916
rect 5964 29426 6020 29428
rect 5964 29374 5966 29426
rect 5966 29374 6018 29426
rect 6018 29374 6020 29426
rect 5964 29372 6020 29374
rect 5852 28924 5908 28980
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 6300 30044 6356 30100
rect 6412 29820 6468 29876
rect 6524 32508 6580 32564
rect 7308 38556 7364 38612
rect 6860 38444 6916 38500
rect 7084 38274 7140 38276
rect 7084 38222 7086 38274
rect 7086 38222 7138 38274
rect 7138 38222 7140 38274
rect 7084 38220 7140 38222
rect 6860 37100 6916 37156
rect 6860 36706 6916 36708
rect 6860 36654 6862 36706
rect 6862 36654 6914 36706
rect 6914 36654 6916 36706
rect 6860 36652 6916 36654
rect 7196 36706 7252 36708
rect 7196 36654 7198 36706
rect 7198 36654 7250 36706
rect 7250 36654 7252 36706
rect 7196 36652 7252 36654
rect 7532 38780 7588 38836
rect 7308 36540 7364 36596
rect 6972 36092 7028 36148
rect 7980 39452 8036 39508
rect 8204 39506 8260 39508
rect 8204 39454 8206 39506
rect 8206 39454 8258 39506
rect 8258 39454 8260 39506
rect 8204 39452 8260 39454
rect 7980 39004 8036 39060
rect 8204 38834 8260 38836
rect 8204 38782 8206 38834
rect 8206 38782 8258 38834
rect 8258 38782 8260 38834
rect 8204 38780 8260 38782
rect 7868 38668 7924 38724
rect 7756 38162 7812 38164
rect 7756 38110 7758 38162
rect 7758 38110 7810 38162
rect 7810 38110 7812 38162
rect 7756 38108 7812 38110
rect 8428 38668 8484 38724
rect 8540 39116 8596 39172
rect 8204 38050 8260 38052
rect 8204 37998 8206 38050
rect 8206 37998 8258 38050
rect 8258 37998 8260 38050
rect 8204 37996 8260 37998
rect 9324 41970 9380 41972
rect 9324 41918 9326 41970
rect 9326 41918 9378 41970
rect 9378 41918 9380 41970
rect 9324 41916 9380 41918
rect 9996 53730 10052 53732
rect 9996 53678 9998 53730
rect 9998 53678 10050 53730
rect 10050 53678 10052 53730
rect 9996 53676 10052 53678
rect 9772 51772 9828 51828
rect 10108 52556 10164 52612
rect 9996 51996 10052 52052
rect 10108 51884 10164 51940
rect 9884 50764 9940 50820
rect 9772 49756 9828 49812
rect 9772 49196 9828 49252
rect 9772 49026 9828 49028
rect 9772 48974 9774 49026
rect 9774 48974 9826 49026
rect 9826 48974 9828 49026
rect 9772 48972 9828 48974
rect 10108 49196 10164 49252
rect 10108 48636 10164 48692
rect 9884 48524 9940 48580
rect 9660 47404 9716 47460
rect 9772 48412 9828 48468
rect 10108 48188 10164 48244
rect 9884 47852 9940 47908
rect 10108 47570 10164 47572
rect 10108 47518 10110 47570
rect 10110 47518 10162 47570
rect 10162 47518 10164 47570
rect 10108 47516 10164 47518
rect 9884 47068 9940 47124
rect 10332 54684 10388 54740
rect 11452 56812 11508 56868
rect 11900 56812 11956 56868
rect 11676 56588 11732 56644
rect 10780 56476 10836 56532
rect 10668 55692 10724 55748
rect 10668 54572 10724 54628
rect 10556 54236 10612 54292
rect 10332 53452 10388 53508
rect 10668 53452 10724 53508
rect 11004 55916 11060 55972
rect 11564 55858 11620 55860
rect 11564 55806 11566 55858
rect 11566 55806 11618 55858
rect 11618 55806 11620 55858
rect 11564 55804 11620 55806
rect 11900 56588 11956 56644
rect 12348 56252 12404 56308
rect 13244 56700 13300 56756
rect 13468 56700 13524 56756
rect 13244 56252 13300 56308
rect 11788 55692 11844 55748
rect 11900 55298 11956 55300
rect 11900 55246 11902 55298
rect 11902 55246 11954 55298
rect 11954 55246 11956 55298
rect 11900 55244 11956 55246
rect 11452 54684 11508 54740
rect 10892 54460 10948 54516
rect 11004 54572 11060 54628
rect 11900 54572 11956 54628
rect 11004 53618 11060 53620
rect 11004 53566 11006 53618
rect 11006 53566 11058 53618
rect 11058 53566 11060 53618
rect 11004 53564 11060 53566
rect 11340 53564 11396 53620
rect 10780 53340 10836 53396
rect 10444 53228 10500 53284
rect 10332 49138 10388 49140
rect 10332 49086 10334 49138
rect 10334 49086 10386 49138
rect 10386 49086 10388 49138
rect 10332 49084 10388 49086
rect 10332 48636 10388 48692
rect 10332 46956 10388 47012
rect 9772 45836 9828 45892
rect 9884 45612 9940 45668
rect 9548 44604 9604 44660
rect 9996 45276 10052 45332
rect 9548 43820 9604 43876
rect 9548 43596 9604 43652
rect 9884 44994 9940 44996
rect 9884 44942 9886 44994
rect 9886 44942 9938 44994
rect 9938 44942 9940 44994
rect 9884 44940 9940 44942
rect 9884 44380 9940 44436
rect 9660 43484 9716 43540
rect 9772 44044 9828 44100
rect 9660 43036 9716 43092
rect 9660 42812 9716 42868
rect 10220 45276 10276 45332
rect 9996 43932 10052 43988
rect 9884 43596 9940 43652
rect 9996 43036 10052 43092
rect 9100 40908 9156 40964
rect 9324 41186 9380 41188
rect 9324 41134 9326 41186
rect 9326 41134 9378 41186
rect 9378 41134 9380 41186
rect 9324 41132 9380 41134
rect 9548 42140 9604 42196
rect 8316 37548 8372 37604
rect 8204 37212 8260 37268
rect 8540 37548 8596 37604
rect 7868 36876 7924 36932
rect 7756 36764 7812 36820
rect 7420 36092 7476 36148
rect 8092 36764 8148 36820
rect 8204 36988 8260 37044
rect 8316 36594 8372 36596
rect 8316 36542 8318 36594
rect 8318 36542 8370 36594
rect 8370 36542 8372 36594
rect 8316 36540 8372 36542
rect 8204 36370 8260 36372
rect 8204 36318 8206 36370
rect 8206 36318 8258 36370
rect 8258 36318 8260 36370
rect 8204 36316 8260 36318
rect 7196 35308 7252 35364
rect 7868 35420 7924 35476
rect 7420 35308 7476 35364
rect 7084 33346 7140 33348
rect 7084 33294 7086 33346
rect 7086 33294 7138 33346
rect 7138 33294 7140 33346
rect 7084 33292 7140 33294
rect 6860 32844 6916 32900
rect 6636 30604 6692 30660
rect 6636 30210 6692 30212
rect 6636 30158 6638 30210
rect 6638 30158 6690 30210
rect 6690 30158 6692 30210
rect 6636 30156 6692 30158
rect 6076 28700 6132 28756
rect 6636 28812 6692 28868
rect 5516 27580 5572 27636
rect 5740 27468 5796 27524
rect 5404 25788 5460 25844
rect 5628 25788 5684 25844
rect 5292 25564 5348 25620
rect 3804 25114 3860 25116
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4012 25060 4068 25062
rect 5180 25452 5236 25508
rect 3948 24556 4004 24612
rect 3948 24220 4004 24276
rect 3724 24162 3780 24164
rect 3724 24110 3726 24162
rect 3726 24110 3778 24162
rect 3778 24110 3780 24162
rect 3724 24108 3780 24110
rect 3836 23938 3892 23940
rect 3836 23886 3838 23938
rect 3838 23886 3890 23938
rect 3890 23886 3892 23938
rect 3836 23884 3892 23886
rect 3612 23548 3668 23604
rect 2716 20300 2772 20356
rect 2828 20748 2884 20804
rect 2716 20130 2772 20132
rect 2716 20078 2718 20130
rect 2718 20078 2770 20130
rect 2770 20078 2772 20130
rect 2716 20076 2772 20078
rect 2716 18732 2772 18788
rect 2716 16940 2772 16996
rect 3804 23546 3860 23548
rect 3276 23436 3332 23492
rect 3388 22930 3444 22932
rect 3388 22878 3390 22930
rect 3390 22878 3442 22930
rect 3442 22878 3444 22930
rect 3388 22876 3444 22878
rect 3388 22540 3444 22596
rect 3388 21868 3444 21924
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 5628 25340 5684 25396
rect 5292 25004 5348 25060
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4844 24332 4900 24388
rect 3612 23324 3668 23380
rect 4060 23266 4116 23268
rect 4060 23214 4062 23266
rect 4062 23214 4114 23266
rect 4114 23214 4116 23266
rect 4060 23212 4116 23214
rect 3724 22316 3780 22372
rect 4172 22930 4228 22932
rect 4172 22878 4174 22930
rect 4174 22878 4226 22930
rect 4226 22878 4228 22930
rect 4172 22876 4228 22878
rect 4732 23436 4788 23492
rect 5068 24108 5124 24164
rect 5516 25228 5572 25284
rect 5628 24780 5684 24836
rect 5516 24610 5572 24612
rect 5516 24558 5518 24610
rect 5518 24558 5570 24610
rect 5570 24558 5572 24610
rect 5516 24556 5572 24558
rect 5404 24108 5460 24164
rect 5068 23772 5124 23828
rect 4844 23100 4900 23156
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 4844 22652 4900 22708
rect 3948 22316 4004 22372
rect 3500 21084 3556 21140
rect 4956 22370 5012 22372
rect 4956 22318 4958 22370
rect 4958 22318 5010 22370
rect 5010 22318 5012 22370
rect 4956 22316 5012 22318
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 4172 21756 4228 21812
rect 3164 20636 3220 20692
rect 4060 21084 4116 21140
rect 4284 21698 4340 21700
rect 4284 21646 4286 21698
rect 4286 21646 4338 21698
rect 4338 21646 4340 21698
rect 4284 21644 4340 21646
rect 5068 21868 5124 21924
rect 5180 23154 5236 23156
rect 5180 23102 5182 23154
rect 5182 23102 5234 23154
rect 5234 23102 5236 23154
rect 5180 23100 5236 23102
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4672 21140 4728 21142
rect 4732 20914 4788 20916
rect 4732 20862 4734 20914
rect 4734 20862 4786 20914
rect 4786 20862 4788 20914
rect 4732 20860 4788 20862
rect 3276 20412 3332 20468
rect 3164 18338 3220 18340
rect 3164 18286 3166 18338
rect 3166 18286 3218 18338
rect 3218 18286 3220 18338
rect 3164 18284 3220 18286
rect 2716 15426 2772 15428
rect 2716 15374 2718 15426
rect 2718 15374 2770 15426
rect 2770 15374 2772 15426
rect 2716 15372 2772 15374
rect 2828 15820 2884 15876
rect 2156 14028 2212 14084
rect 2716 14028 2772 14084
rect 2380 13244 2436 13300
rect 2268 13186 2324 13188
rect 2268 13134 2270 13186
rect 2270 13134 2322 13186
rect 2322 13134 2324 13186
rect 2268 13132 2324 13134
rect 2268 12572 2324 12628
rect 2156 12348 2212 12404
rect 1932 10444 1988 10500
rect 1820 10220 1876 10276
rect 1708 9100 1764 9156
rect 2604 13522 2660 13524
rect 2604 13470 2606 13522
rect 2606 13470 2658 13522
rect 2658 13470 2660 13522
rect 2604 13468 2660 13470
rect 2492 12908 2548 12964
rect 2380 10220 2436 10276
rect 2492 11340 2548 11396
rect 1596 8316 1652 8372
rect 2156 9772 2212 9828
rect 1484 6860 1540 6916
rect 1596 7980 1652 8036
rect 1372 6300 1428 6356
rect 1372 6076 1428 6132
rect 1596 5964 1652 6020
rect 1708 8092 1764 8148
rect 1708 5180 1764 5236
rect 1820 7980 1876 8036
rect 2044 8482 2100 8484
rect 2044 8430 2046 8482
rect 2046 8430 2098 8482
rect 2098 8430 2100 8482
rect 2044 8428 2100 8430
rect 2044 8204 2100 8260
rect 1932 6802 1988 6804
rect 1932 6750 1934 6802
rect 1934 6750 1986 6802
rect 1986 6750 1988 6802
rect 1932 6748 1988 6750
rect 1820 4226 1876 4228
rect 1820 4174 1822 4226
rect 1822 4174 1874 4226
rect 1874 4174 1876 4226
rect 1820 4172 1876 4174
rect 1372 4060 1428 4116
rect 1372 3778 1428 3780
rect 1372 3726 1374 3778
rect 1374 3726 1426 3778
rect 1426 3726 1428 3778
rect 1372 3724 1428 3726
rect 1596 3554 1652 3556
rect 1596 3502 1598 3554
rect 1598 3502 1650 3554
rect 1650 3502 1652 3554
rect 1596 3500 1652 3502
rect 2268 7420 2324 7476
rect 2492 9826 2548 9828
rect 2492 9774 2494 9826
rect 2494 9774 2546 9826
rect 2546 9774 2548 9826
rect 2492 9772 2548 9774
rect 2380 6412 2436 6468
rect 2492 9548 2548 9604
rect 2380 5852 2436 5908
rect 2492 5292 2548 5348
rect 2268 4172 2324 4228
rect 2380 4844 2436 4900
rect 2380 4060 2436 4116
rect 2380 3554 2436 3556
rect 2380 3502 2382 3554
rect 2382 3502 2434 3554
rect 2434 3502 2436 3554
rect 2380 3500 2436 3502
rect 2268 2716 2324 2772
rect 1372 1708 1428 1764
rect 1932 1708 1988 1764
rect 2044 1932 2100 1988
rect 1148 1484 1204 1540
rect 1036 1202 1092 1204
rect 1036 1150 1038 1202
rect 1038 1150 1090 1202
rect 1090 1150 1092 1202
rect 1036 1148 1092 1150
rect 1596 1484 1652 1540
rect 1372 1090 1428 1092
rect 1372 1038 1374 1090
rect 1374 1038 1426 1090
rect 1426 1038 1428 1090
rect 1372 1036 1428 1038
rect 1820 1202 1876 1204
rect 1820 1150 1822 1202
rect 1822 1150 1874 1202
rect 1874 1150 1876 1202
rect 1820 1148 1876 1150
rect 2828 12012 2884 12068
rect 3164 16492 3220 16548
rect 3052 15372 3108 15428
rect 3052 14028 3108 14084
rect 3388 18508 3444 18564
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3612 20076 3668 20132
rect 3948 19964 4004 20020
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 4396 19964 4452 20020
rect 4956 20412 5012 20468
rect 4844 19964 4900 20020
rect 4396 19740 4452 19796
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 5180 21532 5236 21588
rect 5292 23772 5348 23828
rect 5628 23884 5684 23940
rect 5404 21756 5460 21812
rect 5180 21084 5236 21140
rect 4284 18844 4340 18900
rect 4620 18732 4676 18788
rect 4172 18508 4228 18564
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 5292 20972 5348 21028
rect 5516 20802 5572 20804
rect 5516 20750 5518 20802
rect 5518 20750 5570 20802
rect 5570 20750 5572 20802
rect 5516 20748 5572 20750
rect 4464 18058 4520 18060
rect 3612 17836 3668 17892
rect 4284 17948 4340 18004
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 3948 17666 4004 17668
rect 3948 17614 3950 17666
rect 3950 17614 4002 17666
rect 4002 17614 4004 17666
rect 3948 17612 4004 17614
rect 3612 17500 3668 17556
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 5068 17948 5124 18004
rect 4396 17388 4452 17444
rect 4732 17388 4788 17444
rect 4284 17164 4340 17220
rect 3388 16716 3444 16772
rect 3724 16492 3780 16548
rect 4172 16658 4228 16660
rect 4172 16606 4174 16658
rect 4174 16606 4226 16658
rect 4226 16606 4228 16658
rect 4172 16604 4228 16606
rect 4060 16492 4116 16548
rect 4464 16490 4520 16492
rect 3388 16380 3444 16436
rect 3612 16380 3668 16436
rect 3276 15820 3332 15876
rect 3164 15260 3220 15316
rect 3052 13468 3108 13524
rect 2940 11004 2996 11060
rect 2716 9548 2772 9604
rect 2716 8540 2772 8596
rect 2828 7644 2884 7700
rect 2828 6018 2884 6020
rect 2828 5966 2830 6018
rect 2830 5966 2882 6018
rect 2882 5966 2884 6018
rect 2828 5964 2884 5966
rect 3052 8930 3108 8932
rect 3052 8878 3054 8930
rect 3054 8878 3106 8930
rect 3106 8878 3108 8930
rect 3052 8876 3108 8878
rect 3052 8428 3108 8484
rect 3276 14700 3332 14756
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 4172 16380 4228 16436
rect 3500 15708 3556 15764
rect 4060 16098 4116 16100
rect 4060 16046 4062 16098
rect 4062 16046 4114 16098
rect 4114 16046 4116 16098
rect 4060 16044 4116 16046
rect 3612 15596 3668 15652
rect 3804 15706 3860 15708
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 4172 15484 4228 15540
rect 3612 15260 3668 15316
rect 3948 15202 4004 15204
rect 3948 15150 3950 15202
rect 3950 15150 4002 15202
rect 4002 15150 4004 15202
rect 3948 15148 4004 15150
rect 4060 14924 4116 14980
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 4620 14754 4676 14756
rect 4620 14702 4622 14754
rect 4622 14702 4674 14754
rect 4674 14702 4676 14754
rect 4620 14700 4676 14702
rect 4956 16098 5012 16100
rect 4956 16046 4958 16098
rect 4958 16046 5010 16098
rect 5010 16046 5012 16098
rect 4956 16044 5012 16046
rect 4956 15820 5012 15876
rect 5404 17948 5460 18004
rect 6076 28140 6132 28196
rect 5964 27634 6020 27636
rect 5964 27582 5966 27634
rect 5966 27582 6018 27634
rect 6018 27582 6020 27634
rect 5964 27580 6020 27582
rect 5852 26236 5908 26292
rect 5852 25116 5908 25172
rect 6188 27580 6244 27636
rect 6188 26348 6244 26404
rect 6300 27132 6356 27188
rect 6412 27020 6468 27076
rect 6636 26796 6692 26852
rect 6748 28588 6804 28644
rect 6076 25900 6132 25956
rect 6076 25340 6132 25396
rect 6188 24780 6244 24836
rect 6300 25564 6356 25620
rect 6412 25004 6468 25060
rect 6076 24162 6132 24164
rect 6076 24110 6078 24162
rect 6078 24110 6130 24162
rect 6130 24110 6132 24162
rect 6076 24108 6132 24110
rect 5964 23772 6020 23828
rect 5852 21420 5908 21476
rect 7756 34914 7812 34916
rect 7756 34862 7758 34914
rect 7758 34862 7810 34914
rect 7810 34862 7812 34914
rect 7756 34860 7812 34862
rect 7532 33404 7588 33460
rect 6860 27804 6916 27860
rect 7308 31836 7364 31892
rect 6860 27244 6916 27300
rect 7196 30940 7252 30996
rect 6972 27074 7028 27076
rect 6972 27022 6974 27074
rect 6974 27022 7026 27074
rect 7026 27022 7028 27074
rect 6972 27020 7028 27022
rect 7084 30156 7140 30212
rect 6860 26684 6916 26740
rect 7196 27356 7252 27412
rect 7756 33740 7812 33796
rect 7756 32284 7812 32340
rect 7644 32172 7700 32228
rect 8092 35026 8148 35028
rect 8092 34974 8094 35026
rect 8094 34974 8146 35026
rect 8146 34974 8148 35026
rect 8092 34972 8148 34974
rect 7980 34748 8036 34804
rect 8092 34076 8148 34132
rect 8428 34524 8484 34580
rect 8428 33964 8484 34020
rect 8428 33068 8484 33124
rect 7980 32786 8036 32788
rect 7980 32734 7982 32786
rect 7982 32734 8034 32786
rect 8034 32734 8036 32786
rect 7980 32732 8036 32734
rect 8204 32284 8260 32340
rect 8428 32396 8484 32452
rect 7868 32060 7924 32116
rect 7420 30156 7476 30212
rect 7644 31500 7700 31556
rect 7420 29820 7476 29876
rect 7980 31836 8036 31892
rect 7980 30604 8036 30660
rect 7868 30380 7924 30436
rect 7756 30210 7812 30212
rect 7756 30158 7758 30210
rect 7758 30158 7810 30210
rect 7810 30158 7812 30210
rect 7756 30156 7812 30158
rect 7868 29820 7924 29876
rect 8204 31388 8260 31444
rect 8316 31500 8372 31556
rect 8652 35868 8708 35924
rect 8652 33740 8708 33796
rect 8876 39788 8932 39844
rect 10668 53228 10724 53284
rect 10556 52668 10612 52724
rect 10556 51548 10612 51604
rect 11004 52780 11060 52836
rect 10668 51212 10724 51268
rect 10556 48972 10612 49028
rect 10668 49756 10724 49812
rect 11900 54348 11956 54404
rect 12460 55020 12516 55076
rect 12796 55020 12852 55076
rect 12124 54908 12180 54964
rect 11788 53004 11844 53060
rect 12012 53676 12068 53732
rect 11676 52780 11732 52836
rect 11004 49644 11060 49700
rect 11116 51996 11172 52052
rect 12684 54124 12740 54180
rect 12460 53730 12516 53732
rect 12460 53678 12462 53730
rect 12462 53678 12514 53730
rect 12514 53678 12516 53730
rect 12460 53676 12516 53678
rect 12684 53676 12740 53732
rect 12348 52892 12404 52948
rect 13020 54684 13076 54740
rect 13132 54572 13188 54628
rect 11788 52108 11844 52164
rect 11452 51436 11508 51492
rect 11340 50594 11396 50596
rect 11340 50542 11342 50594
rect 11342 50542 11394 50594
rect 11394 50542 11396 50594
rect 11340 50540 11396 50542
rect 11340 50316 11396 50372
rect 11116 48636 11172 48692
rect 11340 49532 11396 49588
rect 10668 47964 10724 48020
rect 10556 46562 10612 46564
rect 10556 46510 10558 46562
rect 10558 46510 10610 46562
rect 10610 46510 10612 46562
rect 10556 46508 10612 46510
rect 10668 46396 10724 46452
rect 11004 48188 11060 48244
rect 11228 48242 11284 48244
rect 11228 48190 11230 48242
rect 11230 48190 11282 48242
rect 11282 48190 11284 48242
rect 11228 48188 11284 48190
rect 11676 51996 11732 52052
rect 11564 48524 11620 48580
rect 11676 50876 11732 50932
rect 11116 47740 11172 47796
rect 11228 47628 11284 47684
rect 11452 47628 11508 47684
rect 11788 49810 11844 49812
rect 11788 49758 11790 49810
rect 11790 49758 11842 49810
rect 11842 49758 11844 49810
rect 11788 49756 11844 49758
rect 11004 46396 11060 46452
rect 11004 45890 11060 45892
rect 11004 45838 11006 45890
rect 11006 45838 11058 45890
rect 11058 45838 11060 45890
rect 11004 45836 11060 45838
rect 10668 45666 10724 45668
rect 10668 45614 10670 45666
rect 10670 45614 10722 45666
rect 10722 45614 10724 45666
rect 10668 45612 10724 45614
rect 10332 44828 10388 44884
rect 10332 44044 10388 44100
rect 10108 42476 10164 42532
rect 10220 43260 10276 43316
rect 9660 41746 9716 41748
rect 9660 41694 9662 41746
rect 9662 41694 9714 41746
rect 9714 41694 9716 41746
rect 9660 41692 9716 41694
rect 9660 41244 9716 41300
rect 9324 40348 9380 40404
rect 8988 38556 9044 38612
rect 8876 38162 8932 38164
rect 8876 38110 8878 38162
rect 8878 38110 8930 38162
rect 8930 38110 8932 38162
rect 8876 38108 8932 38110
rect 9212 38722 9268 38724
rect 9212 38670 9214 38722
rect 9214 38670 9266 38722
rect 9266 38670 9268 38722
rect 9212 38668 9268 38670
rect 8876 37548 8932 37604
rect 9212 38108 9268 38164
rect 9324 38050 9380 38052
rect 9324 37998 9326 38050
rect 9326 37998 9378 38050
rect 9378 37998 9380 38050
rect 9324 37996 9380 37998
rect 8876 36316 8932 36372
rect 9772 41186 9828 41188
rect 9772 41134 9774 41186
rect 9774 41134 9826 41186
rect 9826 41134 9828 41186
rect 9772 41132 9828 41134
rect 9772 39676 9828 39732
rect 9884 38892 9940 38948
rect 9772 38668 9828 38724
rect 9548 38444 9604 38500
rect 9660 37548 9716 37604
rect 8988 35980 9044 36036
rect 8988 35586 9044 35588
rect 8988 35534 8990 35586
rect 8990 35534 9042 35586
rect 9042 35534 9044 35586
rect 8988 35532 9044 35534
rect 8764 34412 8820 34468
rect 8876 32844 8932 32900
rect 8988 32508 9044 32564
rect 8764 32172 8820 32228
rect 8540 31276 8596 31332
rect 8540 30994 8596 30996
rect 8540 30942 8542 30994
rect 8542 30942 8594 30994
rect 8594 30942 8596 30994
rect 8540 30940 8596 30942
rect 8876 31276 8932 31332
rect 8428 30604 8484 30660
rect 8204 30098 8260 30100
rect 8204 30046 8206 30098
rect 8206 30046 8258 30098
rect 8258 30046 8260 30098
rect 8204 30044 8260 30046
rect 8316 29986 8372 29988
rect 8316 29934 8318 29986
rect 8318 29934 8370 29986
rect 8370 29934 8372 29986
rect 8316 29932 8372 29934
rect 8092 29820 8148 29876
rect 7420 28924 7476 28980
rect 7532 28476 7588 28532
rect 8204 28642 8260 28644
rect 8204 28590 8206 28642
rect 8206 28590 8258 28642
rect 8258 28590 8260 28642
rect 8204 28588 8260 28590
rect 7980 28140 8036 28196
rect 7868 27916 7924 27972
rect 7756 27804 7812 27860
rect 7980 27468 8036 27524
rect 7980 27186 8036 27188
rect 7980 27134 7982 27186
rect 7982 27134 8034 27186
rect 8034 27134 8036 27186
rect 7980 27132 8036 27134
rect 7868 27020 7924 27076
rect 7756 26796 7812 26852
rect 7308 26684 7364 26740
rect 7644 26684 7700 26740
rect 7196 26124 7252 26180
rect 7084 25900 7140 25956
rect 6972 25618 7028 25620
rect 6972 25566 6974 25618
rect 6974 25566 7026 25618
rect 7026 25566 7028 25618
rect 6972 25564 7028 25566
rect 6860 24834 6916 24836
rect 6860 24782 6862 24834
rect 6862 24782 6914 24834
rect 6914 24782 6916 24834
rect 6860 24780 6916 24782
rect 6524 24108 6580 24164
rect 6748 23660 6804 23716
rect 6860 23548 6916 23604
rect 6412 23212 6468 23268
rect 6972 23212 7028 23268
rect 6188 21532 6244 21588
rect 6524 23100 6580 23156
rect 6748 21474 6804 21476
rect 6748 21422 6750 21474
rect 6750 21422 6802 21474
rect 6802 21422 6804 21474
rect 6748 21420 6804 21422
rect 7420 26124 7476 26180
rect 7308 25788 7364 25844
rect 7756 25788 7812 25844
rect 7868 26460 7924 26516
rect 9884 37212 9940 37268
rect 9324 36876 9380 36932
rect 9212 36706 9268 36708
rect 9212 36654 9214 36706
rect 9214 36654 9266 36706
rect 9266 36654 9268 36706
rect 9212 36652 9268 36654
rect 9660 37042 9716 37044
rect 9660 36990 9662 37042
rect 9662 36990 9714 37042
rect 9714 36990 9716 37042
rect 9660 36988 9716 36990
rect 9772 36876 9828 36932
rect 9660 36764 9716 36820
rect 9436 36428 9492 36484
rect 9436 35868 9492 35924
rect 9548 36316 9604 36372
rect 9324 34748 9380 34804
rect 9212 32732 9268 32788
rect 9212 32562 9268 32564
rect 9212 32510 9214 32562
rect 9214 32510 9266 32562
rect 9266 32510 9268 32562
rect 9212 32508 9268 32510
rect 9212 32172 9268 32228
rect 9436 32450 9492 32452
rect 9436 32398 9438 32450
rect 9438 32398 9490 32450
rect 9490 32398 9492 32450
rect 9436 32396 9492 32398
rect 9324 31836 9380 31892
rect 9772 34188 9828 34244
rect 10668 44380 10724 44436
rect 10780 44044 10836 44100
rect 10892 45500 10948 45556
rect 10668 43932 10724 43988
rect 11788 46396 11844 46452
rect 11340 44716 11396 44772
rect 11116 43932 11172 43988
rect 10780 43650 10836 43652
rect 10780 43598 10782 43650
rect 10782 43598 10834 43650
rect 10834 43598 10836 43650
rect 10780 43596 10836 43598
rect 11004 43596 11060 43652
rect 11340 43650 11396 43652
rect 11340 43598 11342 43650
rect 11342 43598 11394 43650
rect 11394 43598 11396 43650
rect 11340 43596 11396 43598
rect 10444 43372 10500 43428
rect 10556 43484 10612 43540
rect 11676 45164 11732 45220
rect 11564 44994 11620 44996
rect 11564 44942 11566 44994
rect 11566 44942 11618 44994
rect 11618 44942 11620 44994
rect 11564 44940 11620 44942
rect 11564 44716 11620 44772
rect 12012 51996 12068 52052
rect 12124 51490 12180 51492
rect 12124 51438 12126 51490
rect 12126 51438 12178 51490
rect 12178 51438 12180 51490
rect 12124 51436 12180 51438
rect 12460 52162 12516 52164
rect 12460 52110 12462 52162
rect 12462 52110 12514 52162
rect 12514 52110 12516 52162
rect 12460 52108 12516 52110
rect 12908 52108 12964 52164
rect 12348 51324 12404 51380
rect 12684 51660 12740 51716
rect 12460 51212 12516 51268
rect 12796 51266 12852 51268
rect 12796 51214 12798 51266
rect 12798 51214 12850 51266
rect 12850 51214 12852 51266
rect 12796 51212 12852 51214
rect 12236 51154 12292 51156
rect 12236 51102 12238 51154
rect 12238 51102 12290 51154
rect 12290 51102 12292 51154
rect 12236 51100 12292 51102
rect 12684 50988 12740 51044
rect 12460 50876 12516 50932
rect 12348 50818 12404 50820
rect 12348 50766 12350 50818
rect 12350 50766 12402 50818
rect 12402 50766 12404 50818
rect 12348 50764 12404 50766
rect 12012 50652 12068 50708
rect 12236 49980 12292 50036
rect 12460 50540 12516 50596
rect 12236 49698 12292 49700
rect 12236 49646 12238 49698
rect 12238 49646 12290 49698
rect 12290 49646 12292 49698
rect 12236 49644 12292 49646
rect 12012 49532 12068 49588
rect 11900 45164 11956 45220
rect 12012 47404 12068 47460
rect 11676 44268 11732 44324
rect 11452 43484 11508 43540
rect 11228 43426 11284 43428
rect 11228 43374 11230 43426
rect 11230 43374 11282 43426
rect 11282 43374 11284 43426
rect 11228 43372 11284 43374
rect 11564 43260 11620 43316
rect 10556 42476 10612 42532
rect 10444 42028 10500 42084
rect 10332 41804 10388 41860
rect 10332 41298 10388 41300
rect 10332 41246 10334 41298
rect 10334 41246 10386 41298
rect 10386 41246 10388 41298
rect 10332 41244 10388 41246
rect 10220 40460 10276 40516
rect 10332 41020 10388 41076
rect 9996 36876 10052 36932
rect 10108 39788 10164 39844
rect 10332 38834 10388 38836
rect 10332 38782 10334 38834
rect 10334 38782 10386 38834
rect 10386 38782 10388 38834
rect 10332 38780 10388 38782
rect 10892 42252 10948 42308
rect 11788 42588 11844 42644
rect 11004 41916 11060 41972
rect 11116 42252 11172 42308
rect 10668 41244 10724 41300
rect 10668 39676 10724 39732
rect 10892 40124 10948 40180
rect 10108 36764 10164 36820
rect 10780 38668 10836 38724
rect 10108 36370 10164 36372
rect 10108 36318 10110 36370
rect 10110 36318 10162 36370
rect 10162 36318 10164 36370
rect 10108 36316 10164 36318
rect 10556 38050 10612 38052
rect 10556 37998 10558 38050
rect 10558 37998 10610 38050
rect 10610 37998 10612 38050
rect 10556 37996 10612 37998
rect 10332 37266 10388 37268
rect 10332 37214 10334 37266
rect 10334 37214 10386 37266
rect 10386 37214 10388 37266
rect 10332 37212 10388 37214
rect 10444 36988 10500 37044
rect 10444 36092 10500 36148
rect 10556 35756 10612 35812
rect 9884 33740 9940 33796
rect 9996 34802 10052 34804
rect 9996 34750 9998 34802
rect 9998 34750 10050 34802
rect 10050 34750 10052 34802
rect 9996 34748 10052 34750
rect 11788 42028 11844 42084
rect 11340 41580 11396 41636
rect 11340 40908 11396 40964
rect 12124 47292 12180 47348
rect 12124 46284 12180 46340
rect 12460 46396 12516 46452
rect 12124 44994 12180 44996
rect 12124 44942 12126 44994
rect 12126 44942 12178 44994
rect 12178 44942 12180 44994
rect 12124 44940 12180 44942
rect 12460 45836 12516 45892
rect 12348 44716 12404 44772
rect 12236 43932 12292 43988
rect 12236 43372 12292 43428
rect 12124 43314 12180 43316
rect 12124 43262 12126 43314
rect 12126 43262 12178 43314
rect 12178 43262 12180 43314
rect 12124 43260 12180 43262
rect 12124 42700 12180 42756
rect 12236 42642 12292 42644
rect 12236 42590 12238 42642
rect 12238 42590 12290 42642
rect 12290 42590 12292 42642
rect 12236 42588 12292 42590
rect 12124 42476 12180 42532
rect 12012 42028 12068 42084
rect 12348 42028 12404 42084
rect 12124 41970 12180 41972
rect 12124 41918 12126 41970
rect 12126 41918 12178 41970
rect 12178 41918 12180 41970
rect 12124 41916 12180 41918
rect 12012 41580 12068 41636
rect 13244 53900 13300 53956
rect 13356 53004 13412 53060
rect 13020 51996 13076 52052
rect 13132 52332 13188 52388
rect 13244 52220 13300 52276
rect 13244 51884 13300 51940
rect 14140 57036 14196 57092
rect 13692 54796 13748 54852
rect 13804 55244 13860 55300
rect 13692 53564 13748 53620
rect 14588 56028 14644 56084
rect 14140 54290 14196 54292
rect 14140 54238 14142 54290
rect 14142 54238 14194 54290
rect 14194 54238 14196 54290
rect 14140 54236 14196 54238
rect 14028 53340 14084 53396
rect 13916 53116 13972 53172
rect 13580 52722 13636 52724
rect 13580 52670 13582 52722
rect 13582 52670 13634 52722
rect 13634 52670 13636 52722
rect 13580 52668 13636 52670
rect 14140 52668 14196 52724
rect 13580 51212 13636 51268
rect 13468 51100 13524 51156
rect 13468 49644 13524 49700
rect 13580 49586 13636 49588
rect 13580 49534 13582 49586
rect 13582 49534 13634 49586
rect 13634 49534 13636 49586
rect 13580 49532 13636 49534
rect 12684 48412 12740 48468
rect 12796 48748 12852 48804
rect 12684 47516 12740 47572
rect 13020 47458 13076 47460
rect 13020 47406 13022 47458
rect 13022 47406 13074 47458
rect 13074 47406 13076 47458
rect 13020 47404 13076 47406
rect 12908 46508 12964 46564
rect 13804 51324 13860 51380
rect 15036 55916 15092 55972
rect 14476 55410 14532 55412
rect 14476 55358 14478 55410
rect 14478 55358 14530 55410
rect 14530 55358 14532 55410
rect 14476 55356 14532 55358
rect 14924 54572 14980 54628
rect 14924 54348 14980 54404
rect 15372 55244 15428 55300
rect 15484 54572 15540 54628
rect 15820 55410 15876 55412
rect 15820 55358 15822 55410
rect 15822 55358 15874 55410
rect 15874 55358 15876 55410
rect 15820 55356 15876 55358
rect 15596 55020 15652 55076
rect 15148 54290 15204 54292
rect 15148 54238 15150 54290
rect 15150 54238 15202 54290
rect 15202 54238 15204 54290
rect 15148 54236 15204 54238
rect 14476 54124 14532 54180
rect 15036 53676 15092 53732
rect 14364 52556 14420 52612
rect 14252 51884 14308 51940
rect 14476 52220 14532 52276
rect 13804 50652 13860 50708
rect 14140 50540 14196 50596
rect 15148 53004 15204 53060
rect 14700 51660 14756 51716
rect 15148 52556 15204 52612
rect 15260 52668 15316 52724
rect 15484 52556 15540 52612
rect 16044 54572 16100 54628
rect 15820 54290 15876 54292
rect 15820 54238 15822 54290
rect 15822 54238 15874 54290
rect 15874 54238 15876 54290
rect 15820 54236 15876 54238
rect 15932 53900 15988 53956
rect 15708 53676 15764 53732
rect 15820 53452 15876 53508
rect 15708 53058 15764 53060
rect 15708 53006 15710 53058
rect 15710 53006 15762 53058
rect 15762 53006 15764 53058
rect 15708 53004 15764 53006
rect 16828 56364 16884 56420
rect 16828 55970 16884 55972
rect 16828 55918 16830 55970
rect 16830 55918 16882 55970
rect 16882 55918 16884 55970
rect 16828 55916 16884 55918
rect 16380 54908 16436 54964
rect 17164 55858 17220 55860
rect 17164 55806 17166 55858
rect 17166 55806 17218 55858
rect 17218 55806 17220 55858
rect 17164 55804 17220 55806
rect 16716 55020 16772 55076
rect 17164 55020 17220 55076
rect 16828 54908 16884 54964
rect 16492 54796 16548 54852
rect 16380 54572 16436 54628
rect 18620 56700 18676 56756
rect 18844 56700 18900 56756
rect 18172 56588 18228 56644
rect 17724 56476 17780 56532
rect 18620 56476 18676 56532
rect 17612 56364 17668 56420
rect 17500 55410 17556 55412
rect 17500 55358 17502 55410
rect 17502 55358 17554 55410
rect 17554 55358 17556 55410
rect 17500 55356 17556 55358
rect 18172 56028 18228 56084
rect 17948 55468 18004 55524
rect 17612 55244 17668 55300
rect 17836 55244 17892 55300
rect 17388 55020 17444 55076
rect 17276 54572 17332 54628
rect 18732 56252 18788 56308
rect 18508 55020 18564 55076
rect 18284 54460 18340 54516
rect 18508 54402 18564 54404
rect 18508 54350 18510 54402
rect 18510 54350 18562 54402
rect 18562 54350 18564 54402
rect 18508 54348 18564 54350
rect 16268 54236 16324 54292
rect 16940 53452 16996 53508
rect 16492 53116 16548 53172
rect 16044 52946 16100 52948
rect 16044 52894 16046 52946
rect 16046 52894 16098 52946
rect 16098 52894 16100 52946
rect 16044 52892 16100 52894
rect 15932 52780 15988 52836
rect 15148 52162 15204 52164
rect 15148 52110 15150 52162
rect 15150 52110 15202 52162
rect 15202 52110 15204 52162
rect 15148 52108 15204 52110
rect 15932 52162 15988 52164
rect 15932 52110 15934 52162
rect 15934 52110 15986 52162
rect 15986 52110 15988 52162
rect 15932 52108 15988 52110
rect 15708 51436 15764 51492
rect 15036 51378 15092 51380
rect 15036 51326 15038 51378
rect 15038 51326 15090 51378
rect 15090 51326 15092 51378
rect 15036 51324 15092 51326
rect 14588 50652 14644 50708
rect 14476 50594 14532 50596
rect 14476 50542 14478 50594
rect 14478 50542 14530 50594
rect 14530 50542 14532 50594
rect 14476 50540 14532 50542
rect 14140 49868 14196 49924
rect 13692 48188 13748 48244
rect 13692 48018 13748 48020
rect 13692 47966 13694 48018
rect 13694 47966 13746 48018
rect 13746 47966 13748 48018
rect 13692 47964 13748 47966
rect 13356 47516 13412 47572
rect 13468 47852 13524 47908
rect 13468 47292 13524 47348
rect 13692 47068 13748 47124
rect 13132 45836 13188 45892
rect 13132 45666 13188 45668
rect 13132 45614 13134 45666
rect 13134 45614 13186 45666
rect 13186 45614 13188 45666
rect 13132 45612 13188 45614
rect 13244 45106 13300 45108
rect 13244 45054 13246 45106
rect 13246 45054 13298 45106
rect 13298 45054 13300 45106
rect 13244 45052 13300 45054
rect 12796 44716 12852 44772
rect 12684 43708 12740 43764
rect 12684 43260 12740 43316
rect 13580 46562 13636 46564
rect 13580 46510 13582 46562
rect 13582 46510 13634 46562
rect 13634 46510 13636 46562
rect 13580 46508 13636 46510
rect 14028 47852 14084 47908
rect 13916 47740 13972 47796
rect 13804 46732 13860 46788
rect 13804 46284 13860 46340
rect 13356 44716 13412 44772
rect 13132 44380 13188 44436
rect 12796 42140 12852 42196
rect 12908 42028 12964 42084
rect 13020 41804 13076 41860
rect 12796 41468 12852 41524
rect 12796 41132 12852 41188
rect 12236 40684 12292 40740
rect 11900 39676 11956 39732
rect 11788 39228 11844 39284
rect 11900 39116 11956 39172
rect 11788 39058 11844 39060
rect 11788 39006 11790 39058
rect 11790 39006 11842 39058
rect 11842 39006 11844 39058
rect 11788 39004 11844 39006
rect 11004 38668 11060 38724
rect 11004 38162 11060 38164
rect 11004 38110 11006 38162
rect 11006 38110 11058 38162
rect 11058 38110 11060 38162
rect 11004 38108 11060 38110
rect 12124 38274 12180 38276
rect 12124 38222 12126 38274
rect 12126 38222 12178 38274
rect 12178 38222 12180 38274
rect 12124 38220 12180 38222
rect 11564 38108 11620 38164
rect 11340 37772 11396 37828
rect 11228 37548 11284 37604
rect 11004 36482 11060 36484
rect 11004 36430 11006 36482
rect 11006 36430 11058 36482
rect 11058 36430 11060 36482
rect 11004 36428 11060 36430
rect 10556 34242 10612 34244
rect 10556 34190 10558 34242
rect 10558 34190 10610 34242
rect 10610 34190 10612 34242
rect 10556 34188 10612 34190
rect 11340 36764 11396 36820
rect 11116 35308 11172 35364
rect 9996 33852 10052 33908
rect 9884 33458 9940 33460
rect 9884 33406 9886 33458
rect 9886 33406 9938 33458
rect 9938 33406 9940 33458
rect 9884 33404 9940 33406
rect 9884 32732 9940 32788
rect 9772 32396 9828 32452
rect 10556 32956 10612 33012
rect 10332 32060 10388 32116
rect 10780 33516 10836 33572
rect 11004 34076 11060 34132
rect 11004 33906 11060 33908
rect 11004 33854 11006 33906
rect 11006 33854 11058 33906
rect 11058 33854 11060 33906
rect 11004 33852 11060 33854
rect 9660 31836 9716 31892
rect 9212 30940 9268 30996
rect 9548 31388 9604 31444
rect 8764 30604 8820 30660
rect 8764 29708 8820 29764
rect 8988 30044 9044 30100
rect 8988 29372 9044 29428
rect 9436 30492 9492 30548
rect 9324 30434 9380 30436
rect 9324 30382 9326 30434
rect 9326 30382 9378 30434
rect 9378 30382 9380 30434
rect 9324 30380 9380 30382
rect 9996 31388 10052 31444
rect 9884 30994 9940 30996
rect 9884 30942 9886 30994
rect 9886 30942 9938 30994
rect 9938 30942 9940 30994
rect 9884 30940 9940 30942
rect 9772 30210 9828 30212
rect 9772 30158 9774 30210
rect 9774 30158 9826 30210
rect 9826 30158 9828 30210
rect 9772 30156 9828 30158
rect 9660 29820 9716 29876
rect 8764 28700 8820 28756
rect 9884 29426 9940 29428
rect 9884 29374 9886 29426
rect 9886 29374 9938 29426
rect 9938 29374 9940 29426
rect 9884 29372 9940 29374
rect 8876 27916 8932 27972
rect 9100 28252 9156 28308
rect 8540 27746 8596 27748
rect 8540 27694 8542 27746
rect 8542 27694 8594 27746
rect 8594 27694 8596 27746
rect 8540 27692 8596 27694
rect 8876 27746 8932 27748
rect 8876 27694 8878 27746
rect 8878 27694 8930 27746
rect 8930 27694 8932 27746
rect 8876 27692 8932 27694
rect 8428 27580 8484 27636
rect 8988 27132 9044 27188
rect 8428 26460 8484 26516
rect 8092 26236 8148 26292
rect 8316 26236 8372 26292
rect 7420 25506 7476 25508
rect 7420 25454 7422 25506
rect 7422 25454 7474 25506
rect 7474 25454 7476 25506
rect 7420 25452 7476 25454
rect 7532 25394 7588 25396
rect 7532 25342 7534 25394
rect 7534 25342 7586 25394
rect 7586 25342 7588 25394
rect 7532 25340 7588 25342
rect 7868 25618 7924 25620
rect 7868 25566 7870 25618
rect 7870 25566 7922 25618
rect 7922 25566 7924 25618
rect 7868 25564 7924 25566
rect 7756 25228 7812 25284
rect 7644 24722 7700 24724
rect 7644 24670 7646 24722
rect 7646 24670 7698 24722
rect 7698 24670 7700 24722
rect 7644 24668 7700 24670
rect 7756 24556 7812 24612
rect 7308 23660 7364 23716
rect 7420 23884 7476 23940
rect 7868 23884 7924 23940
rect 7756 23548 7812 23604
rect 7868 23660 7924 23716
rect 7420 23100 7476 23156
rect 7196 22764 7252 22820
rect 7980 23100 8036 23156
rect 8204 25900 8260 25956
rect 8764 26124 8820 26180
rect 8988 26124 9044 26180
rect 8764 25452 8820 25508
rect 7532 22540 7588 22596
rect 6972 21308 7028 21364
rect 7084 21980 7140 22036
rect 5964 20412 6020 20468
rect 6300 20412 6356 20468
rect 6524 20748 6580 20804
rect 6188 20188 6244 20244
rect 5740 20018 5796 20020
rect 5740 19966 5742 20018
rect 5742 19966 5794 20018
rect 5794 19966 5796 20018
rect 5740 19964 5796 19966
rect 5852 19628 5908 19684
rect 5852 19404 5908 19460
rect 5964 19292 6020 19348
rect 6076 19180 6132 19236
rect 6300 19964 6356 20020
rect 5852 18508 5908 18564
rect 5628 18060 5684 18116
rect 5740 17890 5796 17892
rect 5740 17838 5742 17890
rect 5742 17838 5794 17890
rect 5794 17838 5796 17890
rect 5740 17836 5796 17838
rect 5404 16994 5460 16996
rect 5404 16942 5406 16994
rect 5406 16942 5458 16994
rect 5458 16942 5460 16994
rect 5404 16940 5460 16942
rect 5628 17724 5684 17780
rect 5852 17612 5908 17668
rect 5516 16380 5572 16436
rect 5516 15372 5572 15428
rect 5740 15596 5796 15652
rect 5180 15260 5236 15316
rect 5292 15202 5348 15204
rect 5292 15150 5294 15202
rect 5294 15150 5346 15202
rect 5346 15150 5348 15202
rect 5292 15148 5348 15150
rect 5180 14700 5236 14756
rect 5292 14924 5348 14980
rect 6076 18732 6132 18788
rect 6188 18396 6244 18452
rect 5964 16940 6020 16996
rect 6412 18508 6468 18564
rect 5964 16604 6020 16660
rect 5964 15596 6020 15652
rect 4956 14476 5012 14532
rect 3836 14252 3892 14308
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 3500 13916 3556 13972
rect 4172 14028 4228 14084
rect 3948 13132 4004 13188
rect 3500 13074 3556 13076
rect 3500 13022 3502 13074
rect 3502 13022 3554 13074
rect 3554 13022 3556 13074
rect 3500 13020 3556 13022
rect 3388 12460 3444 12516
rect 3276 12236 3332 12292
rect 3276 11900 3332 11956
rect 4844 14252 4900 14308
rect 4732 14140 4788 14196
rect 5628 14476 5684 14532
rect 5180 14252 5236 14308
rect 4732 13580 4788 13636
rect 5180 14028 5236 14084
rect 5404 14028 5460 14084
rect 5292 13468 5348 13524
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 5068 13356 5124 13412
rect 4620 13020 4676 13076
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4508 12572 4564 12628
rect 4012 12516 4068 12518
rect 4396 12460 4452 12516
rect 3612 11900 3668 11956
rect 3724 12124 3780 12180
rect 3500 11788 3556 11844
rect 3388 10386 3444 10388
rect 3388 10334 3390 10386
rect 3390 10334 3442 10386
rect 3442 10334 3444 10386
rect 3388 10332 3444 10334
rect 3724 11228 3780 11284
rect 4172 12012 4228 12068
rect 4508 12236 4564 12292
rect 4956 12290 5012 12292
rect 4956 12238 4958 12290
rect 4958 12238 5010 12290
rect 5010 12238 5012 12290
rect 4956 12236 5012 12238
rect 5852 14530 5908 14532
rect 5852 14478 5854 14530
rect 5854 14478 5906 14530
rect 5906 14478 5908 14530
rect 5852 14476 5908 14478
rect 6076 16044 6132 16100
rect 6076 14924 6132 14980
rect 6076 14642 6132 14644
rect 6076 14590 6078 14642
rect 6078 14590 6130 14642
rect 6130 14590 6132 14642
rect 6076 14588 6132 14590
rect 6076 14252 6132 14308
rect 5740 12460 5796 12516
rect 5180 12124 5236 12180
rect 5628 12124 5684 12180
rect 4844 12012 4900 12068
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4172 11228 4228 11284
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4396 11004 4452 11060
rect 4012 10948 4068 10950
rect 4172 10892 4228 10948
rect 3612 10610 3668 10612
rect 3612 10558 3614 10610
rect 3614 10558 3666 10610
rect 3666 10558 3668 10610
rect 3612 10556 3668 10558
rect 4172 10220 4228 10276
rect 3388 9884 3444 9940
rect 3500 8876 3556 8932
rect 3948 9826 4004 9828
rect 3948 9774 3950 9826
rect 3950 9774 4002 9826
rect 4002 9774 4004 9826
rect 3948 9772 4004 9774
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 3612 8764 3668 8820
rect 3948 8876 4004 8932
rect 3612 8370 3668 8372
rect 3612 8318 3614 8370
rect 3614 8318 3666 8370
rect 3666 8318 3668 8370
rect 3612 8316 3668 8318
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4732 9938 4788 9940
rect 4732 9886 4734 9938
rect 4734 9886 4786 9938
rect 4786 9886 4788 9938
rect 4732 9884 4788 9886
rect 4284 9548 4340 9604
rect 4396 9324 4452 9380
rect 4284 8876 4340 8932
rect 4284 8540 4340 8596
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 4508 8258 4564 8260
rect 4508 8206 4510 8258
rect 4510 8206 4562 8258
rect 4562 8206 4564 8258
rect 4508 8204 4564 8206
rect 3388 7980 3444 8036
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4956 11564 5012 11620
rect 5180 11564 5236 11620
rect 5068 10556 5124 10612
rect 5180 11340 5236 11396
rect 3164 7698 3220 7700
rect 3164 7646 3166 7698
rect 3166 7646 3218 7698
rect 3218 7646 3220 7698
rect 3164 7644 3220 7646
rect 5068 10386 5124 10388
rect 5068 10334 5070 10386
rect 5070 10334 5122 10386
rect 5122 10334 5124 10386
rect 5068 10332 5124 10334
rect 6300 16380 6356 16436
rect 6300 16098 6356 16100
rect 6300 16046 6302 16098
rect 6302 16046 6354 16098
rect 6354 16046 6356 16098
rect 6300 16044 6356 16046
rect 6188 13468 6244 13524
rect 6188 13020 6244 13076
rect 6524 18450 6580 18452
rect 6524 18398 6526 18450
rect 6526 18398 6578 18450
rect 6578 18398 6580 18450
rect 6524 18396 6580 18398
rect 6636 19964 6692 20020
rect 6636 18172 6692 18228
rect 6524 17164 6580 17220
rect 8428 25228 8484 25284
rect 9212 25228 9268 25284
rect 8988 24162 9044 24164
rect 8988 24110 8990 24162
rect 8990 24110 9042 24162
rect 9042 24110 9044 24162
rect 8988 24108 9044 24110
rect 9324 23938 9380 23940
rect 9324 23886 9326 23938
rect 9326 23886 9378 23938
rect 9378 23886 9380 23938
rect 9324 23884 9380 23886
rect 9324 23660 9380 23716
rect 8092 22652 8148 22708
rect 7196 21308 7252 21364
rect 7532 21586 7588 21588
rect 7532 21534 7534 21586
rect 7534 21534 7586 21586
rect 7586 21534 7588 21586
rect 7532 21532 7588 21534
rect 7196 19740 7252 19796
rect 7196 19180 7252 19236
rect 6972 17666 7028 17668
rect 6972 17614 6974 17666
rect 6974 17614 7026 17666
rect 7026 17614 7028 17666
rect 6972 17612 7028 17614
rect 6972 17276 7028 17332
rect 7084 17052 7140 17108
rect 6860 16322 6916 16324
rect 6860 16270 6862 16322
rect 6862 16270 6914 16322
rect 6914 16270 6916 16322
rect 6860 16268 6916 16270
rect 7308 18450 7364 18452
rect 7308 18398 7310 18450
rect 7310 18398 7362 18450
rect 7362 18398 7364 18450
rect 7308 18396 7364 18398
rect 7756 21756 7812 21812
rect 7868 21420 7924 21476
rect 8316 21868 8372 21924
rect 8204 21644 8260 21700
rect 8092 21308 8148 21364
rect 8092 20636 8148 20692
rect 7756 19740 7812 19796
rect 7532 17612 7588 17668
rect 7644 19068 7700 19124
rect 7532 16716 7588 16772
rect 7420 16658 7476 16660
rect 7420 16606 7422 16658
rect 7422 16606 7474 16658
rect 7474 16606 7476 16658
rect 7420 16604 7476 16606
rect 7420 16322 7476 16324
rect 7420 16270 7422 16322
rect 7422 16270 7474 16322
rect 7474 16270 7476 16322
rect 7420 16268 7476 16270
rect 7756 16828 7812 16884
rect 7868 18060 7924 18116
rect 6524 15372 6580 15428
rect 6636 15314 6692 15316
rect 6636 15262 6638 15314
rect 6638 15262 6690 15314
rect 6690 15262 6692 15314
rect 6636 15260 6692 15262
rect 6748 15090 6804 15092
rect 6748 15038 6750 15090
rect 6750 15038 6802 15090
rect 6802 15038 6804 15090
rect 6748 15036 6804 15038
rect 7308 16044 7364 16100
rect 6860 14924 6916 14980
rect 7084 14924 7140 14980
rect 6636 14588 6692 14644
rect 6636 13580 6692 13636
rect 6748 13692 6804 13748
rect 7196 14588 7252 14644
rect 7084 14252 7140 14308
rect 8204 19234 8260 19236
rect 8204 19182 8206 19234
rect 8206 19182 8258 19234
rect 8258 19182 8260 19234
rect 8204 19180 8260 19182
rect 8204 18508 8260 18564
rect 7980 17164 8036 17220
rect 7868 14588 7924 14644
rect 7980 16940 8036 16996
rect 8092 15596 8148 15652
rect 7084 13692 7140 13748
rect 6748 13356 6804 13412
rect 6636 13244 6692 13300
rect 6972 13132 7028 13188
rect 6300 12460 6356 12516
rect 5852 12012 5908 12068
rect 5964 11676 6020 11732
rect 5292 11228 5348 11284
rect 5852 11506 5908 11508
rect 5852 11454 5854 11506
rect 5854 11454 5906 11506
rect 5906 11454 5908 11506
rect 6524 12012 6580 12068
rect 5852 11452 5908 11454
rect 6300 11900 6356 11956
rect 6748 12908 6804 12964
rect 6300 11452 6356 11508
rect 5628 11004 5684 11060
rect 5628 10780 5684 10836
rect 5292 10556 5348 10612
rect 5516 10610 5572 10612
rect 5516 10558 5518 10610
rect 5518 10558 5570 10610
rect 5570 10558 5572 10610
rect 5516 10556 5572 10558
rect 5292 10386 5348 10388
rect 5292 10334 5294 10386
rect 5294 10334 5346 10386
rect 5346 10334 5348 10386
rect 5292 10332 5348 10334
rect 5292 10108 5348 10164
rect 5292 9826 5348 9828
rect 5292 9774 5294 9826
rect 5294 9774 5346 9826
rect 5346 9774 5348 9826
rect 5292 9772 5348 9774
rect 5180 8876 5236 8932
rect 5292 8652 5348 8708
rect 5292 8316 5348 8372
rect 5180 8258 5236 8260
rect 5180 8206 5182 8258
rect 5182 8206 5234 8258
rect 5234 8206 5236 8258
rect 5180 8204 5236 8206
rect 3612 7362 3668 7364
rect 3612 7310 3614 7362
rect 3614 7310 3666 7362
rect 3666 7310 3668 7362
rect 3612 7308 3668 7310
rect 3388 6972 3444 7028
rect 3948 7474 4004 7476
rect 3948 7422 3950 7474
rect 3950 7422 4002 7474
rect 4002 7422 4004 7474
rect 3948 7420 4004 7422
rect 4172 7308 4228 7364
rect 5964 10610 6020 10612
rect 5964 10558 5966 10610
rect 5966 10558 6018 10610
rect 6018 10558 6020 10610
rect 5964 10556 6020 10558
rect 6076 10444 6132 10500
rect 5852 8876 5908 8932
rect 6300 10780 6356 10836
rect 6076 10220 6132 10276
rect 6300 10220 6356 10276
rect 5628 8428 5684 8484
rect 5740 8764 5796 8820
rect 4396 7362 4452 7364
rect 4396 7310 4398 7362
rect 4398 7310 4450 7362
rect 4450 7310 4452 7362
rect 4396 7308 4452 7310
rect 5516 8204 5572 8260
rect 4284 7084 4340 7140
rect 4844 7196 4900 7252
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 4172 6412 4228 6468
rect 3388 6300 3444 6356
rect 2716 5122 2772 5124
rect 2716 5070 2718 5122
rect 2718 5070 2770 5122
rect 2770 5070 2772 5122
rect 2716 5068 2772 5070
rect 2940 4956 2996 5012
rect 2604 4508 2660 4564
rect 2940 4562 2996 4564
rect 2940 4510 2942 4562
rect 2942 4510 2994 4562
rect 2994 4510 2996 4562
rect 2940 4508 2996 4510
rect 2716 4060 2772 4116
rect 3276 4284 3332 4340
rect 3804 6298 3860 6300
rect 3500 6188 3556 6244
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 4060 5852 4116 5908
rect 3836 5682 3892 5684
rect 3836 5630 3838 5682
rect 3838 5630 3890 5682
rect 3890 5630 3892 5682
rect 3836 5628 3892 5630
rect 3612 5122 3668 5124
rect 3612 5070 3614 5122
rect 3614 5070 3666 5122
rect 3666 5070 3668 5122
rect 3612 5068 3668 5070
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 3948 4508 4004 4564
rect 3724 4338 3780 4340
rect 3724 4286 3726 4338
rect 3726 4286 3778 4338
rect 3778 4286 3780 4338
rect 3724 4284 3780 4286
rect 3500 3948 3556 4004
rect 4620 6690 4676 6692
rect 4620 6638 4622 6690
rect 4622 6638 4674 6690
rect 4674 6638 4676 6690
rect 4620 6636 4676 6638
rect 4956 7084 5012 7140
rect 4284 6300 4340 6356
rect 4844 5964 4900 6020
rect 4464 5514 4520 5516
rect 4284 5404 4340 5460
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4396 4620 4452 4676
rect 4620 4396 4676 4452
rect 4508 4284 4564 4340
rect 5628 7474 5684 7476
rect 5628 7422 5630 7474
rect 5630 7422 5682 7474
rect 5682 7422 5684 7474
rect 5628 7420 5684 7422
rect 5404 7084 5460 7140
rect 5628 7084 5684 7140
rect 5292 6972 5348 7028
rect 5516 6524 5572 6580
rect 5180 6412 5236 6468
rect 5292 6300 5348 6356
rect 5180 5740 5236 5796
rect 5180 5516 5236 5572
rect 5628 6300 5684 6356
rect 6076 8764 6132 8820
rect 5964 8204 6020 8260
rect 5852 6412 5908 6468
rect 6636 11564 6692 11620
rect 6636 10444 6692 10500
rect 6412 9772 6468 9828
rect 6300 8428 6356 8484
rect 6972 12124 7028 12180
rect 7196 12460 7252 12516
rect 6748 9772 6804 9828
rect 6972 11506 7028 11508
rect 6972 11454 6974 11506
rect 6974 11454 7026 11506
rect 7026 11454 7028 11506
rect 6972 11452 7028 11454
rect 6860 10556 6916 10612
rect 7084 10780 7140 10836
rect 6972 9548 7028 9604
rect 6972 9212 7028 9268
rect 6636 9100 6692 9156
rect 6636 8428 6692 8484
rect 6748 8876 6804 8932
rect 6524 8316 6580 8372
rect 6300 7644 6356 7700
rect 5964 5852 6020 5908
rect 6188 6300 6244 6356
rect 5852 5740 5908 5796
rect 5516 5068 5572 5124
rect 4172 3948 4228 4004
rect 3500 3388 3556 3444
rect 3276 3276 3332 3332
rect 2716 2380 2772 2436
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 3388 2828 3444 2884
rect 3724 2770 3780 2772
rect 3724 2718 3726 2770
rect 3726 2718 3778 2770
rect 3778 2718 3780 2770
rect 3724 2716 3780 2718
rect 3164 2156 3220 2212
rect 3276 2044 3332 2100
rect 2604 1260 2660 1316
rect 2940 1372 2996 1428
rect 2044 588 2100 644
rect 2492 588 2548 644
rect 4060 2268 4116 2324
rect 3612 1820 3668 1876
rect 3388 1596 3444 1652
rect 3276 476 3332 532
rect 3388 1148 3444 1204
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 5068 3388 5124 3444
rect 4508 2940 4564 2996
rect 4508 2716 4564 2772
rect 5068 2716 5124 2772
rect 4284 2380 4340 2436
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 5068 2268 5124 2324
rect 4732 2098 4788 2100
rect 4732 2046 4734 2098
rect 4734 2046 4786 2098
rect 4786 2046 4788 2098
rect 4732 2044 4788 2046
rect 4396 1484 4452 1540
rect 3500 924 3556 980
rect 4508 1820 4564 1876
rect 4844 1202 4900 1204
rect 4844 1150 4846 1202
rect 4846 1150 4898 1202
rect 4898 1150 4900 1202
rect 4844 1148 4900 1150
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 5180 2156 5236 2212
rect 5180 978 5236 980
rect 5180 926 5182 978
rect 5182 926 5234 978
rect 5234 926 5236 978
rect 5180 924 5236 926
rect 5180 700 5236 756
rect 5740 5068 5796 5124
rect 5628 4732 5684 4788
rect 5628 3836 5684 3892
rect 5964 3052 6020 3108
rect 6412 7532 6468 7588
rect 6412 6860 6468 6916
rect 6412 6412 6468 6468
rect 6636 6524 6692 6580
rect 6636 6300 6692 6356
rect 6412 6076 6468 6132
rect 6300 4844 6356 4900
rect 6748 5516 6804 5572
rect 6636 5404 6692 5460
rect 7868 13916 7924 13972
rect 7420 13746 7476 13748
rect 7420 13694 7422 13746
rect 7422 13694 7474 13746
rect 7474 13694 7476 13746
rect 7420 13692 7476 13694
rect 7756 13132 7812 13188
rect 8092 14812 8148 14868
rect 8540 23042 8596 23044
rect 8540 22990 8542 23042
rect 8542 22990 8594 23042
rect 8594 22990 8596 23042
rect 8540 22988 8596 22990
rect 9212 23436 9268 23492
rect 8540 17106 8596 17108
rect 8540 17054 8542 17106
rect 8542 17054 8594 17106
rect 8594 17054 8596 17106
rect 8540 17052 8596 17054
rect 8316 14028 8372 14084
rect 8428 14588 8484 14644
rect 8204 13746 8260 13748
rect 8204 13694 8206 13746
rect 8206 13694 8258 13746
rect 8258 13694 8260 13746
rect 8204 13692 8260 13694
rect 8428 13468 8484 13524
rect 8316 13244 8372 13300
rect 7532 12962 7588 12964
rect 7532 12910 7534 12962
rect 7534 12910 7586 12962
rect 7586 12910 7588 12962
rect 7532 12908 7588 12910
rect 7420 12348 7476 12404
rect 7644 12012 7700 12068
rect 7644 10610 7700 10612
rect 7644 10558 7646 10610
rect 7646 10558 7698 10610
rect 7698 10558 7700 10610
rect 7644 10556 7700 10558
rect 7644 10332 7700 10388
rect 7420 9826 7476 9828
rect 7420 9774 7422 9826
rect 7422 9774 7474 9826
rect 7474 9774 7476 9826
rect 7420 9772 7476 9774
rect 7308 9042 7364 9044
rect 7308 8990 7310 9042
rect 7310 8990 7362 9042
rect 7362 8990 7364 9042
rect 7308 8988 7364 8990
rect 7420 8818 7476 8820
rect 7420 8766 7422 8818
rect 7422 8766 7474 8818
rect 7474 8766 7476 8818
rect 7420 8764 7476 8766
rect 6972 8204 7028 8260
rect 7196 6972 7252 7028
rect 6972 6524 7028 6580
rect 7084 6748 7140 6804
rect 6860 5404 6916 5460
rect 6972 6300 7028 6356
rect 6300 4226 6356 4228
rect 6300 4174 6302 4226
rect 6302 4174 6354 4226
rect 6354 4174 6356 4226
rect 6300 4172 6356 4174
rect 6524 3948 6580 4004
rect 6412 2210 6468 2212
rect 6412 2158 6414 2210
rect 6414 2158 6466 2210
rect 6466 2158 6468 2210
rect 6412 2156 6468 2158
rect 6188 2044 6244 2100
rect 6076 1596 6132 1652
rect 5404 364 5460 420
rect 5628 1148 5684 1204
rect 7308 6412 7364 6468
rect 8092 13020 8148 13076
rect 8204 11788 8260 11844
rect 8204 11618 8260 11620
rect 8204 11566 8206 11618
rect 8206 11566 8258 11618
rect 8258 11566 8260 11618
rect 8204 11564 8260 11566
rect 8092 10220 8148 10276
rect 8204 11228 8260 11284
rect 8764 21586 8820 21588
rect 8764 21534 8766 21586
rect 8766 21534 8818 21586
rect 8818 21534 8820 21586
rect 8764 21532 8820 21534
rect 9212 21308 9268 21364
rect 9884 28476 9940 28532
rect 10220 30940 10276 30996
rect 10332 31612 10388 31668
rect 10332 30380 10388 30436
rect 10220 30210 10276 30212
rect 10220 30158 10222 30210
rect 10222 30158 10274 30210
rect 10274 30158 10276 30210
rect 10220 30156 10276 30158
rect 10332 30044 10388 30100
rect 10332 28530 10388 28532
rect 10332 28478 10334 28530
rect 10334 28478 10386 28530
rect 10386 28478 10388 28530
rect 10332 28476 10388 28478
rect 9996 28252 10052 28308
rect 10108 28364 10164 28420
rect 9660 27468 9716 27524
rect 9548 27020 9604 27076
rect 9548 26684 9604 26740
rect 9772 26514 9828 26516
rect 9772 26462 9774 26514
rect 9774 26462 9826 26514
rect 9826 26462 9828 26514
rect 9772 26460 9828 26462
rect 9660 26290 9716 26292
rect 9660 26238 9662 26290
rect 9662 26238 9714 26290
rect 9714 26238 9716 26290
rect 9660 26236 9716 26238
rect 9772 26178 9828 26180
rect 9772 26126 9774 26178
rect 9774 26126 9826 26178
rect 9826 26126 9828 26178
rect 9772 26124 9828 26126
rect 9548 23548 9604 23604
rect 9884 25228 9940 25284
rect 10108 27298 10164 27300
rect 10108 27246 10110 27298
rect 10110 27246 10162 27298
rect 10162 27246 10164 27298
rect 10108 27244 10164 27246
rect 9996 25452 10052 25508
rect 9772 24780 9828 24836
rect 10332 27692 10388 27748
rect 10108 25900 10164 25956
rect 9772 24220 9828 24276
rect 9772 23154 9828 23156
rect 9772 23102 9774 23154
rect 9774 23102 9826 23154
rect 9826 23102 9828 23154
rect 9772 23100 9828 23102
rect 9884 22988 9940 23044
rect 9996 23660 10052 23716
rect 9436 21980 9492 22036
rect 9548 21532 9604 21588
rect 9548 21084 9604 21140
rect 9660 22652 9716 22708
rect 8764 20748 8820 20804
rect 9212 20636 9268 20692
rect 9324 20748 9380 20804
rect 8988 18060 9044 18116
rect 8876 17836 8932 17892
rect 8652 12796 8708 12852
rect 8764 17612 8820 17668
rect 9212 20076 9268 20132
rect 9212 19458 9268 19460
rect 9212 19406 9214 19458
rect 9214 19406 9266 19458
rect 9266 19406 9268 19458
rect 9212 19404 9268 19406
rect 10332 26178 10388 26180
rect 10332 26126 10334 26178
rect 10334 26126 10386 26178
rect 10386 26126 10388 26178
rect 10332 26124 10388 26126
rect 10220 25004 10276 25060
rect 10892 32060 10948 32116
rect 11004 33068 11060 33124
rect 10780 31948 10836 32004
rect 10668 30044 10724 30100
rect 10780 31276 10836 31332
rect 10556 29932 10612 29988
rect 10892 30380 10948 30436
rect 10892 29820 10948 29876
rect 10780 28924 10836 28980
rect 10892 28812 10948 28868
rect 10668 28252 10724 28308
rect 10668 27074 10724 27076
rect 10668 27022 10670 27074
rect 10670 27022 10722 27074
rect 10722 27022 10724 27074
rect 10668 27020 10724 27022
rect 10892 28252 10948 28308
rect 10780 27244 10836 27300
rect 10780 26908 10836 26964
rect 10892 27580 10948 27636
rect 10444 23772 10500 23828
rect 10220 22652 10276 22708
rect 9884 22092 9940 22148
rect 9772 21586 9828 21588
rect 9772 21534 9774 21586
rect 9774 21534 9826 21586
rect 9826 21534 9828 21586
rect 9772 21532 9828 21534
rect 9660 20860 9716 20916
rect 9436 19964 9492 20020
rect 9772 20636 9828 20692
rect 9884 19852 9940 19908
rect 9996 21980 10052 22036
rect 9772 19740 9828 19796
rect 9324 18450 9380 18452
rect 9324 18398 9326 18450
rect 9326 18398 9378 18450
rect 9378 18398 9380 18450
rect 9324 18396 9380 18398
rect 9100 17666 9156 17668
rect 9100 17614 9102 17666
rect 9102 17614 9154 17666
rect 9154 17614 9156 17666
rect 9100 17612 9156 17614
rect 8764 17276 8820 17332
rect 8540 12684 8596 12740
rect 8652 12460 8708 12516
rect 8428 11228 8484 11284
rect 8316 10556 8372 10612
rect 8428 10892 8484 10948
rect 8204 9996 8260 10052
rect 7868 9548 7924 9604
rect 7756 9100 7812 9156
rect 7868 8876 7924 8932
rect 7756 7868 7812 7924
rect 7644 7250 7700 7252
rect 7644 7198 7646 7250
rect 7646 7198 7698 7250
rect 7698 7198 7700 7250
rect 7644 7196 7700 7198
rect 8316 9548 8372 9604
rect 8540 10610 8596 10612
rect 8540 10558 8542 10610
rect 8542 10558 8594 10610
rect 8594 10558 8596 10610
rect 8540 10556 8596 10558
rect 8652 9884 8708 9940
rect 8652 8930 8708 8932
rect 8652 8878 8654 8930
rect 8654 8878 8706 8930
rect 8706 8878 8708 8930
rect 8652 8876 8708 8878
rect 8428 8764 8484 8820
rect 8652 8204 8708 8260
rect 8428 7644 8484 7700
rect 7980 6860 8036 6916
rect 8316 7196 8372 7252
rect 7868 6524 7924 6580
rect 7196 5740 7252 5796
rect 7084 5180 7140 5236
rect 6972 4226 7028 4228
rect 6972 4174 6974 4226
rect 6974 4174 7026 4226
rect 7026 4174 7028 4226
rect 6972 4172 7028 4174
rect 7420 5794 7476 5796
rect 7420 5742 7422 5794
rect 7422 5742 7474 5794
rect 7474 5742 7476 5794
rect 7420 5740 7476 5742
rect 7308 5068 7364 5124
rect 7308 4732 7364 4788
rect 7644 5516 7700 5572
rect 8092 5404 8148 5460
rect 8204 6860 8260 6916
rect 7980 5346 8036 5348
rect 7980 5294 7982 5346
rect 7982 5294 8034 5346
rect 8034 5294 8036 5346
rect 7980 5292 8036 5294
rect 7980 5122 8036 5124
rect 7980 5070 7982 5122
rect 7982 5070 8034 5122
rect 8034 5070 8036 5122
rect 7980 5068 8036 5070
rect 7308 4172 7364 4228
rect 7756 4620 7812 4676
rect 7196 3500 7252 3556
rect 6636 2716 6692 2772
rect 6860 2658 6916 2660
rect 6860 2606 6862 2658
rect 6862 2606 6914 2658
rect 6914 2606 6916 2658
rect 6860 2604 6916 2606
rect 6636 2044 6692 2100
rect 7308 2604 7364 2660
rect 7308 2156 7364 2212
rect 7196 1596 7252 1652
rect 6972 1484 7028 1540
rect 6860 1148 6916 1204
rect 7532 4226 7588 4228
rect 7532 4174 7534 4226
rect 7534 4174 7586 4226
rect 7586 4174 7588 4226
rect 7532 4172 7588 4174
rect 7420 1596 7476 1652
rect 7532 3948 7588 4004
rect 7644 3666 7700 3668
rect 7644 3614 7646 3666
rect 7646 3614 7698 3666
rect 7698 3614 7700 3666
rect 7644 3612 7700 3614
rect 7868 3724 7924 3780
rect 8092 4172 8148 4228
rect 8316 4060 8372 4116
rect 8092 3948 8148 4004
rect 7532 700 7588 756
rect 7308 252 7364 308
rect 7196 140 7252 196
rect 7756 252 7812 308
rect 7980 3164 8036 3220
rect 8092 2770 8148 2772
rect 8092 2718 8094 2770
rect 8094 2718 8146 2770
rect 8146 2718 8148 2770
rect 8092 2716 8148 2718
rect 8652 7586 8708 7588
rect 8652 7534 8654 7586
rect 8654 7534 8706 7586
rect 8706 7534 8708 7586
rect 8652 7532 8708 7534
rect 9324 17388 9380 17444
rect 8988 16994 9044 16996
rect 8988 16942 8990 16994
rect 8990 16942 9042 16994
rect 9042 16942 9044 16994
rect 8988 16940 9044 16942
rect 8876 16828 8932 16884
rect 8988 16380 9044 16436
rect 9660 18732 9716 18788
rect 9436 16268 9492 16324
rect 9548 18060 9604 18116
rect 9772 18172 9828 18228
rect 9884 19292 9940 19348
rect 9996 18732 10052 18788
rect 10556 26684 10612 26740
rect 10556 21980 10612 22036
rect 10668 26460 10724 26516
rect 10780 25900 10836 25956
rect 10556 21698 10612 21700
rect 10556 21646 10558 21698
rect 10558 21646 10610 21698
rect 10610 21646 10612 21698
rect 10556 21644 10612 21646
rect 10780 23100 10836 23156
rect 10668 20914 10724 20916
rect 10668 20862 10670 20914
rect 10670 20862 10722 20914
rect 10722 20862 10724 20914
rect 10668 20860 10724 20862
rect 10556 20412 10612 20468
rect 10892 22652 10948 22708
rect 11340 32956 11396 33012
rect 11452 34860 11508 34916
rect 11452 32562 11508 32564
rect 11452 32510 11454 32562
rect 11454 32510 11506 32562
rect 11506 32510 11508 32562
rect 11452 32508 11508 32510
rect 11228 29372 11284 29428
rect 11452 28924 11508 28980
rect 11340 28252 11396 28308
rect 11452 27020 11508 27076
rect 11004 22316 11060 22372
rect 11116 23884 11172 23940
rect 11340 25228 11396 25284
rect 11228 22988 11284 23044
rect 11340 22370 11396 22372
rect 11340 22318 11342 22370
rect 11342 22318 11394 22370
rect 11394 22318 11396 22370
rect 11340 22316 11396 22318
rect 11116 21756 11172 21812
rect 10780 20412 10836 20468
rect 10892 21532 10948 21588
rect 10332 19794 10388 19796
rect 10332 19742 10334 19794
rect 10334 19742 10386 19794
rect 10386 19742 10388 19794
rect 10332 19740 10388 19742
rect 10220 19068 10276 19124
rect 9212 15932 9268 15988
rect 9100 15596 9156 15652
rect 8988 15260 9044 15316
rect 8876 14754 8932 14756
rect 8876 14702 8878 14754
rect 8878 14702 8930 14754
rect 8930 14702 8932 14754
rect 8876 14700 8932 14702
rect 9324 15484 9380 15540
rect 9436 15036 9492 15092
rect 9660 16940 9716 16996
rect 9996 18338 10052 18340
rect 9996 18286 9998 18338
rect 9998 18286 10050 18338
rect 10050 18286 10052 18338
rect 9996 18284 10052 18286
rect 9996 16828 10052 16884
rect 9996 16492 10052 16548
rect 10108 16098 10164 16100
rect 10108 16046 10110 16098
rect 10110 16046 10162 16098
rect 10162 16046 10164 16098
rect 10108 16044 10164 16046
rect 9996 15372 10052 15428
rect 9660 15202 9716 15204
rect 9660 15150 9662 15202
rect 9662 15150 9714 15202
rect 9714 15150 9716 15202
rect 9660 15148 9716 15150
rect 9772 15036 9828 15092
rect 9548 14364 9604 14420
rect 9436 13244 9492 13300
rect 8988 13074 9044 13076
rect 8988 13022 8990 13074
rect 8990 13022 9042 13074
rect 9042 13022 9044 13074
rect 8988 13020 9044 13022
rect 9100 12962 9156 12964
rect 9100 12910 9102 12962
rect 9102 12910 9154 12962
rect 9154 12910 9156 12962
rect 9100 12908 9156 12910
rect 8988 12460 9044 12516
rect 9548 11788 9604 11844
rect 9324 11564 9380 11620
rect 9884 14642 9940 14644
rect 9884 14590 9886 14642
rect 9886 14590 9938 14642
rect 9938 14590 9940 14642
rect 9884 14588 9940 14590
rect 10108 15484 10164 15540
rect 10780 19906 10836 19908
rect 10780 19854 10782 19906
rect 10782 19854 10834 19906
rect 10834 19854 10836 19906
rect 10780 19852 10836 19854
rect 10780 19346 10836 19348
rect 10780 19294 10782 19346
rect 10782 19294 10834 19346
rect 10834 19294 10836 19346
rect 10780 19292 10836 19294
rect 10668 19068 10724 19124
rect 10332 17164 10388 17220
rect 10556 18396 10612 18452
rect 11900 35756 11956 35812
rect 12460 40684 12516 40740
rect 12684 40460 12740 40516
rect 12460 39116 12516 39172
rect 12572 39228 12628 39284
rect 12348 36988 12404 37044
rect 12460 38892 12516 38948
rect 12684 38834 12740 38836
rect 12684 38782 12686 38834
rect 12686 38782 12738 38834
rect 12738 38782 12740 38834
rect 12684 38780 12740 38782
rect 12908 38780 12964 38836
rect 13356 44268 13412 44324
rect 13244 43538 13300 43540
rect 13244 43486 13246 43538
rect 13246 43486 13298 43538
rect 13298 43486 13300 43538
rect 13244 43484 13300 43486
rect 13244 43260 13300 43316
rect 13468 42028 13524 42084
rect 13468 41804 13524 41860
rect 13356 40684 13412 40740
rect 13804 44098 13860 44100
rect 13804 44046 13806 44098
rect 13806 44046 13858 44098
rect 13858 44046 13860 44098
rect 13804 44044 13860 44046
rect 13580 40460 13636 40516
rect 14028 45890 14084 45892
rect 14028 45838 14030 45890
rect 14030 45838 14082 45890
rect 14082 45838 14084 45890
rect 14028 45836 14084 45838
rect 14028 45276 14084 45332
rect 14476 48524 14532 48580
rect 13916 43372 13972 43428
rect 14252 47964 14308 48020
rect 14252 44940 14308 44996
rect 13692 41020 13748 41076
rect 13468 40348 13524 40404
rect 13580 40290 13636 40292
rect 13580 40238 13582 40290
rect 13582 40238 13634 40290
rect 13634 40238 13636 40290
rect 13580 40236 13636 40238
rect 13356 39788 13412 39844
rect 13244 39116 13300 39172
rect 12684 36988 12740 37044
rect 12572 36764 12628 36820
rect 12124 35756 12180 35812
rect 12348 36092 12404 36148
rect 12348 34972 12404 35028
rect 12012 34524 12068 34580
rect 12124 33516 12180 33572
rect 11900 32508 11956 32564
rect 12012 32844 12068 32900
rect 11900 31948 11956 32004
rect 12012 31724 12068 31780
rect 12236 32396 12292 32452
rect 12236 31612 12292 31668
rect 12348 31724 12404 31780
rect 12124 31388 12180 31444
rect 12236 30268 12292 30324
rect 11788 29596 11844 29652
rect 11676 29426 11732 29428
rect 11676 29374 11678 29426
rect 11678 29374 11730 29426
rect 11730 29374 11732 29426
rect 11676 29372 11732 29374
rect 12236 29314 12292 29316
rect 12236 29262 12238 29314
rect 12238 29262 12290 29314
rect 12290 29262 12292 29314
rect 12236 29260 12292 29262
rect 11676 27468 11732 27524
rect 12572 31948 12628 32004
rect 12572 31500 12628 31556
rect 12796 35644 12852 35700
rect 13244 37100 13300 37156
rect 13020 35196 13076 35252
rect 13020 34914 13076 34916
rect 13020 34862 13022 34914
rect 13022 34862 13074 34914
rect 13074 34862 13076 34914
rect 13020 34860 13076 34862
rect 12908 33068 12964 33124
rect 13468 39452 13524 39508
rect 13356 36652 13412 36708
rect 13580 38444 13636 38500
rect 13916 41692 13972 41748
rect 13916 40684 13972 40740
rect 13916 40124 13972 40180
rect 13692 38108 13748 38164
rect 13804 38332 13860 38388
rect 13804 37212 13860 37268
rect 13580 36540 13636 36596
rect 13244 35420 13300 35476
rect 13468 36316 13524 36372
rect 13468 34636 13524 34692
rect 13244 33516 13300 33572
rect 13132 31724 13188 31780
rect 13244 33068 13300 33124
rect 12684 31388 12740 31444
rect 13020 31276 13076 31332
rect 12684 30322 12740 30324
rect 12684 30270 12686 30322
rect 12686 30270 12738 30322
rect 12738 30270 12740 30322
rect 12684 30268 12740 30270
rect 12460 29596 12516 29652
rect 12908 29650 12964 29652
rect 12908 29598 12910 29650
rect 12910 29598 12962 29650
rect 12962 29598 12964 29650
rect 12908 29596 12964 29598
rect 13132 30882 13188 30884
rect 13132 30830 13134 30882
rect 13134 30830 13186 30882
rect 13186 30830 13188 30882
rect 13132 30828 13188 30830
rect 12348 29148 12404 29204
rect 12348 28588 12404 28644
rect 12572 28642 12628 28644
rect 12572 28590 12574 28642
rect 12574 28590 12626 28642
rect 12626 28590 12628 28642
rect 12572 28588 12628 28590
rect 12348 28140 12404 28196
rect 12796 28252 12852 28308
rect 12124 27746 12180 27748
rect 12124 27694 12126 27746
rect 12126 27694 12178 27746
rect 12178 27694 12180 27746
rect 12124 27692 12180 27694
rect 11900 27356 11956 27412
rect 12236 27244 12292 27300
rect 11900 27186 11956 27188
rect 11900 27134 11902 27186
rect 11902 27134 11954 27186
rect 11954 27134 11956 27186
rect 11900 27132 11956 27134
rect 12460 27186 12516 27188
rect 12460 27134 12462 27186
rect 12462 27134 12514 27186
rect 12514 27134 12516 27186
rect 12460 27132 12516 27134
rect 11676 26796 11732 26852
rect 12124 26796 12180 26852
rect 11676 25900 11732 25956
rect 11900 25788 11956 25844
rect 11788 25452 11844 25508
rect 11788 24780 11844 24836
rect 11676 24050 11732 24052
rect 11676 23998 11678 24050
rect 11678 23998 11730 24050
rect 11730 23998 11732 24050
rect 11676 23996 11732 23998
rect 11452 21196 11508 21252
rect 11788 22540 11844 22596
rect 11340 20914 11396 20916
rect 11340 20862 11342 20914
rect 11342 20862 11394 20914
rect 11394 20862 11396 20914
rect 11340 20860 11396 20862
rect 11116 20802 11172 20804
rect 11116 20750 11118 20802
rect 11118 20750 11170 20802
rect 11170 20750 11172 20802
rect 11116 20748 11172 20750
rect 11228 20690 11284 20692
rect 11228 20638 11230 20690
rect 11230 20638 11282 20690
rect 11282 20638 11284 20690
rect 11228 20636 11284 20638
rect 11116 19906 11172 19908
rect 11116 19854 11118 19906
rect 11118 19854 11170 19906
rect 11170 19854 11172 19906
rect 11116 19852 11172 19854
rect 11452 20412 11508 20468
rect 11004 19794 11060 19796
rect 11004 19742 11006 19794
rect 11006 19742 11058 19794
rect 11058 19742 11060 19794
rect 11004 19740 11060 19742
rect 11004 19404 11060 19460
rect 11004 18284 11060 18340
rect 10892 18060 10948 18116
rect 11228 18396 11284 18452
rect 11340 18508 11396 18564
rect 10668 17442 10724 17444
rect 10668 17390 10670 17442
rect 10670 17390 10722 17442
rect 10722 17390 10724 17442
rect 10668 17388 10724 17390
rect 10556 16940 10612 16996
rect 10668 16492 10724 16548
rect 10332 16322 10388 16324
rect 10332 16270 10334 16322
rect 10334 16270 10386 16322
rect 10386 16270 10388 16322
rect 10332 16268 10388 16270
rect 10556 16268 10612 16324
rect 10556 15820 10612 15876
rect 10220 15372 10276 15428
rect 10556 15426 10612 15428
rect 10556 15374 10558 15426
rect 10558 15374 10610 15426
rect 10610 15374 10612 15426
rect 10556 15372 10612 15374
rect 9660 11564 9716 11620
rect 9212 11452 9268 11508
rect 9100 11170 9156 11172
rect 9100 11118 9102 11170
rect 9102 11118 9154 11170
rect 9154 11118 9156 11170
rect 9100 11116 9156 11118
rect 9100 10892 9156 10948
rect 8876 10668 8932 10724
rect 9212 9996 9268 10052
rect 9772 10668 9828 10724
rect 10220 13132 10276 13188
rect 11228 17276 11284 17332
rect 11004 16380 11060 16436
rect 11116 16156 11172 16212
rect 10892 15202 10948 15204
rect 10892 15150 10894 15202
rect 10894 15150 10946 15202
rect 10946 15150 10948 15202
rect 10892 15148 10948 15150
rect 10332 11452 10388 11508
rect 10444 13692 10500 13748
rect 10332 10556 10388 10612
rect 10556 13132 10612 13188
rect 10556 10780 10612 10836
rect 9772 10386 9828 10388
rect 9772 10334 9774 10386
rect 9774 10334 9826 10386
rect 9826 10334 9828 10386
rect 9772 10332 9828 10334
rect 9996 10332 10052 10388
rect 9660 10220 9716 10276
rect 9548 10108 9604 10164
rect 9324 9884 9380 9940
rect 9884 9938 9940 9940
rect 9884 9886 9886 9938
rect 9886 9886 9938 9938
rect 9938 9886 9940 9938
rect 9884 9884 9940 9886
rect 9100 9212 9156 9268
rect 9660 9324 9716 9380
rect 9548 9212 9604 9268
rect 9324 8652 9380 8708
rect 9548 8258 9604 8260
rect 9548 8206 9550 8258
rect 9550 8206 9602 8258
rect 9602 8206 9604 8258
rect 9548 8204 9604 8206
rect 9100 7868 9156 7924
rect 8988 7196 9044 7252
rect 9324 7196 9380 7252
rect 8876 6860 8932 6916
rect 9100 6802 9156 6804
rect 9100 6750 9102 6802
rect 9102 6750 9154 6802
rect 9154 6750 9156 6802
rect 9100 6748 9156 6750
rect 8876 6690 8932 6692
rect 8876 6638 8878 6690
rect 8878 6638 8930 6690
rect 8930 6638 8932 6690
rect 8876 6636 8932 6638
rect 9212 6690 9268 6692
rect 9212 6638 9214 6690
rect 9214 6638 9266 6690
rect 9266 6638 9268 6690
rect 9212 6636 9268 6638
rect 9100 6524 9156 6580
rect 8540 5906 8596 5908
rect 8540 5854 8542 5906
rect 8542 5854 8594 5906
rect 8594 5854 8596 5906
rect 8540 5852 8596 5854
rect 8540 5068 8596 5124
rect 8764 5794 8820 5796
rect 8764 5742 8766 5794
rect 8766 5742 8818 5794
rect 8818 5742 8820 5794
rect 8764 5740 8820 5742
rect 9212 5404 9268 5460
rect 9884 9212 9940 9268
rect 9884 8092 9940 8148
rect 10108 9212 10164 9268
rect 9660 5740 9716 5796
rect 9436 5292 9492 5348
rect 8988 4956 9044 5012
rect 8876 4844 8932 4900
rect 8876 4508 8932 4564
rect 10108 7532 10164 7588
rect 9996 7474 10052 7476
rect 9996 7422 9998 7474
rect 9998 7422 10050 7474
rect 10050 7422 10052 7474
rect 9996 7420 10052 7422
rect 9884 6300 9940 6356
rect 10108 5180 10164 5236
rect 9772 5068 9828 5124
rect 9548 4284 9604 4340
rect 9772 3778 9828 3780
rect 9772 3726 9774 3778
rect 9774 3726 9826 3778
rect 9826 3726 9828 3778
rect 9772 3724 9828 3726
rect 9212 3388 9268 3444
rect 9324 3164 9380 3220
rect 8652 2716 8708 2772
rect 8876 2770 8932 2772
rect 8876 2718 8878 2770
rect 8878 2718 8930 2770
rect 8930 2718 8932 2770
rect 8876 2716 8932 2718
rect 8540 2268 8596 2324
rect 8540 2044 8596 2100
rect 8204 1986 8260 1988
rect 8204 1934 8206 1986
rect 8206 1934 8258 1986
rect 8258 1934 8260 1986
rect 8204 1932 8260 1934
rect 7980 1596 8036 1652
rect 8316 1596 8372 1652
rect 8092 978 8148 980
rect 8092 926 8094 978
rect 8094 926 8146 978
rect 8146 926 8148 978
rect 8092 924 8148 926
rect 7980 252 8036 308
rect 10108 3500 10164 3556
rect 10332 8258 10388 8260
rect 10332 8206 10334 8258
rect 10334 8206 10386 8258
rect 10386 8206 10388 8258
rect 10332 8204 10388 8206
rect 10332 6578 10388 6580
rect 10332 6526 10334 6578
rect 10334 6526 10386 6578
rect 10386 6526 10388 6578
rect 10332 6524 10388 6526
rect 9660 2604 9716 2660
rect 9660 2210 9716 2212
rect 9660 2158 9662 2210
rect 9662 2158 9714 2210
rect 9714 2158 9716 2210
rect 9660 2156 9716 2158
rect 9324 1932 9380 1988
rect 9660 1932 9716 1988
rect 9212 1596 9268 1652
rect 8764 1484 8820 1540
rect 8540 1148 8596 1204
rect 8764 1148 8820 1204
rect 9884 1260 9940 1316
rect 9996 924 10052 980
rect 10332 5740 10388 5796
rect 11004 13692 11060 13748
rect 12012 25506 12068 25508
rect 12012 25454 12014 25506
rect 12014 25454 12066 25506
rect 12066 25454 12068 25506
rect 12012 25452 12068 25454
rect 12684 26236 12740 26292
rect 13020 28252 13076 28308
rect 13020 28028 13076 28084
rect 13468 32396 13524 32452
rect 13244 28476 13300 28532
rect 13356 30828 13412 30884
rect 13916 35698 13972 35700
rect 13916 35646 13918 35698
rect 13918 35646 13970 35698
rect 13970 35646 13972 35698
rect 13916 35644 13972 35646
rect 13692 34690 13748 34692
rect 13692 34638 13694 34690
rect 13694 34638 13746 34690
rect 13746 34638 13748 34690
rect 13692 34636 13748 34638
rect 13916 34636 13972 34692
rect 14364 47292 14420 47348
rect 14812 49868 14868 49924
rect 14700 49810 14756 49812
rect 14700 49758 14702 49810
rect 14702 49758 14754 49810
rect 14754 49758 14756 49810
rect 14700 49756 14756 49758
rect 15148 51100 15204 51156
rect 15260 50594 15316 50596
rect 15260 50542 15262 50594
rect 15262 50542 15314 50594
rect 15314 50542 15316 50594
rect 15260 50540 15316 50542
rect 16828 52220 16884 52276
rect 16156 51436 16212 51492
rect 16940 51996 16996 52052
rect 16044 51324 16100 51380
rect 16268 50652 16324 50708
rect 15708 50540 15764 50596
rect 15036 49868 15092 49924
rect 15148 49698 15204 49700
rect 15148 49646 15150 49698
rect 15150 49646 15202 49698
rect 15202 49646 15204 49698
rect 15148 49644 15204 49646
rect 15148 49420 15204 49476
rect 14924 48914 14980 48916
rect 14924 48862 14926 48914
rect 14926 48862 14978 48914
rect 14978 48862 14980 48914
rect 14924 48860 14980 48862
rect 15260 48354 15316 48356
rect 15260 48302 15262 48354
rect 15262 48302 15314 48354
rect 15314 48302 15316 48354
rect 15260 48300 15316 48302
rect 14812 47852 14868 47908
rect 14700 47458 14756 47460
rect 14700 47406 14702 47458
rect 14702 47406 14754 47458
rect 14754 47406 14756 47458
rect 14700 47404 14756 47406
rect 14588 47068 14644 47124
rect 14588 46732 14644 46788
rect 14476 45164 14532 45220
rect 14140 40684 14196 40740
rect 14252 40236 14308 40292
rect 14700 45164 14756 45220
rect 14812 45057 14814 45108
rect 14814 45057 14866 45108
rect 14866 45057 14868 45108
rect 14812 45052 14868 45057
rect 15260 47292 15316 47348
rect 15036 46732 15092 46788
rect 15260 46620 15316 46676
rect 15036 44882 15092 44884
rect 15036 44830 15038 44882
rect 15038 44830 15090 44882
rect 15090 44830 15092 44882
rect 15036 44828 15092 44830
rect 14588 42588 14644 42644
rect 15148 44268 15204 44324
rect 15148 43820 15204 43876
rect 15148 43484 15204 43540
rect 14924 42588 14980 42644
rect 14924 42364 14980 42420
rect 14924 42028 14980 42084
rect 14812 41970 14868 41972
rect 14812 41918 14814 41970
rect 14814 41918 14866 41970
rect 14866 41918 14868 41970
rect 14812 41916 14868 41918
rect 14700 41804 14756 41860
rect 14812 41298 14868 41300
rect 14812 41246 14814 41298
rect 14814 41246 14866 41298
rect 14866 41246 14868 41298
rect 14812 41244 14868 41246
rect 14588 40460 14644 40516
rect 14476 40402 14532 40404
rect 14476 40350 14478 40402
rect 14478 40350 14530 40402
rect 14530 40350 14532 40402
rect 14476 40348 14532 40350
rect 15820 50316 15876 50372
rect 15708 49980 15764 50036
rect 15484 49810 15540 49812
rect 15484 49758 15486 49810
rect 15486 49758 15538 49810
rect 15538 49758 15540 49810
rect 15484 49756 15540 49758
rect 15708 49756 15764 49812
rect 15932 49810 15988 49812
rect 15932 49758 15934 49810
rect 15934 49758 15986 49810
rect 15986 49758 15988 49810
rect 15932 49756 15988 49758
rect 16044 48972 16100 49028
rect 15932 48748 15988 48804
rect 16044 48412 16100 48468
rect 15708 47852 15764 47908
rect 15820 48300 15876 48356
rect 15484 46674 15540 46676
rect 15484 46622 15486 46674
rect 15486 46622 15538 46674
rect 15538 46622 15540 46674
rect 15484 46620 15540 46622
rect 15372 43820 15428 43876
rect 15484 45724 15540 45780
rect 15372 43538 15428 43540
rect 15372 43486 15374 43538
rect 15374 43486 15426 43538
rect 15426 43486 15428 43538
rect 15372 43484 15428 43486
rect 15708 46620 15764 46676
rect 16940 51212 16996 51268
rect 16828 51100 16884 51156
rect 18396 54124 18452 54180
rect 19292 56140 19348 56196
rect 19068 55916 19124 55972
rect 19180 55580 19236 55636
rect 18732 54124 18788 54180
rect 18396 53788 18452 53844
rect 18620 53788 18676 53844
rect 17388 53340 17444 53396
rect 17724 52946 17780 52948
rect 17724 52894 17726 52946
rect 17726 52894 17778 52946
rect 17778 52894 17780 52946
rect 17724 52892 17780 52894
rect 17948 52892 18004 52948
rect 17948 52668 18004 52724
rect 17276 52108 17332 52164
rect 17164 51436 17220 51492
rect 17164 50764 17220 50820
rect 16492 50316 16548 50372
rect 16940 50428 16996 50484
rect 16940 49980 16996 50036
rect 17052 50204 17108 50260
rect 16828 49868 16884 49924
rect 16380 48300 16436 48356
rect 16492 49644 16548 49700
rect 15932 47852 15988 47908
rect 15932 47068 15988 47124
rect 17164 49196 17220 49252
rect 17612 51212 17668 51268
rect 17836 51266 17892 51268
rect 17836 51214 17838 51266
rect 17838 51214 17890 51266
rect 17890 51214 17892 51266
rect 17836 51212 17892 51214
rect 17500 50876 17556 50932
rect 17500 50540 17556 50596
rect 17724 50876 17780 50932
rect 17276 49026 17332 49028
rect 17276 48974 17278 49026
rect 17278 48974 17330 49026
rect 17330 48974 17332 49026
rect 17276 48972 17332 48974
rect 17052 48860 17108 48916
rect 16828 47964 16884 48020
rect 16268 47852 16324 47908
rect 16716 47852 16772 47908
rect 16156 47346 16212 47348
rect 16156 47294 16158 47346
rect 16158 47294 16210 47346
rect 16210 47294 16212 47346
rect 16156 47292 16212 47294
rect 16044 46508 16100 46564
rect 15932 46396 15988 46452
rect 16156 45388 16212 45444
rect 16044 45106 16100 45108
rect 16044 45054 16046 45106
rect 16046 45054 16098 45106
rect 16098 45054 16100 45106
rect 16044 45052 16100 45054
rect 15484 42812 15540 42868
rect 15820 42140 15876 42196
rect 15484 41916 15540 41972
rect 15260 41244 15316 41300
rect 15596 41244 15652 41300
rect 15708 40348 15764 40404
rect 14140 39676 14196 39732
rect 14252 39564 14308 39620
rect 14140 39452 14196 39508
rect 14252 38444 14308 38500
rect 14588 38780 14644 38836
rect 14476 38332 14532 38388
rect 14476 37548 14532 37604
rect 14476 37154 14532 37156
rect 14476 37102 14478 37154
rect 14478 37102 14530 37154
rect 14530 37102 14532 37154
rect 14476 37100 14532 37102
rect 14476 36764 14532 36820
rect 14364 35586 14420 35588
rect 14364 35534 14366 35586
rect 14366 35534 14418 35586
rect 14418 35534 14420 35586
rect 14364 35532 14420 35534
rect 14140 34636 14196 34692
rect 14140 34188 14196 34244
rect 15820 40124 15876 40180
rect 15260 39452 15316 39508
rect 14924 39116 14980 39172
rect 14812 38220 14868 38276
rect 14812 37212 14868 37268
rect 14924 38780 14980 38836
rect 16044 43596 16100 43652
rect 16604 47404 16660 47460
rect 16492 47068 16548 47124
rect 17276 48242 17332 48244
rect 17276 48190 17278 48242
rect 17278 48190 17330 48242
rect 17330 48190 17332 48242
rect 17276 48188 17332 48190
rect 16716 46620 16772 46676
rect 16716 46396 16772 46452
rect 16156 44044 16212 44100
rect 16044 43426 16100 43428
rect 16044 43374 16046 43426
rect 16046 43374 16098 43426
rect 16098 43374 16100 43426
rect 16044 43372 16100 43374
rect 16044 42642 16100 42644
rect 16044 42590 16046 42642
rect 16046 42590 16098 42642
rect 16098 42590 16100 42642
rect 16044 42588 16100 42590
rect 16044 42364 16100 42420
rect 16380 43820 16436 43876
rect 16940 47068 16996 47124
rect 16940 46844 16996 46900
rect 16940 46060 16996 46116
rect 17164 47570 17220 47572
rect 17164 47518 17166 47570
rect 17166 47518 17218 47570
rect 17218 47518 17220 47570
rect 17164 47516 17220 47518
rect 17276 47458 17332 47460
rect 17276 47406 17278 47458
rect 17278 47406 17330 47458
rect 17330 47406 17332 47458
rect 17276 47404 17332 47406
rect 17276 46844 17332 46900
rect 17052 45836 17108 45892
rect 16940 45778 16996 45780
rect 16940 45726 16942 45778
rect 16942 45726 16994 45778
rect 16994 45726 16996 45778
rect 16940 45724 16996 45726
rect 16940 45388 16996 45444
rect 17052 44716 17108 44772
rect 17276 44716 17332 44772
rect 16828 43820 16884 43876
rect 16492 43426 16548 43428
rect 16492 43374 16494 43426
rect 16494 43374 16546 43426
rect 16546 43374 16548 43426
rect 16492 43372 16548 43374
rect 16268 42252 16324 42308
rect 16044 41580 16100 41636
rect 16828 42252 16884 42308
rect 16492 41692 16548 41748
rect 16044 41298 16100 41300
rect 16044 41246 16046 41298
rect 16046 41246 16098 41298
rect 16098 41246 16100 41298
rect 16044 41244 16100 41246
rect 16156 40124 16212 40180
rect 16268 39676 16324 39732
rect 16044 39506 16100 39508
rect 16044 39454 16046 39506
rect 16046 39454 16098 39506
rect 16098 39454 16100 39506
rect 16044 39452 16100 39454
rect 15820 39116 15876 39172
rect 15260 38332 15316 38388
rect 15036 37772 15092 37828
rect 15036 37100 15092 37156
rect 14924 36594 14980 36596
rect 14924 36542 14926 36594
rect 14926 36542 14978 36594
rect 14978 36542 14980 36594
rect 14924 36540 14980 36542
rect 14700 36428 14756 36484
rect 14924 36204 14980 36260
rect 14588 35420 14644 35476
rect 14028 33740 14084 33796
rect 13916 33570 13972 33572
rect 13916 33518 13918 33570
rect 13918 33518 13970 33570
rect 13970 33518 13972 33570
rect 13916 33516 13972 33518
rect 13804 33404 13860 33460
rect 13916 32338 13972 32340
rect 13916 32286 13918 32338
rect 13918 32286 13970 32338
rect 13970 32286 13972 32338
rect 13916 32284 13972 32286
rect 13916 31724 13972 31780
rect 13804 30434 13860 30436
rect 13804 30382 13806 30434
rect 13806 30382 13858 30434
rect 13858 30382 13860 30434
rect 13804 30380 13860 30382
rect 13580 29932 13636 29988
rect 13468 29596 13524 29652
rect 13692 29820 13748 29876
rect 13692 29596 13748 29652
rect 13356 28028 13412 28084
rect 13132 27804 13188 27860
rect 13020 27746 13076 27748
rect 13020 27694 13022 27746
rect 13022 27694 13074 27746
rect 13074 27694 13076 27746
rect 13020 27692 13076 27694
rect 12908 27020 12964 27076
rect 13020 27356 13076 27412
rect 12908 26796 12964 26852
rect 12572 26124 12628 26180
rect 12460 25340 12516 25396
rect 11900 21420 11956 21476
rect 12236 24780 12292 24836
rect 12124 22370 12180 22372
rect 12124 22318 12126 22370
rect 12126 22318 12178 22370
rect 12178 22318 12180 22370
rect 12124 22316 12180 22318
rect 12124 21810 12180 21812
rect 12124 21758 12126 21810
rect 12126 21758 12178 21810
rect 12178 21758 12180 21810
rect 12124 21756 12180 21758
rect 12012 21644 12068 21700
rect 11788 20636 11844 20692
rect 11900 20412 11956 20468
rect 11788 19906 11844 19908
rect 11788 19854 11790 19906
rect 11790 19854 11842 19906
rect 11842 19854 11844 19906
rect 11788 19852 11844 19854
rect 11452 18060 11508 18116
rect 11452 17890 11508 17892
rect 11452 17838 11454 17890
rect 11454 17838 11506 17890
rect 11506 17838 11508 17890
rect 11452 17836 11508 17838
rect 11116 13468 11172 13524
rect 11228 13804 11284 13860
rect 11004 13244 11060 13300
rect 10892 12962 10948 12964
rect 10892 12910 10894 12962
rect 10894 12910 10946 12962
rect 10946 12910 10948 12962
rect 10892 12908 10948 12910
rect 10892 10834 10948 10836
rect 10892 10782 10894 10834
rect 10894 10782 10946 10834
rect 10946 10782 10948 10834
rect 10892 10780 10948 10782
rect 11340 13132 11396 13188
rect 11116 11788 11172 11844
rect 11564 11564 11620 11620
rect 11116 11394 11172 11396
rect 11116 11342 11118 11394
rect 11118 11342 11170 11394
rect 11170 11342 11172 11394
rect 11116 11340 11172 11342
rect 11004 10556 11060 10612
rect 11116 10780 11172 10836
rect 11004 10050 11060 10052
rect 11004 9998 11006 10050
rect 11006 9998 11058 10050
rect 11058 9998 11060 10050
rect 11004 9996 11060 9998
rect 10780 9884 10836 9940
rect 11004 9324 11060 9380
rect 11004 8764 11060 8820
rect 10892 8258 10948 8260
rect 10892 8206 10894 8258
rect 10894 8206 10946 8258
rect 10946 8206 10948 8258
rect 10892 8204 10948 8206
rect 10668 8092 10724 8148
rect 10556 7868 10612 7924
rect 10556 7420 10612 7476
rect 10668 6412 10724 6468
rect 10780 6860 10836 6916
rect 10780 6188 10836 6244
rect 10892 5906 10948 5908
rect 10892 5854 10894 5906
rect 10894 5854 10946 5906
rect 10946 5854 10948 5906
rect 10892 5852 10948 5854
rect 10892 5292 10948 5348
rect 10780 5068 10836 5124
rect 10556 4956 10612 5012
rect 10444 4562 10500 4564
rect 10444 4510 10446 4562
rect 10446 4510 10498 4562
rect 10498 4510 10500 4562
rect 10444 4508 10500 4510
rect 10668 4172 10724 4228
rect 11452 10722 11508 10724
rect 11452 10670 11454 10722
rect 11454 10670 11506 10722
rect 11506 10670 11508 10722
rect 11452 10668 11508 10670
rect 12012 19794 12068 19796
rect 12012 19742 12014 19794
rect 12014 19742 12066 19794
rect 12066 19742 12068 19794
rect 12012 19740 12068 19742
rect 12348 22540 12404 22596
rect 12348 22092 12404 22148
rect 12236 19852 12292 19908
rect 12012 19404 12068 19460
rect 12796 25788 12852 25844
rect 12572 23660 12628 23716
rect 12572 23436 12628 23492
rect 12684 24220 12740 24276
rect 13692 28476 13748 28532
rect 13244 26796 13300 26852
rect 13244 26290 13300 26292
rect 13244 26238 13246 26290
rect 13246 26238 13298 26290
rect 13298 26238 13300 26290
rect 13244 26236 13300 26238
rect 13580 27020 13636 27076
rect 13916 29036 13972 29092
rect 14476 32396 14532 32452
rect 14924 35644 14980 35700
rect 14700 35196 14756 35252
rect 14812 35026 14868 35028
rect 14812 34974 14814 35026
rect 14814 34974 14866 35026
rect 14866 34974 14868 35026
rect 14812 34972 14868 34974
rect 15148 36988 15204 37044
rect 15372 37996 15428 38052
rect 15260 36092 15316 36148
rect 14812 34130 14868 34132
rect 14812 34078 14814 34130
rect 14814 34078 14866 34130
rect 14866 34078 14868 34130
rect 14812 34076 14868 34078
rect 15820 37772 15876 37828
rect 15484 37042 15540 37044
rect 15484 36990 15486 37042
rect 15486 36990 15538 37042
rect 15538 36990 15540 37042
rect 15484 36988 15540 36990
rect 16044 37826 16100 37828
rect 16044 37774 16046 37826
rect 16046 37774 16098 37826
rect 16098 37774 16100 37826
rect 16044 37772 16100 37774
rect 15932 37266 15988 37268
rect 15932 37214 15934 37266
rect 15934 37214 15986 37266
rect 15986 37214 15988 37266
rect 15932 37212 15988 37214
rect 15596 36316 15652 36372
rect 15820 36204 15876 36260
rect 15820 35644 15876 35700
rect 15596 35532 15652 35588
rect 14700 32508 14756 32564
rect 14588 31276 14644 31332
rect 15372 34914 15428 34916
rect 15372 34862 15374 34914
rect 15374 34862 15426 34914
rect 15426 34862 15428 34914
rect 15372 34860 15428 34862
rect 15372 34636 15428 34692
rect 16268 38332 16324 38388
rect 16156 35084 16212 35140
rect 15708 34524 15764 34580
rect 15596 33852 15652 33908
rect 15372 33404 15428 33460
rect 14924 33346 14980 33348
rect 14924 33294 14926 33346
rect 14926 33294 14978 33346
rect 14978 33294 14980 33346
rect 14924 33292 14980 33294
rect 15148 33292 15204 33348
rect 15036 32562 15092 32564
rect 15036 32510 15038 32562
rect 15038 32510 15090 32562
rect 15090 32510 15092 32562
rect 15036 32508 15092 32510
rect 14924 31890 14980 31892
rect 14924 31838 14926 31890
rect 14926 31838 14978 31890
rect 14978 31838 14980 31890
rect 14924 31836 14980 31838
rect 14140 30940 14196 30996
rect 14588 30380 14644 30436
rect 14476 30210 14532 30212
rect 14476 30158 14478 30210
rect 14478 30158 14530 30210
rect 14530 30158 14532 30210
rect 14476 30156 14532 30158
rect 14364 29932 14420 29988
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 13916 27298 13972 27300
rect 13916 27246 13918 27298
rect 13918 27246 13970 27298
rect 13970 27246 13972 27298
rect 13916 27244 13972 27246
rect 13580 26572 13636 26628
rect 13580 26124 13636 26180
rect 13132 26066 13188 26068
rect 13132 26014 13134 26066
rect 13134 26014 13186 26066
rect 13186 26014 13188 26066
rect 13132 26012 13188 26014
rect 13468 25788 13524 25844
rect 13356 25564 13412 25620
rect 13244 25340 13300 25396
rect 13132 25228 13188 25284
rect 12796 22092 12852 22148
rect 12796 21196 12852 21252
rect 13132 21756 13188 21812
rect 13020 21196 13076 21252
rect 12684 20636 12740 20692
rect 12684 20188 12740 20244
rect 12796 19234 12852 19236
rect 12796 19182 12798 19234
rect 12798 19182 12850 19234
rect 12850 19182 12852 19234
rect 12796 19180 12852 19182
rect 12684 18508 12740 18564
rect 12348 18172 12404 18228
rect 11900 16156 11956 16212
rect 12012 17724 12068 17780
rect 12236 17666 12292 17668
rect 12236 17614 12238 17666
rect 12238 17614 12290 17666
rect 12290 17614 12292 17666
rect 12236 17612 12292 17614
rect 11788 12348 11844 12404
rect 12348 15372 12404 15428
rect 12124 15202 12180 15204
rect 12124 15150 12126 15202
rect 12126 15150 12178 15202
rect 12178 15150 12180 15202
rect 12124 15148 12180 15150
rect 12348 14924 12404 14980
rect 12124 14530 12180 14532
rect 12124 14478 12126 14530
rect 12126 14478 12178 14530
rect 12178 14478 12180 14530
rect 12124 14476 12180 14478
rect 12124 13970 12180 13972
rect 12124 13918 12126 13970
rect 12126 13918 12178 13970
rect 12178 13918 12180 13970
rect 12124 13916 12180 13918
rect 12908 18396 12964 18452
rect 13468 23772 13524 23828
rect 13692 23772 13748 23828
rect 13692 23324 13748 23380
rect 13804 23436 13860 23492
rect 13804 23212 13860 23268
rect 13804 22428 13860 22484
rect 13692 22316 13748 22372
rect 13804 21980 13860 22036
rect 14476 29820 14532 29876
rect 14588 30044 14644 30100
rect 14476 29148 14532 29204
rect 14252 27692 14308 27748
rect 14364 25900 14420 25956
rect 14364 25564 14420 25620
rect 14252 24332 14308 24388
rect 14140 23436 14196 23492
rect 13916 21756 13972 21812
rect 14700 29260 14756 29316
rect 14588 27858 14644 27860
rect 14588 27806 14590 27858
rect 14590 27806 14642 27858
rect 14642 27806 14644 27858
rect 14588 27804 14644 27806
rect 14700 25564 14756 25620
rect 14924 30492 14980 30548
rect 15260 32956 15316 33012
rect 15260 32732 15316 32788
rect 15036 28252 15092 28308
rect 15260 30156 15316 30212
rect 15260 28588 15316 28644
rect 15484 32732 15540 32788
rect 15484 32284 15540 32340
rect 15372 28476 15428 28532
rect 15484 31836 15540 31892
rect 15148 27746 15204 27748
rect 15148 27694 15150 27746
rect 15150 27694 15202 27746
rect 15202 27694 15204 27746
rect 15148 27692 15204 27694
rect 15036 26796 15092 26852
rect 14588 24332 14644 24388
rect 14700 23884 14756 23940
rect 14476 23436 14532 23492
rect 14476 23266 14532 23268
rect 14476 23214 14478 23266
rect 14478 23214 14530 23266
rect 14530 23214 14532 23266
rect 14476 23212 14532 23214
rect 14812 22370 14868 22372
rect 14812 22318 14814 22370
rect 14814 22318 14866 22370
rect 14866 22318 14868 22370
rect 14812 22316 14868 22318
rect 14252 21756 14308 21812
rect 13804 21644 13860 21700
rect 13580 20524 13636 20580
rect 14140 20188 14196 20244
rect 13580 19906 13636 19908
rect 13580 19854 13582 19906
rect 13582 19854 13634 19906
rect 13634 19854 13636 19906
rect 13580 19852 13636 19854
rect 13020 19180 13076 19236
rect 13356 19458 13412 19460
rect 13356 19406 13358 19458
rect 13358 19406 13410 19458
rect 13410 19406 13412 19458
rect 13356 19404 13412 19406
rect 13468 19346 13524 19348
rect 13468 19294 13470 19346
rect 13470 19294 13522 19346
rect 13522 19294 13524 19346
rect 13468 19292 13524 19294
rect 13244 18396 13300 18452
rect 13020 18172 13076 18228
rect 12796 17388 12852 17444
rect 13020 17724 13076 17780
rect 13244 17164 13300 17220
rect 13356 17612 13412 17668
rect 13580 17164 13636 17220
rect 13468 16716 13524 16772
rect 13916 16940 13972 16996
rect 13804 16770 13860 16772
rect 13804 16718 13806 16770
rect 13806 16718 13858 16770
rect 13858 16718 13860 16770
rect 13804 16716 13860 16718
rect 13804 16380 13860 16436
rect 13244 15708 13300 15764
rect 12908 15260 12964 15316
rect 12908 14924 12964 14980
rect 12796 14700 12852 14756
rect 12572 14476 12628 14532
rect 12908 14530 12964 14532
rect 12908 14478 12910 14530
rect 12910 14478 12962 14530
rect 12962 14478 12964 14530
rect 12908 14476 12964 14478
rect 12572 14252 12628 14308
rect 12460 13132 12516 13188
rect 12236 12348 12292 12404
rect 11676 11452 11732 11508
rect 12012 11788 12068 11844
rect 11564 10610 11620 10612
rect 11564 10558 11566 10610
rect 11566 10558 11618 10610
rect 11618 10558 11620 10610
rect 11564 10556 11620 10558
rect 11676 11228 11732 11284
rect 11564 10108 11620 10164
rect 11452 9996 11508 10052
rect 11340 9884 11396 9940
rect 11452 9714 11508 9716
rect 11452 9662 11454 9714
rect 11454 9662 11506 9714
rect 11506 9662 11508 9714
rect 11452 9660 11508 9662
rect 11900 11452 11956 11508
rect 11788 10386 11844 10388
rect 11788 10334 11790 10386
rect 11790 10334 11842 10386
rect 11842 10334 11844 10386
rect 11788 10332 11844 10334
rect 12236 11228 12292 11284
rect 12348 11900 12404 11956
rect 12124 11116 12180 11172
rect 12348 10892 12404 10948
rect 12460 10668 12516 10724
rect 12348 10556 12404 10612
rect 13020 13916 13076 13972
rect 13244 14812 13300 14868
rect 13244 14364 13300 14420
rect 13468 15596 13524 15652
rect 13580 15708 13636 15764
rect 13580 15484 13636 15540
rect 13580 15314 13636 15316
rect 13580 15262 13582 15314
rect 13582 15262 13634 15314
rect 13634 15262 13636 15314
rect 13580 15260 13636 15262
rect 13804 14588 13860 14644
rect 13580 14140 13636 14196
rect 13692 14476 13748 14532
rect 13580 13970 13636 13972
rect 13580 13918 13582 13970
rect 13582 13918 13634 13970
rect 13634 13918 13636 13970
rect 13580 13916 13636 13918
rect 13132 12962 13188 12964
rect 13132 12910 13134 12962
rect 13134 12910 13186 12962
rect 13186 12910 13188 12962
rect 13132 12908 13188 12910
rect 13020 12572 13076 12628
rect 13244 12572 13300 12628
rect 13356 13692 13412 13748
rect 13020 12124 13076 12180
rect 13132 11676 13188 11732
rect 12908 10444 12964 10500
rect 12572 10332 12628 10388
rect 12236 9938 12292 9940
rect 12236 9886 12238 9938
rect 12238 9886 12290 9938
rect 12290 9886 12292 9938
rect 12236 9884 12292 9886
rect 11900 9548 11956 9604
rect 12796 9938 12852 9940
rect 12796 9886 12798 9938
rect 12798 9886 12850 9938
rect 12850 9886 12852 9938
rect 12796 9884 12852 9886
rect 13132 9660 13188 9716
rect 13244 10556 13300 10612
rect 11788 9324 11844 9380
rect 12572 9548 12628 9604
rect 11116 7084 11172 7140
rect 11228 6748 11284 6804
rect 11564 8092 11620 8148
rect 11116 6412 11172 6468
rect 11116 6188 11172 6244
rect 11116 5068 11172 5124
rect 11788 7980 11844 8036
rect 11788 7756 11844 7812
rect 11900 8204 11956 8260
rect 11676 7420 11732 7476
rect 12012 7532 12068 7588
rect 11900 7474 11956 7476
rect 11900 7422 11902 7474
rect 11902 7422 11954 7474
rect 11954 7422 11956 7474
rect 11900 7420 11956 7422
rect 11788 6636 11844 6692
rect 11452 6524 11508 6580
rect 11900 6524 11956 6580
rect 11676 6412 11732 6468
rect 11788 5964 11844 6020
rect 11564 4396 11620 4452
rect 11228 3836 11284 3892
rect 11116 3778 11172 3780
rect 11116 3726 11118 3778
rect 11118 3726 11170 3778
rect 11170 3726 11172 3778
rect 11116 3724 11172 3726
rect 12236 7868 12292 7924
rect 12236 6300 12292 6356
rect 12348 7420 12404 7476
rect 12572 8370 12628 8372
rect 12572 8318 12574 8370
rect 12574 8318 12626 8370
rect 12626 8318 12628 8370
rect 12572 8316 12628 8318
rect 12460 7084 12516 7140
rect 12124 6188 12180 6244
rect 12012 6018 12068 6020
rect 12012 5966 12014 6018
rect 12014 5966 12066 6018
rect 12066 5966 12068 6018
rect 12012 5964 12068 5966
rect 12236 5964 12292 6020
rect 12236 5180 12292 5236
rect 11900 5122 11956 5124
rect 11900 5070 11902 5122
rect 11902 5070 11954 5122
rect 11954 5070 11956 5122
rect 11900 5068 11956 5070
rect 11900 4114 11956 4116
rect 11900 4062 11902 4114
rect 11902 4062 11954 4114
rect 11954 4062 11956 4114
rect 11900 4060 11956 4062
rect 13244 9324 13300 9380
rect 13356 11228 13412 11284
rect 13580 13692 13636 13748
rect 13356 10108 13412 10164
rect 13468 10332 13524 10388
rect 12796 8428 12852 8484
rect 13244 8428 13300 8484
rect 13132 7644 13188 7700
rect 13244 7084 13300 7140
rect 12908 6018 12964 6020
rect 12908 5966 12910 6018
rect 12910 5966 12962 6018
rect 12962 5966 12964 6018
rect 12908 5964 12964 5966
rect 12348 5068 12404 5124
rect 12460 5292 12516 5348
rect 11228 2770 11284 2772
rect 11228 2718 11230 2770
rect 11230 2718 11282 2770
rect 11282 2718 11284 2770
rect 11228 2716 11284 2718
rect 12236 2716 12292 2772
rect 12348 4844 12404 4900
rect 10444 1148 10500 1204
rect 10556 1932 10612 1988
rect 10332 140 10388 196
rect 11564 1820 11620 1876
rect 11452 1596 11508 1652
rect 11676 1596 11732 1652
rect 11004 1484 11060 1540
rect 10892 700 10948 756
rect 11228 1090 11284 1092
rect 11228 1038 11230 1090
rect 11230 1038 11282 1090
rect 11282 1038 11284 1090
rect 11228 1036 11284 1038
rect 12236 2156 12292 2212
rect 13580 9772 13636 9828
rect 13692 12908 13748 12964
rect 13580 8540 13636 8596
rect 14028 16098 14084 16100
rect 14028 16046 14030 16098
rect 14030 16046 14082 16098
rect 14082 16046 14084 16098
rect 14028 16044 14084 16046
rect 13916 13132 13972 13188
rect 14252 15708 14308 15764
rect 15372 26236 15428 26292
rect 15148 25004 15204 25060
rect 15260 26012 15316 26068
rect 15036 23212 15092 23268
rect 14812 20914 14868 20916
rect 14812 20862 14814 20914
rect 14814 20862 14866 20914
rect 14866 20862 14868 20914
rect 14812 20860 14868 20862
rect 14588 20748 14644 20804
rect 14476 20076 14532 20132
rect 14476 19234 14532 19236
rect 14476 19182 14478 19234
rect 14478 19182 14530 19234
rect 14530 19182 14532 19234
rect 14476 19180 14532 19182
rect 14812 20018 14868 20020
rect 14812 19966 14814 20018
rect 14814 19966 14866 20018
rect 14866 19966 14868 20018
rect 14812 19964 14868 19966
rect 15596 30156 15652 30212
rect 15596 28642 15652 28644
rect 15596 28590 15598 28642
rect 15598 28590 15650 28642
rect 15650 28590 15652 28642
rect 15596 28588 15652 28590
rect 16268 37660 16324 37716
rect 16044 33516 16100 33572
rect 16044 33180 16100 33236
rect 15820 32562 15876 32564
rect 15820 32510 15822 32562
rect 15822 32510 15874 32562
rect 15874 32510 15876 32562
rect 15820 32508 15876 32510
rect 16044 32396 16100 32452
rect 16268 32562 16324 32564
rect 16268 32510 16270 32562
rect 16270 32510 16322 32562
rect 16322 32510 16324 32562
rect 16268 32508 16324 32510
rect 15596 25116 15652 25172
rect 15708 24498 15764 24500
rect 15708 24446 15710 24498
rect 15710 24446 15762 24498
rect 15762 24446 15764 24498
rect 15708 24444 15764 24446
rect 16940 41468 16996 41524
rect 16828 40962 16884 40964
rect 16828 40910 16830 40962
rect 16830 40910 16882 40962
rect 16882 40910 16884 40962
rect 16828 40908 16884 40910
rect 16604 40236 16660 40292
rect 16604 39116 16660 39172
rect 16604 38892 16660 38948
rect 16940 39788 16996 39844
rect 16492 34524 16548 34580
rect 16828 39452 16884 39508
rect 16828 36988 16884 37044
rect 17276 43932 17332 43988
rect 17164 43596 17220 43652
rect 17388 43260 17444 43316
rect 17836 50652 17892 50708
rect 17836 50428 17892 50484
rect 18172 51660 18228 51716
rect 18284 51436 18340 51492
rect 18396 51996 18452 52052
rect 18508 52220 18564 52276
rect 20412 56476 20468 56532
rect 19964 55916 20020 55972
rect 20412 55970 20468 55972
rect 20412 55918 20414 55970
rect 20414 55918 20466 55970
rect 20466 55918 20468 55970
rect 20412 55916 20468 55918
rect 19516 55858 19572 55860
rect 19516 55806 19518 55858
rect 19518 55806 19570 55858
rect 19570 55806 19572 55858
rect 19516 55804 19572 55806
rect 20860 56028 20916 56084
rect 19516 55410 19572 55412
rect 19516 55358 19518 55410
rect 19518 55358 19570 55410
rect 19570 55358 19572 55410
rect 19516 55356 19572 55358
rect 20860 55410 20916 55412
rect 20860 55358 20862 55410
rect 20862 55358 20914 55410
rect 20914 55358 20916 55410
rect 20860 55356 20916 55358
rect 19404 55244 19460 55300
rect 18956 54348 19012 54404
rect 20076 54908 20132 54964
rect 19740 54796 19796 54852
rect 19292 54124 19348 54180
rect 19516 54012 19572 54068
rect 19964 54012 20020 54068
rect 20300 54796 20356 54852
rect 21644 56364 21700 56420
rect 22204 56700 22260 56756
rect 21980 55970 22036 55972
rect 21980 55918 21982 55970
rect 21982 55918 22034 55970
rect 22034 55918 22036 55970
rect 21980 55916 22036 55918
rect 20860 54124 20916 54180
rect 18844 53452 18900 53508
rect 19292 52722 19348 52724
rect 19292 52670 19294 52722
rect 19294 52670 19346 52722
rect 19346 52670 19348 52722
rect 19292 52668 19348 52670
rect 19516 52668 19572 52724
rect 18732 52556 18788 52612
rect 19404 52556 19460 52612
rect 18956 52274 19012 52276
rect 18956 52222 18958 52274
rect 18958 52222 19010 52274
rect 19010 52222 19012 52274
rect 18956 52220 19012 52222
rect 19180 52162 19236 52164
rect 19180 52110 19182 52162
rect 19182 52110 19234 52162
rect 19234 52110 19236 52162
rect 19180 52108 19236 52110
rect 19404 52108 19460 52164
rect 19516 51996 19572 52052
rect 18620 51772 18676 51828
rect 19516 51772 19572 51828
rect 18508 51436 18564 51492
rect 17948 49420 18004 49476
rect 18172 50540 18228 50596
rect 17948 49196 18004 49252
rect 17612 48188 17668 48244
rect 17724 48524 17780 48580
rect 17836 47404 17892 47460
rect 17500 45388 17556 45444
rect 17388 41298 17444 41300
rect 17388 41246 17390 41298
rect 17390 41246 17442 41298
rect 17442 41246 17444 41298
rect 17388 41244 17444 41246
rect 17164 40962 17220 40964
rect 17164 40910 17166 40962
rect 17166 40910 17218 40962
rect 17218 40910 17220 40962
rect 17164 40908 17220 40910
rect 18172 48636 18228 48692
rect 18620 51100 18676 51156
rect 18844 50876 18900 50932
rect 19292 50652 19348 50708
rect 18396 49196 18452 49252
rect 18396 47628 18452 47684
rect 18508 48412 18564 48468
rect 18284 47292 18340 47348
rect 17948 46060 18004 46116
rect 17836 44380 17892 44436
rect 18172 46396 18228 46452
rect 18732 49868 18788 49924
rect 19180 49810 19236 49812
rect 19180 49758 19182 49810
rect 19182 49758 19234 49810
rect 19234 49758 19236 49810
rect 19180 49756 19236 49758
rect 19068 49644 19124 49700
rect 18844 48972 18900 49028
rect 19180 49138 19236 49140
rect 19180 49086 19182 49138
rect 19182 49086 19234 49138
rect 19234 49086 19236 49138
rect 19180 49084 19236 49086
rect 18284 46284 18340 46340
rect 18508 46114 18564 46116
rect 18508 46062 18510 46114
rect 18510 46062 18562 46114
rect 18562 46062 18564 46114
rect 18508 46060 18564 46062
rect 18172 45724 18228 45780
rect 18284 44604 18340 44660
rect 18396 44492 18452 44548
rect 17612 41970 17668 41972
rect 17612 41918 17614 41970
rect 17614 41918 17666 41970
rect 17666 41918 17668 41970
rect 17612 41916 17668 41918
rect 17724 41244 17780 41300
rect 18060 42866 18116 42868
rect 18060 42814 18062 42866
rect 18062 42814 18114 42866
rect 18114 42814 18116 42866
rect 18060 42812 18116 42814
rect 17836 40908 17892 40964
rect 17164 37660 17220 37716
rect 16828 36092 16884 36148
rect 17388 37100 17444 37156
rect 18060 37548 18116 37604
rect 17612 37266 17668 37268
rect 17612 37214 17614 37266
rect 17614 37214 17666 37266
rect 17666 37214 17668 37266
rect 17612 37212 17668 37214
rect 17500 36764 17556 36820
rect 17836 36764 17892 36820
rect 16828 35084 16884 35140
rect 16604 32508 16660 32564
rect 16716 34636 16772 34692
rect 16492 32338 16548 32340
rect 16492 32286 16494 32338
rect 16494 32286 16546 32338
rect 16546 32286 16548 32338
rect 16492 32284 16548 32286
rect 16716 31836 16772 31892
rect 15932 30604 15988 30660
rect 16044 30210 16100 30212
rect 16044 30158 16046 30210
rect 16046 30158 16098 30210
rect 16098 30158 16100 30210
rect 16044 30156 16100 30158
rect 15932 28924 15988 28980
rect 15932 28588 15988 28644
rect 16492 29036 16548 29092
rect 16380 28812 16436 28868
rect 16268 28252 16324 28308
rect 16492 28364 16548 28420
rect 16044 27692 16100 27748
rect 16044 26460 16100 26516
rect 16380 27132 16436 27188
rect 16044 25676 16100 25732
rect 15932 23714 15988 23716
rect 15932 23662 15934 23714
rect 15934 23662 15986 23714
rect 15986 23662 15988 23714
rect 15932 23660 15988 23662
rect 15148 22988 15204 23044
rect 15484 23042 15540 23044
rect 15484 22990 15486 23042
rect 15486 22990 15538 23042
rect 15538 22990 15540 23042
rect 15484 22988 15540 22990
rect 15260 22930 15316 22932
rect 15260 22878 15262 22930
rect 15262 22878 15314 22930
rect 15314 22878 15316 22930
rect 15260 22876 15316 22878
rect 15372 22316 15428 22372
rect 15372 19852 15428 19908
rect 15484 19964 15540 20020
rect 14924 18508 14980 18564
rect 15036 18450 15092 18452
rect 15036 18398 15038 18450
rect 15038 18398 15090 18450
rect 15090 18398 15092 18450
rect 15036 18396 15092 18398
rect 14924 17948 14980 18004
rect 14812 17836 14868 17892
rect 14364 15484 14420 15540
rect 14476 17666 14532 17668
rect 14476 17614 14478 17666
rect 14478 17614 14530 17666
rect 14530 17614 14532 17666
rect 14476 17612 14532 17614
rect 14364 15148 14420 15204
rect 14700 16380 14756 16436
rect 14700 16156 14756 16212
rect 15260 17388 15316 17444
rect 14924 17164 14980 17220
rect 15484 17106 15540 17108
rect 15484 17054 15486 17106
rect 15486 17054 15538 17106
rect 15538 17054 15540 17106
rect 15484 17052 15540 17054
rect 15372 16882 15428 16884
rect 15372 16830 15374 16882
rect 15374 16830 15426 16882
rect 15426 16830 15428 16882
rect 15372 16828 15428 16830
rect 15708 22316 15764 22372
rect 15820 21756 15876 21812
rect 15820 21586 15876 21588
rect 15820 21534 15822 21586
rect 15822 21534 15874 21586
rect 15874 21534 15876 21586
rect 15820 21532 15876 21534
rect 15708 21196 15764 21252
rect 15820 20412 15876 20468
rect 16156 25564 16212 25620
rect 17276 35644 17332 35700
rect 17164 35196 17220 35252
rect 17052 34130 17108 34132
rect 17052 34078 17054 34130
rect 17054 34078 17106 34130
rect 17106 34078 17108 34130
rect 17052 34076 17108 34078
rect 17164 33740 17220 33796
rect 16940 32450 16996 32452
rect 16940 32398 16942 32450
rect 16942 32398 16994 32450
rect 16994 32398 16996 32450
rect 16940 32396 16996 32398
rect 16828 30828 16884 30884
rect 16940 31276 16996 31332
rect 16716 30380 16772 30436
rect 16828 29148 16884 29204
rect 16940 29820 16996 29876
rect 16716 29036 16772 29092
rect 16940 27916 16996 27972
rect 16604 27580 16660 27636
rect 16604 27132 16660 27188
rect 17388 35532 17444 35588
rect 17612 33740 17668 33796
rect 17388 32396 17444 32452
rect 17500 32060 17556 32116
rect 17836 31724 17892 31780
rect 17948 36092 18004 36148
rect 18060 35532 18116 35588
rect 18060 34972 18116 35028
rect 18060 34188 18116 34244
rect 17836 31276 17892 31332
rect 17724 30940 17780 30996
rect 17164 30156 17220 30212
rect 17276 30380 17332 30436
rect 17164 28476 17220 28532
rect 17164 27132 17220 27188
rect 17388 29820 17444 29876
rect 17388 28140 17444 28196
rect 17500 27970 17556 27972
rect 17500 27918 17502 27970
rect 17502 27918 17554 27970
rect 17554 27918 17556 27970
rect 17500 27916 17556 27918
rect 17612 27020 17668 27076
rect 17388 26796 17444 26852
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 16604 26012 16660 26068
rect 16492 25452 16548 25508
rect 16828 25900 16884 25956
rect 16380 25004 16436 25060
rect 16492 25116 16548 25172
rect 16268 24444 16324 24500
rect 16828 24668 16884 24724
rect 16268 22204 16324 22260
rect 16156 21756 16212 21812
rect 16268 21644 16324 21700
rect 17052 25676 17108 25732
rect 17052 24444 17108 24500
rect 17164 25452 17220 25508
rect 16492 23100 16548 23156
rect 16156 20412 16212 20468
rect 16044 19458 16100 19460
rect 16044 19406 16046 19458
rect 16046 19406 16098 19458
rect 16098 19406 16100 19458
rect 16044 19404 16100 19406
rect 16268 19516 16324 19572
rect 16380 21084 16436 21140
rect 16268 18732 16324 18788
rect 16268 18508 16324 18564
rect 15932 17836 15988 17892
rect 16268 18172 16324 18228
rect 16044 17666 16100 17668
rect 16044 17614 16046 17666
rect 16046 17614 16098 17666
rect 16098 17614 16100 17666
rect 16044 17612 16100 17614
rect 16156 17500 16212 17556
rect 15596 16716 15652 16772
rect 15260 16604 15316 16660
rect 16044 16210 16100 16212
rect 16044 16158 16046 16210
rect 16046 16158 16098 16210
rect 16098 16158 16100 16210
rect 16044 16156 16100 16158
rect 15596 15820 15652 15876
rect 14364 14364 14420 14420
rect 14476 13132 14532 13188
rect 14140 12236 14196 12292
rect 13916 11788 13972 11844
rect 13916 11170 13972 11172
rect 13916 11118 13918 11170
rect 13918 11118 13970 11170
rect 13970 11118 13972 11170
rect 13916 11116 13972 11118
rect 13804 10780 13860 10836
rect 13804 9772 13860 9828
rect 14028 10108 14084 10164
rect 14924 15148 14980 15204
rect 14924 14924 14980 14980
rect 15036 14140 15092 14196
rect 14700 12124 14756 12180
rect 14364 11228 14420 11284
rect 14588 11228 14644 11284
rect 14364 10892 14420 10948
rect 16156 15148 16212 15204
rect 15708 14364 15764 14420
rect 15820 14700 15876 14756
rect 15596 13916 15652 13972
rect 15036 11564 15092 11620
rect 15148 13468 15204 13524
rect 15036 11340 15092 11396
rect 15260 13132 15316 13188
rect 15372 13244 15428 13300
rect 15484 13186 15540 13188
rect 15484 13134 15486 13186
rect 15486 13134 15538 13186
rect 15538 13134 15540 13186
rect 15484 13132 15540 13134
rect 15260 11676 15316 11732
rect 15596 11788 15652 11844
rect 15372 11564 15428 11620
rect 15708 11676 15764 11732
rect 15596 11564 15652 11620
rect 14924 10780 14980 10836
rect 15484 10780 15540 10836
rect 14700 10668 14756 10724
rect 14588 10610 14644 10612
rect 14588 10558 14590 10610
rect 14590 10558 14642 10610
rect 14642 10558 14644 10610
rect 14588 10556 14644 10558
rect 14924 10556 14980 10612
rect 14476 10444 14532 10500
rect 14140 8988 14196 9044
rect 13580 7420 13636 7476
rect 13580 6860 13636 6916
rect 13804 6860 13860 6916
rect 12908 5180 12964 5236
rect 12684 5122 12740 5124
rect 12684 5070 12686 5122
rect 12686 5070 12738 5122
rect 12738 5070 12740 5122
rect 12684 5068 12740 5070
rect 13132 5122 13188 5124
rect 13132 5070 13134 5122
rect 13134 5070 13186 5122
rect 13186 5070 13188 5122
rect 13132 5068 13188 5070
rect 14028 7250 14084 7252
rect 14028 7198 14030 7250
rect 14030 7198 14082 7250
rect 14082 7198 14084 7250
rect 14028 7196 14084 7198
rect 14252 8428 14308 8484
rect 14252 7362 14308 7364
rect 14252 7310 14254 7362
rect 14254 7310 14306 7362
rect 14306 7310 14308 7362
rect 14252 7308 14308 7310
rect 15708 10610 15764 10612
rect 15708 10558 15710 10610
rect 15710 10558 15762 10610
rect 15762 10558 15764 10610
rect 15708 10556 15764 10558
rect 15484 10444 15540 10500
rect 14588 9772 14644 9828
rect 14700 9042 14756 9044
rect 14700 8990 14702 9042
rect 14702 8990 14754 9042
rect 14754 8990 14756 9042
rect 14700 8988 14756 8990
rect 15372 10332 15428 10388
rect 15260 9996 15316 10052
rect 14924 8316 14980 8372
rect 14700 8258 14756 8260
rect 14700 8206 14702 8258
rect 14702 8206 14754 8258
rect 14754 8206 14756 8258
rect 14700 8204 14756 8206
rect 14588 8092 14644 8148
rect 14924 7756 14980 7812
rect 14476 7308 14532 7364
rect 14812 7532 14868 7588
rect 14364 6972 14420 7028
rect 14476 7084 14532 7140
rect 14588 6802 14644 6804
rect 14588 6750 14590 6802
rect 14590 6750 14642 6802
rect 14642 6750 14644 6802
rect 14588 6748 14644 6750
rect 15596 10050 15652 10052
rect 15596 9998 15598 10050
rect 15598 9998 15650 10050
rect 15650 9998 15652 10050
rect 15596 9996 15652 9998
rect 16492 20412 16548 20468
rect 16492 19852 16548 19908
rect 17052 23436 17108 23492
rect 16828 22652 16884 22708
rect 17052 22876 17108 22932
rect 16940 22316 16996 22372
rect 16828 20748 16884 20804
rect 16716 19852 16772 19908
rect 16604 19516 16660 19572
rect 16492 16770 16548 16772
rect 16492 16718 16494 16770
rect 16494 16718 16546 16770
rect 16546 16718 16548 16770
rect 16492 16716 16548 16718
rect 16492 16156 16548 16212
rect 16492 15260 16548 15316
rect 16828 19404 16884 19460
rect 17612 26572 17668 26628
rect 17948 31164 18004 31220
rect 17836 29426 17892 29428
rect 17836 29374 17838 29426
rect 17838 29374 17890 29426
rect 17890 29374 17892 29426
rect 17836 29372 17892 29374
rect 17948 27916 18004 27972
rect 17948 27634 18004 27636
rect 17948 27582 17950 27634
rect 17950 27582 18002 27634
rect 18002 27582 18004 27634
rect 17948 27580 18004 27582
rect 18060 27020 18116 27076
rect 18284 42588 18340 42644
rect 19180 48018 19236 48020
rect 19180 47966 19182 48018
rect 19182 47966 19234 48018
rect 19234 47966 19236 48018
rect 19180 47964 19236 47966
rect 19068 47852 19124 47908
rect 19068 47068 19124 47124
rect 18956 46956 19012 47012
rect 19740 52556 19796 52612
rect 19740 51660 19796 51716
rect 19964 53228 20020 53284
rect 20076 53170 20132 53172
rect 20076 53118 20078 53170
rect 20078 53118 20130 53170
rect 20130 53118 20132 53170
rect 20076 53116 20132 53118
rect 20188 52892 20244 52948
rect 19964 51772 20020 51828
rect 19628 51212 19684 51268
rect 19964 50988 20020 51044
rect 19516 50540 19572 50596
rect 20076 50316 20132 50372
rect 19964 50092 20020 50148
rect 20524 53900 20580 53956
rect 21196 54460 21252 54516
rect 21756 55580 21812 55636
rect 22652 55970 22708 55972
rect 22652 55918 22654 55970
rect 22654 55918 22706 55970
rect 22706 55918 22708 55970
rect 22652 55916 22708 55918
rect 23100 55916 23156 55972
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 24444 56476 24500 56532
rect 22540 55804 22596 55860
rect 24892 56812 24948 56868
rect 24556 56252 24612 56308
rect 22988 55858 23044 55860
rect 22988 55806 22990 55858
rect 22990 55806 23042 55858
rect 23042 55806 23044 55858
rect 22988 55804 23044 55806
rect 25340 56924 25396 56980
rect 25116 56364 25172 56420
rect 25788 55970 25844 55972
rect 25788 55918 25790 55970
rect 25790 55918 25842 55970
rect 25842 55918 25844 55970
rect 25788 55916 25844 55918
rect 21756 55298 21812 55300
rect 21756 55246 21758 55298
rect 21758 55246 21810 55298
rect 21810 55246 21812 55298
rect 21756 55244 21812 55246
rect 21756 54684 21812 54740
rect 23212 55468 23268 55524
rect 22540 55298 22596 55300
rect 22540 55246 22542 55298
rect 22542 55246 22594 55298
rect 22594 55246 22596 55298
rect 22540 55244 22596 55246
rect 22876 55020 22932 55076
rect 21196 53618 21252 53620
rect 21196 53566 21198 53618
rect 21198 53566 21250 53618
rect 21250 53566 21252 53618
rect 21196 53564 21252 53566
rect 21532 53564 21588 53620
rect 21644 52946 21700 52948
rect 21644 52894 21646 52946
rect 21646 52894 21698 52946
rect 21698 52894 21700 52946
rect 21644 52892 21700 52894
rect 20636 52332 20692 52388
rect 20860 52274 20916 52276
rect 20860 52222 20862 52274
rect 20862 52222 20914 52274
rect 20914 52222 20916 52274
rect 20860 52220 20916 52222
rect 20524 51884 20580 51940
rect 20636 51996 20692 52052
rect 20636 51378 20692 51380
rect 20636 51326 20638 51378
rect 20638 51326 20690 51378
rect 20690 51326 20692 51378
rect 20636 51324 20692 51326
rect 21532 52162 21588 52164
rect 21532 52110 21534 52162
rect 21534 52110 21586 52162
rect 21586 52110 21588 52162
rect 21532 52108 21588 52110
rect 21420 51996 21476 52052
rect 20748 51212 20804 51268
rect 20188 50204 20244 50260
rect 20076 49756 20132 49812
rect 19740 49644 19796 49700
rect 19964 49698 20020 49700
rect 19964 49646 19966 49698
rect 19966 49646 20018 49698
rect 20018 49646 20020 49698
rect 19964 49644 20020 49646
rect 19628 49196 19684 49252
rect 19404 47404 19460 47460
rect 19404 47068 19460 47124
rect 18620 44380 18676 44436
rect 18956 46060 19012 46116
rect 19404 46172 19460 46228
rect 19068 45612 19124 45668
rect 19292 44492 19348 44548
rect 19068 44044 19124 44100
rect 18732 41804 18788 41860
rect 19068 41970 19124 41972
rect 19068 41918 19070 41970
rect 19070 41918 19122 41970
rect 19122 41918 19124 41970
rect 19068 41916 19124 41918
rect 18508 41244 18564 41300
rect 18620 40908 18676 40964
rect 18284 37660 18340 37716
rect 18508 38556 18564 38612
rect 18396 37548 18452 37604
rect 18284 36988 18340 37044
rect 18284 31778 18340 31780
rect 18284 31726 18286 31778
rect 18286 31726 18338 31778
rect 18338 31726 18340 31778
rect 18284 31724 18340 31726
rect 18508 37100 18564 37156
rect 18508 36092 18564 36148
rect 18844 41020 18900 41076
rect 19292 41244 19348 41300
rect 18956 40796 19012 40852
rect 18844 40684 18900 40740
rect 19180 40348 19236 40404
rect 18844 40290 18900 40292
rect 18844 40238 18846 40290
rect 18846 40238 18898 40290
rect 18898 40238 18900 40290
rect 18844 40236 18900 40238
rect 19068 40012 19124 40068
rect 18844 39730 18900 39732
rect 18844 39678 18846 39730
rect 18846 39678 18898 39730
rect 18898 39678 18900 39730
rect 18844 39676 18900 39678
rect 18844 38722 18900 38724
rect 18844 38670 18846 38722
rect 18846 38670 18898 38722
rect 18898 38670 18900 38722
rect 18844 38668 18900 38670
rect 18844 36876 18900 36932
rect 18620 35308 18676 35364
rect 18508 35196 18564 35252
rect 19292 38556 19348 38612
rect 19180 37324 19236 37380
rect 20188 49196 20244 49252
rect 19740 48748 19796 48804
rect 19964 48412 20020 48468
rect 19852 48018 19908 48020
rect 19852 47966 19854 48018
rect 19854 47966 19906 48018
rect 19906 47966 19908 48018
rect 19852 47964 19908 47966
rect 19740 47180 19796 47236
rect 19852 47516 19908 47572
rect 19964 47404 20020 47460
rect 20076 47180 20132 47236
rect 20076 46844 20132 46900
rect 19964 46060 20020 46116
rect 20076 46396 20132 46452
rect 19628 44044 19684 44100
rect 19740 45836 19796 45892
rect 19516 41468 19572 41524
rect 19628 43484 19684 43540
rect 19964 44716 20020 44772
rect 19852 43538 19908 43540
rect 19852 43486 19854 43538
rect 19854 43486 19906 43538
rect 19906 43486 19908 43538
rect 19852 43484 19908 43486
rect 20300 48802 20356 48804
rect 20300 48750 20302 48802
rect 20302 48750 20354 48802
rect 20354 48750 20356 48802
rect 20300 48748 20356 48750
rect 20300 47570 20356 47572
rect 20300 47518 20302 47570
rect 20302 47518 20354 47570
rect 20354 47518 20356 47570
rect 20300 47516 20356 47518
rect 20300 46732 20356 46788
rect 20076 44210 20132 44212
rect 20076 44158 20078 44210
rect 20078 44158 20130 44210
rect 20130 44158 20132 44210
rect 20076 44156 20132 44158
rect 19964 43372 20020 43428
rect 19740 43036 19796 43092
rect 20188 43036 20244 43092
rect 19628 42588 19684 42644
rect 19516 41020 19572 41076
rect 19516 40348 19572 40404
rect 19740 42252 19796 42308
rect 19740 40236 19796 40292
rect 20188 41916 20244 41972
rect 19964 40402 20020 40404
rect 19964 40350 19966 40402
rect 19966 40350 20018 40402
rect 20018 40350 20020 40402
rect 19964 40348 20020 40350
rect 19852 40012 19908 40068
rect 20076 40012 20132 40068
rect 20524 50204 20580 50260
rect 20748 48914 20804 48916
rect 20748 48862 20750 48914
rect 20750 48862 20802 48914
rect 20802 48862 20804 48914
rect 20748 48860 20804 48862
rect 20636 48636 20692 48692
rect 21084 50988 21140 51044
rect 21084 50540 21140 50596
rect 21084 49922 21140 49924
rect 21084 49870 21086 49922
rect 21086 49870 21138 49922
rect 21138 49870 21140 49922
rect 21084 49868 21140 49870
rect 20972 48860 21028 48916
rect 20524 47292 20580 47348
rect 20748 47180 20804 47236
rect 20748 46898 20804 46900
rect 20748 46846 20750 46898
rect 20750 46846 20802 46898
rect 20802 46846 20804 46898
rect 20748 46844 20804 46846
rect 20860 46674 20916 46676
rect 20860 46622 20862 46674
rect 20862 46622 20914 46674
rect 20914 46622 20916 46674
rect 20860 46620 20916 46622
rect 20748 46562 20804 46564
rect 20748 46510 20750 46562
rect 20750 46510 20802 46562
rect 20802 46510 20804 46562
rect 20748 46508 20804 46510
rect 20524 45724 20580 45780
rect 20524 44268 20580 44324
rect 20636 44828 20692 44884
rect 20412 43372 20468 43428
rect 20636 43708 20692 43764
rect 20524 42588 20580 42644
rect 20748 43484 20804 43540
rect 21084 48748 21140 48804
rect 21532 51772 21588 51828
rect 21532 50988 21588 51044
rect 21532 49756 21588 49812
rect 21420 49420 21476 49476
rect 22428 54402 22484 54404
rect 22428 54350 22430 54402
rect 22430 54350 22482 54402
rect 22482 54350 22484 54402
rect 22428 54348 22484 54350
rect 22092 54012 22148 54068
rect 21980 53788 22036 53844
rect 22092 53730 22148 53732
rect 22092 53678 22094 53730
rect 22094 53678 22146 53730
rect 22146 53678 22148 53730
rect 22092 53676 22148 53678
rect 22092 53452 22148 53508
rect 21980 52834 22036 52836
rect 21980 52782 21982 52834
rect 21982 52782 22034 52834
rect 22034 52782 22036 52834
rect 21980 52780 22036 52782
rect 21756 51548 21812 51604
rect 21868 51490 21924 51492
rect 21868 51438 21870 51490
rect 21870 51438 21922 51490
rect 21922 51438 21924 51490
rect 21868 51436 21924 51438
rect 21756 51324 21812 51380
rect 21756 50876 21812 50932
rect 21756 50706 21812 50708
rect 21756 50654 21758 50706
rect 21758 50654 21810 50706
rect 21810 50654 21812 50706
rect 21756 50652 21812 50654
rect 21644 49308 21700 49364
rect 21868 48972 21924 49028
rect 22428 53452 22484 53508
rect 23100 54290 23156 54292
rect 23100 54238 23102 54290
rect 23102 54238 23154 54290
rect 23154 54238 23156 54290
rect 23100 54236 23156 54238
rect 22764 53452 22820 53508
rect 23100 53900 23156 53956
rect 22652 52892 22708 52948
rect 22428 52780 22484 52836
rect 22316 52722 22372 52724
rect 22316 52670 22318 52722
rect 22318 52670 22370 52722
rect 22370 52670 22372 52722
rect 22316 52668 22372 52670
rect 22092 52332 22148 52388
rect 22764 52386 22820 52388
rect 22764 52334 22766 52386
rect 22766 52334 22818 52386
rect 22818 52334 22820 52386
rect 22764 52332 22820 52334
rect 22316 51436 22372 51492
rect 22316 50764 22372 50820
rect 22764 51100 22820 51156
rect 22764 50876 22820 50932
rect 21980 48860 22036 48916
rect 21980 48412 22036 48468
rect 21420 47068 21476 47124
rect 21868 47404 21924 47460
rect 21644 47292 21700 47348
rect 22092 48130 22148 48132
rect 22092 48078 22094 48130
rect 22094 48078 22146 48130
rect 22146 48078 22148 48130
rect 22092 48076 22148 48078
rect 22764 49084 22820 49140
rect 22652 48748 22708 48804
rect 22316 47180 22372 47236
rect 20636 42364 20692 42420
rect 20860 42700 20916 42756
rect 20860 41916 20916 41972
rect 20972 41580 21028 41636
rect 20972 40012 21028 40068
rect 21084 40236 21140 40292
rect 19628 37884 19684 37940
rect 19404 37100 19460 37156
rect 19740 36482 19796 36484
rect 19740 36430 19742 36482
rect 19742 36430 19794 36482
rect 19794 36430 19796 36482
rect 19740 36428 19796 36430
rect 19404 36092 19460 36148
rect 18620 35084 18676 35140
rect 19180 35084 19236 35140
rect 18620 34130 18676 34132
rect 18620 34078 18622 34130
rect 18622 34078 18674 34130
rect 18674 34078 18676 34130
rect 18620 34076 18676 34078
rect 19068 34690 19124 34692
rect 19068 34638 19070 34690
rect 19070 34638 19122 34690
rect 19122 34638 19124 34690
rect 19068 34636 19124 34638
rect 19068 34412 19124 34468
rect 19964 37996 20020 38052
rect 19404 35084 19460 35140
rect 19740 35308 19796 35364
rect 20412 34972 20468 35028
rect 19628 34636 19684 34692
rect 19852 34802 19908 34804
rect 19852 34750 19854 34802
rect 19854 34750 19906 34802
rect 19906 34750 19908 34802
rect 19852 34748 19908 34750
rect 19516 34412 19572 34468
rect 18844 34076 18900 34132
rect 18508 34018 18564 34020
rect 18508 33966 18510 34018
rect 18510 33966 18562 34018
rect 18562 33966 18564 34018
rect 18508 33964 18564 33966
rect 19628 34130 19684 34132
rect 19628 34078 19630 34130
rect 19630 34078 19682 34130
rect 19682 34078 19684 34130
rect 19628 34076 19684 34078
rect 19516 33458 19572 33460
rect 19516 33406 19518 33458
rect 19518 33406 19570 33458
rect 19570 33406 19572 33458
rect 19516 33404 19572 33406
rect 18620 32732 18676 32788
rect 18508 32562 18564 32564
rect 18508 32510 18510 32562
rect 18510 32510 18562 32562
rect 18562 32510 18564 32562
rect 18508 32508 18564 32510
rect 18396 30940 18452 30996
rect 18508 30380 18564 30436
rect 18172 28924 18228 28980
rect 18844 32620 18900 32676
rect 18620 28924 18676 28980
rect 18732 31612 18788 31668
rect 18508 28866 18564 28868
rect 18508 28814 18510 28866
rect 18510 28814 18562 28866
rect 18562 28814 18564 28866
rect 18508 28812 18564 28814
rect 19516 32508 19572 32564
rect 18844 31164 18900 31220
rect 19180 31500 19236 31556
rect 18844 30994 18900 30996
rect 18844 30942 18846 30994
rect 18846 30942 18898 30994
rect 18898 30942 18900 30994
rect 18844 30940 18900 30942
rect 18508 28588 18564 28644
rect 18844 30492 18900 30548
rect 18508 27804 18564 27860
rect 18396 27356 18452 27412
rect 18284 27020 18340 27076
rect 18396 26908 18452 26964
rect 17612 26178 17668 26180
rect 17612 26126 17614 26178
rect 17614 26126 17666 26178
rect 17666 26126 17668 26178
rect 17612 26124 17668 26126
rect 17500 26066 17556 26068
rect 17500 26014 17502 26066
rect 17502 26014 17554 26066
rect 17554 26014 17556 26066
rect 17500 26012 17556 26014
rect 17724 25618 17780 25620
rect 17724 25566 17726 25618
rect 17726 25566 17778 25618
rect 17778 25566 17780 25618
rect 17724 25564 17780 25566
rect 17500 25452 17556 25508
rect 17276 23660 17332 23716
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 17388 22652 17444 22708
rect 17164 21756 17220 21812
rect 17836 23324 17892 23380
rect 18172 23660 18228 23716
rect 18060 23436 18116 23492
rect 18060 23154 18116 23156
rect 18060 23102 18062 23154
rect 18062 23102 18114 23154
rect 18114 23102 18116 23154
rect 18060 23100 18116 23102
rect 17612 22652 17668 22708
rect 17500 21756 17556 21812
rect 17388 21308 17444 21364
rect 17276 20412 17332 20468
rect 17164 20076 17220 20132
rect 17164 19404 17220 19460
rect 17164 18450 17220 18452
rect 17164 18398 17166 18450
rect 17166 18398 17218 18450
rect 17218 18398 17220 18450
rect 17164 18396 17220 18398
rect 16940 17778 16996 17780
rect 16940 17726 16942 17778
rect 16942 17726 16994 17778
rect 16994 17726 16996 17778
rect 16940 17724 16996 17726
rect 16828 17164 16884 17220
rect 16716 16828 16772 16884
rect 17164 17052 17220 17108
rect 16940 16044 16996 16100
rect 17052 16716 17108 16772
rect 16604 15148 16660 15204
rect 16716 15932 16772 15988
rect 16380 14252 16436 14308
rect 15932 12124 15988 12180
rect 17052 15484 17108 15540
rect 17164 15314 17220 15316
rect 17164 15262 17166 15314
rect 17166 15262 17218 15314
rect 17218 15262 17220 15314
rect 17164 15260 17220 15262
rect 16828 13916 16884 13972
rect 17612 21362 17668 21364
rect 17612 21310 17614 21362
rect 17614 21310 17666 21362
rect 17666 21310 17668 21362
rect 17612 21308 17668 21310
rect 18060 22652 18116 22708
rect 17948 22258 18004 22260
rect 17948 22206 17950 22258
rect 17950 22206 18002 22258
rect 18002 22206 18004 22258
rect 17948 22204 18004 22206
rect 18060 21420 18116 21476
rect 17948 21308 18004 21364
rect 17612 20076 17668 20132
rect 17836 20802 17892 20804
rect 17836 20750 17838 20802
rect 17838 20750 17890 20802
rect 17890 20750 17892 20802
rect 17836 20748 17892 20750
rect 18172 20914 18228 20916
rect 18172 20862 18174 20914
rect 18174 20862 18226 20914
rect 18226 20862 18228 20914
rect 18172 20860 18228 20862
rect 17948 20524 18004 20580
rect 18060 20018 18116 20020
rect 18060 19966 18062 20018
rect 18062 19966 18114 20018
rect 18114 19966 18116 20018
rect 18060 19964 18116 19966
rect 18060 19516 18116 19572
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 17948 18172 18004 18228
rect 17388 16268 17444 16324
rect 17500 14924 17556 14980
rect 17500 14140 17556 14196
rect 16492 12684 16548 12740
rect 16156 11788 16212 11844
rect 16156 11116 16212 11172
rect 16380 11340 16436 11396
rect 16268 11004 16324 11060
rect 16044 9996 16100 10052
rect 16604 11116 16660 11172
rect 16716 10780 16772 10836
rect 16828 10556 16884 10612
rect 16940 11116 16996 11172
rect 16716 10444 16772 10500
rect 17388 13916 17444 13972
rect 17500 12908 17556 12964
rect 17724 17106 17780 17108
rect 17724 17054 17726 17106
rect 17726 17054 17778 17106
rect 17778 17054 17780 17106
rect 17724 17052 17780 17054
rect 17836 16604 17892 16660
rect 17836 16044 17892 16100
rect 18172 15986 18228 15988
rect 18172 15934 18174 15986
rect 18174 15934 18226 15986
rect 18226 15934 18228 15986
rect 18172 15932 18228 15934
rect 18172 15260 18228 15316
rect 17948 15148 18004 15204
rect 17724 14476 17780 14532
rect 17388 11340 17444 11396
rect 17500 10892 17556 10948
rect 17276 10780 17332 10836
rect 16492 9996 16548 10052
rect 16156 9938 16212 9940
rect 16156 9886 16158 9938
rect 16158 9886 16210 9938
rect 16210 9886 16212 9938
rect 16156 9884 16212 9886
rect 15820 9436 15876 9492
rect 15708 8764 15764 8820
rect 15596 8204 15652 8260
rect 14700 6524 14756 6580
rect 14252 6412 14308 6468
rect 13916 5068 13972 5124
rect 13580 5010 13636 5012
rect 13580 4958 13582 5010
rect 13582 4958 13634 5010
rect 13634 4958 13636 5010
rect 13580 4956 13636 4958
rect 13020 4508 13076 4564
rect 12908 4396 12964 4452
rect 13020 3778 13076 3780
rect 13020 3726 13022 3778
rect 13022 3726 13074 3778
rect 13074 3726 13076 3778
rect 13020 3724 13076 3726
rect 12684 3666 12740 3668
rect 12684 3614 12686 3666
rect 12686 3614 12738 3666
rect 12738 3614 12740 3666
rect 12684 3612 12740 3614
rect 13468 4284 13524 4340
rect 13356 4226 13412 4228
rect 13356 4174 13358 4226
rect 13358 4174 13410 4226
rect 13410 4174 13412 4226
rect 13356 4172 13412 4174
rect 13580 4172 13636 4228
rect 13916 4172 13972 4228
rect 14140 5180 14196 5236
rect 14028 3948 14084 4004
rect 14252 3724 14308 3780
rect 14476 6018 14532 6020
rect 14476 5966 14478 6018
rect 14478 5966 14530 6018
rect 14530 5966 14532 6018
rect 14476 5964 14532 5966
rect 13020 3052 13076 3108
rect 12796 2546 12852 2548
rect 12796 2494 12798 2546
rect 12798 2494 12850 2546
rect 12850 2494 12852 2546
rect 12796 2492 12852 2494
rect 13580 2716 13636 2772
rect 12348 1932 12404 1988
rect 12908 1986 12964 1988
rect 12908 1934 12910 1986
rect 12910 1934 12962 1986
rect 12962 1934 12964 1986
rect 12908 1932 12964 1934
rect 13468 1708 13524 1764
rect 12348 1596 12404 1652
rect 11564 812 11620 868
rect 11900 700 11956 756
rect 13244 1596 13300 1652
rect 12796 1260 12852 1316
rect 12572 1202 12628 1204
rect 12572 1150 12574 1202
rect 12574 1150 12626 1202
rect 12626 1150 12628 1202
rect 12572 1148 12628 1150
rect 7644 28 7700 84
rect 13804 2882 13860 2884
rect 13804 2830 13806 2882
rect 13806 2830 13858 2882
rect 13858 2830 13860 2882
rect 13804 2828 13860 2830
rect 13916 2380 13972 2436
rect 14252 3276 14308 3332
rect 14252 2380 14308 2436
rect 14252 1932 14308 1988
rect 14588 5794 14644 5796
rect 14588 5742 14590 5794
rect 14590 5742 14642 5794
rect 14642 5742 14644 5794
rect 14588 5740 14644 5742
rect 14588 5516 14644 5572
rect 14924 5516 14980 5572
rect 14476 5180 14532 5236
rect 14700 4844 14756 4900
rect 14588 4562 14644 4564
rect 14588 4510 14590 4562
rect 14590 4510 14642 4562
rect 14642 4510 14644 4562
rect 14588 4508 14644 4510
rect 14476 2828 14532 2884
rect 15260 6802 15316 6804
rect 15260 6750 15262 6802
rect 15262 6750 15314 6802
rect 15314 6750 15316 6802
rect 15260 6748 15316 6750
rect 15148 4956 15204 5012
rect 15260 6300 15316 6356
rect 16044 9660 16100 9716
rect 16044 9324 16100 9380
rect 16268 9548 16324 9604
rect 16268 9324 16324 9380
rect 16828 9826 16884 9828
rect 16828 9774 16830 9826
rect 16830 9774 16882 9826
rect 16882 9774 16884 9826
rect 16828 9772 16884 9774
rect 16940 9660 16996 9716
rect 16604 9324 16660 9380
rect 16716 9042 16772 9044
rect 16716 8990 16718 9042
rect 16718 8990 16770 9042
rect 16770 8990 16772 9042
rect 16716 8988 16772 8990
rect 16940 8370 16996 8372
rect 16940 8318 16942 8370
rect 16942 8318 16994 8370
rect 16994 8318 16996 8370
rect 16940 8316 16996 8318
rect 16268 8204 16324 8260
rect 16156 7420 16212 7476
rect 17276 9772 17332 9828
rect 17052 7756 17108 7812
rect 16716 7532 16772 7588
rect 15820 7308 15876 7364
rect 16492 7308 16548 7364
rect 15932 6972 15988 7028
rect 16268 7196 16324 7252
rect 15932 6802 15988 6804
rect 15932 6750 15934 6802
rect 15934 6750 15986 6802
rect 15986 6750 15988 6802
rect 15932 6748 15988 6750
rect 15708 6690 15764 6692
rect 15708 6638 15710 6690
rect 15710 6638 15762 6690
rect 15762 6638 15764 6690
rect 15708 6636 15764 6638
rect 15596 6300 15652 6356
rect 15932 6300 15988 6356
rect 15484 5964 15540 6020
rect 15820 5964 15876 6020
rect 15932 5794 15988 5796
rect 15932 5742 15934 5794
rect 15934 5742 15986 5794
rect 15986 5742 15988 5794
rect 15932 5740 15988 5742
rect 16268 5964 16324 6020
rect 16156 5068 16212 5124
rect 16604 6636 16660 6692
rect 16716 6076 16772 6132
rect 17052 6690 17108 6692
rect 17052 6638 17054 6690
rect 17054 6638 17106 6690
rect 17106 6638 17108 6690
rect 17052 6636 17108 6638
rect 17164 6524 17220 6580
rect 15260 4732 15316 4788
rect 14924 4060 14980 4116
rect 14924 3666 14980 3668
rect 14924 3614 14926 3666
rect 14926 3614 14978 3666
rect 14978 3614 14980 3666
rect 14924 3612 14980 3614
rect 16604 4732 16660 4788
rect 16268 4508 16324 4564
rect 15932 4338 15988 4340
rect 15932 4286 15934 4338
rect 15934 4286 15986 4338
rect 15986 4286 15988 4338
rect 15932 4284 15988 4286
rect 16828 4508 16884 4564
rect 16940 4956 16996 5012
rect 15932 3724 15988 3780
rect 16156 3500 16212 3556
rect 16268 4060 16324 4116
rect 14700 3164 14756 3220
rect 15820 3276 15876 3332
rect 14700 2604 14756 2660
rect 15596 2716 15652 2772
rect 15260 2268 15316 2324
rect 14924 2210 14980 2212
rect 14924 2158 14926 2210
rect 14926 2158 14978 2210
rect 14978 2158 14980 2210
rect 14924 2156 14980 2158
rect 16156 2940 16212 2996
rect 14588 2098 14644 2100
rect 14588 2046 14590 2098
rect 14590 2046 14642 2098
rect 14642 2046 14644 2098
rect 14588 2044 14644 2046
rect 16828 3948 16884 4004
rect 16716 3724 16772 3780
rect 16604 3554 16660 3556
rect 16604 3502 16606 3554
rect 16606 3502 16658 3554
rect 16658 3502 16660 3554
rect 16604 3500 16660 3502
rect 16492 3388 16548 3444
rect 14364 1708 14420 1764
rect 16044 1762 16100 1764
rect 16044 1710 16046 1762
rect 16046 1710 16098 1762
rect 16098 1710 16100 1762
rect 16044 1708 16100 1710
rect 14588 1596 14644 1652
rect 14140 924 14196 980
rect 13692 812 13748 868
rect 15036 1596 15092 1652
rect 15932 1596 15988 1652
rect 15484 1202 15540 1204
rect 15484 1150 15486 1202
rect 15486 1150 15538 1202
rect 15538 1150 15540 1202
rect 15484 1148 15540 1150
rect 15148 700 15204 756
rect 15484 700 15540 756
rect 16380 1596 16436 1652
rect 16268 476 16324 532
rect 17500 9042 17556 9044
rect 17500 8990 17502 9042
rect 17502 8990 17554 9042
rect 17554 8990 17556 9042
rect 17500 8988 17556 8990
rect 17388 8258 17444 8260
rect 17388 8206 17390 8258
rect 17390 8206 17442 8258
rect 17442 8206 17444 8258
rect 17388 8204 17444 8206
rect 17388 7362 17444 7364
rect 17388 7310 17390 7362
rect 17390 7310 17442 7362
rect 17442 7310 17444 7362
rect 17388 7308 17444 7310
rect 17836 13244 17892 13300
rect 17948 11228 18004 11284
rect 18172 14476 18228 14532
rect 17724 11116 17780 11172
rect 17836 10610 17892 10612
rect 17836 10558 17838 10610
rect 17838 10558 17890 10610
rect 17890 10558 17892 10610
rect 17836 10556 17892 10558
rect 18060 9996 18116 10052
rect 17724 9938 17780 9940
rect 17724 9886 17726 9938
rect 17726 9886 17778 9938
rect 17778 9886 17780 9938
rect 17724 9884 17780 9886
rect 17836 9660 17892 9716
rect 18508 25676 18564 25732
rect 18732 27074 18788 27076
rect 18732 27022 18734 27074
rect 18734 27022 18786 27074
rect 18786 27022 18788 27074
rect 18732 27020 18788 27022
rect 19068 30434 19124 30436
rect 19068 30382 19070 30434
rect 19070 30382 19122 30434
rect 19122 30382 19124 30434
rect 19068 30380 19124 30382
rect 18956 30268 19012 30324
rect 19628 30828 19684 30884
rect 19964 34076 20020 34132
rect 19852 33740 19908 33796
rect 21084 37548 21140 37604
rect 22092 46562 22148 46564
rect 22092 46510 22094 46562
rect 22094 46510 22146 46562
rect 22146 46510 22148 46562
rect 22092 46508 22148 46510
rect 21756 46114 21812 46116
rect 21756 46062 21758 46114
rect 21758 46062 21810 46114
rect 21810 46062 21812 46114
rect 21756 46060 21812 46062
rect 21980 46060 22036 46116
rect 21644 45612 21700 45668
rect 21980 45612 22036 45668
rect 21644 45052 21700 45108
rect 21644 43372 21700 43428
rect 21756 43260 21812 43316
rect 21868 43484 21924 43540
rect 21756 43036 21812 43092
rect 21420 40348 21476 40404
rect 21644 40572 21700 40628
rect 21308 38946 21364 38948
rect 21308 38894 21310 38946
rect 21310 38894 21362 38946
rect 21362 38894 21364 38946
rect 21308 38892 21364 38894
rect 21644 38722 21700 38724
rect 21644 38670 21646 38722
rect 21646 38670 21698 38722
rect 21698 38670 21700 38722
rect 21644 38668 21700 38670
rect 21308 36988 21364 37044
rect 20972 36764 21028 36820
rect 20636 35084 20692 35140
rect 21084 36092 21140 36148
rect 20524 34860 20580 34916
rect 20972 34972 21028 35028
rect 20748 34802 20804 34804
rect 20748 34750 20750 34802
rect 20750 34750 20802 34802
rect 20802 34750 20804 34802
rect 20748 34748 20804 34750
rect 20524 34130 20580 34132
rect 20524 34078 20526 34130
rect 20526 34078 20578 34130
rect 20578 34078 20580 34130
rect 20524 34076 20580 34078
rect 20860 34130 20916 34132
rect 20860 34078 20862 34130
rect 20862 34078 20914 34130
rect 20914 34078 20916 34130
rect 20860 34076 20916 34078
rect 20748 34018 20804 34020
rect 20748 33966 20750 34018
rect 20750 33966 20802 34018
rect 20802 33966 20804 34018
rect 20748 33964 20804 33966
rect 20188 33740 20244 33796
rect 20636 33740 20692 33796
rect 19964 33346 20020 33348
rect 19964 33294 19966 33346
rect 19966 33294 20018 33346
rect 20018 33294 20020 33346
rect 19964 33292 20020 33294
rect 21084 33292 21140 33348
rect 20748 33068 20804 33124
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 19852 30604 19908 30660
rect 19740 30268 19796 30324
rect 19964 30380 20020 30436
rect 19628 30156 19684 30212
rect 19180 29932 19236 29988
rect 19516 29932 19572 29988
rect 19180 29426 19236 29428
rect 19180 29374 19182 29426
rect 19182 29374 19234 29426
rect 19234 29374 19236 29426
rect 19180 29372 19236 29374
rect 20076 30828 20132 30884
rect 19852 30044 19908 30100
rect 19068 29314 19124 29316
rect 19068 29262 19070 29314
rect 19070 29262 19122 29314
rect 19122 29262 19124 29314
rect 19068 29260 19124 29262
rect 19180 29148 19236 29204
rect 19068 28866 19124 28868
rect 19068 28814 19070 28866
rect 19070 28814 19122 28866
rect 19122 28814 19124 28866
rect 19068 28812 19124 28814
rect 19852 29148 19908 29204
rect 19516 28588 19572 28644
rect 19292 28530 19348 28532
rect 19292 28478 19294 28530
rect 19294 28478 19346 28530
rect 19346 28478 19348 28530
rect 19292 28476 19348 28478
rect 19180 27916 19236 27972
rect 19068 27858 19124 27860
rect 19068 27806 19070 27858
rect 19070 27806 19122 27858
rect 19122 27806 19124 27858
rect 19068 27804 19124 27806
rect 19404 27916 19460 27972
rect 19628 27858 19684 27860
rect 19628 27806 19630 27858
rect 19630 27806 19682 27858
rect 19682 27806 19684 27858
rect 19628 27804 19684 27806
rect 19404 27580 19460 27636
rect 20076 29036 20132 29092
rect 20748 31500 20804 31556
rect 21420 35084 21476 35140
rect 21420 32620 21476 32676
rect 20636 31276 20692 31332
rect 20524 31164 20580 31220
rect 21308 32450 21364 32452
rect 21308 32398 21310 32450
rect 21310 32398 21362 32450
rect 21362 32398 21364 32450
rect 21308 32396 21364 32398
rect 21196 31948 21252 32004
rect 20860 31106 20916 31108
rect 20860 31054 20862 31106
rect 20862 31054 20914 31106
rect 20914 31054 20916 31106
rect 20860 31052 20916 31054
rect 20300 30828 20356 30884
rect 20412 29932 20468 29988
rect 20076 28476 20132 28532
rect 21420 31164 21476 31220
rect 20972 30210 21028 30212
rect 20972 30158 20974 30210
rect 20974 30158 21026 30210
rect 21026 30158 21028 30210
rect 20972 30156 21028 30158
rect 21196 30156 21252 30212
rect 21196 29932 21252 29988
rect 20636 29314 20692 29316
rect 20636 29262 20638 29314
rect 20638 29262 20690 29314
rect 20690 29262 20692 29314
rect 20636 29260 20692 29262
rect 20748 28812 20804 28868
rect 20636 28754 20692 28756
rect 20636 28702 20638 28754
rect 20638 28702 20690 28754
rect 20690 28702 20692 28754
rect 20636 28700 20692 28702
rect 20860 28588 20916 28644
rect 20972 28700 21028 28756
rect 20524 28476 20580 28532
rect 20076 27468 20132 27524
rect 18956 27132 19012 27188
rect 19180 27020 19236 27076
rect 18956 25340 19012 25396
rect 18844 24892 18900 24948
rect 19852 27132 19908 27188
rect 19740 26348 19796 26404
rect 19404 25340 19460 25396
rect 19516 26012 19572 26068
rect 19180 23884 19236 23940
rect 18396 22652 18452 22708
rect 18396 22204 18452 22260
rect 18508 21756 18564 21812
rect 18844 23100 18900 23156
rect 18620 20412 18676 20468
rect 18732 22988 18788 23044
rect 18508 20188 18564 20244
rect 18844 21362 18900 21364
rect 18844 21310 18846 21362
rect 18846 21310 18898 21362
rect 18898 21310 18900 21362
rect 18844 21308 18900 21310
rect 18844 20636 18900 20692
rect 18508 19628 18564 19684
rect 18396 19404 18452 19460
rect 18396 17164 18452 17220
rect 18732 17276 18788 17332
rect 18508 16210 18564 16212
rect 18508 16158 18510 16210
rect 18510 16158 18562 16210
rect 18562 16158 18564 16210
rect 18508 16156 18564 16158
rect 18956 19852 19012 19908
rect 18956 19292 19012 19348
rect 18956 17836 19012 17892
rect 18956 16828 19012 16884
rect 18956 15372 19012 15428
rect 19292 24332 19348 24388
rect 19404 23378 19460 23380
rect 19404 23326 19406 23378
rect 19406 23326 19458 23378
rect 19458 23326 19460 23378
rect 19404 23324 19460 23326
rect 19404 23100 19460 23156
rect 19740 26012 19796 26068
rect 19740 25506 19796 25508
rect 19740 25454 19742 25506
rect 19742 25454 19794 25506
rect 19794 25454 19796 25506
rect 19740 25452 19796 25454
rect 19628 24722 19684 24724
rect 19628 24670 19630 24722
rect 19630 24670 19682 24722
rect 19682 24670 19684 24722
rect 19628 24668 19684 24670
rect 19740 24444 19796 24500
rect 19740 23938 19796 23940
rect 19740 23886 19742 23938
rect 19742 23886 19794 23938
rect 19794 23886 19796 23938
rect 19740 23884 19796 23886
rect 19740 23100 19796 23156
rect 19628 22428 19684 22484
rect 19740 22876 19796 22932
rect 19516 22370 19572 22372
rect 19516 22318 19518 22370
rect 19518 22318 19570 22370
rect 19570 22318 19572 22370
rect 19516 22316 19572 22318
rect 19292 19404 19348 19460
rect 19404 19292 19460 19348
rect 19180 17836 19236 17892
rect 19292 17164 19348 17220
rect 19404 18060 19460 18116
rect 19628 20076 19684 20132
rect 18956 14812 19012 14868
rect 18396 14476 18452 14532
rect 18508 13522 18564 13524
rect 18508 13470 18510 13522
rect 18510 13470 18562 13522
rect 18562 13470 18564 13522
rect 18508 13468 18564 13470
rect 18620 13020 18676 13076
rect 18508 12348 18564 12404
rect 18396 12178 18452 12180
rect 18396 12126 18398 12178
rect 18398 12126 18450 12178
rect 18450 12126 18452 12178
rect 18396 12124 18452 12126
rect 18508 11116 18564 11172
rect 18508 10610 18564 10612
rect 18508 10558 18510 10610
rect 18510 10558 18562 10610
rect 18562 10558 18564 10610
rect 18508 10556 18564 10558
rect 18060 8428 18116 8484
rect 18396 9212 18452 9268
rect 17948 8204 18004 8260
rect 17612 8092 17668 8148
rect 18060 8092 18116 8148
rect 17612 7756 17668 7812
rect 17948 7084 18004 7140
rect 18060 6802 18116 6804
rect 18060 6750 18062 6802
rect 18062 6750 18114 6802
rect 18114 6750 18116 6802
rect 18060 6748 18116 6750
rect 17948 6076 18004 6132
rect 17500 4732 17556 4788
rect 17052 4060 17108 4116
rect 16716 2658 16772 2660
rect 16716 2606 16718 2658
rect 16718 2606 16770 2658
rect 16770 2606 16772 2658
rect 16716 2604 16772 2606
rect 19068 13468 19124 13524
rect 18956 12850 19012 12852
rect 18956 12798 18958 12850
rect 18958 12798 19010 12850
rect 19010 12798 19012 12850
rect 18956 12796 19012 12798
rect 19292 13580 19348 13636
rect 19516 17052 19572 17108
rect 19964 25564 20020 25620
rect 19964 24668 20020 24724
rect 19964 22876 20020 22932
rect 21196 28588 21252 28644
rect 21980 42252 22036 42308
rect 22204 44156 22260 44212
rect 21980 41970 22036 41972
rect 21980 41918 21982 41970
rect 21982 41918 22034 41970
rect 22034 41918 22036 41970
rect 21980 41916 22036 41918
rect 21980 41692 22036 41748
rect 22092 41298 22148 41300
rect 22092 41246 22094 41298
rect 22094 41246 22146 41298
rect 22146 41246 22148 41298
rect 22092 41244 22148 41246
rect 21980 40684 22036 40740
rect 22092 40348 22148 40404
rect 22540 48300 22596 48356
rect 22540 46508 22596 46564
rect 22764 47628 22820 47684
rect 22764 46844 22820 46900
rect 22764 45890 22820 45892
rect 22764 45838 22766 45890
rect 22766 45838 22818 45890
rect 22818 45838 22820 45890
rect 22764 45836 22820 45838
rect 22652 45388 22708 45444
rect 22540 44994 22596 44996
rect 22540 44942 22542 44994
rect 22542 44942 22594 44994
rect 22594 44942 22596 44994
rect 22540 44940 22596 44942
rect 22428 44604 22484 44660
rect 22428 44156 22484 44212
rect 22540 44380 22596 44436
rect 22316 42252 22372 42308
rect 22428 43708 22484 43764
rect 22316 41916 22372 41972
rect 22764 44268 22820 44324
rect 22652 43314 22708 43316
rect 22652 43262 22654 43314
rect 22654 43262 22706 43314
rect 22706 43262 22708 43314
rect 22652 43260 22708 43262
rect 22540 41970 22596 41972
rect 22540 41918 22542 41970
rect 22542 41918 22594 41970
rect 22594 41918 22596 41970
rect 22540 41916 22596 41918
rect 22764 41244 22820 41300
rect 22428 40460 22484 40516
rect 22764 40460 22820 40516
rect 22652 40236 22708 40292
rect 22988 53730 23044 53732
rect 22988 53678 22990 53730
rect 22990 53678 23042 53730
rect 23042 53678 23044 53730
rect 22988 53676 23044 53678
rect 23100 53228 23156 53284
rect 23100 51324 23156 51380
rect 23100 50988 23156 51044
rect 23548 55410 23604 55412
rect 23548 55358 23550 55410
rect 23550 55358 23602 55410
rect 23602 55358 23604 55410
rect 23548 55356 23604 55358
rect 23436 54290 23492 54292
rect 23436 54238 23438 54290
rect 23438 54238 23490 54290
rect 23490 54238 23492 54290
rect 23436 54236 23492 54238
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 23772 54684 23828 54740
rect 23884 54290 23940 54292
rect 23884 54238 23886 54290
rect 23886 54238 23938 54290
rect 23938 54238 23940 54290
rect 23884 54236 23940 54238
rect 23324 53564 23380 53620
rect 24108 53788 24164 53844
rect 23212 49196 23268 49252
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 24780 55132 24836 55188
rect 24556 54572 24612 54628
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 24220 53564 24276 53620
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 24220 53340 24276 53396
rect 24108 53116 24164 53172
rect 23548 52444 23604 52500
rect 23660 52892 23716 52948
rect 23660 52220 23716 52276
rect 23884 52274 23940 52276
rect 23884 52222 23886 52274
rect 23886 52222 23938 52274
rect 23938 52222 23940 52274
rect 23884 52220 23940 52222
rect 24220 52892 24276 52948
rect 24220 52108 24276 52164
rect 24668 53730 24724 53732
rect 24668 53678 24670 53730
rect 24670 53678 24722 53730
rect 24722 53678 24724 53730
rect 24668 53676 24724 53678
rect 24780 53116 24836 53172
rect 25340 55804 25396 55860
rect 25116 53340 25172 53396
rect 25340 54124 25396 54180
rect 24892 53004 24948 53060
rect 24668 52780 24724 52836
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 25004 52892 25060 52948
rect 25676 54460 25732 54516
rect 25564 54124 25620 54180
rect 26124 55580 26180 55636
rect 26684 56812 26740 56868
rect 27132 56028 27188 56084
rect 26908 55916 26964 55972
rect 26460 55858 26516 55860
rect 26460 55806 26462 55858
rect 26462 55806 26514 55858
rect 26514 55806 26516 55858
rect 26460 55804 26516 55806
rect 26236 55468 26292 55524
rect 26124 54348 26180 54404
rect 25788 53788 25844 53844
rect 25452 53730 25508 53732
rect 25452 53678 25454 53730
rect 25454 53678 25506 53730
rect 25506 53678 25508 53730
rect 25452 53676 25508 53678
rect 25676 53676 25732 53732
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 24012 51716 24068 51718
rect 23772 51548 23828 51604
rect 23436 50988 23492 51044
rect 23996 51548 24052 51604
rect 24332 51266 24388 51268
rect 24332 51214 24334 51266
rect 24334 51214 24386 51266
rect 24386 51214 24388 51266
rect 24332 51212 24388 51214
rect 25340 52722 25396 52724
rect 25340 52670 25342 52722
rect 25342 52670 25394 52722
rect 25394 52670 25396 52722
rect 25340 52668 25396 52670
rect 25228 52220 25284 52276
rect 25004 51548 25060 51604
rect 24668 51378 24724 51380
rect 24668 51326 24670 51378
rect 24670 51326 24722 51378
rect 24722 51326 24724 51378
rect 24668 51324 24724 51326
rect 25004 51324 25060 51380
rect 24108 50988 24164 51044
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 24108 50764 24164 50820
rect 25004 50652 25060 50708
rect 24332 50428 24388 50484
rect 23436 50204 23492 50260
rect 23436 49980 23492 50036
rect 23436 49532 23492 49588
rect 23660 50204 23716 50260
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 24220 50092 24276 50148
rect 23996 49980 24052 50036
rect 23548 49420 23604 49476
rect 24556 50482 24612 50484
rect 24556 50430 24558 50482
rect 24558 50430 24610 50482
rect 24610 50430 24612 50482
rect 24556 50428 24612 50430
rect 24220 49420 24276 49476
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 23324 48412 23380 48468
rect 23436 49084 23492 49140
rect 23324 47628 23380 47684
rect 23324 46898 23380 46900
rect 23324 46846 23326 46898
rect 23326 46846 23378 46898
rect 23378 46846 23380 46898
rect 23324 46844 23380 46846
rect 22988 41132 23044 41188
rect 23100 40348 23156 40404
rect 21756 37884 21812 37940
rect 21868 36764 21924 36820
rect 21756 36316 21812 36372
rect 21868 35532 21924 35588
rect 21644 35084 21700 35140
rect 21756 34076 21812 34132
rect 21644 33964 21700 34020
rect 21868 33628 21924 33684
rect 21756 33346 21812 33348
rect 21756 33294 21758 33346
rect 21758 33294 21810 33346
rect 21810 33294 21812 33346
rect 21756 33292 21812 33294
rect 21532 30828 21588 30884
rect 21644 32620 21700 32676
rect 22316 37884 22372 37940
rect 22092 36482 22148 36484
rect 22092 36430 22094 36482
rect 22094 36430 22146 36482
rect 22146 36430 22148 36482
rect 22092 36428 22148 36430
rect 22204 36316 22260 36372
rect 22092 35586 22148 35588
rect 22092 35534 22094 35586
rect 22094 35534 22146 35586
rect 22146 35534 22148 35586
rect 22092 35532 22148 35534
rect 22204 35026 22260 35028
rect 22204 34974 22206 35026
rect 22206 34974 22258 35026
rect 22258 34974 22260 35026
rect 22204 34972 22260 34974
rect 21868 32620 21924 32676
rect 21980 33180 22036 33236
rect 21980 31836 22036 31892
rect 21644 30604 21700 30660
rect 21756 31052 21812 31108
rect 21420 29820 21476 29876
rect 21644 30380 21700 30436
rect 21308 28476 21364 28532
rect 20636 27858 20692 27860
rect 20636 27806 20638 27858
rect 20638 27806 20690 27858
rect 20690 27806 20692 27858
rect 20636 27804 20692 27806
rect 20524 27356 20580 27412
rect 20524 27132 20580 27188
rect 20972 27356 21028 27412
rect 20524 26908 20580 26964
rect 20524 26684 20580 26740
rect 20972 26684 21028 26740
rect 20860 26460 20916 26516
rect 20412 25676 20468 25732
rect 21308 27468 21364 27524
rect 21308 27132 21364 27188
rect 21196 26460 21252 26516
rect 21308 26796 21364 26852
rect 21196 26236 21252 26292
rect 20636 25676 20692 25732
rect 20636 25506 20692 25508
rect 20636 25454 20638 25506
rect 20638 25454 20690 25506
rect 20690 25454 20692 25506
rect 20636 25452 20692 25454
rect 20524 25340 20580 25396
rect 20524 24892 20580 24948
rect 20524 23100 20580 23156
rect 19852 20748 19908 20804
rect 19964 20412 20020 20468
rect 19740 19516 19796 19572
rect 20300 19458 20356 19460
rect 20300 19406 20302 19458
rect 20302 19406 20354 19458
rect 20354 19406 20356 19458
rect 20300 19404 20356 19406
rect 20076 19234 20132 19236
rect 20076 19182 20078 19234
rect 20078 19182 20130 19234
rect 20130 19182 20132 19234
rect 20076 19180 20132 19182
rect 20524 22428 20580 22484
rect 21308 25900 21364 25956
rect 20972 25564 21028 25620
rect 21196 25564 21252 25620
rect 21084 25452 21140 25508
rect 21644 30156 21700 30212
rect 22540 39900 22596 39956
rect 22540 39618 22596 39620
rect 22540 39566 22542 39618
rect 22542 39566 22594 39618
rect 22594 39566 22596 39618
rect 22540 39564 22596 39566
rect 22876 37884 22932 37940
rect 22540 37154 22596 37156
rect 22540 37102 22542 37154
rect 22542 37102 22594 37154
rect 22594 37102 22596 37154
rect 22540 37100 22596 37102
rect 22428 35644 22484 35700
rect 22764 36988 22820 37044
rect 22652 33516 22708 33572
rect 22316 32732 22372 32788
rect 22540 33292 22596 33348
rect 22428 31836 22484 31892
rect 22092 30940 22148 30996
rect 22428 31218 22484 31220
rect 22428 31166 22430 31218
rect 22430 31166 22482 31218
rect 22482 31166 22484 31218
rect 22428 31164 22484 31166
rect 22316 30044 22372 30100
rect 21868 29484 21924 29540
rect 21532 27356 21588 27412
rect 21532 27132 21588 27188
rect 22092 29314 22148 29316
rect 22092 29262 22094 29314
rect 22094 29262 22146 29314
rect 22146 29262 22148 29314
rect 22092 29260 22148 29262
rect 22204 28700 22260 28756
rect 22092 28642 22148 28644
rect 22092 28590 22094 28642
rect 22094 28590 22146 28642
rect 22146 28590 22148 28642
rect 22092 28588 22148 28590
rect 21756 27468 21812 27524
rect 21756 26684 21812 26740
rect 21868 27132 21924 27188
rect 21644 26290 21700 26292
rect 21644 26238 21646 26290
rect 21646 26238 21698 26290
rect 21698 26238 21700 26290
rect 21644 26236 21700 26238
rect 21196 24332 21252 24388
rect 21644 24556 21700 24612
rect 21308 24220 21364 24276
rect 21644 24332 21700 24388
rect 20860 23996 20916 24052
rect 21420 24050 21476 24052
rect 21420 23998 21422 24050
rect 21422 23998 21474 24050
rect 21474 23998 21476 24050
rect 21420 23996 21476 23998
rect 21868 26348 21924 26404
rect 22092 27916 22148 27972
rect 22652 31052 22708 31108
rect 22652 30492 22708 30548
rect 22316 28140 22372 28196
rect 22316 27356 22372 27412
rect 22204 25900 22260 25956
rect 22316 25788 22372 25844
rect 22540 24892 22596 24948
rect 22652 25116 22708 25172
rect 20748 23100 20804 23156
rect 21084 23772 21140 23828
rect 20748 22876 20804 22932
rect 20972 22594 21028 22596
rect 20972 22542 20974 22594
rect 20974 22542 21026 22594
rect 21026 22542 21028 22594
rect 20972 22540 21028 22542
rect 20748 22204 20804 22260
rect 20524 21196 20580 21252
rect 20972 21532 21028 21588
rect 21308 23772 21364 23828
rect 21868 23772 21924 23828
rect 21196 23660 21252 23716
rect 21532 23660 21588 23716
rect 21308 23436 21364 23492
rect 21868 23324 21924 23380
rect 22092 23436 22148 23492
rect 21532 22652 21588 22708
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 21420 21196 21476 21252
rect 20748 20412 20804 20468
rect 20860 20636 20916 20692
rect 20748 19346 20804 19348
rect 20748 19294 20750 19346
rect 20750 19294 20802 19346
rect 20802 19294 20804 19346
rect 20748 19292 20804 19294
rect 20412 18732 20468 18788
rect 20412 18508 20468 18564
rect 20300 18396 20356 18452
rect 20188 17890 20244 17892
rect 20188 17838 20190 17890
rect 20190 17838 20242 17890
rect 20242 17838 20244 17890
rect 20188 17836 20244 17838
rect 20076 17164 20132 17220
rect 19628 16268 19684 16324
rect 19964 16828 20020 16884
rect 19740 16098 19796 16100
rect 19740 16046 19742 16098
rect 19742 16046 19794 16098
rect 19794 16046 19796 16098
rect 19740 16044 19796 16046
rect 19852 15708 19908 15764
rect 19740 14812 19796 14868
rect 19404 13020 19460 13076
rect 19516 14028 19572 14084
rect 19068 12124 19124 12180
rect 19180 12066 19236 12068
rect 19180 12014 19182 12066
rect 19182 12014 19234 12066
rect 19234 12014 19236 12066
rect 19180 12012 19236 12014
rect 18732 11564 18788 11620
rect 18844 11676 18900 11732
rect 19180 11340 19236 11396
rect 19180 11116 19236 11172
rect 18956 10556 19012 10612
rect 18732 9714 18788 9716
rect 18732 9662 18734 9714
rect 18734 9662 18786 9714
rect 18786 9662 18788 9714
rect 18732 9660 18788 9662
rect 18620 8988 18676 9044
rect 17612 3500 17668 3556
rect 17276 2882 17332 2884
rect 17276 2830 17278 2882
rect 17278 2830 17330 2882
rect 17330 2830 17332 2882
rect 17276 2828 17332 2830
rect 17500 2828 17556 2884
rect 17164 2604 17220 2660
rect 16716 1148 16772 1204
rect 16828 1596 16884 1652
rect 17276 1596 17332 1652
rect 17724 2546 17780 2548
rect 17724 2494 17726 2546
rect 17726 2494 17778 2546
rect 17778 2494 17780 2546
rect 17724 2492 17780 2494
rect 17612 2268 17668 2324
rect 17724 2098 17780 2100
rect 17724 2046 17726 2098
rect 17726 2046 17778 2098
rect 17778 2046 17780 2098
rect 17724 2044 17780 2046
rect 18844 8988 18900 9044
rect 18396 8428 18452 8484
rect 18620 8316 18676 8372
rect 18620 6636 18676 6692
rect 19068 10108 19124 10164
rect 19068 9324 19124 9380
rect 19180 9660 19236 9716
rect 19180 8428 19236 8484
rect 19068 8258 19124 8260
rect 19068 8206 19070 8258
rect 19070 8206 19122 8258
rect 19122 8206 19124 8258
rect 19068 8204 19124 8206
rect 18396 5852 18452 5908
rect 18508 6300 18564 6356
rect 19516 11676 19572 11732
rect 20188 16492 20244 16548
rect 20412 17836 20468 17892
rect 21084 20636 21140 20692
rect 20524 16098 20580 16100
rect 20524 16046 20526 16098
rect 20526 16046 20578 16098
rect 20578 16046 20580 16098
rect 20524 16044 20580 16046
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 21532 19964 21588 20020
rect 21308 19516 21364 19572
rect 21532 19516 21588 19572
rect 21420 19180 21476 19236
rect 21980 22428 22036 22484
rect 21868 20524 21924 20580
rect 21756 19180 21812 19236
rect 21532 18172 21588 18228
rect 21308 17612 21364 17668
rect 21196 17554 21252 17556
rect 21196 17502 21198 17554
rect 21198 17502 21250 17554
rect 21250 17502 21252 17554
rect 21196 17500 21252 17502
rect 20860 17164 20916 17220
rect 21756 17164 21812 17220
rect 21308 16828 21364 16884
rect 21196 16322 21252 16324
rect 21196 16270 21198 16322
rect 21198 16270 21250 16322
rect 21250 16270 21252 16322
rect 21196 16268 21252 16270
rect 20412 15932 20468 15988
rect 20076 14812 20132 14868
rect 21532 16492 21588 16548
rect 20972 14812 21028 14868
rect 21084 15148 21140 15204
rect 19852 14252 19908 14308
rect 19740 13692 19796 13748
rect 19740 13522 19796 13524
rect 19740 13470 19742 13522
rect 19742 13470 19794 13522
rect 19794 13470 19796 13522
rect 19740 13468 19796 13470
rect 20636 14476 20692 14532
rect 20188 13132 20244 13188
rect 20188 12962 20244 12964
rect 20188 12910 20190 12962
rect 20190 12910 20242 12962
rect 20242 12910 20244 12962
rect 20188 12908 20244 12910
rect 20748 13468 20804 13524
rect 20972 14028 21028 14084
rect 21084 13468 21140 13524
rect 19852 12178 19908 12180
rect 19852 12126 19854 12178
rect 19854 12126 19906 12178
rect 19906 12126 19908 12178
rect 19852 12124 19908 12126
rect 20076 12178 20132 12180
rect 20076 12126 20078 12178
rect 20078 12126 20130 12178
rect 20130 12126 20132 12178
rect 20076 12124 20132 12126
rect 19740 11676 19796 11732
rect 20300 12012 20356 12068
rect 20188 11618 20244 11620
rect 20188 11566 20190 11618
rect 20190 11566 20242 11618
rect 20242 11566 20244 11618
rect 20188 11564 20244 11566
rect 19628 11452 19684 11508
rect 19404 9996 19460 10052
rect 19292 7756 19348 7812
rect 19292 7420 19348 7476
rect 19964 10780 20020 10836
rect 20076 10892 20132 10948
rect 19964 8316 20020 8372
rect 19180 6690 19236 6692
rect 19180 6638 19182 6690
rect 19182 6638 19234 6690
rect 19234 6638 19236 6690
rect 19180 6636 19236 6638
rect 19852 7420 19908 7476
rect 19516 6524 19572 6580
rect 19852 6636 19908 6692
rect 18396 4956 18452 5012
rect 18284 4396 18340 4452
rect 18172 3554 18228 3556
rect 18172 3502 18174 3554
rect 18174 3502 18226 3554
rect 18226 3502 18228 3554
rect 18172 3500 18228 3502
rect 17948 2828 18004 2884
rect 18060 2604 18116 2660
rect 18396 4284 18452 4340
rect 18956 6076 19012 6132
rect 18508 3500 18564 3556
rect 18620 5180 18676 5236
rect 20076 8092 20132 8148
rect 20188 9996 20244 10052
rect 20188 7308 20244 7364
rect 20076 7196 20132 7252
rect 20188 6636 20244 6692
rect 18956 4732 19012 4788
rect 18508 3276 18564 3332
rect 18060 2044 18116 2100
rect 18284 2098 18340 2100
rect 18284 2046 18286 2098
rect 18286 2046 18338 2098
rect 18338 2046 18340 2098
rect 18284 2044 18340 2046
rect 17948 1986 18004 1988
rect 17948 1934 17950 1986
rect 17950 1934 18002 1986
rect 18002 1934 18004 1986
rect 17948 1932 18004 1934
rect 18060 1708 18116 1764
rect 18172 1596 18228 1652
rect 19628 5516 19684 5572
rect 19180 5068 19236 5124
rect 19740 5122 19796 5124
rect 19740 5070 19742 5122
rect 19742 5070 19794 5122
rect 19794 5070 19796 5122
rect 19740 5068 19796 5070
rect 18956 4172 19012 4228
rect 18732 3666 18788 3668
rect 18732 3614 18734 3666
rect 18734 3614 18786 3666
rect 18786 3614 18788 3666
rect 18732 3612 18788 3614
rect 18844 3388 18900 3444
rect 19628 3724 19684 3780
rect 18956 3052 19012 3108
rect 18620 2828 18676 2884
rect 19068 2716 19124 2772
rect 18620 2380 18676 2436
rect 18844 2380 18900 2436
rect 18732 1986 18788 1988
rect 18732 1934 18734 1986
rect 18734 1934 18786 1986
rect 18786 1934 18788 1986
rect 18732 1932 18788 1934
rect 19516 2770 19572 2772
rect 19516 2718 19518 2770
rect 19518 2718 19570 2770
rect 19570 2718 19572 2770
rect 19516 2716 19572 2718
rect 19292 2210 19348 2212
rect 19292 2158 19294 2210
rect 19294 2158 19346 2210
rect 19346 2158 19348 2210
rect 19292 2156 19348 2158
rect 19180 1932 19236 1988
rect 19516 1932 19572 1988
rect 19964 5516 20020 5572
rect 20972 13020 21028 13076
rect 20860 12796 20916 12852
rect 20748 11452 20804 11508
rect 20972 12012 21028 12068
rect 21756 16268 21812 16324
rect 21532 15596 21588 15652
rect 21644 16044 21700 16100
rect 21308 15484 21364 15540
rect 21756 15596 21812 15652
rect 21868 15484 21924 15540
rect 21756 14812 21812 14868
rect 21308 14530 21364 14532
rect 21308 14478 21310 14530
rect 21310 14478 21362 14530
rect 21362 14478 21364 14530
rect 21308 14476 21364 14478
rect 21420 13746 21476 13748
rect 21420 13694 21422 13746
rect 21422 13694 21474 13746
rect 21474 13694 21476 13746
rect 21420 13692 21476 13694
rect 20860 11116 20916 11172
rect 20524 8370 20580 8372
rect 20524 8318 20526 8370
rect 20526 8318 20578 8370
rect 20578 8318 20580 8370
rect 20524 8316 20580 8318
rect 20636 7756 20692 7812
rect 20636 6636 20692 6692
rect 20972 10722 21028 10724
rect 20972 10670 20974 10722
rect 20974 10670 21026 10722
rect 21026 10670 21028 10722
rect 20972 10668 21028 10670
rect 21196 10556 21252 10612
rect 21308 12908 21364 12964
rect 21532 12962 21588 12964
rect 21532 12910 21534 12962
rect 21534 12910 21586 12962
rect 21586 12910 21588 12962
rect 21532 12908 21588 12910
rect 21308 11676 21364 11732
rect 21308 11228 21364 11284
rect 20972 8258 21028 8260
rect 20972 8206 20974 8258
rect 20974 8206 21026 8258
rect 21026 8206 21028 8258
rect 20972 8204 21028 8206
rect 21420 12796 21476 12852
rect 21420 10668 21476 10724
rect 21532 12460 21588 12516
rect 21644 12124 21700 12180
rect 21868 13692 21924 13748
rect 22316 23324 22372 23380
rect 22540 23100 22596 23156
rect 22764 24892 22820 24948
rect 22764 24668 22820 24724
rect 22764 23548 22820 23604
rect 22764 22652 22820 22708
rect 22204 21756 22260 21812
rect 23100 36988 23156 37044
rect 22988 36316 23044 36372
rect 22988 35532 23044 35588
rect 23100 35420 23156 35476
rect 23100 30994 23156 30996
rect 23100 30942 23102 30994
rect 23102 30942 23154 30994
rect 23154 30942 23156 30994
rect 23100 30940 23156 30942
rect 22988 27356 23044 27412
rect 22988 27132 23044 27188
rect 23100 29260 23156 29316
rect 22988 26124 23044 26180
rect 23100 24332 23156 24388
rect 22988 23660 23044 23716
rect 23100 23154 23156 23156
rect 23100 23102 23102 23154
rect 23102 23102 23154 23154
rect 23154 23102 23156 23154
rect 23100 23100 23156 23102
rect 22988 22370 23044 22372
rect 22988 22318 22990 22370
rect 22990 22318 23042 22370
rect 23042 22318 23044 22370
rect 22988 22316 23044 22318
rect 23660 49084 23716 49140
rect 23548 48412 23604 48468
rect 23548 46508 23604 46564
rect 23772 48748 23828 48804
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 24012 48580 24068 48582
rect 24220 48636 24276 48692
rect 24220 47740 24276 47796
rect 24332 48130 24388 48132
rect 24332 48078 24334 48130
rect 24334 48078 24386 48130
rect 24386 48078 24388 48130
rect 24332 48076 24388 48078
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 24444 47180 24500 47236
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 24220 46956 24276 47012
rect 24444 46620 24500 46676
rect 25004 50092 25060 50148
rect 25788 53618 25844 53620
rect 25788 53566 25790 53618
rect 25790 53566 25842 53618
rect 25842 53566 25844 53618
rect 25788 53564 25844 53566
rect 26572 54460 26628 54516
rect 26348 53900 26404 53956
rect 26460 54348 26516 54404
rect 26348 53730 26404 53732
rect 26348 53678 26350 53730
rect 26350 53678 26402 53730
rect 26402 53678 26404 53730
rect 26348 53676 26404 53678
rect 26236 53228 26292 53284
rect 26124 53116 26180 53172
rect 25900 52892 25956 52948
rect 26908 55298 26964 55300
rect 26908 55246 26910 55298
rect 26910 55246 26962 55298
rect 26962 55246 26964 55298
rect 26908 55244 26964 55246
rect 27468 55804 27524 55860
rect 27132 54796 27188 54852
rect 27244 54290 27300 54292
rect 27244 54238 27246 54290
rect 27246 54238 27298 54290
rect 27298 54238 27300 54290
rect 27244 54236 27300 54238
rect 26572 53116 26628 53172
rect 26348 52780 26404 52836
rect 25676 52444 25732 52500
rect 25116 49250 25172 49252
rect 25116 49198 25118 49250
rect 25118 49198 25170 49250
rect 25170 49198 25172 49250
rect 25116 49196 25172 49198
rect 25004 49084 25060 49140
rect 25004 47458 25060 47460
rect 25004 47406 25006 47458
rect 25006 47406 25058 47458
rect 25058 47406 25060 47458
rect 25004 47404 25060 47406
rect 24668 46396 24724 46452
rect 23884 46284 23940 46340
rect 24464 46282 24520 46284
rect 23660 46172 23716 46228
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 25004 46284 25060 46340
rect 23884 45890 23940 45892
rect 23884 45838 23886 45890
rect 23886 45838 23938 45890
rect 23938 45838 23940 45890
rect 23884 45836 23940 45838
rect 23660 45500 23716 45556
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 24332 45388 24388 45444
rect 23772 45164 23828 45220
rect 24668 45106 24724 45108
rect 24668 45054 24670 45106
rect 24670 45054 24722 45106
rect 24722 45054 24724 45106
rect 24668 45052 24724 45054
rect 24444 44940 24500 44996
rect 23660 44716 23716 44772
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 23996 44044 24052 44100
rect 24220 44044 24276 44100
rect 23436 43036 23492 43092
rect 23548 43932 23604 43988
rect 23324 41916 23380 41972
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 24220 43820 24276 43876
rect 24780 44268 24836 44324
rect 24780 44044 24836 44100
rect 24892 43932 24948 43988
rect 25004 43538 25060 43540
rect 25004 43486 25006 43538
rect 25006 43486 25058 43538
rect 25058 43486 25060 43538
rect 25004 43484 25060 43486
rect 23772 43036 23828 43092
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 24332 43372 24388 43428
rect 24332 43036 24388 43092
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 25340 50652 25396 50708
rect 25564 51212 25620 51268
rect 25564 50204 25620 50260
rect 25452 48802 25508 48804
rect 25452 48750 25454 48802
rect 25454 48750 25506 48802
rect 25506 48750 25508 48802
rect 25452 48748 25508 48750
rect 25900 52386 25956 52388
rect 25900 52334 25902 52386
rect 25902 52334 25954 52386
rect 25954 52334 25956 52386
rect 25900 52332 25956 52334
rect 26236 52108 26292 52164
rect 25900 50876 25956 50932
rect 25900 50428 25956 50484
rect 25564 48412 25620 48468
rect 25676 48972 25732 49028
rect 25564 48018 25620 48020
rect 25564 47966 25566 48018
rect 25566 47966 25618 48018
rect 25618 47966 25620 48018
rect 25564 47964 25620 47966
rect 25340 47570 25396 47572
rect 25340 47518 25342 47570
rect 25342 47518 25394 47570
rect 25394 47518 25396 47570
rect 25340 47516 25396 47518
rect 25340 46172 25396 46228
rect 25340 45724 25396 45780
rect 25900 48972 25956 49028
rect 25452 45164 25508 45220
rect 25228 44882 25284 44884
rect 25228 44830 25230 44882
rect 25230 44830 25282 44882
rect 25282 44830 25284 44882
rect 25228 44828 25284 44830
rect 25228 44604 25284 44660
rect 24220 42028 24276 42084
rect 25228 42364 25284 42420
rect 24780 41692 24836 41748
rect 25004 41916 25060 41972
rect 23548 41580 23604 41636
rect 24220 41580 24276 41636
rect 23884 41468 23940 41524
rect 23660 41186 23716 41188
rect 23660 41134 23662 41186
rect 23662 41134 23714 41186
rect 23714 41134 23716 41186
rect 23660 41132 23716 41134
rect 23436 40402 23492 40404
rect 23436 40350 23438 40402
rect 23438 40350 23490 40402
rect 23490 40350 23492 40402
rect 23436 40348 23492 40350
rect 23548 40236 23604 40292
rect 23436 40012 23492 40068
rect 23324 38668 23380 38724
rect 23324 38108 23380 38164
rect 23324 35980 23380 36036
rect 23324 35532 23380 35588
rect 23548 39116 23604 39172
rect 23548 38946 23604 38948
rect 23548 38894 23550 38946
rect 23550 38894 23602 38946
rect 23602 38894 23604 38946
rect 23548 38892 23604 38894
rect 23548 38050 23604 38052
rect 23548 37998 23550 38050
rect 23550 37998 23602 38050
rect 23602 37998 23604 38050
rect 23548 37996 23604 37998
rect 23436 33964 23492 34020
rect 23884 40908 23940 40964
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 23772 40460 23828 40516
rect 23772 39452 23828 39508
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 24444 40796 24500 40852
rect 25228 41132 25284 41188
rect 25676 46284 25732 46340
rect 25564 44268 25620 44324
rect 25900 44156 25956 44212
rect 25676 43426 25732 43428
rect 25676 43374 25678 43426
rect 25678 43374 25730 43426
rect 25730 43374 25732 43426
rect 25676 43372 25732 43374
rect 25900 41746 25956 41748
rect 25900 41694 25902 41746
rect 25902 41694 25954 41746
rect 25954 41694 25956 41746
rect 25900 41692 25956 41694
rect 25116 40348 25172 40404
rect 24220 40124 24276 40180
rect 24892 40236 24948 40292
rect 24464 40010 24520 40012
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 24108 39452 24164 39508
rect 24332 39564 24388 39620
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 24012 39172 24068 39174
rect 23772 38780 23828 38836
rect 23996 38780 24052 38836
rect 23996 38556 24052 38612
rect 23772 38444 23828 38500
rect 23884 38162 23940 38164
rect 23884 38110 23886 38162
rect 23886 38110 23938 38162
rect 23938 38110 23940 38162
rect 23884 38108 23940 38110
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24332 37660 24388 37716
rect 24012 37604 24068 37606
rect 24220 37548 24276 37604
rect 24220 37154 24276 37156
rect 24220 37102 24222 37154
rect 24222 37102 24274 37154
rect 24274 37102 24276 37154
rect 24220 37100 24276 37102
rect 23772 36764 23828 36820
rect 24556 37884 24612 37940
rect 25228 39676 25284 39732
rect 25340 40908 25396 40964
rect 25116 38892 25172 38948
rect 24892 37548 24948 37604
rect 24556 37100 24612 37156
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 23548 36428 23604 36484
rect 25116 37212 25172 37268
rect 24892 36428 24948 36484
rect 23324 30156 23380 30212
rect 23436 29484 23492 29540
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 23324 25116 23380 25172
rect 23436 26124 23492 26180
rect 23324 23212 23380 23268
rect 25228 38108 25284 38164
rect 23660 36204 23716 36260
rect 24892 36204 24948 36260
rect 25228 36092 25284 36148
rect 23804 36090 23860 36092
rect 23660 35980 23716 36036
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 24892 35980 24948 36036
rect 23772 35532 23828 35588
rect 23772 35196 23828 35252
rect 23772 34860 23828 34916
rect 24444 35474 24500 35476
rect 24444 35422 24446 35474
rect 24446 35422 24498 35474
rect 24498 35422 24500 35474
rect 24444 35420 24500 35422
rect 24668 35420 24724 35476
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 23884 34636 23940 34692
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 24556 34524 24612 34580
rect 23884 33852 23940 33908
rect 24108 33906 24164 33908
rect 24108 33854 24110 33906
rect 24110 33854 24162 33906
rect 24162 33854 24164 33906
rect 24108 33852 24164 33854
rect 25116 35308 25172 35364
rect 25116 34748 25172 34804
rect 26124 50540 26180 50596
rect 26348 51378 26404 51380
rect 26348 51326 26350 51378
rect 26350 51326 26402 51378
rect 26402 51326 26404 51378
rect 26348 51324 26404 51326
rect 26460 51660 26516 51716
rect 26796 53452 26852 53508
rect 27132 53788 27188 53844
rect 26908 52892 26964 52948
rect 27020 52668 27076 52724
rect 26908 52556 26964 52612
rect 26908 52332 26964 52388
rect 26796 51660 26852 51716
rect 26236 49138 26292 49140
rect 26236 49086 26238 49138
rect 26238 49086 26290 49138
rect 26290 49086 26292 49138
rect 26236 49084 26292 49086
rect 26236 46956 26292 47012
rect 26236 46284 26292 46340
rect 26460 49868 26516 49924
rect 26460 49532 26516 49588
rect 26684 49308 26740 49364
rect 26796 49196 26852 49252
rect 26684 48636 26740 48692
rect 26348 46060 26404 46116
rect 26460 48300 26516 48356
rect 26572 48130 26628 48132
rect 26572 48078 26574 48130
rect 26574 48078 26626 48130
rect 26626 48078 26628 48130
rect 26572 48076 26628 48078
rect 26684 47346 26740 47348
rect 26684 47294 26686 47346
rect 26686 47294 26738 47346
rect 26738 47294 26740 47346
rect 26684 47292 26740 47294
rect 26684 47068 26740 47124
rect 26796 46844 26852 46900
rect 26124 44492 26180 44548
rect 25676 39340 25732 39396
rect 25676 39004 25732 39060
rect 25452 38444 25508 38500
rect 25452 37324 25508 37380
rect 25676 37266 25732 37268
rect 25676 37214 25678 37266
rect 25678 37214 25730 37266
rect 25730 37214 25732 37266
rect 25676 37212 25732 37214
rect 25564 36988 25620 37044
rect 25340 34748 25396 34804
rect 25452 36876 25508 36932
rect 25564 35474 25620 35476
rect 25564 35422 25566 35474
rect 25566 35422 25618 35474
rect 25618 35422 25620 35474
rect 25564 35420 25620 35422
rect 25676 34860 25732 34916
rect 24332 33740 24388 33796
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 23884 33404 23940 33460
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 24220 32956 24276 33012
rect 23884 32060 23940 32116
rect 23884 31778 23940 31780
rect 23884 31726 23886 31778
rect 23886 31726 23938 31778
rect 23938 31726 23940 31778
rect 23884 31724 23940 31726
rect 23660 31276 23716 31332
rect 23804 31386 23860 31388
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23884 30994 23940 30996
rect 23884 30942 23886 30994
rect 23886 30942 23938 30994
rect 23938 30942 23940 30994
rect 23884 30940 23940 30942
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 23660 29036 23716 29092
rect 23660 28700 23716 28756
rect 23996 29538 24052 29540
rect 23996 29486 23998 29538
rect 23998 29486 24050 29538
rect 24050 29486 24052 29538
rect 23996 29484 24052 29486
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24556 31948 24612 32004
rect 24668 31666 24724 31668
rect 24668 31614 24670 31666
rect 24670 31614 24722 31666
rect 24722 31614 24724 31666
rect 24668 31612 24724 31614
rect 24556 31164 24612 31220
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 24332 30156 24388 30212
rect 24444 29314 24500 29316
rect 24444 29262 24446 29314
rect 24446 29262 24498 29314
rect 24498 29262 24500 29314
rect 24444 29260 24500 29262
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 24332 28476 24388 28532
rect 25116 33516 25172 33572
rect 25116 33292 25172 33348
rect 25452 33068 25508 33124
rect 25004 32956 25060 33012
rect 25340 32956 25396 33012
rect 25004 32172 25060 32228
rect 25228 31890 25284 31892
rect 25228 31838 25230 31890
rect 25230 31838 25282 31890
rect 25282 31838 25284 31890
rect 25228 31836 25284 31838
rect 25228 30994 25284 30996
rect 25228 30942 25230 30994
rect 25230 30942 25282 30994
rect 25282 30942 25284 30994
rect 25228 30940 25284 30942
rect 25116 30882 25172 30884
rect 25116 30830 25118 30882
rect 25118 30830 25170 30882
rect 25170 30830 25172 30882
rect 25116 30828 25172 30830
rect 25116 29036 25172 29092
rect 25116 28700 25172 28756
rect 24892 28476 24948 28532
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24220 28252 24276 28308
rect 25676 31948 25732 32004
rect 25564 30828 25620 30884
rect 25676 30268 25732 30324
rect 25452 30156 25508 30212
rect 25676 30098 25732 30100
rect 25676 30046 25678 30098
rect 25678 30046 25730 30098
rect 25730 30046 25732 30098
rect 25676 30044 25732 30046
rect 24012 28196 24068 28198
rect 24780 28028 24836 28084
rect 24220 27858 24276 27860
rect 24220 27806 24222 27858
rect 24222 27806 24274 27858
rect 24274 27806 24276 27858
rect 24220 27804 24276 27806
rect 24780 27692 24836 27748
rect 25676 28812 25732 28868
rect 23884 27356 23940 27412
rect 24220 27468 24276 27524
rect 23660 26908 23716 26964
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 24464 27466 24520 27468
rect 24332 27356 24388 27412
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24892 27468 24948 27524
rect 25116 27244 25172 27300
rect 24220 26572 24276 26628
rect 25004 27132 25060 27188
rect 25116 26796 25172 26852
rect 25564 27020 25620 27076
rect 24220 26124 24276 26180
rect 24444 26124 24500 26180
rect 25004 26178 25060 26180
rect 25004 26126 25006 26178
rect 25006 26126 25058 26178
rect 25058 26126 25060 26178
rect 25004 26124 25060 26126
rect 24332 25788 24388 25844
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 24780 25730 24836 25732
rect 24780 25678 24782 25730
rect 24782 25678 24834 25730
rect 24834 25678 24836 25730
rect 24780 25676 24836 25678
rect 23548 25004 23604 25060
rect 23548 24220 23604 24276
rect 23548 23042 23604 23044
rect 23548 22990 23550 23042
rect 23550 22990 23602 23042
rect 23602 22990 23604 23042
rect 23548 22988 23604 22990
rect 22316 20690 22372 20692
rect 22316 20638 22318 20690
rect 22318 20638 22370 20690
rect 22370 20638 22372 20690
rect 22316 20636 22372 20638
rect 22204 20524 22260 20580
rect 22652 20524 22708 20580
rect 22428 19964 22484 20020
rect 22204 16604 22260 16660
rect 22316 19852 22372 19908
rect 22092 14364 22148 14420
rect 22092 13468 22148 13524
rect 21980 12066 22036 12068
rect 21980 12014 21982 12066
rect 21982 12014 22034 12066
rect 22034 12014 22036 12066
rect 21980 12012 22036 12014
rect 21756 11116 21812 11172
rect 21980 11788 22036 11844
rect 21868 10892 21924 10948
rect 21868 9996 21924 10052
rect 21532 9884 21588 9940
rect 21756 9884 21812 9940
rect 20972 7474 21028 7476
rect 20972 7422 20974 7474
rect 20974 7422 21026 7474
rect 21026 7422 21028 7474
rect 20972 7420 21028 7422
rect 20860 7084 20916 7140
rect 21644 7250 21700 7252
rect 21644 7198 21646 7250
rect 21646 7198 21698 7250
rect 21698 7198 21700 7250
rect 21644 7196 21700 7198
rect 20412 5964 20468 6020
rect 20972 5516 21028 5572
rect 20860 5404 20916 5460
rect 20300 5068 20356 5124
rect 20524 5122 20580 5124
rect 20524 5070 20526 5122
rect 20526 5070 20578 5122
rect 20578 5070 20580 5122
rect 20524 5068 20580 5070
rect 19964 4338 20020 4340
rect 19964 4286 19966 4338
rect 19966 4286 20018 4338
rect 20018 4286 20020 4338
rect 19964 4284 20020 4286
rect 20748 4620 20804 4676
rect 20636 4338 20692 4340
rect 20636 4286 20638 4338
rect 20638 4286 20690 4338
rect 20690 4286 20692 4338
rect 20636 4284 20692 4286
rect 20188 4060 20244 4116
rect 19852 3666 19908 3668
rect 19852 3614 19854 3666
rect 19854 3614 19906 3666
rect 19906 3614 19908 3666
rect 19852 3612 19908 3614
rect 19964 2658 20020 2660
rect 19964 2606 19966 2658
rect 19966 2606 20018 2658
rect 20018 2606 20020 2658
rect 19964 2604 20020 2606
rect 20076 2546 20132 2548
rect 20076 2494 20078 2546
rect 20078 2494 20130 2546
rect 20130 2494 20132 2546
rect 20076 2492 20132 2494
rect 19852 2380 19908 2436
rect 19852 1986 19908 1988
rect 19852 1934 19854 1986
rect 19854 1934 19906 1986
rect 19906 1934 19908 1986
rect 19852 1932 19908 1934
rect 19516 1372 19572 1428
rect 18732 1148 18788 1204
rect 18508 924 18564 980
rect 19068 364 19124 420
rect 20972 5180 21028 5236
rect 21084 4732 21140 4788
rect 22764 18060 22820 18116
rect 22316 16044 22372 16100
rect 22428 16828 22484 16884
rect 23100 21308 23156 21364
rect 23100 20860 23156 20916
rect 23212 20636 23268 20692
rect 23100 19906 23156 19908
rect 23100 19854 23102 19906
rect 23102 19854 23154 19906
rect 23154 19854 23156 19906
rect 23100 19852 23156 19854
rect 23436 21980 23492 22036
rect 23548 21474 23604 21476
rect 23548 21422 23550 21474
rect 23550 21422 23602 21474
rect 23602 21422 23604 21474
rect 23548 21420 23604 21422
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 24444 25116 24500 25172
rect 24444 24668 24500 24724
rect 24556 24556 24612 24612
rect 24464 24330 24520 24332
rect 24220 24220 24276 24276
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 23884 23938 23940 23940
rect 23884 23886 23886 23938
rect 23886 23886 23938 23938
rect 23938 23886 23940 23938
rect 23884 23884 23940 23886
rect 23804 23546 23860 23548
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 24556 23996 24612 24052
rect 24556 23772 24612 23828
rect 24220 23436 24276 23492
rect 23884 23154 23940 23156
rect 23884 23102 23886 23154
rect 23886 23102 23938 23154
rect 23938 23102 23940 23154
rect 23884 23100 23940 23102
rect 24220 23100 24276 23156
rect 24220 22876 24276 22932
rect 25004 25340 25060 25396
rect 25228 25506 25284 25508
rect 25228 25454 25230 25506
rect 25230 25454 25282 25506
rect 25282 25454 25284 25506
rect 25228 25452 25284 25454
rect 25116 23324 25172 23380
rect 25228 25116 25284 25172
rect 25004 23212 25060 23268
rect 25340 24668 25396 24724
rect 25564 23548 25620 23604
rect 25676 23660 25732 23716
rect 24892 22988 24948 23044
rect 24780 22876 24836 22932
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 24332 22540 24388 22596
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 24556 21980 24612 22036
rect 25228 22876 25284 22932
rect 24556 21532 24612 21588
rect 24780 21586 24836 21588
rect 24780 21534 24782 21586
rect 24782 21534 24834 21586
rect 24834 21534 24836 21586
rect 24780 21532 24836 21534
rect 24892 21420 24948 21476
rect 24332 21196 24388 21252
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 23660 20748 23716 20804
rect 23884 20802 23940 20804
rect 23884 20750 23886 20802
rect 23886 20750 23938 20802
rect 23938 20750 23940 20802
rect 23884 20748 23940 20750
rect 24556 20690 24612 20692
rect 24556 20638 24558 20690
rect 24558 20638 24610 20690
rect 24610 20638 24612 20690
rect 24556 20636 24612 20638
rect 23436 20300 23492 20356
rect 23436 20018 23492 20020
rect 23436 19966 23438 20018
rect 23438 19966 23490 20018
rect 23490 19966 23492 20018
rect 23436 19964 23492 19966
rect 23100 18284 23156 18340
rect 22988 16828 23044 16884
rect 23324 16882 23380 16884
rect 23324 16830 23326 16882
rect 23326 16830 23378 16882
rect 23378 16830 23380 16882
rect 23324 16828 23380 16830
rect 23324 16492 23380 16548
rect 23548 17948 23604 18004
rect 23100 16156 23156 16212
rect 22428 15538 22484 15540
rect 22428 15486 22430 15538
rect 22430 15486 22482 15538
rect 22482 15486 22484 15538
rect 22428 15484 22484 15486
rect 22204 11676 22260 11732
rect 22316 14476 22372 14532
rect 22204 11452 22260 11508
rect 22204 10892 22260 10948
rect 22204 10668 22260 10724
rect 22316 10444 22372 10500
rect 22428 12908 22484 12964
rect 22316 9042 22372 9044
rect 22316 8990 22318 9042
rect 22318 8990 22370 9042
rect 22370 8990 22372 9042
rect 22316 8988 22372 8990
rect 22316 8204 22372 8260
rect 21756 6524 21812 6580
rect 21980 6748 22036 6804
rect 21420 5740 21476 5796
rect 21420 5122 21476 5124
rect 21420 5070 21422 5122
rect 21422 5070 21474 5122
rect 21474 5070 21476 5122
rect 21420 5068 21476 5070
rect 21868 5852 21924 5908
rect 21756 5516 21812 5572
rect 21532 4620 21588 4676
rect 21644 5404 21700 5460
rect 21532 4396 21588 4452
rect 20860 3388 20916 3444
rect 20300 2828 20356 2884
rect 21084 3442 21140 3444
rect 21084 3390 21086 3442
rect 21086 3390 21138 3442
rect 21138 3390 21140 3442
rect 21084 3388 21140 3390
rect 21196 2770 21252 2772
rect 21196 2718 21198 2770
rect 21198 2718 21250 2770
rect 21250 2718 21252 2770
rect 21196 2716 21252 2718
rect 21196 2492 21252 2548
rect 20748 2380 20804 2436
rect 20412 1596 20468 1652
rect 20860 1484 20916 1540
rect 20636 476 20692 532
rect 21756 4732 21812 4788
rect 21644 3778 21700 3780
rect 21644 3726 21646 3778
rect 21646 3726 21698 3778
rect 21698 3726 21700 3778
rect 21644 3724 21700 3726
rect 21756 3666 21812 3668
rect 21756 3614 21758 3666
rect 21758 3614 21810 3666
rect 21810 3614 21812 3666
rect 21756 3612 21812 3614
rect 22092 4338 22148 4340
rect 22092 4286 22094 4338
rect 22094 4286 22146 4338
rect 22146 4286 22148 4338
rect 22092 4284 22148 4286
rect 22652 12908 22708 12964
rect 22652 12460 22708 12516
rect 22540 12012 22596 12068
rect 22764 11788 22820 11844
rect 22876 15708 22932 15764
rect 23100 15708 23156 15764
rect 22988 15596 23044 15652
rect 23212 15148 23268 15204
rect 23100 13580 23156 13636
rect 22988 13132 23044 13188
rect 23212 13074 23268 13076
rect 23212 13022 23214 13074
rect 23214 13022 23266 13074
rect 23266 13022 23268 13074
rect 23212 13020 23268 13022
rect 23100 12178 23156 12180
rect 23100 12126 23102 12178
rect 23102 12126 23154 12178
rect 23154 12126 23156 12178
rect 23100 12124 23156 12126
rect 23548 16156 23604 16212
rect 23436 15820 23492 15876
rect 23436 13020 23492 13076
rect 23548 15708 23604 15764
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 24780 20636 24836 20692
rect 24892 20524 24948 20580
rect 24556 20412 24612 20468
rect 24220 20300 24276 20356
rect 24220 19852 24276 19908
rect 24108 19516 24164 19572
rect 24220 19628 24276 19684
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24220 18844 24276 18900
rect 24332 19180 24388 19236
rect 24012 18788 24068 18790
rect 24220 17388 24276 17444
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 23772 17052 23828 17108
rect 24108 16882 24164 16884
rect 24108 16830 24110 16882
rect 24110 16830 24162 16882
rect 24162 16830 24164 16882
rect 24108 16828 24164 16830
rect 24108 16380 24164 16436
rect 24108 15932 24164 15988
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 23660 13244 23716 13300
rect 23772 13132 23828 13188
rect 25116 20524 25172 20580
rect 25116 19852 25172 19908
rect 24892 18396 24948 18452
rect 25004 18732 25060 18788
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 24892 18060 24948 18116
rect 24668 16828 24724 16884
rect 24780 17276 24836 17332
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 24892 16156 24948 16212
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 25116 17612 25172 17668
rect 26124 43932 26180 43988
rect 26348 43538 26404 43540
rect 26348 43486 26350 43538
rect 26350 43486 26402 43538
rect 26402 43486 26404 43538
rect 26348 43484 26404 43486
rect 26460 43036 26516 43092
rect 26348 42700 26404 42756
rect 27020 45052 27076 45108
rect 26908 43708 26964 43764
rect 26460 42252 26516 42308
rect 26236 41580 26292 41636
rect 26348 41804 26404 41860
rect 26236 41132 26292 41188
rect 26236 40908 26292 40964
rect 26236 40402 26292 40404
rect 26236 40350 26238 40402
rect 26238 40350 26290 40402
rect 26290 40350 26292 40402
rect 26236 40348 26292 40350
rect 26572 41244 26628 41300
rect 26236 39676 26292 39732
rect 26236 39116 26292 39172
rect 26236 38834 26292 38836
rect 26236 38782 26238 38834
rect 26238 38782 26290 38834
rect 26290 38782 26292 38834
rect 26236 38780 26292 38782
rect 26012 37548 26068 37604
rect 26236 38332 26292 38388
rect 26012 37100 26068 37156
rect 26124 35698 26180 35700
rect 26124 35646 26126 35698
rect 26126 35646 26178 35698
rect 26178 35646 26180 35698
rect 26124 35644 26180 35646
rect 26012 35532 26068 35588
rect 26124 33292 26180 33348
rect 26012 31612 26068 31668
rect 26460 39506 26516 39508
rect 26460 39454 26462 39506
rect 26462 39454 26514 39506
rect 26514 39454 26516 39506
rect 26460 39452 26516 39454
rect 26684 40178 26740 40180
rect 26684 40126 26686 40178
rect 26686 40126 26738 40178
rect 26738 40126 26740 40178
rect 26684 40124 26740 40126
rect 26796 39900 26852 39956
rect 26684 39452 26740 39508
rect 26460 39116 26516 39172
rect 26684 39116 26740 39172
rect 26460 37100 26516 37156
rect 26796 36482 26852 36484
rect 26796 36430 26798 36482
rect 26798 36430 26850 36482
rect 26850 36430 26852 36482
rect 26796 36428 26852 36430
rect 26908 37660 26964 37716
rect 26684 36092 26740 36148
rect 26684 34188 26740 34244
rect 26796 34076 26852 34132
rect 26236 32060 26292 32116
rect 26124 31388 26180 31444
rect 26124 31164 26180 31220
rect 26572 32060 26628 32116
rect 26012 28812 26068 28868
rect 26012 28530 26068 28532
rect 26012 28478 26014 28530
rect 26014 28478 26066 28530
rect 26066 28478 26068 28530
rect 26012 28476 26068 28478
rect 25900 25676 25956 25732
rect 25900 23892 25902 23940
rect 25902 23892 25954 23940
rect 25954 23892 25956 23940
rect 25900 23884 25956 23892
rect 25788 22652 25844 22708
rect 26236 29538 26292 29540
rect 26236 29486 26238 29538
rect 26238 29486 26290 29538
rect 26290 29486 26292 29538
rect 26236 29484 26292 29486
rect 27804 56252 27860 56308
rect 27580 55468 27636 55524
rect 27692 55580 27748 55636
rect 27580 54460 27636 54516
rect 27468 54236 27524 54292
rect 27468 53788 27524 53844
rect 27356 53452 27412 53508
rect 27356 53058 27412 53060
rect 27356 53006 27358 53058
rect 27358 53006 27410 53058
rect 27410 53006 27412 53058
rect 27356 53004 27412 53006
rect 27916 55858 27972 55860
rect 27916 55806 27918 55858
rect 27918 55806 27970 55858
rect 27970 55806 27972 55858
rect 27916 55804 27972 55806
rect 28252 56588 28308 56644
rect 28028 55468 28084 55524
rect 28140 56140 28196 56196
rect 28588 54684 28644 54740
rect 29260 55580 29316 55636
rect 28812 55132 28868 55188
rect 28700 54572 28756 54628
rect 27916 54290 27972 54292
rect 27916 54238 27918 54290
rect 27918 54238 27970 54290
rect 27970 54238 27972 54290
rect 27916 54236 27972 54238
rect 27804 54012 27860 54068
rect 27804 53730 27860 53732
rect 27804 53678 27806 53730
rect 27806 53678 27858 53730
rect 27858 53678 27860 53730
rect 27804 53676 27860 53678
rect 27692 53564 27748 53620
rect 27580 52780 27636 52836
rect 27916 53228 27972 53284
rect 27244 51884 27300 51940
rect 27356 52556 27412 52612
rect 27804 52444 27860 52500
rect 27692 51436 27748 51492
rect 27692 51100 27748 51156
rect 27804 50988 27860 51044
rect 27580 50876 27636 50932
rect 27356 48972 27412 49028
rect 27468 50652 27524 50708
rect 27692 49138 27748 49140
rect 27692 49086 27694 49138
rect 27694 49086 27746 49138
rect 27746 49086 27748 49138
rect 27692 49084 27748 49086
rect 27580 48860 27636 48916
rect 27692 48748 27748 48804
rect 27244 47964 27300 48020
rect 27804 47516 27860 47572
rect 27356 47404 27412 47460
rect 27580 47458 27636 47460
rect 27580 47406 27582 47458
rect 27582 47406 27634 47458
rect 27634 47406 27636 47458
rect 27580 47404 27636 47406
rect 28028 49532 28084 49588
rect 28252 52892 28308 52948
rect 28252 49420 28308 49476
rect 28924 54460 28980 54516
rect 28476 54124 28532 54180
rect 28476 53900 28532 53956
rect 28476 53228 28532 53284
rect 28700 53340 28756 53396
rect 28588 53004 28644 53060
rect 28588 52108 28644 52164
rect 28700 52332 28756 52388
rect 29148 54908 29204 54964
rect 29148 54738 29204 54740
rect 29148 54686 29150 54738
rect 29150 54686 29202 54738
rect 29202 54686 29204 54738
rect 29148 54684 29204 54686
rect 29036 52668 29092 52724
rect 28700 51602 28756 51604
rect 28700 51550 28702 51602
rect 28702 51550 28754 51602
rect 28754 51550 28756 51602
rect 28700 51548 28756 51550
rect 28588 51436 28644 51492
rect 28588 50988 28644 51044
rect 29036 51660 29092 51716
rect 29372 55468 29428 55524
rect 29484 56140 29540 56196
rect 29596 55858 29652 55860
rect 29596 55806 29598 55858
rect 29598 55806 29650 55858
rect 29650 55806 29652 55858
rect 29596 55804 29652 55806
rect 30604 57036 30660 57092
rect 30268 56028 30324 56084
rect 30380 56476 30436 56532
rect 29932 55970 29988 55972
rect 29932 55918 29934 55970
rect 29934 55918 29986 55970
rect 29986 55918 29988 55970
rect 29932 55916 29988 55918
rect 30268 55858 30324 55860
rect 30268 55806 30270 55858
rect 30270 55806 30322 55858
rect 30322 55806 30324 55858
rect 30268 55804 30324 55806
rect 29820 55692 29876 55748
rect 29484 55356 29540 55412
rect 29820 55410 29876 55412
rect 29820 55358 29822 55410
rect 29822 55358 29874 55410
rect 29874 55358 29876 55410
rect 29820 55356 29876 55358
rect 29596 55298 29652 55300
rect 29596 55246 29598 55298
rect 29598 55246 29650 55298
rect 29650 55246 29652 55298
rect 29596 55244 29652 55246
rect 30268 54684 30324 54740
rect 29260 53676 29316 53732
rect 29372 54572 29428 54628
rect 29372 52892 29428 52948
rect 29484 52444 29540 52500
rect 29372 52108 29428 52164
rect 29148 51266 29204 51268
rect 29148 51214 29150 51266
rect 29150 51214 29202 51266
rect 29202 51214 29204 51266
rect 29148 51212 29204 51214
rect 29484 51996 29540 52052
rect 29260 50988 29316 51044
rect 29484 51100 29540 51156
rect 29372 50876 29428 50932
rect 28700 50204 28756 50260
rect 28140 48076 28196 48132
rect 28924 49980 28980 50036
rect 27468 46956 27524 47012
rect 27468 45836 27524 45892
rect 27244 44322 27300 44324
rect 27244 44270 27246 44322
rect 27246 44270 27298 44322
rect 27298 44270 27300 44322
rect 27244 44268 27300 44270
rect 28140 47628 28196 47684
rect 28252 47516 28308 47572
rect 28476 48972 28532 49028
rect 28140 46844 28196 46900
rect 28420 46844 28476 46900
rect 28700 47292 28756 47348
rect 29036 48860 29092 48916
rect 29372 48748 29428 48804
rect 29820 52892 29876 52948
rect 30156 52444 30212 52500
rect 29820 50652 29876 50708
rect 29932 52332 29988 52388
rect 29708 49868 29764 49924
rect 29820 50316 29876 50372
rect 29596 49698 29652 49700
rect 29596 49646 29598 49698
rect 29598 49646 29650 49698
rect 29650 49646 29652 49698
rect 29596 49644 29652 49646
rect 29708 48636 29764 48692
rect 29820 47516 29876 47572
rect 29708 47458 29764 47460
rect 29708 47406 29710 47458
rect 29710 47406 29762 47458
rect 29762 47406 29764 47458
rect 29708 47404 29764 47406
rect 30268 52108 30324 52164
rect 30492 56140 30548 56196
rect 30492 55410 30548 55412
rect 30492 55358 30494 55410
rect 30494 55358 30546 55410
rect 30546 55358 30548 55410
rect 30492 55356 30548 55358
rect 30940 55692 30996 55748
rect 30716 55468 30772 55524
rect 31388 56812 31444 56868
rect 30828 55244 30884 55300
rect 31164 55298 31220 55300
rect 31164 55246 31166 55298
rect 31166 55246 31218 55298
rect 31218 55246 31220 55298
rect 31164 55244 31220 55246
rect 30604 52444 30660 52500
rect 30380 50876 30436 50932
rect 30492 50764 30548 50820
rect 30044 50540 30100 50596
rect 30268 50594 30324 50596
rect 30268 50542 30270 50594
rect 30270 50542 30322 50594
rect 30322 50542 30324 50594
rect 30268 50540 30324 50542
rect 30380 49868 30436 49924
rect 30268 49810 30324 49812
rect 30268 49758 30270 49810
rect 30270 49758 30322 49810
rect 30322 49758 30324 49810
rect 30268 49756 30324 49758
rect 30604 50540 30660 50596
rect 31276 54572 31332 54628
rect 32060 57148 32116 57204
rect 31612 56252 31668 56308
rect 31724 56700 31780 56756
rect 31500 56140 31556 56196
rect 31836 56476 31892 56532
rect 31724 55858 31780 55860
rect 31724 55806 31726 55858
rect 31726 55806 31778 55858
rect 31778 55806 31780 55858
rect 31724 55804 31780 55806
rect 32508 56028 32564 56084
rect 32732 55970 32788 55972
rect 32732 55918 32734 55970
rect 32734 55918 32786 55970
rect 32786 55918 32788 55970
rect 32732 55916 32788 55918
rect 31948 53900 32004 53956
rect 31276 53788 31332 53844
rect 30828 53564 30884 53620
rect 31164 53452 31220 53508
rect 30940 52834 30996 52836
rect 30940 52782 30942 52834
rect 30942 52782 30994 52834
rect 30994 52782 30996 52834
rect 30940 52780 30996 52782
rect 30828 52108 30884 52164
rect 30828 50594 30884 50596
rect 30828 50542 30830 50594
rect 30830 50542 30882 50594
rect 30882 50542 30884 50594
rect 30828 50540 30884 50542
rect 31052 52162 31108 52164
rect 31052 52110 31054 52162
rect 31054 52110 31106 52162
rect 31106 52110 31108 52162
rect 31052 52108 31108 52110
rect 31164 51378 31220 51380
rect 31164 51326 31166 51378
rect 31166 51326 31218 51378
rect 31218 51326 31220 51378
rect 31164 51324 31220 51326
rect 31276 50092 31332 50148
rect 31500 53730 31556 53732
rect 31500 53678 31502 53730
rect 31502 53678 31554 53730
rect 31554 53678 31556 53730
rect 31500 53676 31556 53678
rect 31724 53676 31780 53732
rect 31500 53452 31556 53508
rect 31836 53116 31892 53172
rect 31500 52668 31556 52724
rect 31500 52274 31556 52276
rect 31500 52222 31502 52274
rect 31502 52222 31554 52274
rect 31554 52222 31556 52274
rect 31500 52220 31556 52222
rect 32172 53564 32228 53620
rect 32060 53170 32116 53172
rect 32060 53118 32062 53170
rect 32062 53118 32114 53170
rect 32114 53118 32116 53170
rect 32060 53116 32116 53118
rect 31612 50652 31668 50708
rect 31388 49980 31444 50036
rect 30940 49868 30996 49924
rect 30828 49250 30884 49252
rect 30828 49198 30830 49250
rect 30830 49198 30882 49250
rect 30882 49198 30884 49250
rect 30828 49196 30884 49198
rect 30492 49026 30548 49028
rect 30492 48974 30494 49026
rect 30494 48974 30546 49026
rect 30546 48974 30548 49026
rect 30492 48972 30548 48974
rect 30156 48300 30212 48356
rect 29036 46956 29092 47012
rect 28588 46508 28644 46564
rect 27692 46060 27748 46116
rect 27580 44716 27636 44772
rect 27468 43484 27524 43540
rect 27244 43372 27300 43428
rect 28028 46172 28084 46228
rect 27916 46114 27972 46116
rect 27916 46062 27918 46114
rect 27918 46062 27970 46114
rect 27970 46062 27972 46114
rect 27916 46060 27972 46062
rect 28588 45948 28644 46004
rect 28364 45890 28420 45892
rect 28364 45838 28366 45890
rect 28366 45838 28418 45890
rect 28418 45838 28420 45890
rect 28364 45836 28420 45838
rect 28700 45276 28756 45332
rect 28812 46508 28868 46564
rect 28700 45052 28756 45108
rect 27916 44604 27972 44660
rect 27804 44268 27860 44324
rect 28252 43484 28308 43540
rect 27916 43036 27972 43092
rect 27244 42028 27300 42084
rect 27692 42252 27748 42308
rect 28140 41580 28196 41636
rect 27468 40124 27524 40180
rect 27244 39618 27300 39620
rect 27244 39566 27246 39618
rect 27246 39566 27298 39618
rect 27298 39566 27300 39618
rect 27244 39564 27300 39566
rect 27132 37324 27188 37380
rect 27244 37266 27300 37268
rect 27244 37214 27246 37266
rect 27246 37214 27298 37266
rect 27298 37214 27300 37266
rect 27244 37212 27300 37214
rect 27020 37100 27076 37156
rect 27804 38610 27860 38612
rect 27804 38558 27806 38610
rect 27806 38558 27858 38610
rect 27858 38558 27860 38610
rect 27804 38556 27860 38558
rect 28028 40124 28084 40180
rect 28140 38444 28196 38500
rect 27916 37996 27972 38052
rect 28476 44322 28532 44324
rect 28476 44270 28478 44322
rect 28478 44270 28530 44322
rect 28530 44270 28532 44322
rect 28476 44268 28532 44270
rect 28700 43932 28756 43988
rect 28588 43372 28644 43428
rect 28476 42588 28532 42644
rect 28476 41580 28532 41636
rect 28700 42754 28756 42756
rect 28700 42702 28702 42754
rect 28702 42702 28754 42754
rect 28754 42702 28756 42754
rect 28700 42700 28756 42702
rect 28700 42028 28756 42084
rect 30044 47068 30100 47124
rect 29148 46508 29204 46564
rect 28812 41468 28868 41524
rect 29036 45836 29092 45892
rect 29036 45276 29092 45332
rect 28588 40124 28644 40180
rect 28700 40684 28756 40740
rect 28700 40460 28756 40516
rect 28700 39116 28756 39172
rect 27468 36428 27524 36484
rect 27244 34636 27300 34692
rect 27020 33852 27076 33908
rect 27132 33740 27188 33796
rect 27580 35196 27636 35252
rect 27580 33852 27636 33908
rect 27580 33628 27636 33684
rect 28028 34914 28084 34916
rect 28028 34862 28030 34914
rect 28030 34862 28082 34914
rect 28082 34862 28084 34914
rect 28028 34860 28084 34862
rect 27580 32844 27636 32900
rect 28924 41020 28980 41076
rect 29708 46450 29764 46452
rect 29708 46398 29710 46450
rect 29710 46398 29762 46450
rect 29762 46398 29764 46450
rect 29708 46396 29764 46398
rect 29932 46284 29988 46340
rect 29596 44828 29652 44884
rect 29148 44156 29204 44212
rect 29148 42476 29204 42532
rect 29372 43260 29428 43316
rect 29596 43260 29652 43316
rect 29484 43036 29540 43092
rect 29372 42028 29428 42084
rect 29036 39116 29092 39172
rect 28588 38780 28644 38836
rect 28476 37378 28532 37380
rect 28476 37326 28478 37378
rect 28478 37326 28530 37378
rect 28530 37326 28532 37378
rect 28476 37324 28532 37326
rect 28364 37212 28420 37268
rect 28252 33628 28308 33684
rect 27468 32396 27524 32452
rect 28140 32396 28196 32452
rect 27356 32284 27412 32340
rect 26908 31778 26964 31780
rect 26908 31726 26910 31778
rect 26910 31726 26962 31778
rect 26962 31726 26964 31778
rect 26908 31724 26964 31726
rect 26908 31164 26964 31220
rect 26796 31052 26852 31108
rect 26684 30380 26740 30436
rect 26684 29260 26740 29316
rect 26460 28866 26516 28868
rect 26460 28814 26462 28866
rect 26462 28814 26514 28866
rect 26514 28814 26516 28866
rect 26460 28812 26516 28814
rect 26124 27132 26180 27188
rect 26236 28476 26292 28532
rect 26236 28140 26292 28196
rect 26460 27916 26516 27972
rect 26348 27244 26404 27300
rect 26348 26908 26404 26964
rect 26124 25116 26180 25172
rect 26236 25340 26292 25396
rect 26124 24668 26180 24724
rect 26124 23212 26180 23268
rect 26012 22316 26068 22372
rect 26572 27186 26628 27188
rect 26572 27134 26574 27186
rect 26574 27134 26626 27186
rect 26626 27134 26628 27186
rect 26572 27132 26628 27134
rect 26572 26178 26628 26180
rect 26572 26126 26574 26178
rect 26574 26126 26626 26178
rect 26626 26126 26628 26178
rect 26572 26124 26628 26126
rect 27468 30994 27524 30996
rect 27468 30942 27470 30994
rect 27470 30942 27522 30994
rect 27522 30942 27524 30994
rect 27468 30940 27524 30942
rect 27804 30770 27860 30772
rect 27804 30718 27806 30770
rect 27806 30718 27858 30770
rect 27858 30718 27860 30770
rect 27804 30716 27860 30718
rect 27692 30604 27748 30660
rect 28028 30940 28084 30996
rect 27020 30268 27076 30324
rect 27804 30156 27860 30212
rect 27020 28028 27076 28084
rect 27244 30044 27300 30100
rect 26908 27468 26964 27524
rect 26908 27074 26964 27076
rect 26908 27022 26910 27074
rect 26910 27022 26962 27074
rect 26962 27022 26964 27074
rect 26908 27020 26964 27022
rect 27132 27468 27188 27524
rect 26684 25452 26740 25508
rect 26796 25676 26852 25732
rect 26460 24220 26516 24276
rect 26684 24498 26740 24500
rect 26684 24446 26686 24498
rect 26686 24446 26738 24498
rect 26738 24446 26740 24498
rect 26684 24444 26740 24446
rect 26348 23938 26404 23940
rect 26348 23886 26350 23938
rect 26350 23886 26402 23938
rect 26402 23886 26404 23938
rect 26348 23884 26404 23886
rect 25452 21756 25508 21812
rect 25340 21420 25396 21476
rect 25676 21308 25732 21364
rect 25564 21196 25620 21252
rect 25340 20860 25396 20916
rect 25452 19964 25508 20020
rect 25564 20076 25620 20132
rect 25340 19852 25396 19908
rect 25340 19628 25396 19684
rect 25564 19068 25620 19124
rect 25452 18508 25508 18564
rect 26124 21420 26180 21476
rect 26124 20802 26180 20804
rect 26124 20750 26126 20802
rect 26126 20750 26178 20802
rect 26178 20750 26180 20802
rect 26124 20748 26180 20750
rect 25788 20300 25844 20356
rect 26684 23436 26740 23492
rect 26684 22988 26740 23044
rect 26460 21756 26516 21812
rect 26796 21980 26852 22036
rect 26684 21084 26740 21140
rect 26236 20018 26292 20020
rect 26236 19966 26238 20018
rect 26238 19966 26290 20018
rect 26290 19966 26292 20018
rect 26236 19964 26292 19966
rect 26236 19740 26292 19796
rect 26348 19292 26404 19348
rect 26684 20636 26740 20692
rect 26572 19852 26628 19908
rect 26236 19180 26292 19236
rect 26460 19234 26516 19236
rect 26460 19182 26462 19234
rect 26462 19182 26514 19234
rect 26514 19182 26516 19234
rect 26460 19180 26516 19182
rect 26348 18732 26404 18788
rect 26236 18450 26292 18452
rect 26236 18398 26238 18450
rect 26238 18398 26290 18450
rect 26290 18398 26292 18450
rect 26236 18396 26292 18398
rect 26124 18284 26180 18340
rect 25228 16882 25284 16884
rect 25228 16830 25230 16882
rect 25230 16830 25282 16882
rect 25282 16830 25284 16882
rect 25228 16828 25284 16830
rect 25116 15820 25172 15876
rect 24332 14364 24388 14420
rect 25116 14476 25172 14532
rect 24892 14028 24948 14084
rect 24892 13692 24948 13748
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24220 12572 24276 12628
rect 24444 12572 24500 12628
rect 24012 12516 24068 12518
rect 23324 12012 23380 12068
rect 22876 11564 22932 11620
rect 23100 11900 23156 11956
rect 22540 10892 22596 10948
rect 22540 10444 22596 10500
rect 22988 10498 23044 10500
rect 22988 10446 22990 10498
rect 22990 10446 23042 10498
rect 23042 10446 23044 10498
rect 22988 10444 23044 10446
rect 22988 10220 23044 10276
rect 22764 10050 22820 10052
rect 22764 9998 22766 10050
rect 22766 9998 22818 10050
rect 22818 9998 22820 10050
rect 22764 9996 22820 9998
rect 22764 8092 22820 8148
rect 22876 6972 22932 7028
rect 22316 5068 22372 5124
rect 22876 5740 22932 5796
rect 22764 5122 22820 5124
rect 22764 5070 22766 5122
rect 22766 5070 22818 5122
rect 22818 5070 22820 5122
rect 22764 5068 22820 5070
rect 21532 3276 21588 3332
rect 21420 2716 21476 2772
rect 21308 2268 21364 2324
rect 21420 2380 21476 2436
rect 21420 1708 21476 1764
rect 21980 1708 22036 1764
rect 22204 3276 22260 3332
rect 22652 4114 22708 4116
rect 22652 4062 22654 4114
rect 22654 4062 22706 4114
rect 22706 4062 22708 4114
rect 22652 4060 22708 4062
rect 22764 3948 22820 4004
rect 22652 3836 22708 3892
rect 23548 12066 23604 12068
rect 23548 12014 23550 12066
rect 23550 12014 23602 12066
rect 23602 12014 23604 12066
rect 23548 12012 23604 12014
rect 23436 11452 23492 11508
rect 23324 10892 23380 10948
rect 23436 10444 23492 10500
rect 23100 9212 23156 9268
rect 23436 8988 23492 9044
rect 23324 7532 23380 7588
rect 23884 12178 23940 12180
rect 23884 12126 23886 12178
rect 23886 12126 23938 12178
rect 23938 12126 23940 12178
rect 23884 12124 23940 12126
rect 23996 12012 24052 12068
rect 23772 11788 23828 11844
rect 23772 11116 23828 11172
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23884 10556 23940 10612
rect 23996 10386 24052 10388
rect 23996 10334 23998 10386
rect 23998 10334 24050 10386
rect 24050 10334 24052 10386
rect 23996 10332 24052 10334
rect 23804 9434 23860 9436
rect 23660 9324 23716 9380
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 23660 8988 23716 9044
rect 23884 8204 23940 8260
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 23548 6748 23604 6804
rect 23436 6578 23492 6580
rect 23436 6526 23438 6578
rect 23438 6526 23490 6578
rect 23490 6526 23492 6578
rect 23436 6524 23492 6526
rect 23100 6076 23156 6132
rect 22876 3164 22932 3220
rect 23996 6524 24052 6580
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 24332 11564 24388 11620
rect 24444 10610 24500 10612
rect 24444 10558 24446 10610
rect 24446 10558 24498 10610
rect 24498 10558 24500 10610
rect 24444 10556 24500 10558
rect 25004 10610 25060 10612
rect 25004 10558 25006 10610
rect 25006 10558 25058 10610
rect 25058 10558 25060 10610
rect 25004 10556 25060 10558
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24332 9660 24388 9716
rect 24332 9324 24388 9380
rect 25228 14252 25284 14308
rect 25228 13692 25284 13748
rect 25228 12460 25284 12516
rect 25228 12236 25284 12292
rect 24332 8540 24388 8596
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24332 8204 24388 8260
rect 24668 7644 24724 7700
rect 24668 7308 24724 7364
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 24332 6636 24388 6692
rect 24332 6300 24388 6356
rect 25004 8204 25060 8260
rect 24444 6188 24500 6244
rect 23660 5404 23716 5460
rect 24220 5906 24276 5908
rect 24220 5854 24222 5906
rect 24222 5854 24274 5906
rect 24274 5854 24276 5906
rect 24220 5852 24276 5854
rect 24892 6690 24948 6692
rect 24892 6638 24894 6690
rect 24894 6638 24946 6690
rect 24946 6638 24948 6690
rect 24892 6636 24948 6638
rect 24668 6018 24724 6020
rect 24668 5966 24670 6018
rect 24670 5966 24722 6018
rect 24722 5966 24724 6018
rect 24668 5964 24724 5966
rect 24556 5740 24612 5796
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24220 4620 24276 4676
rect 23660 4284 23716 4340
rect 23884 4284 23940 4340
rect 23996 4114 24052 4116
rect 23996 4062 23998 4114
rect 23998 4062 24050 4114
rect 24050 4062 24052 4114
rect 23996 4060 24052 4062
rect 23884 3948 23940 4004
rect 23548 3724 23604 3780
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 25116 6972 25172 7028
rect 25116 6748 25172 6804
rect 25228 6636 25284 6692
rect 25004 5906 25060 5908
rect 25004 5854 25006 5906
rect 25006 5854 25058 5906
rect 25058 5854 25060 5906
rect 25004 5852 25060 5854
rect 24220 3500 24276 3556
rect 23436 3164 23492 3220
rect 23548 3052 23604 3108
rect 22428 2770 22484 2772
rect 22428 2718 22430 2770
rect 22430 2718 22482 2770
rect 22482 2718 22484 2770
rect 22428 2716 22484 2718
rect 23100 2658 23156 2660
rect 23100 2606 23102 2658
rect 23102 2606 23154 2658
rect 23154 2606 23156 2658
rect 23100 2604 23156 2606
rect 22540 2044 22596 2100
rect 22652 2156 22708 2212
rect 23100 1932 23156 1988
rect 21756 1596 21812 1652
rect 21644 1372 21700 1428
rect 21308 700 21364 756
rect 21420 588 21476 644
rect 22316 1090 22372 1092
rect 22316 1038 22318 1090
rect 22318 1038 22370 1090
rect 22370 1038 22372 1090
rect 22316 1036 22372 1038
rect 22652 700 22708 756
rect 22764 364 22820 420
rect 23100 924 23156 980
rect 23436 2658 23492 2660
rect 23436 2606 23438 2658
rect 23438 2606 23490 2658
rect 23490 2606 23492 2658
rect 23436 2604 23492 2606
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 24332 3164 24388 3220
rect 23884 2716 23940 2772
rect 24108 2492 24164 2548
rect 23772 2380 23828 2436
rect 24444 2546 24500 2548
rect 24444 2494 24446 2546
rect 24446 2494 24498 2546
rect 24498 2494 24500 2546
rect 24444 2492 24500 2494
rect 23548 2268 23604 2324
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24892 2268 24948 2324
rect 23548 1596 23604 1652
rect 23324 978 23380 980
rect 23324 926 23326 978
rect 23326 926 23378 978
rect 23378 926 23380 978
rect 23324 924 23380 926
rect 23212 252 23268 308
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24332 1484 24388 1540
rect 25228 6076 25284 6132
rect 25228 5516 25284 5572
rect 25788 16882 25844 16884
rect 25788 16830 25790 16882
rect 25790 16830 25842 16882
rect 25842 16830 25844 16882
rect 25788 16828 25844 16830
rect 26236 17666 26292 17668
rect 26236 17614 26238 17666
rect 26238 17614 26290 17666
rect 26290 17614 26292 17666
rect 26236 17612 26292 17614
rect 25900 16268 25956 16324
rect 26124 16492 26180 16548
rect 26124 16268 26180 16324
rect 25676 14476 25732 14532
rect 25900 14364 25956 14420
rect 25452 13522 25508 13524
rect 25452 13470 25454 13522
rect 25454 13470 25506 13522
rect 25506 13470 25508 13522
rect 25452 13468 25508 13470
rect 25564 12460 25620 12516
rect 25452 12124 25508 12180
rect 25564 11788 25620 11844
rect 25452 11340 25508 11396
rect 25452 10668 25508 10724
rect 25900 13580 25956 13636
rect 26236 13580 26292 13636
rect 25788 13356 25844 13412
rect 26124 13468 26180 13524
rect 25788 13186 25844 13188
rect 25788 13134 25790 13186
rect 25790 13134 25842 13186
rect 25842 13134 25844 13186
rect 25788 13132 25844 13134
rect 25900 12572 25956 12628
rect 25676 10556 25732 10612
rect 25788 11116 25844 11172
rect 25788 10332 25844 10388
rect 25452 8316 25508 8372
rect 25452 8092 25508 8148
rect 25676 7980 25732 8036
rect 25452 7756 25508 7812
rect 25452 6412 25508 6468
rect 26236 12850 26292 12852
rect 26236 12798 26238 12850
rect 26238 12798 26290 12850
rect 26290 12798 26292 12850
rect 26236 12796 26292 12798
rect 26124 12460 26180 12516
rect 26012 10892 26068 10948
rect 26012 10332 26068 10388
rect 26460 17164 26516 17220
rect 26460 14028 26516 14084
rect 26684 20076 26740 20132
rect 26908 23436 26964 23492
rect 26796 18732 26852 18788
rect 26796 18172 26852 18228
rect 26684 16268 26740 16324
rect 26796 16156 26852 16212
rect 26684 15932 26740 15988
rect 26908 15932 26964 15988
rect 26348 12124 26404 12180
rect 26572 11676 26628 11732
rect 26572 11228 26628 11284
rect 26684 12124 26740 12180
rect 26796 11394 26852 11396
rect 26796 11342 26798 11394
rect 26798 11342 26850 11394
rect 26850 11342 26852 11394
rect 26796 11340 26852 11342
rect 26348 10780 26404 10836
rect 26124 8316 26180 8372
rect 26012 8258 26068 8260
rect 26012 8206 26014 8258
rect 26014 8206 26066 8258
rect 26066 8206 26068 8258
rect 26012 8204 26068 8206
rect 25900 7980 25956 8036
rect 26124 7644 26180 7700
rect 25900 6690 25956 6692
rect 25900 6638 25902 6690
rect 25902 6638 25954 6690
rect 25954 6638 25956 6690
rect 25900 6636 25956 6638
rect 25564 5516 25620 5572
rect 25116 5180 25172 5236
rect 25900 5404 25956 5460
rect 26572 10780 26628 10836
rect 26348 8316 26404 8372
rect 26460 10556 26516 10612
rect 26572 10444 26628 10500
rect 26684 8652 26740 8708
rect 26460 7084 26516 7140
rect 26236 6412 26292 6468
rect 26460 6412 26516 6468
rect 26348 5964 26404 6020
rect 26684 7644 26740 7700
rect 27020 14140 27076 14196
rect 27020 12796 27076 12852
rect 27020 11676 27076 11732
rect 27916 30098 27972 30100
rect 27916 30046 27918 30098
rect 27918 30046 27970 30098
rect 27970 30046 27972 30098
rect 27916 30044 27972 30046
rect 27916 29484 27972 29540
rect 27580 28754 27636 28756
rect 27580 28702 27582 28754
rect 27582 28702 27634 28754
rect 27634 28702 27636 28754
rect 27580 28700 27636 28702
rect 27580 28028 27636 28084
rect 28140 28028 28196 28084
rect 27916 27746 27972 27748
rect 27916 27694 27918 27746
rect 27918 27694 27970 27746
rect 27970 27694 27972 27746
rect 27916 27692 27972 27694
rect 27356 26908 27412 26964
rect 27356 24556 27412 24612
rect 27804 26290 27860 26292
rect 27804 26238 27806 26290
rect 27806 26238 27858 26290
rect 27858 26238 27860 26290
rect 27804 26236 27860 26238
rect 28028 25788 28084 25844
rect 27916 24668 27972 24724
rect 27804 24610 27860 24612
rect 27804 24558 27806 24610
rect 27806 24558 27858 24610
rect 27858 24558 27860 24610
rect 27804 24556 27860 24558
rect 27916 24444 27972 24500
rect 27692 24332 27748 24388
rect 27692 23938 27748 23940
rect 27692 23886 27694 23938
rect 27694 23886 27746 23938
rect 27746 23886 27748 23938
rect 27692 23884 27748 23886
rect 27692 22594 27748 22596
rect 27692 22542 27694 22594
rect 27694 22542 27746 22594
rect 27746 22542 27748 22594
rect 27692 22540 27748 22542
rect 27916 23884 27972 23940
rect 27804 21868 27860 21924
rect 27804 21644 27860 21700
rect 27692 21420 27748 21476
rect 27468 20300 27524 20356
rect 27244 19234 27300 19236
rect 27244 19182 27246 19234
rect 27246 19182 27298 19234
rect 27298 19182 27300 19234
rect 27244 19180 27300 19182
rect 27356 18060 27412 18116
rect 27356 17612 27412 17668
rect 27244 16492 27300 16548
rect 27244 16210 27300 16212
rect 27244 16158 27246 16210
rect 27246 16158 27298 16210
rect 27298 16158 27300 16210
rect 27244 16156 27300 16158
rect 27244 15148 27300 15204
rect 27244 14476 27300 14532
rect 27356 14140 27412 14196
rect 27244 11116 27300 11172
rect 27356 9996 27412 10052
rect 27804 20636 27860 20692
rect 27692 19516 27748 19572
rect 27916 19628 27972 19684
rect 27804 19180 27860 19236
rect 27692 18508 27748 18564
rect 28140 22482 28196 22484
rect 28140 22430 28142 22482
rect 28142 22430 28194 22482
rect 28194 22430 28196 22482
rect 28140 22428 28196 22430
rect 28700 38050 28756 38052
rect 28700 37998 28702 38050
rect 28702 37998 28754 38050
rect 28754 37998 28756 38050
rect 28700 37996 28756 37998
rect 28700 35420 28756 35476
rect 28812 35084 28868 35140
rect 29036 38050 29092 38052
rect 29036 37998 29038 38050
rect 29038 37998 29090 38050
rect 29090 37998 29092 38050
rect 29036 37996 29092 37998
rect 28924 34860 28980 34916
rect 28476 33628 28532 33684
rect 28364 31052 28420 31108
rect 28812 33964 28868 34020
rect 28924 33628 28980 33684
rect 29036 37100 29092 37156
rect 28924 32338 28980 32340
rect 28924 32286 28926 32338
rect 28926 32286 28978 32338
rect 28978 32286 28980 32338
rect 28924 32284 28980 32286
rect 28812 31948 28868 32004
rect 28924 31724 28980 31780
rect 30380 47570 30436 47572
rect 30380 47518 30382 47570
rect 30382 47518 30434 47570
rect 30434 47518 30436 47570
rect 30380 47516 30436 47518
rect 30716 48636 30772 48692
rect 30716 47852 30772 47908
rect 30716 47516 30772 47572
rect 30828 47404 30884 47460
rect 30716 47234 30772 47236
rect 30716 47182 30718 47234
rect 30718 47182 30770 47234
rect 30770 47182 30772 47234
rect 30716 47180 30772 47182
rect 30492 46956 30548 47012
rect 30156 45612 30212 45668
rect 30044 45388 30100 45444
rect 30156 45106 30212 45108
rect 30156 45054 30158 45106
rect 30158 45054 30210 45106
rect 30210 45054 30212 45106
rect 30156 45052 30212 45054
rect 30604 46620 30660 46676
rect 30604 46396 30660 46452
rect 30380 45052 30436 45108
rect 30492 45890 30548 45892
rect 30492 45838 30494 45890
rect 30494 45838 30546 45890
rect 30546 45838 30548 45890
rect 30492 45836 30548 45838
rect 30044 44828 30100 44884
rect 29932 43484 29988 43540
rect 30604 45666 30660 45668
rect 30604 45614 30606 45666
rect 30606 45614 30658 45666
rect 30658 45614 30660 45666
rect 30604 45612 30660 45614
rect 30828 45836 30884 45892
rect 30716 45388 30772 45444
rect 32172 51772 32228 51828
rect 31836 50428 31892 50484
rect 31948 51100 32004 51156
rect 32172 51100 32228 51156
rect 31724 50092 31780 50148
rect 31500 48972 31556 49028
rect 31612 49644 31668 49700
rect 31276 48914 31332 48916
rect 31276 48862 31278 48914
rect 31278 48862 31330 48914
rect 31330 48862 31332 48914
rect 31276 48860 31332 48862
rect 31948 49644 32004 49700
rect 31500 48748 31556 48804
rect 31388 47682 31444 47684
rect 31388 47630 31390 47682
rect 31390 47630 31442 47682
rect 31442 47630 31444 47682
rect 31388 47628 31444 47630
rect 30940 45276 30996 45332
rect 31276 47458 31332 47460
rect 31276 47406 31278 47458
rect 31278 47406 31330 47458
rect 31330 47406 31332 47458
rect 31276 47404 31332 47406
rect 31052 46284 31108 46340
rect 30940 45106 30996 45108
rect 30940 45054 30942 45106
rect 30942 45054 30994 45106
rect 30994 45054 30996 45106
rect 30940 45052 30996 45054
rect 30716 44716 30772 44772
rect 30604 44434 30660 44436
rect 30604 44382 30606 44434
rect 30606 44382 30658 44434
rect 30658 44382 30660 44434
rect 30604 44380 30660 44382
rect 29820 43372 29876 43428
rect 30268 43314 30324 43316
rect 30268 43262 30270 43314
rect 30270 43262 30322 43314
rect 30322 43262 30324 43314
rect 30268 43260 30324 43262
rect 29820 41692 29876 41748
rect 30044 42700 30100 42756
rect 29820 41356 29876 41412
rect 29260 38722 29316 38724
rect 29260 38670 29262 38722
rect 29262 38670 29314 38722
rect 29314 38670 29316 38722
rect 29260 38668 29316 38670
rect 29260 38274 29316 38276
rect 29260 38222 29262 38274
rect 29262 38222 29314 38274
rect 29314 38222 29316 38274
rect 29260 38220 29316 38222
rect 29148 36876 29204 36932
rect 29484 38892 29540 38948
rect 29148 35474 29204 35476
rect 29148 35422 29150 35474
rect 29150 35422 29202 35474
rect 29202 35422 29204 35474
rect 29148 35420 29204 35422
rect 29372 37100 29428 37156
rect 29484 36428 29540 36484
rect 30604 44098 30660 44100
rect 30604 44046 30606 44098
rect 30606 44046 30658 44098
rect 30658 44046 30660 44098
rect 30604 44044 30660 44046
rect 30940 44716 30996 44772
rect 31164 47068 31220 47124
rect 31276 46114 31332 46116
rect 31276 46062 31278 46114
rect 31278 46062 31330 46114
rect 31330 46062 31332 46114
rect 31276 46060 31332 46062
rect 31388 45890 31444 45892
rect 31388 45838 31390 45890
rect 31390 45838 31442 45890
rect 31442 45838 31444 45890
rect 31388 45836 31444 45838
rect 31164 44716 31220 44772
rect 31388 44716 31444 44772
rect 31276 44604 31332 44660
rect 31388 44546 31444 44548
rect 31388 44494 31390 44546
rect 31390 44494 31442 44546
rect 31442 44494 31444 44546
rect 31388 44492 31444 44494
rect 31164 44434 31220 44436
rect 31164 44382 31166 44434
rect 31166 44382 31218 44434
rect 31218 44382 31220 44434
rect 31164 44380 31220 44382
rect 31388 44268 31444 44324
rect 30940 44044 30996 44100
rect 31276 44156 31332 44212
rect 30940 43036 30996 43092
rect 30716 41804 30772 41860
rect 29820 38668 29876 38724
rect 29932 40908 29988 40964
rect 29708 38556 29764 38612
rect 29596 35196 29652 35252
rect 29484 34914 29540 34916
rect 29484 34862 29486 34914
rect 29486 34862 29538 34914
rect 29538 34862 29540 34914
rect 29484 34860 29540 34862
rect 29260 34748 29316 34804
rect 29372 34412 29428 34468
rect 29372 32620 29428 32676
rect 29484 33628 29540 33684
rect 29036 31388 29092 31444
rect 29148 32284 29204 32340
rect 29372 32338 29428 32340
rect 29372 32286 29374 32338
rect 29374 32286 29426 32338
rect 29426 32286 29428 32338
rect 29372 32284 29428 32286
rect 30268 41468 30324 41524
rect 30156 38892 30212 38948
rect 30156 38444 30212 38500
rect 30492 41468 30548 41524
rect 30492 40124 30548 40180
rect 31388 43820 31444 43876
rect 31388 42530 31444 42532
rect 31388 42478 31390 42530
rect 31390 42478 31442 42530
rect 31442 42478 31444 42530
rect 31388 42476 31444 42478
rect 30716 41132 30772 41188
rect 30604 39564 30660 39620
rect 30940 41186 30996 41188
rect 30940 41134 30942 41186
rect 30942 41134 30994 41186
rect 30994 41134 30996 41186
rect 30940 41132 30996 41134
rect 31276 41468 31332 41524
rect 30940 40908 30996 40964
rect 31388 40236 31444 40292
rect 31836 48802 31892 48804
rect 31836 48750 31838 48802
rect 31838 48750 31890 48802
rect 31890 48750 31892 48802
rect 31836 48748 31892 48750
rect 31612 48188 31668 48244
rect 31612 47068 31668 47124
rect 31612 45612 31668 45668
rect 31836 45666 31892 45668
rect 31836 45614 31838 45666
rect 31838 45614 31890 45666
rect 31890 45614 31892 45666
rect 31836 45612 31892 45614
rect 31724 44716 31780 44772
rect 31612 43484 31668 43540
rect 32060 45948 32116 46004
rect 31948 44492 32004 44548
rect 32060 44940 32116 44996
rect 31836 44322 31892 44324
rect 31836 44270 31838 44322
rect 31838 44270 31890 44322
rect 31890 44270 31892 44322
rect 31836 44268 31892 44270
rect 31948 44156 32004 44212
rect 31948 43932 32004 43988
rect 30828 39900 30884 39956
rect 30604 37324 30660 37380
rect 30044 36428 30100 36484
rect 29820 35084 29876 35140
rect 30044 35980 30100 36036
rect 29820 34524 29876 34580
rect 29260 31164 29316 31220
rect 29148 30940 29204 30996
rect 28812 30770 28868 30772
rect 28812 30718 28814 30770
rect 28814 30718 28866 30770
rect 28866 30718 28868 30770
rect 28812 30716 28868 30718
rect 28364 29932 28420 29988
rect 28588 29484 28644 29540
rect 28364 28700 28420 28756
rect 28476 28476 28532 28532
rect 28252 21644 28308 21700
rect 28252 21308 28308 21364
rect 28364 28364 28420 28420
rect 29260 30770 29316 30772
rect 29260 30718 29262 30770
rect 29262 30718 29314 30770
rect 29314 30718 29316 30770
rect 29260 30716 29316 30718
rect 29036 30156 29092 30212
rect 29260 30268 29316 30324
rect 29260 29596 29316 29652
rect 29148 28924 29204 28980
rect 29036 28866 29092 28868
rect 29036 28814 29038 28866
rect 29038 28814 29090 28866
rect 29090 28814 29092 28866
rect 29036 28812 29092 28814
rect 28924 28700 28980 28756
rect 28700 28140 28756 28196
rect 28700 27132 28756 27188
rect 28476 26684 28532 26740
rect 28700 26684 28756 26740
rect 28588 25900 28644 25956
rect 28588 25452 28644 25508
rect 28924 27804 28980 27860
rect 28700 24220 28756 24276
rect 28700 23938 28756 23940
rect 28700 23886 28702 23938
rect 28702 23886 28754 23938
rect 28754 23886 28756 23938
rect 28700 23884 28756 23886
rect 28588 23100 28644 23156
rect 28700 23212 28756 23268
rect 28476 21698 28532 21700
rect 28476 21646 28478 21698
rect 28478 21646 28530 21698
rect 28530 21646 28532 21698
rect 28476 21644 28532 21646
rect 28588 21532 28644 21588
rect 28588 21308 28644 21364
rect 28364 20690 28420 20692
rect 28364 20638 28366 20690
rect 28366 20638 28418 20690
rect 28418 20638 28420 20690
rect 28364 20636 28420 20638
rect 28364 19234 28420 19236
rect 28364 19182 28366 19234
rect 28366 19182 28418 19234
rect 28418 19182 28420 19234
rect 28364 19180 28420 19182
rect 28028 17554 28084 17556
rect 28028 17502 28030 17554
rect 28030 17502 28082 17554
rect 28082 17502 28084 17554
rect 28028 17500 28084 17502
rect 28812 22540 28868 22596
rect 29036 26572 29092 26628
rect 29036 26290 29092 26292
rect 29036 26238 29038 26290
rect 29038 26238 29090 26290
rect 29090 26238 29092 26290
rect 29036 26236 29092 26238
rect 29260 25730 29316 25732
rect 29260 25678 29262 25730
rect 29262 25678 29314 25730
rect 29314 25678 29316 25730
rect 29260 25676 29316 25678
rect 29596 31948 29652 32004
rect 29484 31612 29540 31668
rect 29596 31276 29652 31332
rect 30268 35474 30324 35476
rect 30268 35422 30270 35474
rect 30270 35422 30322 35474
rect 30322 35422 30324 35474
rect 30268 35420 30324 35422
rect 30044 32284 30100 32340
rect 30156 34860 30212 34916
rect 30380 34914 30436 34916
rect 30380 34862 30382 34914
rect 30382 34862 30434 34914
rect 30434 34862 30436 34914
rect 30380 34860 30436 34862
rect 30268 34130 30324 34132
rect 30268 34078 30270 34130
rect 30270 34078 30322 34130
rect 30322 34078 30324 34130
rect 30268 34076 30324 34078
rect 30604 34412 30660 34468
rect 30380 32732 30436 32788
rect 30492 33628 30548 33684
rect 30604 33516 30660 33572
rect 30604 32732 30660 32788
rect 30380 32060 30436 32116
rect 30492 31948 30548 32004
rect 30156 31164 30212 31220
rect 29484 30380 29540 30436
rect 29820 30940 29876 30996
rect 30044 30940 30100 30996
rect 30044 30716 30100 30772
rect 30380 31052 30436 31108
rect 29484 30210 29540 30212
rect 29484 30158 29486 30210
rect 29486 30158 29538 30210
rect 29538 30158 29540 30210
rect 29484 30156 29540 30158
rect 30380 30210 30436 30212
rect 30380 30158 30382 30210
rect 30382 30158 30434 30210
rect 30434 30158 30436 30210
rect 30380 30156 30436 30158
rect 30044 30044 30100 30100
rect 29708 28642 29764 28644
rect 29708 28590 29710 28642
rect 29710 28590 29762 28642
rect 29762 28590 29764 28642
rect 29708 28588 29764 28590
rect 30268 28588 30324 28644
rect 29596 27580 29652 27636
rect 29596 27074 29652 27076
rect 29596 27022 29598 27074
rect 29598 27022 29650 27074
rect 29650 27022 29652 27074
rect 29596 27020 29652 27022
rect 29708 26908 29764 26964
rect 29708 26572 29764 26628
rect 29820 26460 29876 26516
rect 29708 26236 29764 26292
rect 29036 24332 29092 24388
rect 29036 23548 29092 23604
rect 29484 24332 29540 24388
rect 28812 21586 28868 21588
rect 28812 21534 28814 21586
rect 28814 21534 28866 21586
rect 28866 21534 28868 21586
rect 28812 21532 28868 21534
rect 29036 22764 29092 22820
rect 29148 22482 29204 22484
rect 29148 22430 29150 22482
rect 29150 22430 29202 22482
rect 29202 22430 29204 22482
rect 29148 22428 29204 22430
rect 29036 21308 29092 21364
rect 29148 21756 29204 21812
rect 28700 20636 28756 20692
rect 28700 19068 28756 19124
rect 28700 18562 28756 18564
rect 28700 18510 28702 18562
rect 28702 18510 28754 18562
rect 28754 18510 28756 18562
rect 28700 18508 28756 18510
rect 28588 16828 28644 16884
rect 27692 13074 27748 13076
rect 27692 13022 27694 13074
rect 27694 13022 27746 13074
rect 27746 13022 27748 13074
rect 27692 13020 27748 13022
rect 28252 13468 28308 13524
rect 27804 12460 27860 12516
rect 28140 13356 28196 13412
rect 27692 11788 27748 11844
rect 27580 11394 27636 11396
rect 27580 11342 27582 11394
rect 27582 11342 27634 11394
rect 27634 11342 27636 11394
rect 27580 11340 27636 11342
rect 27468 9826 27524 9828
rect 27468 9774 27470 9826
rect 27470 9774 27522 9826
rect 27522 9774 27524 9826
rect 27468 9772 27524 9774
rect 27020 7756 27076 7812
rect 27132 7644 27188 7700
rect 27468 8204 27524 8260
rect 27132 6690 27188 6692
rect 27132 6638 27134 6690
rect 27134 6638 27186 6690
rect 27186 6638 27188 6690
rect 27132 6636 27188 6638
rect 27244 6076 27300 6132
rect 26684 5964 26740 6020
rect 26012 5292 26068 5348
rect 25900 5122 25956 5124
rect 25900 5070 25902 5122
rect 25902 5070 25954 5122
rect 25954 5070 25956 5122
rect 25900 5068 25956 5070
rect 26796 5292 26852 5348
rect 27244 5346 27300 5348
rect 27244 5294 27246 5346
rect 27246 5294 27298 5346
rect 27298 5294 27300 5346
rect 27244 5292 27300 5294
rect 27468 5964 27524 6020
rect 28252 11676 28308 11732
rect 28028 11394 28084 11396
rect 28028 11342 28030 11394
rect 28030 11342 28082 11394
rect 28082 11342 28084 11394
rect 28028 11340 28084 11342
rect 28028 10668 28084 10724
rect 27916 9938 27972 9940
rect 27916 9886 27918 9938
rect 27918 9886 27970 9938
rect 27970 9886 27972 9938
rect 27916 9884 27972 9886
rect 27916 8988 27972 9044
rect 27916 8258 27972 8260
rect 27916 8206 27918 8258
rect 27918 8206 27970 8258
rect 27970 8206 27972 8258
rect 27916 8204 27972 8206
rect 27804 7756 27860 7812
rect 27804 7532 27860 7588
rect 27692 6636 27748 6692
rect 27804 5852 27860 5908
rect 27692 5404 27748 5460
rect 28028 5628 28084 5684
rect 27020 4732 27076 4788
rect 26012 3724 26068 3780
rect 25452 3164 25508 3220
rect 25228 2210 25284 2212
rect 25228 2158 25230 2210
rect 25230 2158 25282 2210
rect 25282 2158 25284 2210
rect 25228 2156 25284 2158
rect 25116 1932 25172 1988
rect 25004 1372 25060 1428
rect 24668 1148 24724 1204
rect 24444 1090 24500 1092
rect 24444 1038 24446 1090
rect 24446 1038 24498 1090
rect 24498 1038 24500 1090
rect 24444 1036 24500 1038
rect 24892 1202 24948 1204
rect 24892 1150 24894 1202
rect 24894 1150 24946 1202
rect 24946 1150 24948 1202
rect 24892 1148 24948 1150
rect 25676 3164 25732 3220
rect 25676 2828 25732 2884
rect 25676 1708 25732 1764
rect 24332 700 24388 756
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 24892 700 24948 756
rect 24892 476 24948 532
rect 13468 28 13524 84
rect 24444 252 24500 308
rect 25116 476 25172 532
rect 25340 588 25396 644
rect 26124 3554 26180 3556
rect 26124 3502 26126 3554
rect 26126 3502 26178 3554
rect 26178 3502 26180 3554
rect 26124 3500 26180 3502
rect 25788 1372 25844 1428
rect 26572 3778 26628 3780
rect 26572 3726 26574 3778
rect 26574 3726 26626 3778
rect 26626 3726 26628 3778
rect 26572 3724 26628 3726
rect 26460 3388 26516 3444
rect 27692 3778 27748 3780
rect 27692 3726 27694 3778
rect 27694 3726 27746 3778
rect 27746 3726 27748 3778
rect 27692 3724 27748 3726
rect 28028 5234 28084 5236
rect 28028 5182 28030 5234
rect 28030 5182 28082 5234
rect 28082 5182 28084 5234
rect 28028 5180 28084 5182
rect 27916 5122 27972 5124
rect 27916 5070 27918 5122
rect 27918 5070 27970 5122
rect 27970 5070 27972 5122
rect 27916 5068 27972 5070
rect 28700 16268 28756 16324
rect 29036 21084 29092 21140
rect 28924 19234 28980 19236
rect 28924 19182 28926 19234
rect 28926 19182 28978 19234
rect 28978 19182 28980 19234
rect 28924 19180 28980 19182
rect 29484 23100 29540 23156
rect 29148 20636 29204 20692
rect 29148 19906 29204 19908
rect 29148 19854 29150 19906
rect 29150 19854 29202 19906
rect 29202 19854 29204 19906
rect 29148 19852 29204 19854
rect 29036 17164 29092 17220
rect 29148 16658 29204 16660
rect 29148 16606 29150 16658
rect 29150 16606 29202 16658
rect 29202 16606 29204 16658
rect 29148 16604 29204 16606
rect 28924 16492 28980 16548
rect 28588 14418 28644 14420
rect 28588 14366 28590 14418
rect 28590 14366 28642 14418
rect 28642 14366 28644 14418
rect 28588 14364 28644 14366
rect 28364 6636 28420 6692
rect 29484 20748 29540 20804
rect 29708 22764 29764 22820
rect 30268 27468 30324 27524
rect 30044 26124 30100 26180
rect 30156 26012 30212 26068
rect 30156 25116 30212 25172
rect 30044 25004 30100 25060
rect 29932 24610 29988 24612
rect 29932 24558 29934 24610
rect 29934 24558 29986 24610
rect 29986 24558 29988 24610
rect 29932 24556 29988 24558
rect 30380 27244 30436 27300
rect 30268 23884 30324 23940
rect 29596 19852 29652 19908
rect 30156 23548 30212 23604
rect 30268 23212 30324 23268
rect 30604 28476 30660 28532
rect 30156 21980 30212 22036
rect 30268 22316 30324 22372
rect 31276 39394 31332 39396
rect 31276 39342 31278 39394
rect 31278 39342 31330 39394
rect 31330 39342 31332 39394
rect 31276 39340 31332 39342
rect 31388 38946 31444 38948
rect 31388 38894 31390 38946
rect 31390 38894 31442 38946
rect 31442 38894 31444 38946
rect 31388 38892 31444 38894
rect 31164 38668 31220 38724
rect 30940 38220 30996 38276
rect 31052 38332 31108 38388
rect 30940 37996 30996 38052
rect 31052 37212 31108 37268
rect 30940 36764 30996 36820
rect 31052 35698 31108 35700
rect 31052 35646 31054 35698
rect 31054 35646 31106 35698
rect 31106 35646 31108 35698
rect 31052 35644 31108 35646
rect 31276 38556 31332 38612
rect 31388 38108 31444 38164
rect 31388 35980 31444 36036
rect 31164 35532 31220 35588
rect 31276 35420 31332 35476
rect 31164 34748 31220 34804
rect 30940 34076 30996 34132
rect 31052 34412 31108 34468
rect 31052 33180 31108 33236
rect 31612 41858 31668 41860
rect 31612 41806 31614 41858
rect 31614 41806 31666 41858
rect 31666 41806 31668 41858
rect 31612 41804 31668 41806
rect 31948 42476 32004 42532
rect 31500 33516 31556 33572
rect 30940 32060 30996 32116
rect 30828 29426 30884 29428
rect 30828 29374 30830 29426
rect 30830 29374 30882 29426
rect 30882 29374 30884 29426
rect 30828 29372 30884 29374
rect 30828 27858 30884 27860
rect 30828 27806 30830 27858
rect 30830 27806 30882 27858
rect 30882 27806 30884 27858
rect 30828 27804 30884 27806
rect 31836 38610 31892 38612
rect 31836 38558 31838 38610
rect 31838 38558 31890 38610
rect 31890 38558 31892 38610
rect 31836 38556 31892 38558
rect 31836 35532 31892 35588
rect 31836 35308 31892 35364
rect 31836 34412 31892 34468
rect 31836 33852 31892 33908
rect 31052 29708 31108 29764
rect 31164 30940 31220 30996
rect 31052 29148 31108 29204
rect 30940 27132 30996 27188
rect 31052 28028 31108 28084
rect 30716 25004 30772 25060
rect 30268 21420 30324 21476
rect 30604 23154 30660 23156
rect 30604 23102 30606 23154
rect 30606 23102 30658 23154
rect 30658 23102 30660 23154
rect 30604 23100 30660 23102
rect 30604 22428 30660 22484
rect 29708 19740 29764 19796
rect 29484 19292 29540 19348
rect 29372 18396 29428 18452
rect 29484 17724 29540 17780
rect 29596 19180 29652 19236
rect 29372 14924 29428 14980
rect 29372 14700 29428 14756
rect 29484 16492 29540 16548
rect 29036 14364 29092 14420
rect 28924 14140 28980 14196
rect 29148 14252 29204 14308
rect 28812 11340 28868 11396
rect 28700 11116 28756 11172
rect 29036 10332 29092 10388
rect 28812 9212 28868 9268
rect 28588 8428 28644 8484
rect 28588 7980 28644 8036
rect 28476 6130 28532 6132
rect 28476 6078 28478 6130
rect 28478 6078 28530 6130
rect 28530 6078 28532 6130
rect 28476 6076 28532 6078
rect 28700 5682 28756 5684
rect 28700 5630 28702 5682
rect 28702 5630 28754 5682
rect 28754 5630 28756 5682
rect 28700 5628 28756 5630
rect 28588 5292 28644 5348
rect 26460 2828 26516 2884
rect 26572 2210 26628 2212
rect 26572 2158 26574 2210
rect 26574 2158 26626 2210
rect 26626 2158 26628 2210
rect 26572 2156 26628 2158
rect 26236 1148 26292 1204
rect 27804 2770 27860 2772
rect 27804 2718 27806 2770
rect 27806 2718 27858 2770
rect 27858 2718 27860 2770
rect 27804 2716 27860 2718
rect 28140 3666 28196 3668
rect 28140 3614 28142 3666
rect 28142 3614 28194 3666
rect 28194 3614 28196 3666
rect 28140 3612 28196 3614
rect 28028 3164 28084 3220
rect 27916 2492 27972 2548
rect 28028 1260 28084 1316
rect 27020 1036 27076 1092
rect 26236 364 26292 420
rect 26460 252 26516 308
rect 26684 924 26740 980
rect 27132 978 27188 980
rect 27132 926 27134 978
rect 27134 926 27186 978
rect 27186 926 27188 978
rect 27132 924 27188 926
rect 28476 3724 28532 3780
rect 29036 4732 29092 4788
rect 29260 13634 29316 13636
rect 29260 13582 29262 13634
rect 29262 13582 29314 13634
rect 29314 13582 29316 13634
rect 29260 13580 29316 13582
rect 29708 18508 29764 18564
rect 29820 20076 29876 20132
rect 29708 17052 29764 17108
rect 29596 16268 29652 16324
rect 29596 14754 29652 14756
rect 29596 14702 29598 14754
rect 29598 14702 29650 14754
rect 29650 14702 29652 14754
rect 29596 14700 29652 14702
rect 29484 14252 29540 14308
rect 30940 26012 30996 26068
rect 31052 23548 31108 23604
rect 31276 29484 31332 29540
rect 31612 31948 31668 32004
rect 31500 30770 31556 30772
rect 31500 30718 31502 30770
rect 31502 30718 31554 30770
rect 31554 30718 31556 30770
rect 31500 30716 31556 30718
rect 31500 30210 31556 30212
rect 31500 30158 31502 30210
rect 31502 30158 31554 30210
rect 31554 30158 31556 30210
rect 31500 30156 31556 30158
rect 33180 56252 33236 56308
rect 33404 56028 33460 56084
rect 32396 55356 32452 55412
rect 32508 55298 32564 55300
rect 32508 55246 32510 55298
rect 32510 55246 32562 55298
rect 32562 55246 32564 55298
rect 32508 55244 32564 55246
rect 32396 54012 32452 54068
rect 32508 53954 32564 53956
rect 32508 53902 32510 53954
rect 32510 53902 32562 53954
rect 32562 53902 32564 53954
rect 32508 53900 32564 53902
rect 32396 53676 32452 53732
rect 32844 54290 32900 54292
rect 32844 54238 32846 54290
rect 32846 54238 32898 54290
rect 32898 54238 32900 54290
rect 32844 54236 32900 54238
rect 32844 54012 32900 54068
rect 32732 53730 32788 53732
rect 32732 53678 32734 53730
rect 32734 53678 32786 53730
rect 32786 53678 32788 53730
rect 32732 53676 32788 53678
rect 32844 53452 32900 53508
rect 32620 52892 32676 52948
rect 32508 52162 32564 52164
rect 32508 52110 32510 52162
rect 32510 52110 32562 52162
rect 32562 52110 32564 52162
rect 32508 52108 32564 52110
rect 32620 51100 32676 51156
rect 33740 55858 33796 55860
rect 33740 55806 33742 55858
rect 33742 55806 33794 55858
rect 33794 55806 33796 55858
rect 33740 55804 33796 55806
rect 33404 55132 33460 55188
rect 33516 55692 33572 55748
rect 33852 55692 33908 55748
rect 33852 55410 33908 55412
rect 33852 55358 33854 55410
rect 33854 55358 33906 55410
rect 33906 55358 33908 55410
rect 33852 55356 33908 55358
rect 33628 55298 33684 55300
rect 33628 55246 33630 55298
rect 33630 55246 33682 55298
rect 33682 55246 33684 55298
rect 33628 55244 33684 55246
rect 34524 57148 34580 57204
rect 34748 56028 34804 56084
rect 34300 55468 34356 55524
rect 33516 54908 33572 54964
rect 34524 55356 34580 55412
rect 33180 54572 33236 54628
rect 33068 53116 33124 53172
rect 33628 53004 33684 53060
rect 33068 52892 33124 52948
rect 33068 52668 33124 52724
rect 32508 50370 32564 50372
rect 32508 50318 32510 50370
rect 32510 50318 32562 50370
rect 32562 50318 32564 50370
rect 32508 50316 32564 50318
rect 32732 50316 32788 50372
rect 32284 50092 32340 50148
rect 32396 49980 32452 50036
rect 32284 49922 32340 49924
rect 32284 49870 32286 49922
rect 32286 49870 32338 49922
rect 32338 49870 32340 49922
rect 32284 49868 32340 49870
rect 32732 49868 32788 49924
rect 33068 52444 33124 52500
rect 33180 52108 33236 52164
rect 34188 53954 34244 53956
rect 34188 53902 34190 53954
rect 34190 53902 34242 53954
rect 34242 53902 34244 53954
rect 34188 53900 34244 53902
rect 33964 53116 34020 53172
rect 34076 53452 34132 53508
rect 33852 52556 33908 52612
rect 33740 52274 33796 52276
rect 33740 52222 33742 52274
rect 33742 52222 33794 52274
rect 33794 52222 33796 52274
rect 33740 52220 33796 52222
rect 33628 51996 33684 52052
rect 32508 48802 32564 48804
rect 32508 48750 32510 48802
rect 32510 48750 32562 48802
rect 32562 48750 32564 48802
rect 32508 48748 32564 48750
rect 32396 47628 32452 47684
rect 32284 47068 32340 47124
rect 32396 45836 32452 45892
rect 32732 47292 32788 47348
rect 33068 50316 33124 50372
rect 33180 51772 33236 51828
rect 32956 49810 33012 49812
rect 32956 49758 32958 49810
rect 32958 49758 33010 49810
rect 33010 49758 33012 49810
rect 32956 49756 33012 49758
rect 32844 47068 32900 47124
rect 33068 47068 33124 47124
rect 35532 56364 35588 56420
rect 35196 55244 35252 55300
rect 36540 56364 36596 56420
rect 35308 55580 35364 55636
rect 34860 53676 34916 53732
rect 35084 54348 35140 54404
rect 35756 55468 35812 55524
rect 35308 53900 35364 53956
rect 35196 53788 35252 53844
rect 34972 53564 35028 53620
rect 35420 53618 35476 53620
rect 35420 53566 35422 53618
rect 35422 53566 35474 53618
rect 35474 53566 35476 53618
rect 35420 53564 35476 53566
rect 34636 53452 34692 53508
rect 34076 51996 34132 52052
rect 33516 51154 33572 51156
rect 33516 51102 33518 51154
rect 33518 51102 33570 51154
rect 33570 51102 33572 51154
rect 33516 51100 33572 51102
rect 34636 52332 34692 52388
rect 34748 52274 34804 52276
rect 34748 52222 34750 52274
rect 34750 52222 34802 52274
rect 34802 52222 34804 52274
rect 34748 52220 34804 52222
rect 33964 50316 34020 50372
rect 33516 48972 33572 49028
rect 33180 47404 33236 47460
rect 32956 46786 33012 46788
rect 32956 46734 32958 46786
rect 32958 46734 33010 46786
rect 33010 46734 33012 46786
rect 32956 46732 33012 46734
rect 32732 46396 32788 46452
rect 32620 46060 32676 46116
rect 32508 45666 32564 45668
rect 32508 45614 32510 45666
rect 32510 45614 32562 45666
rect 32562 45614 32564 45666
rect 32508 45612 32564 45614
rect 32508 44268 32564 44324
rect 32284 43260 32340 43316
rect 33292 48748 33348 48804
rect 33516 48636 33572 48692
rect 33516 48018 33572 48020
rect 33516 47966 33518 48018
rect 33518 47966 33570 48018
rect 33570 47966 33572 48018
rect 33516 47964 33572 47966
rect 34972 51772 35028 51828
rect 34412 49756 34468 49812
rect 34076 49308 34132 49364
rect 34524 49196 34580 49252
rect 33964 48748 34020 48804
rect 34188 48748 34244 48804
rect 34524 48748 34580 48804
rect 34636 49644 34692 49700
rect 34076 48636 34132 48692
rect 34412 48524 34468 48580
rect 33740 47516 33796 47572
rect 33404 46956 33460 47012
rect 33628 46844 33684 46900
rect 32844 44604 32900 44660
rect 32732 43708 32788 43764
rect 32508 43036 32564 43092
rect 32620 41970 32676 41972
rect 32620 41918 32622 41970
rect 32622 41918 32674 41970
rect 32674 41918 32676 41970
rect 32620 41916 32676 41918
rect 32956 42924 33012 42980
rect 32956 41244 33012 41300
rect 32956 40460 33012 40516
rect 32732 40124 32788 40180
rect 32284 40012 32340 40068
rect 33628 45836 33684 45892
rect 33180 45106 33236 45108
rect 33180 45054 33182 45106
rect 33182 45054 33234 45106
rect 33234 45054 33236 45106
rect 33180 45052 33236 45054
rect 33180 44268 33236 44324
rect 33292 45724 33348 45780
rect 34076 45778 34132 45780
rect 34076 45726 34078 45778
rect 34078 45726 34130 45778
rect 34130 45726 34132 45778
rect 34076 45724 34132 45726
rect 33852 45388 33908 45444
rect 33964 45500 34020 45556
rect 33068 40012 33124 40068
rect 33180 43260 33236 43316
rect 33292 41692 33348 41748
rect 33516 43426 33572 43428
rect 33516 43374 33518 43426
rect 33518 43374 33570 43426
rect 33570 43374 33572 43426
rect 33516 43372 33572 43374
rect 34188 45164 34244 45220
rect 34076 44322 34132 44324
rect 34076 44270 34078 44322
rect 34078 44270 34130 44322
rect 34130 44270 34132 44322
rect 34076 44268 34132 44270
rect 33964 43708 34020 43764
rect 33740 43372 33796 43428
rect 33628 42866 33684 42868
rect 33628 42814 33630 42866
rect 33630 42814 33682 42866
rect 33682 42814 33684 42866
rect 33628 42812 33684 42814
rect 33628 41970 33684 41972
rect 33628 41918 33630 41970
rect 33630 41918 33682 41970
rect 33682 41918 33684 41970
rect 33628 41916 33684 41918
rect 33404 41410 33460 41412
rect 33404 41358 33406 41410
rect 33406 41358 33458 41410
rect 33458 41358 33460 41410
rect 33404 41356 33460 41358
rect 33292 40460 33348 40516
rect 33628 40348 33684 40404
rect 33180 38668 33236 38724
rect 33292 40236 33348 40292
rect 32508 36988 32564 37044
rect 33068 37100 33124 37156
rect 32844 36764 32900 36820
rect 32060 34130 32116 34132
rect 32060 34078 32062 34130
rect 32062 34078 32114 34130
rect 32114 34078 32116 34130
rect 32060 34076 32116 34078
rect 31948 33068 32004 33124
rect 32060 31836 32116 31892
rect 32060 31612 32116 31668
rect 32284 34860 32340 34916
rect 32844 34748 32900 34804
rect 32956 36428 33012 36484
rect 32284 34188 32340 34244
rect 32508 34188 32564 34244
rect 32844 33852 32900 33908
rect 33180 36988 33236 37044
rect 33180 36482 33236 36484
rect 33180 36430 33182 36482
rect 33182 36430 33234 36482
rect 33234 36430 33236 36482
rect 33180 36428 33236 36430
rect 33628 39564 33684 39620
rect 33516 38610 33572 38612
rect 33516 38558 33518 38610
rect 33518 38558 33570 38610
rect 33570 38558 33572 38610
rect 33516 38556 33572 38558
rect 33292 36092 33348 36148
rect 33852 43036 33908 43092
rect 33852 40908 33908 40964
rect 34076 41244 34132 41300
rect 33852 40348 33908 40404
rect 33292 35698 33348 35700
rect 33292 35646 33294 35698
rect 33294 35646 33346 35698
rect 33346 35646 33348 35698
rect 33292 35644 33348 35646
rect 33180 35586 33236 35588
rect 33180 35534 33182 35586
rect 33182 35534 33234 35586
rect 33234 35534 33236 35586
rect 33180 35532 33236 35534
rect 33068 33852 33124 33908
rect 33180 34748 33236 34804
rect 32284 30940 32340 30996
rect 32396 31948 32452 32004
rect 32396 31052 32452 31108
rect 31836 29596 31892 29652
rect 31724 28866 31780 28868
rect 31724 28814 31726 28866
rect 31726 28814 31778 28866
rect 31778 28814 31780 28866
rect 31724 28812 31780 28814
rect 31612 28754 31668 28756
rect 31612 28702 31614 28754
rect 31614 28702 31666 28754
rect 31666 28702 31668 28754
rect 31612 28700 31668 28702
rect 31948 28588 32004 28644
rect 31724 27804 31780 27860
rect 31388 27468 31444 27524
rect 31836 27580 31892 27636
rect 31724 27186 31780 27188
rect 31724 27134 31726 27186
rect 31726 27134 31778 27186
rect 31778 27134 31780 27186
rect 31724 27132 31780 27134
rect 31836 27020 31892 27076
rect 31164 22988 31220 23044
rect 31388 26962 31444 26964
rect 31388 26910 31390 26962
rect 31390 26910 31442 26962
rect 31442 26910 31444 26962
rect 31388 26908 31444 26910
rect 31276 26684 31332 26740
rect 31500 26684 31556 26740
rect 31500 25788 31556 25844
rect 31612 26572 31668 26628
rect 31724 25452 31780 25508
rect 31836 25340 31892 25396
rect 31724 25282 31780 25284
rect 31724 25230 31726 25282
rect 31726 25230 31778 25282
rect 31778 25230 31780 25282
rect 31724 25228 31780 25230
rect 31500 24722 31556 24724
rect 31500 24670 31502 24722
rect 31502 24670 31554 24722
rect 31554 24670 31556 24722
rect 31500 24668 31556 24670
rect 31724 24220 31780 24276
rect 31500 23996 31556 24052
rect 31388 23212 31444 23268
rect 31052 22764 31108 22820
rect 30940 21980 30996 22036
rect 30716 21308 30772 21364
rect 30380 20076 30436 20132
rect 29932 19234 29988 19236
rect 29932 19182 29934 19234
rect 29934 19182 29986 19234
rect 29986 19182 29988 19234
rect 29932 19180 29988 19182
rect 30716 19068 30772 19124
rect 30044 18508 30100 18564
rect 29932 16156 29988 16212
rect 29932 13244 29988 13300
rect 30268 18450 30324 18452
rect 30268 18398 30270 18450
rect 30270 18398 30322 18450
rect 30322 18398 30324 18450
rect 30268 18396 30324 18398
rect 30156 17666 30212 17668
rect 30156 17614 30158 17666
rect 30158 17614 30210 17666
rect 30210 17614 30212 17666
rect 30156 17612 30212 17614
rect 30268 17106 30324 17108
rect 30268 17054 30270 17106
rect 30270 17054 30322 17106
rect 30322 17054 30324 17106
rect 30268 17052 30324 17054
rect 30604 16322 30660 16324
rect 30604 16270 30606 16322
rect 30606 16270 30658 16322
rect 30658 16270 30660 16322
rect 30604 16268 30660 16270
rect 30604 16044 30660 16100
rect 30604 15708 30660 15764
rect 30268 15148 30324 15204
rect 30268 14812 30324 14868
rect 30044 14252 30100 14308
rect 29484 11394 29540 11396
rect 29484 11342 29486 11394
rect 29486 11342 29538 11394
rect 29538 11342 29540 11394
rect 29484 11340 29540 11342
rect 29260 10722 29316 10724
rect 29260 10670 29262 10722
rect 29262 10670 29314 10722
rect 29314 10670 29316 10722
rect 29260 10668 29316 10670
rect 29372 6690 29428 6692
rect 29372 6638 29374 6690
rect 29374 6638 29426 6690
rect 29426 6638 29428 6690
rect 29372 6636 29428 6638
rect 29596 10332 29652 10388
rect 30268 14028 30324 14084
rect 30156 13020 30212 13076
rect 30828 18732 30884 18788
rect 30828 18172 30884 18228
rect 30716 12572 30772 12628
rect 30828 17948 30884 18004
rect 30156 11788 30212 11844
rect 30380 11900 30436 11956
rect 30268 11452 30324 11508
rect 30156 11340 30212 11396
rect 30380 10892 30436 10948
rect 30156 10444 30212 10500
rect 30268 10386 30324 10388
rect 30268 10334 30270 10386
rect 30270 10334 30322 10386
rect 30322 10334 30324 10386
rect 30268 10332 30324 10334
rect 29596 9826 29652 9828
rect 29596 9774 29598 9826
rect 29598 9774 29650 9826
rect 29650 9774 29652 9826
rect 29596 9772 29652 9774
rect 29484 6524 29540 6580
rect 29260 5628 29316 5684
rect 30044 9324 30100 9380
rect 30380 8652 30436 8708
rect 30156 7868 30212 7924
rect 30604 8540 30660 8596
rect 30380 7756 30436 7812
rect 30492 8428 30548 8484
rect 30268 7308 30324 7364
rect 30268 6972 30324 7028
rect 30492 6802 30548 6804
rect 30492 6750 30494 6802
rect 30494 6750 30546 6802
rect 30546 6750 30548 6802
rect 30492 6748 30548 6750
rect 30716 7868 30772 7924
rect 29932 5794 29988 5796
rect 29932 5742 29934 5794
rect 29934 5742 29986 5794
rect 29986 5742 29988 5794
rect 29932 5740 29988 5742
rect 30156 5740 30212 5796
rect 29148 4620 29204 4676
rect 28700 3500 28756 3556
rect 28588 3052 28644 3108
rect 29148 3778 29204 3780
rect 29148 3726 29150 3778
rect 29150 3726 29202 3778
rect 29202 3726 29204 3778
rect 29148 3724 29204 3726
rect 29372 4732 29428 4788
rect 30380 4732 30436 4788
rect 29372 3500 29428 3556
rect 29036 2658 29092 2660
rect 29036 2606 29038 2658
rect 29038 2606 29090 2658
rect 29090 2606 29092 2658
rect 29036 2604 29092 2606
rect 28924 2268 28980 2324
rect 28812 1372 28868 1428
rect 29260 3164 29316 3220
rect 29148 1372 29204 1428
rect 28700 1260 28756 1316
rect 29596 2098 29652 2100
rect 29596 2046 29598 2098
rect 29598 2046 29650 2098
rect 29650 2046 29652 2098
rect 29596 2044 29652 2046
rect 30156 3554 30212 3556
rect 30156 3502 30158 3554
rect 30158 3502 30210 3554
rect 30210 3502 30212 3554
rect 30156 3500 30212 3502
rect 29932 3052 29988 3108
rect 29036 1090 29092 1092
rect 29036 1038 29038 1090
rect 29038 1038 29090 1090
rect 29090 1038 29092 1090
rect 29036 1036 29092 1038
rect 27580 476 27636 532
rect 28364 476 28420 532
rect 28924 924 28980 980
rect 28476 252 28532 308
rect 29372 476 29428 532
rect 30268 2380 30324 2436
rect 29932 1484 29988 1540
rect 30604 4450 30660 4452
rect 30604 4398 30606 4450
rect 30606 4398 30658 4450
rect 30658 4398 30660 4450
rect 30604 4396 30660 4398
rect 31164 22370 31220 22372
rect 31164 22318 31166 22370
rect 31166 22318 31218 22370
rect 31218 22318 31220 22370
rect 31164 22316 31220 22318
rect 31276 20802 31332 20804
rect 31276 20750 31278 20802
rect 31278 20750 31330 20802
rect 31330 20750 31332 20802
rect 31276 20748 31332 20750
rect 31052 20018 31108 20020
rect 31052 19966 31054 20018
rect 31054 19966 31106 20018
rect 31106 19966 31108 20018
rect 31052 19964 31108 19966
rect 31276 20076 31332 20132
rect 31052 17666 31108 17668
rect 31052 17614 31054 17666
rect 31054 17614 31106 17666
rect 31106 17614 31108 17666
rect 31052 17612 31108 17614
rect 30940 17052 30996 17108
rect 31164 15932 31220 15988
rect 31276 18284 31332 18340
rect 31164 13020 31220 13076
rect 31724 21644 31780 21700
rect 32732 30994 32788 30996
rect 32732 30942 32734 30994
rect 32734 30942 32786 30994
rect 32786 30942 32788 30994
rect 32732 30940 32788 30942
rect 32060 24556 32116 24612
rect 32732 30716 32788 30772
rect 32060 23436 32116 23492
rect 31612 20578 31668 20580
rect 31612 20526 31614 20578
rect 31614 20526 31666 20578
rect 31666 20526 31668 20578
rect 31612 20524 31668 20526
rect 31500 19964 31556 20020
rect 31500 19794 31556 19796
rect 31500 19742 31502 19794
rect 31502 19742 31554 19794
rect 31554 19742 31556 19794
rect 31500 19740 31556 19742
rect 31612 18732 31668 18788
rect 31388 16380 31444 16436
rect 31500 18284 31556 18340
rect 31836 19068 31892 19124
rect 31724 18060 31780 18116
rect 31276 12124 31332 12180
rect 31388 15820 31444 15876
rect 31276 10610 31332 10612
rect 31276 10558 31278 10610
rect 31278 10558 31330 10610
rect 31330 10558 31332 10610
rect 31276 10556 31332 10558
rect 31724 17612 31780 17668
rect 31836 16828 31892 16884
rect 31948 16492 32004 16548
rect 32060 22540 32116 22596
rect 31500 15260 31556 15316
rect 31612 15932 31668 15988
rect 31948 15596 32004 15652
rect 31724 15260 31780 15316
rect 31612 15148 31668 15204
rect 31388 6636 31444 6692
rect 30828 4284 30884 4340
rect 31276 4396 31332 4452
rect 30380 1932 30436 1988
rect 30492 3164 30548 3220
rect 30268 1596 30324 1652
rect 30044 1372 30100 1428
rect 30156 1202 30212 1204
rect 30156 1150 30158 1202
rect 30158 1150 30210 1202
rect 30210 1150 30212 1202
rect 30156 1148 30212 1150
rect 30380 978 30436 980
rect 30380 926 30382 978
rect 30382 926 30434 978
rect 30434 926 30436 978
rect 30380 924 30436 926
rect 30268 252 30324 308
rect 30716 2492 30772 2548
rect 31164 3554 31220 3556
rect 31164 3502 31166 3554
rect 31166 3502 31218 3554
rect 31218 3502 31220 3554
rect 31164 3500 31220 3502
rect 31164 1708 31220 1764
rect 30492 140 30548 196
rect 30716 700 30772 756
rect 31612 14530 31668 14532
rect 31612 14478 31614 14530
rect 31614 14478 31666 14530
rect 31666 14478 31668 14530
rect 31612 14476 31668 14478
rect 31836 14140 31892 14196
rect 31836 13804 31892 13860
rect 31836 12796 31892 12852
rect 31724 12124 31780 12180
rect 31612 12066 31668 12068
rect 31612 12014 31614 12066
rect 31614 12014 31666 12066
rect 31666 12014 31668 12066
rect 31612 12012 31668 12014
rect 31836 11788 31892 11844
rect 31724 9548 31780 9604
rect 32396 30098 32452 30100
rect 32396 30046 32398 30098
rect 32398 30046 32450 30098
rect 32450 30046 32452 30098
rect 32396 30044 32452 30046
rect 32620 29484 32676 29540
rect 32396 29260 32452 29316
rect 32732 29036 32788 29092
rect 32508 27132 32564 27188
rect 33068 33570 33124 33572
rect 33068 33518 33070 33570
rect 33070 33518 33122 33570
rect 33122 33518 33124 33570
rect 33068 33516 33124 33518
rect 33068 32562 33124 32564
rect 33068 32510 33070 32562
rect 33070 32510 33122 32562
rect 33122 32510 33124 32562
rect 33068 32508 33124 32510
rect 32956 32396 33012 32452
rect 33292 34076 33348 34132
rect 33068 31890 33124 31892
rect 33068 31838 33070 31890
rect 33070 31838 33122 31890
rect 33122 31838 33124 31890
rect 33068 31836 33124 31838
rect 33180 32060 33236 32116
rect 32956 30268 33012 30324
rect 32956 29708 33012 29764
rect 33180 29932 33236 29988
rect 32956 29314 33012 29316
rect 32956 29262 32958 29314
rect 32958 29262 33010 29314
rect 33010 29262 33012 29314
rect 32956 29260 33012 29262
rect 33068 28812 33124 28868
rect 33180 28642 33236 28644
rect 33180 28590 33182 28642
rect 33182 28590 33234 28642
rect 33234 28590 33236 28642
rect 33180 28588 33236 28590
rect 32956 27132 33012 27188
rect 32732 26908 32788 26964
rect 32396 26290 32452 26292
rect 32396 26238 32398 26290
rect 32398 26238 32450 26290
rect 32450 26238 32452 26290
rect 32396 26236 32452 26238
rect 32396 25564 32452 25620
rect 33852 40124 33908 40180
rect 33628 37212 33684 37268
rect 33964 40012 34020 40068
rect 34524 47570 34580 47572
rect 34524 47518 34526 47570
rect 34526 47518 34578 47570
rect 34578 47518 34580 47570
rect 34524 47516 34580 47518
rect 34748 48748 34804 48804
rect 35196 51772 35252 51828
rect 35196 51154 35252 51156
rect 35196 51102 35198 51154
rect 35198 51102 35250 51154
rect 35250 51102 35252 51154
rect 35196 51100 35252 51102
rect 35084 50034 35140 50036
rect 35084 49982 35086 50034
rect 35086 49982 35138 50034
rect 35138 49982 35140 50034
rect 35084 49980 35140 49982
rect 34972 48524 35028 48580
rect 35084 48354 35140 48356
rect 35084 48302 35086 48354
rect 35086 48302 35138 48354
rect 35138 48302 35140 48354
rect 35084 48300 35140 48302
rect 34860 47234 34916 47236
rect 34860 47182 34862 47234
rect 34862 47182 34914 47234
rect 34914 47182 34916 47234
rect 34860 47180 34916 47182
rect 34524 43820 34580 43876
rect 35420 52050 35476 52052
rect 35420 51998 35422 52050
rect 35422 51998 35474 52050
rect 35474 51998 35476 52050
rect 35420 51996 35476 51998
rect 36876 56140 36932 56196
rect 36428 56082 36484 56084
rect 36428 56030 36430 56082
rect 36430 56030 36482 56082
rect 36482 56030 36484 56082
rect 36428 56028 36484 56030
rect 36988 56028 37044 56084
rect 37324 56812 37380 56868
rect 36092 55858 36148 55860
rect 36092 55806 36094 55858
rect 36094 55806 36146 55858
rect 36146 55806 36148 55858
rect 36092 55804 36148 55806
rect 37100 55858 37156 55860
rect 37100 55806 37102 55858
rect 37102 55806 37154 55858
rect 37154 55806 37156 55858
rect 37100 55804 37156 55806
rect 36316 55410 36372 55412
rect 36316 55358 36318 55410
rect 36318 55358 36370 55410
rect 36370 55358 36372 55410
rect 36316 55356 36372 55358
rect 35644 54012 35700 54068
rect 35756 53842 35812 53844
rect 35756 53790 35758 53842
rect 35758 53790 35810 53842
rect 35810 53790 35812 53842
rect 35756 53788 35812 53790
rect 36876 53788 36932 53844
rect 36540 53564 36596 53620
rect 36540 52780 36596 52836
rect 35644 52668 35700 52724
rect 35868 52274 35924 52276
rect 35868 52222 35870 52274
rect 35870 52222 35922 52274
rect 35922 52222 35924 52274
rect 35868 52220 35924 52222
rect 36428 52108 36484 52164
rect 35644 51772 35700 51828
rect 36764 52332 36820 52388
rect 36876 52668 36932 52724
rect 36540 51548 36596 51604
rect 36540 51324 36596 51380
rect 35420 51100 35476 51156
rect 35980 50818 36036 50820
rect 35980 50766 35982 50818
rect 35982 50766 36034 50818
rect 36034 50766 36036 50818
rect 35980 50764 36036 50766
rect 35644 50594 35700 50596
rect 35644 50542 35646 50594
rect 35646 50542 35698 50594
rect 35698 50542 35700 50594
rect 35644 50540 35700 50542
rect 35868 50428 35924 50484
rect 35644 49810 35700 49812
rect 35644 49758 35646 49810
rect 35646 49758 35698 49810
rect 35698 49758 35700 49810
rect 35644 49756 35700 49758
rect 35308 49084 35364 49140
rect 35308 48412 35364 48468
rect 35532 48242 35588 48244
rect 35532 48190 35534 48242
rect 35534 48190 35586 48242
rect 35586 48190 35588 48242
rect 35532 48188 35588 48190
rect 35196 47964 35252 48020
rect 35980 48972 36036 49028
rect 36204 50876 36260 50932
rect 36204 50652 36260 50708
rect 36428 50706 36484 50708
rect 36428 50654 36430 50706
rect 36430 50654 36482 50706
rect 36482 50654 36484 50706
rect 36428 50652 36484 50654
rect 36428 50034 36484 50036
rect 36428 49982 36430 50034
rect 36430 49982 36482 50034
rect 36482 49982 36484 50034
rect 36428 49980 36484 49982
rect 36316 49196 36372 49252
rect 36316 48748 36372 48804
rect 36540 48860 36596 48916
rect 35308 46956 35364 47012
rect 34412 43372 34468 43428
rect 34748 46620 34804 46676
rect 35420 46620 35476 46676
rect 34860 46172 34916 46228
rect 34748 44882 34804 44884
rect 34748 44830 34750 44882
rect 34750 44830 34802 44882
rect 34802 44830 34804 44882
rect 34748 44828 34804 44830
rect 34748 43650 34804 43652
rect 34748 43598 34750 43650
rect 34750 43598 34802 43650
rect 34802 43598 34804 43650
rect 34748 43596 34804 43598
rect 35084 45948 35140 46004
rect 35308 45948 35364 46004
rect 34748 43036 34804 43092
rect 34636 42924 34692 42980
rect 34972 43036 35028 43092
rect 35308 43932 35364 43988
rect 35196 43036 35252 43092
rect 35084 42028 35140 42084
rect 34524 41916 34580 41972
rect 34412 41244 34468 41300
rect 35196 41858 35252 41860
rect 35196 41806 35198 41858
rect 35198 41806 35250 41858
rect 35250 41806 35252 41858
rect 35196 41804 35252 41806
rect 34748 41746 34804 41748
rect 34748 41694 34750 41746
rect 34750 41694 34802 41746
rect 34802 41694 34804 41746
rect 34748 41692 34804 41694
rect 35644 47570 35700 47572
rect 35644 47518 35646 47570
rect 35646 47518 35698 47570
rect 35698 47518 35700 47570
rect 35644 47516 35700 47518
rect 35532 45948 35588 46004
rect 35868 46002 35924 46004
rect 35868 45950 35870 46002
rect 35870 45950 35922 46002
rect 35922 45950 35924 46002
rect 35868 45948 35924 45950
rect 35644 45500 35700 45556
rect 35532 44492 35588 44548
rect 35644 43426 35700 43428
rect 35644 43374 35646 43426
rect 35646 43374 35698 43426
rect 35698 43374 35700 43426
rect 35644 43372 35700 43374
rect 35532 42924 35588 42980
rect 35644 43036 35700 43092
rect 35756 42812 35812 42868
rect 35532 41804 35588 41860
rect 34636 41356 34692 41412
rect 34300 40684 34356 40740
rect 34076 39618 34132 39620
rect 34076 39566 34078 39618
rect 34078 39566 34130 39618
rect 34130 39566 34132 39618
rect 34076 39564 34132 39566
rect 34076 38892 34132 38948
rect 34188 39676 34244 39732
rect 33852 36988 33908 37044
rect 33964 38668 34020 38724
rect 34076 38556 34132 38612
rect 34076 37324 34132 37380
rect 33740 35980 33796 36036
rect 33628 35138 33684 35140
rect 33628 35086 33630 35138
rect 33630 35086 33682 35138
rect 33682 35086 33684 35138
rect 33628 35084 33684 35086
rect 33628 34748 33684 34804
rect 33628 34242 33684 34244
rect 33628 34190 33630 34242
rect 33630 34190 33682 34242
rect 33682 34190 33684 34242
rect 33628 34188 33684 34190
rect 33740 34412 33796 34468
rect 33740 34076 33796 34132
rect 33516 33516 33572 33572
rect 33628 33852 33684 33908
rect 33516 33292 33572 33348
rect 33516 32620 33572 32676
rect 33404 32396 33460 32452
rect 33964 36540 34020 36596
rect 33964 35980 34020 36036
rect 34188 35420 34244 35476
rect 33852 33292 33908 33348
rect 33964 34972 34020 35028
rect 34300 34188 34356 34244
rect 34636 40796 34692 40852
rect 34748 41468 34804 41524
rect 34524 39676 34580 39732
rect 34636 38722 34692 38724
rect 34636 38670 34638 38722
rect 34638 38670 34690 38722
rect 34690 38670 34692 38722
rect 34636 38668 34692 38670
rect 35308 41244 35364 41300
rect 35196 40684 35252 40740
rect 35084 40402 35140 40404
rect 35084 40350 35086 40402
rect 35086 40350 35138 40402
rect 35138 40350 35140 40402
rect 35084 40348 35140 40350
rect 34860 38108 34916 38164
rect 34972 40236 35028 40292
rect 34748 37100 34804 37156
rect 34860 37212 34916 37268
rect 34748 36482 34804 36484
rect 34748 36430 34750 36482
rect 34750 36430 34802 36482
rect 34802 36430 34804 36482
rect 34748 36428 34804 36430
rect 34636 34412 34692 34468
rect 34412 33516 34468 33572
rect 34188 33122 34244 33124
rect 34188 33070 34190 33122
rect 34190 33070 34242 33122
rect 34242 33070 34244 33122
rect 34188 33068 34244 33070
rect 34076 32732 34132 32788
rect 34524 34076 34580 34132
rect 34300 32450 34356 32452
rect 34300 32398 34302 32450
rect 34302 32398 34354 32450
rect 34354 32398 34356 32450
rect 34300 32396 34356 32398
rect 33740 31276 33796 31332
rect 34076 31388 34132 31444
rect 33628 31164 33684 31220
rect 33964 31052 34020 31108
rect 33404 30716 33460 30772
rect 33404 30156 33460 30212
rect 33628 30156 33684 30212
rect 34412 30828 34468 30884
rect 33964 30210 34020 30212
rect 33964 30158 33966 30210
rect 33966 30158 34018 30210
rect 34018 30158 34020 30210
rect 33964 30156 34020 30158
rect 34076 30716 34132 30772
rect 33964 29820 34020 29876
rect 33516 29036 33572 29092
rect 33964 29036 34020 29092
rect 33404 28588 33460 28644
rect 34188 30492 34244 30548
rect 34188 29820 34244 29876
rect 34300 29314 34356 29316
rect 34300 29262 34302 29314
rect 34302 29262 34354 29314
rect 34354 29262 34356 29314
rect 34300 29260 34356 29262
rect 33740 27468 33796 27524
rect 32732 26236 32788 26292
rect 32956 25564 33012 25620
rect 33068 26012 33124 26068
rect 32620 25452 32676 25508
rect 32284 25004 32340 25060
rect 32956 25004 33012 25060
rect 32508 24332 32564 24388
rect 32284 22988 32340 23044
rect 32396 24108 32452 24164
rect 32172 22428 32228 22484
rect 32844 24108 32900 24164
rect 33068 23996 33124 24052
rect 33292 26012 33348 26068
rect 33292 24332 33348 24388
rect 32508 23436 32564 23492
rect 32732 23436 32788 23492
rect 32620 23154 32676 23156
rect 32620 23102 32622 23154
rect 32622 23102 32674 23154
rect 32674 23102 32676 23154
rect 32620 23100 32676 23102
rect 32508 21980 32564 22036
rect 32396 21308 32452 21364
rect 32620 21308 32676 21364
rect 32620 20972 32676 21028
rect 32956 23436 33012 23492
rect 34860 34748 34916 34804
rect 34748 32620 34804 32676
rect 34860 33068 34916 33124
rect 35420 40908 35476 40964
rect 35868 41468 35924 41524
rect 36092 44268 36148 44324
rect 36316 47346 36372 47348
rect 36316 47294 36318 47346
rect 36318 47294 36370 47346
rect 36370 47294 36372 47346
rect 36316 47292 36372 47294
rect 36764 51324 36820 51380
rect 37212 50764 37268 50820
rect 36988 50652 37044 50708
rect 36876 50428 36932 50484
rect 37436 56140 37492 56196
rect 38108 55858 38164 55860
rect 38108 55806 38110 55858
rect 38110 55806 38162 55858
rect 38162 55806 38164 55858
rect 38108 55804 38164 55806
rect 37772 55468 37828 55524
rect 38780 56476 38836 56532
rect 38668 55692 38724 55748
rect 37548 55410 37604 55412
rect 37548 55358 37550 55410
rect 37550 55358 37602 55410
rect 37602 55358 37604 55410
rect 37548 55356 37604 55358
rect 38668 55132 38724 55188
rect 37548 54684 37604 54740
rect 37436 51324 37492 51380
rect 37436 50540 37492 50596
rect 37324 50428 37380 50484
rect 37212 49980 37268 50036
rect 37324 49868 37380 49924
rect 37100 49756 37156 49812
rect 36428 47068 36484 47124
rect 36316 45778 36372 45780
rect 36316 45726 36318 45778
rect 36318 45726 36370 45778
rect 36370 45726 36372 45778
rect 36316 45724 36372 45726
rect 36764 47404 36820 47460
rect 36988 47292 37044 47348
rect 36876 46956 36932 47012
rect 36764 46786 36820 46788
rect 36764 46734 36766 46786
rect 36766 46734 36818 46786
rect 36818 46734 36820 46786
rect 36764 46732 36820 46734
rect 36652 46172 36708 46228
rect 36988 46284 37044 46340
rect 37212 48130 37268 48132
rect 37212 48078 37214 48130
rect 37214 48078 37266 48130
rect 37266 48078 37268 48130
rect 37212 48076 37268 48078
rect 38108 54796 38164 54852
rect 37772 54684 37828 54740
rect 38668 54738 38724 54740
rect 38668 54686 38670 54738
rect 38670 54686 38722 54738
rect 38722 54686 38724 54738
rect 38668 54684 38724 54686
rect 37772 53618 37828 53620
rect 37772 53566 37774 53618
rect 37774 53566 37826 53618
rect 37826 53566 37828 53618
rect 37772 53564 37828 53566
rect 38108 52722 38164 52724
rect 38108 52670 38110 52722
rect 38110 52670 38162 52722
rect 38162 52670 38164 52722
rect 38108 52668 38164 52670
rect 37772 51324 37828 51380
rect 37548 49868 37604 49924
rect 37660 50652 37716 50708
rect 37324 47292 37380 47348
rect 37436 49308 37492 49364
rect 37436 46732 37492 46788
rect 37548 49196 37604 49252
rect 37884 50876 37940 50932
rect 37884 50540 37940 50596
rect 38108 51996 38164 52052
rect 38108 51266 38164 51268
rect 38108 51214 38110 51266
rect 38110 51214 38162 51266
rect 38162 51214 38164 51266
rect 38108 51212 38164 51214
rect 38108 49980 38164 50036
rect 38108 49810 38164 49812
rect 38108 49758 38110 49810
rect 38110 49758 38162 49810
rect 38162 49758 38164 49810
rect 38108 49756 38164 49758
rect 36540 45388 36596 45444
rect 37996 48972 38052 49028
rect 37996 48748 38052 48804
rect 37548 46396 37604 46452
rect 37772 47628 37828 47684
rect 37772 46396 37828 46452
rect 37996 46284 38052 46340
rect 37436 46172 37492 46228
rect 37324 45500 37380 45556
rect 37436 45724 37492 45780
rect 37212 45052 37268 45108
rect 36204 43932 36260 43988
rect 37100 44322 37156 44324
rect 37100 44270 37102 44322
rect 37102 44270 37154 44322
rect 37154 44270 37156 44322
rect 37100 44268 37156 44270
rect 36652 43932 36708 43988
rect 36764 44156 36820 44212
rect 36652 43708 36708 43764
rect 36092 43036 36148 43092
rect 35644 40460 35700 40516
rect 35756 40290 35812 40292
rect 35756 40238 35758 40290
rect 35758 40238 35810 40290
rect 35810 40238 35812 40290
rect 35756 40236 35812 40238
rect 35084 39564 35140 39620
rect 35308 39452 35364 39508
rect 35196 36876 35252 36932
rect 35196 36594 35252 36596
rect 35196 36542 35198 36594
rect 35198 36542 35250 36594
rect 35250 36542 35252 36594
rect 35196 36540 35252 36542
rect 35308 36764 35364 36820
rect 35980 41244 36036 41300
rect 35868 39788 35924 39844
rect 35980 41020 36036 41076
rect 35644 39452 35700 39508
rect 35868 39116 35924 39172
rect 35756 38946 35812 38948
rect 35756 38894 35758 38946
rect 35758 38894 35810 38946
rect 35810 38894 35812 38946
rect 35756 38892 35812 38894
rect 35644 37100 35700 37156
rect 35532 36482 35588 36484
rect 35532 36430 35534 36482
rect 35534 36430 35586 36482
rect 35586 36430 35588 36482
rect 35532 36428 35588 36430
rect 35532 34748 35588 34804
rect 35420 34412 35476 34468
rect 35308 34188 35364 34244
rect 35532 33404 35588 33460
rect 35644 34188 35700 34244
rect 34860 32172 34916 32228
rect 34636 31778 34692 31780
rect 34636 31726 34638 31778
rect 34638 31726 34690 31778
rect 34690 31726 34692 31778
rect 34636 31724 34692 31726
rect 34748 31388 34804 31444
rect 34636 30492 34692 30548
rect 34972 31890 35028 31892
rect 34972 31838 34974 31890
rect 34974 31838 35026 31890
rect 35026 31838 35028 31890
rect 34972 31836 35028 31838
rect 35308 32732 35364 32788
rect 35084 31164 35140 31220
rect 35196 32620 35252 32676
rect 35308 32450 35364 32452
rect 35308 32398 35310 32450
rect 35310 32398 35362 32450
rect 35362 32398 35364 32450
rect 35308 32396 35364 32398
rect 35644 32060 35700 32116
rect 34860 30268 34916 30324
rect 34748 29650 34804 29652
rect 34748 29598 34750 29650
rect 34750 29598 34802 29650
rect 34802 29598 34804 29650
rect 34748 29596 34804 29598
rect 34412 28476 34468 28532
rect 33852 26460 33908 26516
rect 33964 28364 34020 28420
rect 33740 25506 33796 25508
rect 33740 25454 33742 25506
rect 33742 25454 33794 25506
rect 33794 25454 33796 25506
rect 33740 25452 33796 25454
rect 33628 25340 33684 25396
rect 33740 24668 33796 24724
rect 33404 23548 33460 23604
rect 33516 24556 33572 24612
rect 32508 20412 32564 20468
rect 32284 19964 32340 20020
rect 32844 19740 32900 19796
rect 33068 22988 33124 23044
rect 33292 23100 33348 23156
rect 33404 22876 33460 22932
rect 33404 22428 33460 22484
rect 33628 24162 33684 24164
rect 33628 24110 33630 24162
rect 33630 24110 33682 24162
rect 33682 24110 33684 24162
rect 33628 24108 33684 24110
rect 33628 22092 33684 22148
rect 33180 21196 33236 21252
rect 33404 21196 33460 21252
rect 33180 20524 33236 20580
rect 33292 20076 33348 20132
rect 33292 19740 33348 19796
rect 33068 19180 33124 19236
rect 32508 18732 32564 18788
rect 32508 16828 32564 16884
rect 32284 15820 32340 15876
rect 32508 16380 32564 16436
rect 32284 15314 32340 15316
rect 32284 15262 32286 15314
rect 32286 15262 32338 15314
rect 32338 15262 32340 15314
rect 32284 15260 32340 15262
rect 32284 13858 32340 13860
rect 32284 13806 32286 13858
rect 32286 13806 32338 13858
rect 32338 13806 32340 13858
rect 32284 13804 32340 13806
rect 32284 11676 32340 11732
rect 32396 9548 32452 9604
rect 31612 8316 31668 8372
rect 31836 8316 31892 8372
rect 31724 8034 31780 8036
rect 31724 7982 31726 8034
rect 31726 7982 31778 8034
rect 31778 7982 31780 8034
rect 31724 7980 31780 7982
rect 31948 8092 32004 8148
rect 32396 8316 32452 8372
rect 32284 8204 32340 8260
rect 32732 18396 32788 18452
rect 33180 18508 33236 18564
rect 33068 17948 33124 18004
rect 32956 17724 33012 17780
rect 32844 16994 32900 16996
rect 32844 16942 32846 16994
rect 32846 16942 32898 16994
rect 32898 16942 32900 16994
rect 32844 16940 32900 16942
rect 33404 19628 33460 19684
rect 33516 18450 33572 18452
rect 33516 18398 33518 18450
rect 33518 18398 33570 18450
rect 33570 18398 33572 18450
rect 33516 18396 33572 18398
rect 33292 17948 33348 18004
rect 33292 16882 33348 16884
rect 33292 16830 33294 16882
rect 33294 16830 33346 16882
rect 33346 16830 33348 16882
rect 33292 16828 33348 16830
rect 33180 16492 33236 16548
rect 33068 16380 33124 16436
rect 32956 16210 33012 16212
rect 32956 16158 32958 16210
rect 32958 16158 33010 16210
rect 33010 16158 33012 16210
rect 32956 16156 33012 16158
rect 32844 16044 32900 16100
rect 32732 15820 32788 15876
rect 32732 14812 32788 14868
rect 32844 14252 32900 14308
rect 32844 14028 32900 14084
rect 32620 13020 32676 13076
rect 32620 11004 32676 11060
rect 32620 8428 32676 8484
rect 32956 13804 33012 13860
rect 33628 15820 33684 15876
rect 33852 23212 33908 23268
rect 33852 22316 33908 22372
rect 34076 28252 34132 28308
rect 34300 28140 34356 28196
rect 34188 27132 34244 27188
rect 34076 26962 34132 26964
rect 34076 26910 34078 26962
rect 34078 26910 34130 26962
rect 34130 26910 34132 26962
rect 34076 26908 34132 26910
rect 34076 25004 34132 25060
rect 34076 24834 34132 24836
rect 34076 24782 34078 24834
rect 34078 24782 34130 24834
rect 34130 24782 34132 24834
rect 34076 24780 34132 24782
rect 34076 23436 34132 23492
rect 34748 28924 34804 28980
rect 34524 27580 34580 27636
rect 34412 26908 34468 26964
rect 34860 28812 34916 28868
rect 35308 31778 35364 31780
rect 35308 31726 35310 31778
rect 35310 31726 35362 31778
rect 35362 31726 35364 31778
rect 35308 31724 35364 31726
rect 35532 31890 35588 31892
rect 35532 31838 35534 31890
rect 35534 31838 35586 31890
rect 35586 31838 35588 31890
rect 35532 31836 35588 31838
rect 35420 31388 35476 31444
rect 35644 31388 35700 31444
rect 35308 31276 35364 31332
rect 35196 29036 35252 29092
rect 35308 28700 35364 28756
rect 35868 37100 35924 37156
rect 36428 42978 36484 42980
rect 36428 42926 36430 42978
rect 36430 42926 36482 42978
rect 36482 42926 36484 42978
rect 36428 42924 36484 42926
rect 36316 42700 36372 42756
rect 36876 43596 36932 43652
rect 37100 43260 37156 43316
rect 37100 42754 37156 42756
rect 37100 42702 37102 42754
rect 37102 42702 37154 42754
rect 37154 42702 37156 42754
rect 37100 42700 37156 42702
rect 36652 42588 36708 42644
rect 37324 44828 37380 44884
rect 37884 44994 37940 44996
rect 37884 44942 37886 44994
rect 37886 44942 37938 44994
rect 37938 44942 37940 44994
rect 37884 44940 37940 44942
rect 37548 44604 37604 44660
rect 37660 44716 37716 44772
rect 37436 44546 37492 44548
rect 37436 44494 37438 44546
rect 37438 44494 37490 44546
rect 37490 44494 37492 44546
rect 37436 44492 37492 44494
rect 37660 44492 37716 44548
rect 37548 44434 37604 44436
rect 37548 44382 37550 44434
rect 37550 44382 37602 44434
rect 37602 44382 37604 44434
rect 37548 44380 37604 44382
rect 39116 55858 39172 55860
rect 39116 55806 39118 55858
rect 39118 55806 39170 55858
rect 39170 55806 39172 55858
rect 39116 55804 39172 55806
rect 38892 55410 38948 55412
rect 38892 55358 38894 55410
rect 38894 55358 38946 55410
rect 38946 55358 38948 55410
rect 38892 55356 38948 55358
rect 40012 55244 40068 55300
rect 39564 54572 39620 54628
rect 39004 52668 39060 52724
rect 38892 51324 38948 51380
rect 38556 50540 38612 50596
rect 38668 51100 38724 51156
rect 38332 49196 38388 49252
rect 38332 48524 38388 48580
rect 38668 48018 38724 48020
rect 38668 47966 38670 48018
rect 38670 47966 38722 48018
rect 38722 47966 38724 48018
rect 38668 47964 38724 47966
rect 38444 47570 38500 47572
rect 38444 47518 38446 47570
rect 38446 47518 38498 47570
rect 38498 47518 38500 47570
rect 38444 47516 38500 47518
rect 38556 47404 38612 47460
rect 38444 47180 38500 47236
rect 38220 45724 38276 45780
rect 38108 44380 38164 44436
rect 38220 45276 38276 45332
rect 37660 44268 37716 44324
rect 37436 44044 37492 44100
rect 37324 43260 37380 43316
rect 37212 42476 37268 42532
rect 37100 42028 37156 42084
rect 36764 40962 36820 40964
rect 36764 40910 36766 40962
rect 36766 40910 36818 40962
rect 36818 40910 36820 40962
rect 36764 40908 36820 40910
rect 36652 40402 36708 40404
rect 36652 40350 36654 40402
rect 36654 40350 36706 40402
rect 36706 40350 36708 40402
rect 36652 40348 36708 40350
rect 36428 40290 36484 40292
rect 36428 40238 36430 40290
rect 36430 40238 36482 40290
rect 36482 40238 36484 40290
rect 36428 40236 36484 40238
rect 36204 39452 36260 39508
rect 36092 38780 36148 38836
rect 36764 38946 36820 38948
rect 36764 38894 36766 38946
rect 36766 38894 36818 38946
rect 36818 38894 36820 38946
rect 36764 38892 36820 38894
rect 37436 42028 37492 42084
rect 37548 42978 37604 42980
rect 37548 42926 37550 42978
rect 37550 42926 37602 42978
rect 37602 42926 37604 42978
rect 37548 42924 37604 42926
rect 37212 41804 37268 41860
rect 37436 41858 37492 41860
rect 37436 41806 37438 41858
rect 37438 41806 37490 41858
rect 37490 41806 37492 41858
rect 37436 41804 37492 41806
rect 36988 40236 37044 40292
rect 37548 41020 37604 41076
rect 37436 40236 37492 40292
rect 37548 40796 37604 40852
rect 37996 43820 38052 43876
rect 37772 43314 37828 43316
rect 37772 43262 37774 43314
rect 37774 43262 37826 43314
rect 37826 43262 37828 43314
rect 37772 43260 37828 43262
rect 37884 42924 37940 42980
rect 37884 42700 37940 42756
rect 37772 42028 37828 42084
rect 37772 40796 37828 40852
rect 38220 42700 38276 42756
rect 38108 42082 38164 42084
rect 38108 42030 38110 42082
rect 38110 42030 38162 42082
rect 38162 42030 38164 42082
rect 38108 42028 38164 42030
rect 38220 41970 38276 41972
rect 38220 41918 38222 41970
rect 38222 41918 38274 41970
rect 38274 41918 38276 41970
rect 38220 41916 38276 41918
rect 38108 41468 38164 41524
rect 37660 40572 37716 40628
rect 37212 40124 37268 40180
rect 37324 39116 37380 39172
rect 36988 38892 37044 38948
rect 36316 37996 36372 38052
rect 36092 37100 36148 37156
rect 36540 37212 36596 37268
rect 35980 36316 36036 36372
rect 35868 36092 35924 36148
rect 36764 37266 36820 37268
rect 36764 37214 36766 37266
rect 36766 37214 36818 37266
rect 36818 37214 36820 37266
rect 36764 37212 36820 37214
rect 36764 36988 36820 37044
rect 36540 36316 36596 36372
rect 35980 34972 36036 35028
rect 35868 34188 35924 34244
rect 36092 34188 36148 34244
rect 35868 32620 35924 32676
rect 35868 32396 35924 32452
rect 35756 31276 35812 31332
rect 36092 33852 36148 33908
rect 35532 29932 35588 29988
rect 35644 30156 35700 30212
rect 35532 29484 35588 29540
rect 36540 35420 36596 35476
rect 36540 34412 36596 34468
rect 36316 33964 36372 34020
rect 36876 34636 36932 34692
rect 36764 34188 36820 34244
rect 36876 33852 36932 33908
rect 37884 40124 37940 40180
rect 38220 41132 38276 41188
rect 37660 39228 37716 39284
rect 37884 38892 37940 38948
rect 38556 46396 38612 46452
rect 38780 46396 38836 46452
rect 39564 54402 39620 54404
rect 39564 54350 39566 54402
rect 39566 54350 39618 54402
rect 39618 54350 39620 54402
rect 39564 54348 39620 54350
rect 39452 53788 39508 53844
rect 39900 52556 39956 52612
rect 39228 51324 39284 51380
rect 39340 51660 39396 51716
rect 39116 51212 39172 51268
rect 39228 51154 39284 51156
rect 39228 51102 39230 51154
rect 39230 51102 39282 51154
rect 39282 51102 39284 51154
rect 39228 51100 39284 51102
rect 39004 48412 39060 48468
rect 39116 50540 39172 50596
rect 39228 49980 39284 50036
rect 39564 50594 39620 50596
rect 39564 50542 39566 50594
rect 39566 50542 39618 50594
rect 39618 50542 39620 50594
rect 39564 50540 39620 50542
rect 39340 49644 39396 49700
rect 39676 49586 39732 49588
rect 39676 49534 39678 49586
rect 39678 49534 39730 49586
rect 39730 49534 39732 49586
rect 39676 49532 39732 49534
rect 39676 49250 39732 49252
rect 39676 49198 39678 49250
rect 39678 49198 39730 49250
rect 39730 49198 39732 49250
rect 39676 49196 39732 49198
rect 40236 52108 40292 52164
rect 40124 51154 40180 51156
rect 40124 51102 40126 51154
rect 40126 51102 40178 51154
rect 40178 51102 40180 51154
rect 40124 51100 40180 51102
rect 40236 50764 40292 50820
rect 40796 57036 40852 57092
rect 40572 55410 40628 55412
rect 40572 55358 40574 55410
rect 40574 55358 40626 55410
rect 40626 55358 40628 55410
rect 40572 55356 40628 55358
rect 40460 54572 40516 54628
rect 40460 54290 40516 54292
rect 40460 54238 40462 54290
rect 40462 54238 40514 54290
rect 40514 54238 40516 54290
rect 40460 54236 40516 54238
rect 41020 56924 41076 56980
rect 41020 56476 41076 56532
rect 41132 55804 41188 55860
rect 41132 55410 41188 55412
rect 41132 55358 41134 55410
rect 41134 55358 41186 55410
rect 41186 55358 41188 55410
rect 41132 55356 41188 55358
rect 41692 57260 41748 57316
rect 41468 55580 41524 55636
rect 41244 54684 41300 54740
rect 40908 54012 40964 54068
rect 40460 53452 40516 53508
rect 40460 51324 40516 51380
rect 40348 50594 40404 50596
rect 40348 50542 40350 50594
rect 40350 50542 40402 50594
rect 40402 50542 40404 50594
rect 40348 50540 40404 50542
rect 40460 49532 40516 49588
rect 41132 53340 41188 53396
rect 40908 52274 40964 52276
rect 40908 52222 40910 52274
rect 40910 52222 40962 52274
rect 40962 52222 40964 52274
rect 40908 52220 40964 52222
rect 40684 51996 40740 52052
rect 41580 54796 41636 54852
rect 41244 52220 41300 52276
rect 41244 51996 41300 52052
rect 41132 51266 41188 51268
rect 41132 51214 41134 51266
rect 41134 51214 41186 51266
rect 41186 51214 41188 51266
rect 41132 51212 41188 51214
rect 40684 51100 40740 51156
rect 41244 51100 41300 51156
rect 40572 49196 40628 49252
rect 40348 49026 40404 49028
rect 40348 48974 40350 49026
rect 40350 48974 40402 49026
rect 40402 48974 40404 49026
rect 40348 48972 40404 48974
rect 39900 48300 39956 48356
rect 40460 48636 40516 48692
rect 39452 47628 39508 47684
rect 39676 48076 39732 48132
rect 39004 47180 39060 47236
rect 39004 46060 39060 46116
rect 39340 46396 39396 46452
rect 38668 44716 38724 44772
rect 38780 45276 38836 45332
rect 39340 45388 39396 45444
rect 38892 45164 38948 45220
rect 38668 44434 38724 44436
rect 38668 44382 38670 44434
rect 38670 44382 38722 44434
rect 38722 44382 38724 44434
rect 38668 44380 38724 44382
rect 39564 47458 39620 47460
rect 39564 47406 39566 47458
rect 39566 47406 39618 47458
rect 39618 47406 39620 47458
rect 39564 47404 39620 47406
rect 39564 45836 39620 45892
rect 40124 47628 40180 47684
rect 39788 45890 39844 45892
rect 39788 45838 39790 45890
rect 39790 45838 39842 45890
rect 39842 45838 39844 45890
rect 39788 45836 39844 45838
rect 39676 45500 39732 45556
rect 39900 45276 39956 45332
rect 39788 45052 39844 45108
rect 39116 44828 39172 44884
rect 39004 43820 39060 43876
rect 38892 43314 38948 43316
rect 38892 43262 38894 43314
rect 38894 43262 38946 43314
rect 38946 43262 38948 43314
rect 38892 43260 38948 43262
rect 38556 43148 38612 43204
rect 38780 43148 38836 43204
rect 38668 42754 38724 42756
rect 38668 42702 38670 42754
rect 38670 42702 38722 42754
rect 38722 42702 38724 42754
rect 38668 42700 38724 42702
rect 38668 42252 38724 42308
rect 38556 41970 38612 41972
rect 38556 41918 38558 41970
rect 38558 41918 38610 41970
rect 38610 41918 38612 41970
rect 38556 41916 38612 41918
rect 38444 41020 38500 41076
rect 38780 41692 38836 41748
rect 38444 40012 38500 40068
rect 38780 40402 38836 40404
rect 38780 40350 38782 40402
rect 38782 40350 38834 40402
rect 38834 40350 38836 40402
rect 38780 40348 38836 40350
rect 39228 44044 39284 44100
rect 39340 43820 39396 43876
rect 39340 43426 39396 43428
rect 39340 43374 39342 43426
rect 39342 43374 39394 43426
rect 39394 43374 39396 43426
rect 39340 43372 39396 43374
rect 39228 42924 39284 42980
rect 39004 40124 39060 40180
rect 40012 45218 40068 45220
rect 40012 45166 40014 45218
rect 40014 45166 40066 45218
rect 40066 45166 40068 45218
rect 40012 45164 40068 45166
rect 40236 47458 40292 47460
rect 40236 47406 40238 47458
rect 40238 47406 40290 47458
rect 40290 47406 40292 47458
rect 40236 47404 40292 47406
rect 40348 47346 40404 47348
rect 40348 47294 40350 47346
rect 40350 47294 40402 47346
rect 40402 47294 40404 47346
rect 40348 47292 40404 47294
rect 40908 49420 40964 49476
rect 40908 48860 40964 48916
rect 40796 47458 40852 47460
rect 40796 47406 40798 47458
rect 40798 47406 40850 47458
rect 40850 47406 40852 47458
rect 40796 47404 40852 47406
rect 40124 45052 40180 45108
rect 40012 44828 40068 44884
rect 39788 44044 39844 44100
rect 39676 43820 39732 43876
rect 39564 43036 39620 43092
rect 39900 44380 39956 44436
rect 39676 42812 39732 42868
rect 39788 42924 39844 42980
rect 39676 42364 39732 42420
rect 39564 42252 39620 42308
rect 39788 41916 39844 41972
rect 39676 41746 39732 41748
rect 39676 41694 39678 41746
rect 39678 41694 39730 41746
rect 39730 41694 39732 41746
rect 39676 41692 39732 41694
rect 39564 40962 39620 40964
rect 39564 40910 39566 40962
rect 39566 40910 39618 40962
rect 39618 40910 39620 40962
rect 39564 40908 39620 40910
rect 39452 40796 39508 40852
rect 39564 40402 39620 40404
rect 39564 40350 39566 40402
rect 39566 40350 39618 40402
rect 39618 40350 39620 40402
rect 39564 40348 39620 40350
rect 38668 39676 38724 39732
rect 39228 40012 39284 40068
rect 38556 39228 38612 39284
rect 38444 38892 38500 38948
rect 38444 38668 38500 38724
rect 37884 38108 37940 38164
rect 37548 37324 37604 37380
rect 37212 37212 37268 37268
rect 37436 36482 37492 36484
rect 37436 36430 37438 36482
rect 37438 36430 37490 36482
rect 37490 36430 37492 36482
rect 37436 36428 37492 36430
rect 37548 35420 37604 35476
rect 37660 37212 37716 37268
rect 37324 34412 37380 34468
rect 37436 34018 37492 34020
rect 37436 33966 37438 34018
rect 37438 33966 37490 34018
rect 37490 33966 37492 34018
rect 37436 33964 37492 33966
rect 37212 33906 37268 33908
rect 37212 33854 37214 33906
rect 37214 33854 37266 33906
rect 37266 33854 37268 33906
rect 37212 33852 37268 33854
rect 36652 33068 36708 33124
rect 36652 32620 36708 32676
rect 36876 32620 36932 32676
rect 36764 32396 36820 32452
rect 36316 31666 36372 31668
rect 36316 31614 36318 31666
rect 36318 31614 36370 31666
rect 36370 31614 36372 31666
rect 36316 31612 36372 31614
rect 36204 30716 36260 30772
rect 36092 30156 36148 30212
rect 36316 30156 36372 30212
rect 36428 30268 36484 30324
rect 37100 30940 37156 30996
rect 36652 30828 36708 30884
rect 36988 30770 37044 30772
rect 36988 30718 36990 30770
rect 36990 30718 37042 30770
rect 37042 30718 37044 30770
rect 36988 30716 37044 30718
rect 37324 33628 37380 33684
rect 37884 36316 37940 36372
rect 38220 36540 38276 36596
rect 37996 36092 38052 36148
rect 37772 34188 37828 34244
rect 37884 33852 37940 33908
rect 37660 33404 37716 33460
rect 37324 32060 37380 32116
rect 37436 32508 37492 32564
rect 37548 32338 37604 32340
rect 37548 32286 37550 32338
rect 37550 32286 37602 32338
rect 37602 32286 37604 32338
rect 37548 32284 37604 32286
rect 37436 31164 37492 31220
rect 37772 33628 37828 33684
rect 37324 30940 37380 30996
rect 36540 29596 36596 29652
rect 36204 29484 36260 29540
rect 35868 28812 35924 28868
rect 35532 28642 35588 28644
rect 35532 28590 35534 28642
rect 35534 28590 35586 28642
rect 35586 28590 35588 28642
rect 35532 28588 35588 28590
rect 35420 28364 35476 28420
rect 35756 28476 35812 28532
rect 34748 26908 34804 26964
rect 35196 28028 35252 28084
rect 35196 27858 35252 27860
rect 35196 27806 35198 27858
rect 35198 27806 35250 27858
rect 35250 27806 35252 27858
rect 35196 27804 35252 27806
rect 35420 27580 35476 27636
rect 35532 27356 35588 27412
rect 35196 27186 35252 27188
rect 35196 27134 35198 27186
rect 35198 27134 35250 27186
rect 35250 27134 35252 27186
rect 35196 27132 35252 27134
rect 34860 26796 34916 26852
rect 35868 27468 35924 27524
rect 35756 26908 35812 26964
rect 35644 26796 35700 26852
rect 34412 26236 34468 26292
rect 35420 26460 35476 26516
rect 35308 26236 35364 26292
rect 34524 25228 34580 25284
rect 34860 25618 34916 25620
rect 34860 25566 34862 25618
rect 34862 25566 34914 25618
rect 34914 25566 34916 25618
rect 34860 25564 34916 25566
rect 34860 25340 34916 25396
rect 34412 24610 34468 24612
rect 34412 24558 34414 24610
rect 34414 24558 34466 24610
rect 34466 24558 34468 24610
rect 34412 24556 34468 24558
rect 34300 23884 34356 23940
rect 34412 24332 34468 24388
rect 34300 22876 34356 22932
rect 33964 22092 34020 22148
rect 33964 21756 34020 21812
rect 33852 20524 33908 20580
rect 33852 17052 33908 17108
rect 34748 24668 34804 24724
rect 34524 23212 34580 23268
rect 34636 23548 34692 23604
rect 34636 22764 34692 22820
rect 35196 26066 35252 26068
rect 35196 26014 35198 26066
rect 35198 26014 35250 26066
rect 35250 26014 35252 26066
rect 35196 26012 35252 26014
rect 35084 25452 35140 25508
rect 35196 25788 35252 25844
rect 35308 25676 35364 25732
rect 35420 25564 35476 25620
rect 36316 28252 36372 28308
rect 36764 29148 36820 29204
rect 36652 28924 36708 28980
rect 36876 28924 36932 28980
rect 36092 26572 36148 26628
rect 37212 29932 37268 29988
rect 37324 29596 37380 29652
rect 37212 28754 37268 28756
rect 37212 28702 37214 28754
rect 37214 28702 37266 28754
rect 37266 28702 37268 28754
rect 37212 28700 37268 28702
rect 36764 28252 36820 28308
rect 34972 25004 35028 25060
rect 35980 26124 36036 26180
rect 36092 25788 36148 25844
rect 35196 24668 35252 24724
rect 35308 23100 35364 23156
rect 36540 27356 36596 27412
rect 36540 26236 36596 26292
rect 36652 26178 36708 26180
rect 36652 26126 36654 26178
rect 36654 26126 36706 26178
rect 36706 26126 36708 26178
rect 36652 26124 36708 26126
rect 36988 28252 37044 28308
rect 36876 28028 36932 28084
rect 36316 25788 36372 25844
rect 36540 25730 36596 25732
rect 36540 25678 36542 25730
rect 36542 25678 36594 25730
rect 36594 25678 36596 25730
rect 36540 25676 36596 25678
rect 36764 25564 36820 25620
rect 36540 25452 36596 25508
rect 36428 25394 36484 25396
rect 36428 25342 36430 25394
rect 36430 25342 36482 25394
rect 36482 25342 36484 25394
rect 36428 25340 36484 25342
rect 36540 24834 36596 24836
rect 36540 24782 36542 24834
rect 36542 24782 36594 24834
rect 36594 24782 36596 24834
rect 36540 24780 36596 24782
rect 36764 24780 36820 24836
rect 36316 24668 36372 24724
rect 36204 24220 36260 24276
rect 35644 23996 35700 24052
rect 35308 22876 35364 22932
rect 35196 22764 35252 22820
rect 34860 22370 34916 22372
rect 34860 22318 34862 22370
rect 34862 22318 34914 22370
rect 34914 22318 34916 22370
rect 34860 22316 34916 22318
rect 34412 20802 34468 20804
rect 34412 20750 34414 20802
rect 34414 20750 34466 20802
rect 34466 20750 34468 20802
rect 34412 20748 34468 20750
rect 34300 20300 34356 20356
rect 34860 20748 34916 20804
rect 34300 19794 34356 19796
rect 34300 19742 34302 19794
rect 34302 19742 34354 19794
rect 34354 19742 34356 19794
rect 34300 19740 34356 19742
rect 34972 19852 35028 19908
rect 34188 19180 34244 19236
rect 34860 18956 34916 19012
rect 34188 18732 34244 18788
rect 34860 18732 34916 18788
rect 34300 18562 34356 18564
rect 34300 18510 34302 18562
rect 34302 18510 34354 18562
rect 34354 18510 34356 18562
rect 34300 18508 34356 18510
rect 34412 18450 34468 18452
rect 34412 18398 34414 18450
rect 34414 18398 34466 18450
rect 34466 18398 34468 18450
rect 34412 18396 34468 18398
rect 35420 21868 35476 21924
rect 35532 21756 35588 21812
rect 35308 20412 35364 20468
rect 35308 20076 35364 20132
rect 35532 19740 35588 19796
rect 35980 20748 36036 20804
rect 35308 19292 35364 19348
rect 34188 17836 34244 17892
rect 35196 17948 35252 18004
rect 34076 17052 34132 17108
rect 35084 17890 35140 17892
rect 35084 17838 35086 17890
rect 35086 17838 35138 17890
rect 35138 17838 35140 17890
rect 35084 17836 35140 17838
rect 34636 17724 34692 17780
rect 34412 17500 34468 17556
rect 33740 15148 33796 15204
rect 33852 16156 33908 16212
rect 34188 16828 34244 16884
rect 34300 16658 34356 16660
rect 34300 16606 34302 16658
rect 34302 16606 34354 16658
rect 34354 16606 34356 16658
rect 34300 16604 34356 16606
rect 34300 16156 34356 16212
rect 34188 15874 34244 15876
rect 34188 15822 34190 15874
rect 34190 15822 34242 15874
rect 34242 15822 34244 15874
rect 34188 15820 34244 15822
rect 34524 16940 34580 16996
rect 34972 16940 35028 16996
rect 34972 15820 35028 15876
rect 33964 14476 34020 14532
rect 34748 15148 34804 15204
rect 33852 14252 33908 14308
rect 33292 14028 33348 14084
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 33180 13804 33236 13860
rect 33068 12908 33124 12964
rect 33068 12684 33124 12740
rect 32956 12124 33012 12180
rect 33292 13692 33348 13748
rect 34412 13580 34468 13636
rect 34636 13580 34692 13636
rect 33852 12236 33908 12292
rect 33180 10108 33236 10164
rect 33292 10332 33348 10388
rect 33068 9436 33124 9492
rect 33516 10386 33572 10388
rect 33516 10334 33518 10386
rect 33518 10334 33570 10386
rect 33570 10334 33572 10386
rect 33516 10332 33572 10334
rect 33292 9436 33348 9492
rect 32844 9042 32900 9044
rect 32844 8990 32846 9042
rect 32846 8990 32898 9042
rect 32898 8990 32900 9042
rect 32844 8988 32900 8990
rect 32732 8258 32788 8260
rect 32732 8206 32734 8258
rect 32734 8206 32786 8258
rect 32786 8206 32788 8258
rect 32732 8204 32788 8206
rect 32284 7868 32340 7924
rect 32844 7980 32900 8036
rect 32060 7756 32116 7812
rect 31948 7308 32004 7364
rect 31724 6466 31780 6468
rect 31724 6414 31726 6466
rect 31726 6414 31778 6466
rect 31778 6414 31780 6466
rect 31724 6412 31780 6414
rect 31724 4844 31780 4900
rect 31948 4844 32004 4900
rect 32284 5068 32340 5124
rect 32172 4732 32228 4788
rect 31612 4114 31668 4116
rect 31612 4062 31614 4114
rect 31614 4062 31666 4114
rect 31666 4062 31668 4114
rect 31612 4060 31668 4062
rect 32060 3724 32116 3780
rect 31948 2716 32004 2772
rect 31724 2546 31780 2548
rect 31724 2494 31726 2546
rect 31726 2494 31778 2546
rect 31778 2494 31780 2546
rect 31724 2492 31780 2494
rect 31276 1148 31332 1204
rect 31612 1596 31668 1652
rect 31724 1372 31780 1428
rect 32284 4172 32340 4228
rect 32508 7586 32564 7588
rect 32508 7534 32510 7586
rect 32510 7534 32562 7586
rect 32562 7534 32564 7586
rect 32508 7532 32564 7534
rect 32508 7084 32564 7140
rect 32508 6412 32564 6468
rect 32620 5740 32676 5796
rect 32732 5628 32788 5684
rect 32620 4338 32676 4340
rect 32620 4286 32622 4338
rect 32622 4286 32674 4338
rect 32674 4286 32676 4338
rect 32620 4284 32676 4286
rect 33180 8092 33236 8148
rect 33404 8540 33460 8596
rect 33516 8428 33572 8484
rect 33180 7308 33236 7364
rect 33068 6802 33124 6804
rect 33068 6750 33070 6802
rect 33070 6750 33122 6802
rect 33122 6750 33124 6802
rect 33068 6748 33124 6750
rect 33180 6578 33236 6580
rect 33180 6526 33182 6578
rect 33182 6526 33234 6578
rect 33234 6526 33236 6578
rect 33180 6524 33236 6526
rect 32844 5292 32900 5348
rect 32956 6076 33012 6132
rect 32732 4172 32788 4228
rect 32508 4060 32564 4116
rect 32172 2770 32228 2772
rect 32172 2718 32174 2770
rect 32174 2718 32226 2770
rect 32226 2718 32228 2770
rect 32172 2716 32228 2718
rect 32284 3612 32340 3668
rect 32284 2380 32340 2436
rect 32732 3666 32788 3668
rect 32732 3614 32734 3666
rect 32734 3614 32786 3666
rect 32786 3614 32788 3666
rect 32732 3612 32788 3614
rect 33068 5682 33124 5684
rect 33068 5630 33070 5682
rect 33070 5630 33122 5682
rect 33122 5630 33124 5682
rect 33068 5628 33124 5630
rect 33068 5404 33124 5460
rect 33292 6300 33348 6356
rect 33292 5404 33348 5460
rect 33964 12178 34020 12180
rect 33964 12126 33966 12178
rect 33966 12126 34018 12178
rect 34018 12126 34020 12178
rect 33964 12124 34020 12126
rect 34300 10108 34356 10164
rect 34188 8316 34244 8372
rect 33852 7980 33908 8036
rect 33516 7532 33572 7588
rect 33516 6972 33572 7028
rect 33516 6578 33572 6580
rect 33516 6526 33518 6578
rect 33518 6526 33570 6578
rect 33570 6526 33572 6578
rect 33516 6524 33572 6526
rect 34188 6578 34244 6580
rect 34188 6526 34190 6578
rect 34190 6526 34242 6578
rect 34242 6526 34244 6578
rect 34188 6524 34244 6526
rect 34188 6130 34244 6132
rect 34188 6078 34190 6130
rect 34190 6078 34242 6130
rect 34242 6078 34244 6130
rect 34188 6076 34244 6078
rect 34524 11116 34580 11172
rect 34748 11452 34804 11508
rect 34412 9996 34468 10052
rect 34412 9660 34468 9716
rect 34524 10108 34580 10164
rect 34412 8258 34468 8260
rect 34412 8206 34414 8258
rect 34414 8206 34466 8258
rect 34466 8206 34468 8258
rect 34412 8204 34468 8206
rect 34636 9826 34692 9828
rect 34636 9774 34638 9826
rect 34638 9774 34690 9826
rect 34690 9774 34692 9826
rect 34636 9772 34692 9774
rect 34636 8540 34692 8596
rect 34524 6972 34580 7028
rect 34300 5628 34356 5684
rect 34524 6076 34580 6132
rect 33740 5346 33796 5348
rect 33740 5294 33742 5346
rect 33742 5294 33794 5346
rect 33794 5294 33796 5346
rect 33740 5292 33796 5294
rect 34860 14476 34916 14532
rect 34972 14252 35028 14308
rect 35084 12572 35140 12628
rect 34972 12236 35028 12292
rect 34972 11900 35028 11956
rect 35980 18508 36036 18564
rect 35420 18338 35476 18340
rect 35420 18286 35422 18338
rect 35422 18286 35474 18338
rect 35474 18286 35476 18338
rect 35420 18284 35476 18286
rect 35756 18284 35812 18340
rect 35532 16940 35588 16996
rect 35756 15820 35812 15876
rect 36428 23826 36484 23828
rect 36428 23774 36430 23826
rect 36430 23774 36482 23826
rect 36482 23774 36484 23826
rect 36428 23772 36484 23774
rect 36652 23772 36708 23828
rect 36316 23266 36372 23268
rect 36316 23214 36318 23266
rect 36318 23214 36370 23266
rect 36370 23214 36372 23266
rect 36316 23212 36372 23214
rect 36428 22930 36484 22932
rect 36428 22878 36430 22930
rect 36430 22878 36482 22930
rect 36482 22878 36484 22930
rect 36428 22876 36484 22878
rect 36764 23660 36820 23716
rect 36652 23154 36708 23156
rect 36652 23102 36654 23154
rect 36654 23102 36706 23154
rect 36706 23102 36708 23154
rect 36652 23100 36708 23102
rect 36204 21532 36260 21588
rect 36204 20690 36260 20692
rect 36204 20638 36206 20690
rect 36206 20638 36258 20690
rect 36258 20638 36260 20690
rect 36204 20636 36260 20638
rect 36428 21084 36484 21140
rect 37100 27356 37156 27412
rect 36988 25506 37044 25508
rect 36988 25454 36990 25506
rect 36990 25454 37042 25506
rect 37042 25454 37044 25506
rect 36988 25452 37044 25454
rect 36988 24108 37044 24164
rect 36876 23212 36932 23268
rect 37212 26236 37268 26292
rect 38220 34972 38276 35028
rect 38220 34412 38276 34468
rect 38108 34188 38164 34244
rect 38108 33740 38164 33796
rect 38668 38892 38724 38948
rect 39228 39676 39284 39732
rect 39452 40236 39508 40292
rect 38892 37884 38948 37940
rect 38780 35532 38836 35588
rect 39116 35644 39172 35700
rect 38668 35196 38724 35252
rect 38444 35084 38500 35140
rect 38332 34188 38388 34244
rect 38780 34748 38836 34804
rect 38444 33740 38500 33796
rect 38892 34524 38948 34580
rect 39004 34130 39060 34132
rect 39004 34078 39006 34130
rect 39006 34078 39058 34130
rect 39058 34078 39060 34130
rect 39004 34076 39060 34078
rect 39004 33852 39060 33908
rect 38892 33740 38948 33796
rect 37996 32674 38052 32676
rect 37996 32622 37998 32674
rect 37998 32622 38050 32674
rect 38050 32622 38052 32674
rect 37996 32620 38052 32622
rect 37884 31388 37940 31444
rect 37996 31724 38052 31780
rect 37884 31164 37940 31220
rect 37884 30380 37940 30436
rect 37772 29986 37828 29988
rect 37772 29934 37774 29986
rect 37774 29934 37826 29986
rect 37826 29934 37828 29986
rect 37772 29932 37828 29934
rect 37660 29036 37716 29092
rect 37324 25452 37380 25508
rect 37548 25618 37604 25620
rect 37548 25566 37550 25618
rect 37550 25566 37602 25618
rect 37602 25566 37604 25618
rect 37548 25564 37604 25566
rect 37324 24668 37380 24724
rect 37212 23436 37268 23492
rect 37100 23212 37156 23268
rect 37212 23154 37268 23156
rect 37212 23102 37214 23154
rect 37214 23102 37266 23154
rect 37266 23102 37268 23154
rect 37212 23100 37268 23102
rect 37100 22652 37156 22708
rect 37436 23884 37492 23940
rect 37660 24668 37716 24724
rect 37660 24332 37716 24388
rect 37660 23772 37716 23828
rect 37548 22316 37604 22372
rect 37436 22092 37492 22148
rect 36764 21756 36820 21812
rect 36652 21026 36708 21028
rect 36652 20974 36654 21026
rect 36654 20974 36706 21026
rect 36706 20974 36708 21026
rect 36652 20972 36708 20974
rect 36540 20636 36596 20692
rect 36540 18508 36596 18564
rect 36316 18338 36372 18340
rect 36316 18286 36318 18338
rect 36318 18286 36370 18338
rect 36370 18286 36372 18338
rect 36316 18284 36372 18286
rect 36204 16716 36260 16772
rect 36316 17388 36372 17444
rect 35756 15036 35812 15092
rect 35980 15036 36036 15092
rect 36092 14812 36148 14868
rect 35532 14476 35588 14532
rect 35308 14028 35364 14084
rect 35420 14252 35476 14308
rect 35308 11564 35364 11620
rect 35532 13244 35588 13300
rect 35644 11564 35700 11620
rect 35084 9772 35140 9828
rect 34860 7420 34916 7476
rect 34748 6802 34804 6804
rect 34748 6750 34750 6802
rect 34750 6750 34802 6802
rect 34802 6750 34804 6802
rect 34748 6748 34804 6750
rect 35196 6748 35252 6804
rect 34748 6300 34804 6356
rect 35196 6412 35252 6468
rect 36316 13580 36372 13636
rect 36540 15372 36596 15428
rect 37100 20018 37156 20020
rect 37100 19966 37102 20018
rect 37102 19966 37154 20018
rect 37154 19966 37156 20018
rect 37100 19964 37156 19966
rect 36988 19234 37044 19236
rect 36988 19182 36990 19234
rect 36990 19182 37042 19234
rect 37042 19182 37044 19234
rect 36988 19180 37044 19182
rect 36988 18508 37044 18564
rect 37884 28700 37940 28756
rect 37884 26402 37940 26404
rect 37884 26350 37886 26402
rect 37886 26350 37938 26402
rect 37938 26350 37940 26402
rect 37884 26348 37940 26350
rect 37884 24780 37940 24836
rect 38220 32508 38276 32564
rect 39228 35308 39284 35364
rect 39788 39116 39844 39172
rect 39676 38946 39732 38948
rect 39676 38894 39678 38946
rect 39678 38894 39730 38946
rect 39730 38894 39732 38946
rect 39676 38892 39732 38894
rect 40348 46284 40404 46340
rect 40684 45500 40740 45556
rect 40236 44380 40292 44436
rect 40348 43820 40404 43876
rect 40236 43372 40292 43428
rect 40460 43426 40516 43428
rect 40460 43374 40462 43426
rect 40462 43374 40514 43426
rect 40514 43374 40516 43426
rect 40460 43372 40516 43374
rect 40796 44828 40852 44884
rect 41580 53340 41636 53396
rect 41580 52220 41636 52276
rect 42140 56588 42196 56644
rect 42364 56028 42420 56084
rect 41916 55468 41972 55524
rect 41804 54908 41860 54964
rect 41916 54348 41972 54404
rect 42028 54796 42084 54852
rect 43708 57260 43764 57316
rect 43260 56364 43316 56420
rect 43484 56924 43540 56980
rect 42812 55580 42868 55636
rect 42588 55132 42644 55188
rect 42364 54908 42420 54964
rect 42140 54572 42196 54628
rect 41804 54290 41860 54292
rect 41804 54238 41806 54290
rect 41806 54238 41858 54290
rect 41858 54238 41860 54290
rect 41804 54236 41860 54238
rect 42140 53676 42196 53732
rect 41804 52892 41860 52948
rect 41804 52722 41860 52724
rect 41804 52670 41806 52722
rect 41806 52670 41858 52722
rect 41858 52670 41860 52722
rect 41804 52668 41860 52670
rect 41580 50988 41636 51044
rect 41468 50540 41524 50596
rect 41916 51324 41972 51380
rect 41804 49196 41860 49252
rect 42700 54514 42756 54516
rect 42700 54462 42702 54514
rect 42702 54462 42754 54514
rect 42754 54462 42756 54514
rect 42700 54460 42756 54462
rect 42812 54124 42868 54180
rect 42700 53452 42756 53508
rect 42140 51436 42196 51492
rect 42476 51324 42532 51380
rect 42700 51602 42756 51604
rect 42700 51550 42702 51602
rect 42702 51550 42754 51602
rect 42754 51550 42756 51602
rect 42700 51548 42756 51550
rect 43036 54124 43092 54180
rect 44380 56588 44436 56644
rect 43596 56476 43652 56532
rect 45052 56812 45108 56868
rect 45276 56812 45332 56868
rect 45164 56700 45220 56756
rect 43804 56474 43860 56476
rect 43804 56422 43806 56474
rect 43806 56422 43858 56474
rect 43858 56422 43860 56474
rect 43804 56420 43860 56422
rect 43908 56474 43964 56476
rect 43908 56422 43910 56474
rect 43910 56422 43962 56474
rect 43962 56422 43964 56474
rect 43908 56420 43964 56422
rect 44012 56474 44068 56476
rect 44012 56422 44014 56474
rect 44014 56422 44066 56474
rect 44066 56422 44068 56474
rect 44012 56420 44068 56422
rect 44156 56364 44212 56420
rect 43820 56252 43876 56308
rect 44716 56252 44772 56308
rect 44268 56140 44324 56196
rect 44492 55858 44548 55860
rect 44492 55806 44494 55858
rect 44494 55806 44546 55858
rect 44546 55806 44548 55858
rect 44492 55804 44548 55806
rect 44828 55858 44884 55860
rect 44828 55806 44830 55858
rect 44830 55806 44882 55858
rect 44882 55806 44884 55858
rect 44828 55804 44884 55806
rect 44464 55690 44520 55692
rect 43596 55580 43652 55636
rect 44268 55580 44324 55636
rect 44464 55638 44466 55690
rect 44466 55638 44518 55690
rect 44518 55638 44520 55690
rect 44464 55636 44520 55638
rect 44568 55690 44624 55692
rect 44568 55638 44570 55690
rect 44570 55638 44622 55690
rect 44622 55638 44624 55690
rect 44568 55636 44624 55638
rect 44672 55690 44728 55692
rect 44672 55638 44674 55690
rect 44674 55638 44726 55690
rect 44726 55638 44728 55690
rect 44672 55636 44728 55638
rect 45276 56140 45332 56196
rect 45500 56140 45556 56196
rect 45836 56082 45892 56084
rect 45836 56030 45838 56082
rect 45838 56030 45890 56082
rect 45890 56030 45892 56082
rect 45836 56028 45892 56030
rect 43484 55522 43540 55524
rect 43484 55470 43486 55522
rect 43486 55470 43538 55522
rect 43538 55470 43540 55522
rect 43484 55468 43540 55470
rect 44940 55580 44996 55636
rect 43820 55244 43876 55300
rect 44156 55298 44212 55300
rect 44156 55246 44158 55298
rect 44158 55246 44210 55298
rect 44210 55246 44212 55298
rect 44156 55244 44212 55246
rect 44492 55410 44548 55412
rect 44492 55358 44494 55410
rect 44494 55358 44546 55410
rect 44546 55358 44548 55410
rect 44492 55356 44548 55358
rect 46172 57260 46228 57316
rect 46284 56476 46340 56532
rect 45948 55580 46004 55636
rect 44380 55244 44436 55300
rect 43260 55020 43316 55076
rect 43596 54908 43652 54964
rect 43804 54906 43860 54908
rect 43804 54854 43806 54906
rect 43806 54854 43858 54906
rect 43858 54854 43860 54906
rect 43804 54852 43860 54854
rect 43908 54906 43964 54908
rect 43908 54854 43910 54906
rect 43910 54854 43962 54906
rect 43962 54854 43964 54906
rect 43908 54852 43964 54854
rect 44012 54906 44068 54908
rect 44012 54854 44014 54906
rect 44014 54854 44066 54906
rect 44066 54854 44068 54906
rect 44156 54908 44212 54964
rect 44012 54852 44068 54854
rect 44268 54796 44324 54852
rect 43148 53842 43204 53844
rect 43148 53790 43150 53842
rect 43150 53790 43202 53842
rect 43202 53790 43204 53842
rect 43148 53788 43204 53790
rect 43372 53676 43428 53732
rect 43260 53564 43316 53620
rect 42924 53004 42980 53060
rect 43372 52668 43428 52724
rect 43036 52220 43092 52276
rect 44492 54514 44548 54516
rect 44492 54462 44494 54514
rect 44494 54462 44546 54514
rect 44546 54462 44548 54514
rect 44492 54460 44548 54462
rect 44716 54290 44772 54292
rect 44716 54238 44718 54290
rect 44718 54238 44770 54290
rect 44770 54238 44772 54290
rect 44716 54236 44772 54238
rect 44464 54122 44520 54124
rect 44464 54070 44466 54122
rect 44466 54070 44518 54122
rect 44518 54070 44520 54122
rect 44464 54068 44520 54070
rect 44568 54122 44624 54124
rect 44568 54070 44570 54122
rect 44570 54070 44622 54122
rect 44622 54070 44624 54122
rect 44568 54068 44624 54070
rect 44672 54122 44728 54124
rect 44672 54070 44674 54122
rect 44674 54070 44726 54122
rect 44726 54070 44728 54122
rect 44672 54068 44728 54070
rect 45388 54796 45444 54852
rect 45724 54908 45780 54964
rect 44940 54684 44996 54740
rect 46060 55132 46116 55188
rect 45948 54908 46004 54964
rect 46060 54684 46116 54740
rect 45388 54402 45444 54404
rect 45388 54350 45390 54402
rect 45390 54350 45442 54402
rect 45442 54350 45444 54402
rect 45388 54348 45444 54350
rect 44604 53676 44660 53732
rect 43804 53338 43860 53340
rect 43804 53286 43806 53338
rect 43806 53286 43858 53338
rect 43858 53286 43860 53338
rect 43804 53284 43860 53286
rect 43908 53338 43964 53340
rect 43908 53286 43910 53338
rect 43910 53286 43962 53338
rect 43962 53286 43964 53338
rect 43908 53284 43964 53286
rect 44012 53338 44068 53340
rect 44012 53286 44014 53338
rect 44014 53286 44066 53338
rect 44066 53286 44068 53338
rect 44380 53340 44436 53396
rect 44492 53452 44548 53508
rect 44012 53284 44068 53286
rect 43820 53116 43876 53172
rect 43932 52892 43988 52948
rect 44828 53116 44884 53172
rect 44464 52554 44520 52556
rect 44464 52502 44466 52554
rect 44466 52502 44518 52554
rect 44518 52502 44520 52554
rect 44464 52500 44520 52502
rect 44568 52554 44624 52556
rect 44568 52502 44570 52554
rect 44570 52502 44622 52554
rect 44622 52502 44624 52554
rect 44568 52500 44624 52502
rect 44672 52554 44728 52556
rect 44672 52502 44674 52554
rect 44674 52502 44726 52554
rect 44726 52502 44728 52554
rect 44672 52500 44728 52502
rect 44156 52444 44212 52500
rect 43596 52332 43652 52388
rect 43260 52050 43316 52052
rect 43260 51998 43262 52050
rect 43262 51998 43314 52050
rect 43314 51998 43316 52050
rect 43260 51996 43316 51998
rect 43260 51602 43316 51604
rect 43260 51550 43262 51602
rect 43262 51550 43314 51602
rect 43314 51550 43316 51602
rect 43260 51548 43316 51550
rect 42364 49756 42420 49812
rect 42140 49698 42196 49700
rect 42140 49646 42142 49698
rect 42142 49646 42194 49698
rect 42194 49646 42196 49698
rect 42140 49644 42196 49646
rect 41692 48972 41748 49028
rect 41356 48860 41412 48916
rect 41580 48860 41636 48916
rect 41244 48188 41300 48244
rect 41020 48076 41076 48132
rect 41132 46450 41188 46452
rect 41132 46398 41134 46450
rect 41134 46398 41186 46450
rect 41186 46398 41188 46450
rect 41132 46396 41188 46398
rect 41356 47682 41412 47684
rect 41356 47630 41358 47682
rect 41358 47630 41410 47682
rect 41410 47630 41412 47682
rect 41356 47628 41412 47630
rect 41244 46060 41300 46116
rect 41356 45052 41412 45108
rect 41020 44882 41076 44884
rect 41020 44830 41022 44882
rect 41022 44830 41074 44882
rect 41074 44830 41076 44882
rect 41020 44828 41076 44830
rect 41244 44604 41300 44660
rect 40908 44380 40964 44436
rect 41020 43708 41076 43764
rect 40348 41916 40404 41972
rect 40236 41356 40292 41412
rect 40236 40796 40292 40852
rect 40124 40012 40180 40068
rect 40236 39730 40292 39732
rect 40236 39678 40238 39730
rect 40238 39678 40290 39730
rect 40290 39678 40292 39730
rect 40236 39676 40292 39678
rect 39788 38108 39844 38164
rect 39788 37212 39844 37268
rect 39788 35698 39844 35700
rect 39788 35646 39790 35698
rect 39790 35646 39842 35698
rect 39842 35646 39844 35698
rect 39788 35644 39844 35646
rect 40348 38892 40404 38948
rect 40012 38722 40068 38724
rect 40012 38670 40014 38722
rect 40014 38670 40066 38722
rect 40066 38670 40068 38722
rect 40012 38668 40068 38670
rect 40124 37324 40180 37380
rect 39900 35474 39956 35476
rect 39900 35422 39902 35474
rect 39902 35422 39954 35474
rect 39954 35422 39956 35474
rect 39900 35420 39956 35422
rect 39340 33628 39396 33684
rect 39228 32844 39284 32900
rect 39116 32732 39172 32788
rect 38780 32450 38836 32452
rect 38780 32398 38782 32450
rect 38782 32398 38834 32450
rect 38834 32398 38836 32450
rect 38780 32396 38836 32398
rect 38220 32172 38276 32228
rect 38108 31388 38164 31444
rect 38444 31276 38500 31332
rect 38220 30940 38276 30996
rect 38108 30770 38164 30772
rect 38108 30718 38110 30770
rect 38110 30718 38162 30770
rect 38162 30718 38164 30770
rect 38108 30716 38164 30718
rect 38444 30716 38500 30772
rect 38892 31836 38948 31892
rect 39116 32172 39172 32228
rect 38780 31388 38836 31444
rect 38332 29932 38388 29988
rect 39340 31778 39396 31780
rect 39340 31726 39342 31778
rect 39342 31726 39394 31778
rect 39394 31726 39396 31778
rect 39340 31724 39396 31726
rect 39228 30716 39284 30772
rect 38780 29708 38836 29764
rect 38780 29426 38836 29428
rect 38780 29374 38782 29426
rect 38782 29374 38834 29426
rect 38834 29374 38836 29426
rect 38780 29372 38836 29374
rect 38668 28700 38724 28756
rect 38780 28476 38836 28532
rect 38892 28364 38948 28420
rect 38332 27804 38388 27860
rect 38220 27132 38276 27188
rect 38108 26460 38164 26516
rect 38108 26124 38164 26180
rect 37996 24332 38052 24388
rect 37996 24108 38052 24164
rect 37772 21756 37828 21812
rect 38668 27298 38724 27300
rect 38668 27246 38670 27298
rect 38670 27246 38722 27298
rect 38722 27246 38724 27298
rect 38668 27244 38724 27246
rect 38556 26908 38612 26964
rect 38556 26572 38612 26628
rect 38332 26178 38388 26180
rect 38332 26126 38334 26178
rect 38334 26126 38386 26178
rect 38386 26126 38388 26178
rect 38332 26124 38388 26126
rect 38332 25228 38388 25284
rect 38444 23772 38500 23828
rect 37660 20972 37716 21028
rect 37772 21532 37828 21588
rect 38220 21868 38276 21924
rect 37548 20300 37604 20356
rect 37548 19458 37604 19460
rect 37548 19406 37550 19458
rect 37550 19406 37602 19458
rect 37602 19406 37604 19458
rect 37548 19404 37604 19406
rect 37100 18450 37156 18452
rect 37100 18398 37102 18450
rect 37102 18398 37154 18450
rect 37154 18398 37156 18450
rect 37100 18396 37156 18398
rect 37324 18338 37380 18340
rect 37324 18286 37326 18338
rect 37326 18286 37378 18338
rect 37378 18286 37380 18338
rect 37324 18284 37380 18286
rect 37100 17836 37156 17892
rect 37324 17890 37380 17892
rect 37324 17838 37326 17890
rect 37326 17838 37378 17890
rect 37378 17838 37380 17890
rect 37324 17836 37380 17838
rect 36988 16770 37044 16772
rect 36988 16718 36990 16770
rect 36990 16718 37042 16770
rect 37042 16718 37044 16770
rect 36988 16716 37044 16718
rect 37324 16044 37380 16100
rect 37548 18284 37604 18340
rect 37548 16380 37604 16436
rect 37100 15148 37156 15204
rect 36540 13356 36596 13412
rect 36764 13580 36820 13636
rect 36204 12796 36260 12852
rect 36204 12572 36260 12628
rect 35868 11564 35924 11620
rect 35756 10610 35812 10612
rect 35756 10558 35758 10610
rect 35758 10558 35810 10610
rect 35810 10558 35812 10610
rect 35756 10556 35812 10558
rect 35420 10220 35476 10276
rect 36316 11954 36372 11956
rect 36316 11902 36318 11954
rect 36318 11902 36370 11954
rect 36370 11902 36372 11954
rect 36316 11900 36372 11902
rect 35868 9996 35924 10052
rect 35644 9660 35700 9716
rect 35420 8092 35476 8148
rect 36316 9324 36372 9380
rect 35868 7420 35924 7476
rect 35420 6914 35476 6916
rect 35420 6862 35422 6914
rect 35422 6862 35474 6914
rect 35474 6862 35476 6914
rect 35420 6860 35476 6862
rect 35644 6802 35700 6804
rect 35644 6750 35646 6802
rect 35646 6750 35698 6802
rect 35698 6750 35700 6802
rect 35644 6748 35700 6750
rect 35532 6690 35588 6692
rect 35532 6638 35534 6690
rect 35534 6638 35586 6690
rect 35586 6638 35588 6690
rect 35532 6636 35588 6638
rect 35084 5852 35140 5908
rect 35420 5852 35476 5908
rect 34748 5292 34804 5348
rect 35084 5628 35140 5684
rect 33740 4338 33796 4340
rect 33740 4286 33742 4338
rect 33742 4286 33794 4338
rect 33794 4286 33796 4338
rect 33740 4284 33796 4286
rect 32956 2940 33012 2996
rect 33628 3948 33684 4004
rect 32956 2770 33012 2772
rect 32956 2718 32958 2770
rect 32958 2718 33010 2770
rect 33010 2718 33012 2770
rect 32956 2716 33012 2718
rect 33292 2492 33348 2548
rect 32956 2044 33012 2100
rect 32060 476 32116 532
rect 32508 140 32564 196
rect 33852 3724 33908 3780
rect 33740 2770 33796 2772
rect 33740 2718 33742 2770
rect 33742 2718 33794 2770
rect 33794 2718 33796 2770
rect 33740 2716 33796 2718
rect 33964 2268 34020 2324
rect 33852 1820 33908 1876
rect 33404 812 33460 868
rect 33516 252 33572 308
rect 34412 3612 34468 3668
rect 34300 2770 34356 2772
rect 34300 2718 34302 2770
rect 34302 2718 34354 2770
rect 34354 2718 34356 2770
rect 34300 2716 34356 2718
rect 35308 5292 35364 5348
rect 35308 4844 35364 4900
rect 35532 4956 35588 5012
rect 35084 2940 35140 2996
rect 35196 2770 35252 2772
rect 35196 2718 35198 2770
rect 35198 2718 35250 2770
rect 35250 2718 35252 2770
rect 35196 2716 35252 2718
rect 34188 2044 34244 2100
rect 34076 1708 34132 1764
rect 33964 1372 34020 1428
rect 35084 2210 35140 2212
rect 35084 2158 35086 2210
rect 35086 2158 35138 2210
rect 35138 2158 35140 2210
rect 35084 2156 35140 2158
rect 35868 6860 35924 6916
rect 36316 6972 36372 7028
rect 36316 6748 36372 6804
rect 36652 11676 36708 11732
rect 36540 11618 36596 11620
rect 36540 11566 36542 11618
rect 36542 11566 36594 11618
rect 36594 11566 36596 11618
rect 36540 11564 36596 11566
rect 36652 11394 36708 11396
rect 36652 11342 36654 11394
rect 36654 11342 36706 11394
rect 36706 11342 36708 11394
rect 36652 11340 36708 11342
rect 36764 10610 36820 10612
rect 36764 10558 36766 10610
rect 36766 10558 36818 10610
rect 36818 10558 36820 10610
rect 36764 10556 36820 10558
rect 35980 6076 36036 6132
rect 36428 6300 36484 6356
rect 37100 14252 37156 14308
rect 37100 13468 37156 13524
rect 37324 13244 37380 13300
rect 37436 15596 37492 15652
rect 37324 12962 37380 12964
rect 37324 12910 37326 12962
rect 37326 12910 37378 12962
rect 37378 12910 37380 12962
rect 37324 12908 37380 12910
rect 37100 11676 37156 11732
rect 37324 11116 37380 11172
rect 36876 9826 36932 9828
rect 36876 9774 36878 9826
rect 36878 9774 36930 9826
rect 36930 9774 36932 9826
rect 36876 9772 36932 9774
rect 36876 8092 36932 8148
rect 36540 6188 36596 6244
rect 36652 6972 36708 7028
rect 36428 5964 36484 6020
rect 36540 5906 36596 5908
rect 36540 5854 36542 5906
rect 36542 5854 36594 5906
rect 36594 5854 36596 5906
rect 36540 5852 36596 5854
rect 36764 5682 36820 5684
rect 36764 5630 36766 5682
rect 36766 5630 36818 5682
rect 36818 5630 36820 5682
rect 36764 5628 36820 5630
rect 35756 4732 35812 4788
rect 35756 4338 35812 4340
rect 35756 4286 35758 4338
rect 35758 4286 35810 4338
rect 35810 4286 35812 4338
rect 35756 4284 35812 4286
rect 36428 4338 36484 4340
rect 36428 4286 36430 4338
rect 36430 4286 36482 4338
rect 36482 4286 36484 4338
rect 36428 4284 36484 4286
rect 35644 3612 35700 3668
rect 35868 3666 35924 3668
rect 35868 3614 35870 3666
rect 35870 3614 35922 3666
rect 35922 3614 35924 3666
rect 35868 3612 35924 3614
rect 36652 3724 36708 3780
rect 35532 3500 35588 3556
rect 35420 3442 35476 3444
rect 35420 3390 35422 3442
rect 35422 3390 35474 3442
rect 35474 3390 35476 3442
rect 35420 3388 35476 3390
rect 36092 3388 36148 3444
rect 37212 10108 37268 10164
rect 37212 9548 37268 9604
rect 37324 6860 37380 6916
rect 36988 5010 37044 5012
rect 36988 4958 36990 5010
rect 36990 4958 37042 5010
rect 37042 4958 37044 5010
rect 36988 4956 37044 4958
rect 36876 4284 36932 4340
rect 37212 4172 37268 4228
rect 36764 3612 36820 3668
rect 36876 3442 36932 3444
rect 36876 3390 36878 3442
rect 36878 3390 36930 3442
rect 36930 3390 36932 3442
rect 36876 3388 36932 3390
rect 36204 3164 36260 3220
rect 35756 2770 35812 2772
rect 35756 2718 35758 2770
rect 35758 2718 35810 2770
rect 35810 2718 35812 2770
rect 35756 2716 35812 2718
rect 35644 2156 35700 2212
rect 35756 2492 35812 2548
rect 34636 1148 34692 1204
rect 34748 1090 34804 1092
rect 34748 1038 34750 1090
rect 34750 1038 34802 1090
rect 34802 1038 34804 1090
rect 34748 1036 34804 1038
rect 34076 978 34132 980
rect 34076 926 34078 978
rect 34078 926 34130 978
rect 34130 926 34132 978
rect 34076 924 34132 926
rect 34412 700 34468 756
rect 34748 364 34804 420
rect 34300 252 34356 308
rect 35308 1596 35364 1652
rect 35532 1372 35588 1428
rect 36652 2770 36708 2772
rect 36652 2718 36654 2770
rect 36654 2718 36706 2770
rect 36706 2718 36708 2770
rect 36652 2716 36708 2718
rect 36092 2044 36148 2100
rect 35980 476 36036 532
rect 36316 1820 36372 1876
rect 36428 1932 36484 1988
rect 37548 15484 37604 15540
rect 37548 13858 37604 13860
rect 37548 13806 37550 13858
rect 37550 13806 37602 13858
rect 37602 13806 37604 13858
rect 37548 13804 37604 13806
rect 37548 13244 37604 13300
rect 37548 11900 37604 11956
rect 37996 18956 38052 19012
rect 38108 17388 38164 17444
rect 37772 16156 37828 16212
rect 37884 16044 37940 16100
rect 37996 15484 38052 15540
rect 38892 27244 38948 27300
rect 39340 29036 39396 29092
rect 39676 33964 39732 34020
rect 39452 28028 39508 28084
rect 39788 28588 39844 28644
rect 39676 28476 39732 28532
rect 39788 28028 39844 28084
rect 38780 25676 38836 25732
rect 38556 23436 38612 23492
rect 39564 27020 39620 27076
rect 40236 35644 40292 35700
rect 40348 34412 40404 34468
rect 40348 34130 40404 34132
rect 40348 34078 40350 34130
rect 40350 34078 40402 34130
rect 40402 34078 40404 34130
rect 40348 34076 40404 34078
rect 40236 33740 40292 33796
rect 40908 43260 40964 43316
rect 40572 42252 40628 42308
rect 40908 42812 40964 42868
rect 40572 41916 40628 41972
rect 40908 42364 40964 42420
rect 40684 41804 40740 41860
rect 41020 42252 41076 42308
rect 40572 41132 40628 41188
rect 40684 41580 40740 41636
rect 40572 40908 40628 40964
rect 40572 36652 40628 36708
rect 41244 43820 41300 43876
rect 41356 43708 41412 43764
rect 41244 43372 41300 43428
rect 41916 48524 41972 48580
rect 41692 46284 41748 46340
rect 42252 47964 42308 48020
rect 42140 47068 42196 47124
rect 42252 46956 42308 47012
rect 42812 50818 42868 50820
rect 42812 50766 42814 50818
rect 42814 50766 42866 50818
rect 42866 50766 42868 50818
rect 42812 50764 42868 50766
rect 42924 50092 42980 50148
rect 42812 48802 42868 48804
rect 42812 48750 42814 48802
rect 42814 48750 42866 48802
rect 42866 48750 42868 48802
rect 42812 48748 42868 48750
rect 42700 46956 42756 47012
rect 42812 48524 42868 48580
rect 41804 46732 41860 46788
rect 42700 46786 42756 46788
rect 42700 46734 42702 46786
rect 42702 46734 42754 46786
rect 42754 46734 42756 46786
rect 42700 46732 42756 46734
rect 43036 48860 43092 48916
rect 43148 51436 43204 51492
rect 43260 50540 43316 50596
rect 43596 52108 43652 52164
rect 43484 51996 43540 52052
rect 44380 51884 44436 51940
rect 43804 51770 43860 51772
rect 43804 51718 43806 51770
rect 43806 51718 43858 51770
rect 43858 51718 43860 51770
rect 43804 51716 43860 51718
rect 43908 51770 43964 51772
rect 43908 51718 43910 51770
rect 43910 51718 43962 51770
rect 43962 51718 43964 51770
rect 43908 51716 43964 51718
rect 44012 51770 44068 51772
rect 44012 51718 44014 51770
rect 44014 51718 44066 51770
rect 44066 51718 44068 51770
rect 44012 51716 44068 51718
rect 44492 51772 44548 51828
rect 45164 54124 45220 54180
rect 45276 53730 45332 53732
rect 45276 53678 45278 53730
rect 45278 53678 45330 53730
rect 45330 53678 45332 53730
rect 45276 53676 45332 53678
rect 45164 53452 45220 53508
rect 45052 53004 45108 53060
rect 45276 53340 45332 53396
rect 45052 52834 45108 52836
rect 45052 52782 45054 52834
rect 45054 52782 45106 52834
rect 45106 52782 45108 52834
rect 45052 52780 45108 52782
rect 45500 53340 45556 53396
rect 45388 52162 45444 52164
rect 45388 52110 45390 52162
rect 45390 52110 45442 52162
rect 45442 52110 45444 52162
rect 45388 52108 45444 52110
rect 45164 51996 45220 52052
rect 46172 54514 46228 54516
rect 46172 54462 46174 54514
rect 46174 54462 46226 54514
rect 46226 54462 46228 54514
rect 46172 54460 46228 54462
rect 46396 55468 46452 55524
rect 46620 57036 46676 57092
rect 46508 55356 46564 55412
rect 46396 55298 46452 55300
rect 46396 55246 46398 55298
rect 46398 55246 46450 55298
rect 46450 55246 46452 55298
rect 46396 55244 46452 55246
rect 46732 55580 46788 55636
rect 47068 56588 47124 56644
rect 46844 55468 46900 55524
rect 47740 56140 47796 56196
rect 47404 55858 47460 55860
rect 47404 55806 47406 55858
rect 47406 55806 47458 55858
rect 47458 55806 47460 55858
rect 47404 55804 47460 55806
rect 47292 55468 47348 55524
rect 47628 55580 47684 55636
rect 46620 55244 46676 55300
rect 46732 55020 46788 55076
rect 46508 54460 46564 54516
rect 46284 54012 46340 54068
rect 45948 53452 46004 53508
rect 46508 53564 46564 53620
rect 46172 53116 46228 53172
rect 44940 51772 44996 51828
rect 44604 51548 44660 51604
rect 44492 51378 44548 51380
rect 44492 51326 44494 51378
rect 44494 51326 44546 51378
rect 44546 51326 44548 51378
rect 44492 51324 44548 51326
rect 44268 51212 44324 51268
rect 44380 51154 44436 51156
rect 44380 51102 44382 51154
rect 44382 51102 44434 51154
rect 44434 51102 44436 51154
rect 44380 51100 44436 51102
rect 44268 50876 44324 50932
rect 44464 50986 44520 50988
rect 44464 50934 44466 50986
rect 44466 50934 44518 50986
rect 44518 50934 44520 50986
rect 44464 50932 44520 50934
rect 44568 50986 44624 50988
rect 44568 50934 44570 50986
rect 44570 50934 44622 50986
rect 44622 50934 44624 50986
rect 44568 50932 44624 50934
rect 44672 50986 44728 50988
rect 44672 50934 44674 50986
rect 44674 50934 44726 50986
rect 44726 50934 44728 50986
rect 44672 50932 44728 50934
rect 43932 50706 43988 50708
rect 43932 50654 43934 50706
rect 43934 50654 43986 50706
rect 43986 50654 43988 50706
rect 43932 50652 43988 50654
rect 44380 50482 44436 50484
rect 44380 50430 44382 50482
rect 44382 50430 44434 50482
rect 44434 50430 44436 50482
rect 44380 50428 44436 50430
rect 44940 51378 44996 51380
rect 44940 51326 44942 51378
rect 44942 51326 44994 51378
rect 44994 51326 44996 51378
rect 44940 51324 44996 51326
rect 45276 51212 45332 51268
rect 45164 51100 45220 51156
rect 43372 50316 43428 50372
rect 44940 50876 44996 50932
rect 45052 50706 45108 50708
rect 45052 50654 45054 50706
rect 45054 50654 45106 50706
rect 45106 50654 45108 50706
rect 45052 50652 45108 50654
rect 43804 50202 43860 50204
rect 43804 50150 43806 50202
rect 43806 50150 43858 50202
rect 43858 50150 43860 50202
rect 43804 50148 43860 50150
rect 43908 50202 43964 50204
rect 43908 50150 43910 50202
rect 43910 50150 43962 50202
rect 43962 50150 43964 50202
rect 43908 50148 43964 50150
rect 44012 50202 44068 50204
rect 44012 50150 44014 50202
rect 44014 50150 44066 50202
rect 44066 50150 44068 50202
rect 44012 50148 44068 50150
rect 44492 50092 44548 50148
rect 43372 50034 43428 50036
rect 43372 49982 43374 50034
rect 43374 49982 43426 50034
rect 43426 49982 43428 50034
rect 43372 49980 43428 49982
rect 43260 48972 43316 49028
rect 45052 50092 45108 50148
rect 44828 49868 44884 49924
rect 44716 49810 44772 49812
rect 44716 49758 44718 49810
rect 44718 49758 44770 49810
rect 44770 49758 44772 49810
rect 44716 49756 44772 49758
rect 44268 49420 44324 49476
rect 43932 48748 43988 48804
rect 43036 48524 43092 48580
rect 44156 49308 44212 49364
rect 44464 49418 44520 49420
rect 44464 49366 44466 49418
rect 44466 49366 44518 49418
rect 44518 49366 44520 49418
rect 44464 49364 44520 49366
rect 44568 49418 44624 49420
rect 44568 49366 44570 49418
rect 44570 49366 44622 49418
rect 44622 49366 44624 49418
rect 44568 49364 44624 49366
rect 44672 49418 44728 49420
rect 44672 49366 44674 49418
rect 44674 49366 44726 49418
rect 44726 49366 44728 49418
rect 44672 49364 44728 49366
rect 45052 49868 45108 49924
rect 44828 49308 44884 49364
rect 44940 49420 44996 49476
rect 44604 48860 44660 48916
rect 44156 48748 44212 48804
rect 43596 48524 43652 48580
rect 43804 48634 43860 48636
rect 43804 48582 43806 48634
rect 43806 48582 43858 48634
rect 43858 48582 43860 48634
rect 43804 48580 43860 48582
rect 43908 48634 43964 48636
rect 43908 48582 43910 48634
rect 43910 48582 43962 48634
rect 43962 48582 43964 48634
rect 43908 48580 43964 48582
rect 44012 48634 44068 48636
rect 44012 48582 44014 48634
rect 44014 48582 44066 48634
rect 44066 48582 44068 48634
rect 44012 48580 44068 48582
rect 45276 50594 45332 50596
rect 45276 50542 45278 50594
rect 45278 50542 45330 50594
rect 45330 50542 45332 50594
rect 45276 50540 45332 50542
rect 45276 49810 45332 49812
rect 45276 49758 45278 49810
rect 45278 49758 45330 49810
rect 45330 49758 45332 49810
rect 45276 49756 45332 49758
rect 45052 48972 45108 49028
rect 45052 48636 45108 48692
rect 42812 46620 42868 46676
rect 42924 47292 42980 47348
rect 42252 46450 42308 46452
rect 42252 46398 42254 46450
rect 42254 46398 42306 46450
rect 42306 46398 42308 46450
rect 42252 46396 42308 46398
rect 43484 48018 43540 48020
rect 43484 47966 43486 48018
rect 43486 47966 43538 48018
rect 43538 47966 43540 48018
rect 43484 47964 43540 47966
rect 44828 48076 44884 48132
rect 43708 47964 43764 48020
rect 43372 47852 43428 47908
rect 44604 47964 44660 48020
rect 44464 47850 44520 47852
rect 44464 47798 44466 47850
rect 44466 47798 44518 47850
rect 44518 47798 44520 47850
rect 44464 47796 44520 47798
rect 44568 47850 44624 47852
rect 44568 47798 44570 47850
rect 44570 47798 44622 47850
rect 44622 47798 44624 47850
rect 44568 47796 44624 47798
rect 44672 47850 44728 47852
rect 44672 47798 44674 47850
rect 44674 47798 44726 47850
rect 44726 47798 44728 47850
rect 44828 47852 44884 47908
rect 44940 47964 44996 48020
rect 44672 47796 44728 47798
rect 45276 48188 45332 48244
rect 45724 51378 45780 51380
rect 45724 51326 45726 51378
rect 45726 51326 45778 51378
rect 45778 51326 45780 51378
rect 45724 51324 45780 51326
rect 45500 50988 45556 51044
rect 45500 50764 45556 50820
rect 45500 50092 45556 50148
rect 45836 51154 45892 51156
rect 45836 51102 45838 51154
rect 45838 51102 45890 51154
rect 45890 51102 45892 51154
rect 45836 51100 45892 51102
rect 45612 49980 45668 50036
rect 45836 50204 45892 50260
rect 45500 49196 45556 49252
rect 45612 48972 45668 49028
rect 45052 47740 45108 47796
rect 44268 47682 44324 47684
rect 44268 47630 44270 47682
rect 44270 47630 44322 47682
rect 44322 47630 44324 47682
rect 44268 47628 44324 47630
rect 44492 47404 44548 47460
rect 43036 46732 43092 46788
rect 42924 46396 42980 46452
rect 43372 46172 43428 46228
rect 41804 45948 41860 46004
rect 43372 45948 43428 46004
rect 41580 44380 41636 44436
rect 41692 45836 41748 45892
rect 41916 45052 41972 45108
rect 42252 45052 42308 45108
rect 42140 44716 42196 44772
rect 42140 44380 42196 44436
rect 42588 44716 42644 44772
rect 43036 45276 43092 45332
rect 42924 45106 42980 45108
rect 42924 45054 42926 45106
rect 42926 45054 42978 45106
rect 42978 45054 42980 45106
rect 42924 45052 42980 45054
rect 43372 45388 43428 45444
rect 43372 45052 43428 45108
rect 42924 44434 42980 44436
rect 42924 44382 42926 44434
rect 42926 44382 42978 44434
rect 42978 44382 42980 44434
rect 42924 44380 42980 44382
rect 42812 44098 42868 44100
rect 42812 44046 42814 44098
rect 42814 44046 42866 44098
rect 42866 44046 42868 44098
rect 42812 44044 42868 44046
rect 42924 43820 42980 43876
rect 41916 43426 41972 43428
rect 41916 43374 41918 43426
rect 41918 43374 41970 43426
rect 41970 43374 41972 43426
rect 41916 43372 41972 43374
rect 41244 42866 41300 42868
rect 41244 42814 41246 42866
rect 41246 42814 41298 42866
rect 41298 42814 41300 42866
rect 41244 42812 41300 42814
rect 41132 41692 41188 41748
rect 41020 40012 41076 40068
rect 41244 40012 41300 40068
rect 41132 39452 41188 39508
rect 40796 38892 40852 38948
rect 40796 37660 40852 37716
rect 41468 42812 41524 42868
rect 42476 43372 42532 43428
rect 41804 43314 41860 43316
rect 41804 43262 41806 43314
rect 41806 43262 41858 43314
rect 41858 43262 41860 43314
rect 41804 43260 41860 43262
rect 41580 42028 41636 42084
rect 42252 42700 42308 42756
rect 42252 42082 42308 42084
rect 42252 42030 42254 42082
rect 42254 42030 42306 42082
rect 42306 42030 42308 42082
rect 42252 42028 42308 42030
rect 41468 40348 41524 40404
rect 41356 39228 41412 39284
rect 40908 35698 40964 35700
rect 40908 35646 40910 35698
rect 40910 35646 40962 35698
rect 40962 35646 40964 35698
rect 40908 35644 40964 35646
rect 40796 35084 40852 35140
rect 40684 34636 40740 34692
rect 40684 34412 40740 34468
rect 40348 32956 40404 33012
rect 40236 31388 40292 31444
rect 40796 34188 40852 34244
rect 40908 34076 40964 34132
rect 40460 30940 40516 30996
rect 40236 30210 40292 30212
rect 40236 30158 40238 30210
rect 40238 30158 40290 30210
rect 40290 30158 40292 30210
rect 40236 30156 40292 30158
rect 40460 29708 40516 29764
rect 40012 28028 40068 28084
rect 40236 29372 40292 29428
rect 40012 27858 40068 27860
rect 40012 27806 40014 27858
rect 40014 27806 40066 27858
rect 40066 27806 40068 27858
rect 40012 27804 40068 27806
rect 40236 27804 40292 27860
rect 40348 29260 40404 29316
rect 39228 26908 39284 26964
rect 39116 25506 39172 25508
rect 39116 25454 39118 25506
rect 39118 25454 39170 25506
rect 39170 25454 39172 25506
rect 39116 25452 39172 25454
rect 39452 26684 39508 26740
rect 39340 25452 39396 25508
rect 39340 25282 39396 25284
rect 39340 25230 39342 25282
rect 39342 25230 39394 25282
rect 39394 25230 39396 25282
rect 39340 25228 39396 25230
rect 39676 26850 39732 26852
rect 39676 26798 39678 26850
rect 39678 26798 39730 26850
rect 39730 26798 39732 26850
rect 39676 26796 39732 26798
rect 39676 25788 39732 25844
rect 39788 25340 39844 25396
rect 39676 25004 39732 25060
rect 39900 26908 39956 26964
rect 39340 23884 39396 23940
rect 39116 23436 39172 23492
rect 38444 21868 38500 21924
rect 38668 21868 38724 21924
rect 38332 16156 38388 16212
rect 38556 20300 38612 20356
rect 38668 20972 38724 21028
rect 38556 19740 38612 19796
rect 38668 19010 38724 19012
rect 38668 18958 38670 19010
rect 38670 18958 38722 19010
rect 38722 18958 38724 19010
rect 38668 18956 38724 18958
rect 38220 15260 38276 15316
rect 37660 11788 37716 11844
rect 37548 10108 37604 10164
rect 37660 8316 37716 8372
rect 37548 7084 37604 7140
rect 37772 8204 37828 8260
rect 37548 5068 37604 5124
rect 37548 4284 37604 4340
rect 36988 2546 37044 2548
rect 36988 2494 36990 2546
rect 36990 2494 37042 2546
rect 37042 2494 37044 2546
rect 36988 2492 37044 2494
rect 36876 1202 36932 1204
rect 36876 1150 36878 1202
rect 36878 1150 36930 1202
rect 36930 1150 36932 1202
rect 36876 1148 36932 1150
rect 36540 476 36596 532
rect 37436 3276 37492 3332
rect 37660 2940 37716 2996
rect 37324 2770 37380 2772
rect 37324 2718 37326 2770
rect 37326 2718 37378 2770
rect 37378 2718 37380 2770
rect 37324 2716 37380 2718
rect 37548 2210 37604 2212
rect 37548 2158 37550 2210
rect 37550 2158 37602 2210
rect 37602 2158 37604 2210
rect 37548 2156 37604 2158
rect 36764 140 36820 196
rect 37996 14252 38052 14308
rect 38220 14028 38276 14084
rect 37996 13634 38052 13636
rect 37996 13582 37998 13634
rect 37998 13582 38050 13634
rect 38050 13582 38052 13634
rect 37996 13580 38052 13582
rect 38108 12908 38164 12964
rect 37996 11788 38052 11844
rect 38108 11676 38164 11732
rect 38444 15314 38500 15316
rect 38444 15262 38446 15314
rect 38446 15262 38498 15314
rect 38498 15262 38500 15314
rect 38444 15260 38500 15262
rect 39228 22930 39284 22932
rect 39228 22878 39230 22930
rect 39230 22878 39282 22930
rect 39282 22878 39284 22930
rect 39228 22876 39284 22878
rect 39676 24220 39732 24276
rect 40236 27244 40292 27300
rect 40236 27074 40292 27076
rect 40236 27022 40238 27074
rect 40238 27022 40290 27074
rect 40290 27022 40292 27074
rect 40236 27020 40292 27022
rect 40124 26290 40180 26292
rect 40124 26238 40126 26290
rect 40126 26238 40178 26290
rect 40178 26238 40180 26290
rect 40124 26236 40180 26238
rect 40124 25788 40180 25844
rect 40124 25564 40180 25620
rect 40012 23884 40068 23940
rect 40908 33292 40964 33348
rect 41244 36652 41300 36708
rect 41468 38274 41524 38276
rect 41468 38222 41470 38274
rect 41470 38222 41522 38274
rect 41522 38222 41524 38274
rect 41468 38220 41524 38222
rect 41468 37660 41524 37716
rect 41468 37324 41524 37380
rect 41916 41858 41972 41860
rect 41916 41806 41918 41858
rect 41918 41806 41970 41858
rect 41970 41806 41972 41858
rect 41916 41804 41972 41806
rect 42364 41804 42420 41860
rect 42364 41468 42420 41524
rect 42252 41020 42308 41076
rect 42028 40348 42084 40404
rect 41916 39116 41972 39172
rect 43260 44380 43316 44436
rect 43260 43820 43316 43876
rect 43036 43484 43092 43540
rect 42588 41858 42644 41860
rect 42588 41806 42590 41858
rect 42590 41806 42642 41858
rect 42642 41806 42644 41858
rect 42588 41804 42644 41806
rect 42588 41410 42644 41412
rect 42588 41358 42590 41410
rect 42590 41358 42642 41410
rect 42642 41358 42644 41410
rect 42588 41356 42644 41358
rect 43484 44716 43540 44772
rect 43708 47180 43764 47236
rect 43804 47066 43860 47068
rect 43804 47014 43806 47066
rect 43806 47014 43858 47066
rect 43858 47014 43860 47066
rect 43804 47012 43860 47014
rect 43908 47066 43964 47068
rect 43908 47014 43910 47066
rect 43910 47014 43962 47066
rect 43962 47014 43964 47066
rect 43908 47012 43964 47014
rect 44012 47066 44068 47068
rect 44012 47014 44014 47066
rect 44014 47014 44066 47066
rect 44066 47014 44068 47066
rect 44012 47012 44068 47014
rect 44828 47180 44884 47236
rect 45164 47180 45220 47236
rect 43820 46508 43876 46564
rect 43820 45724 43876 45780
rect 43804 45498 43860 45500
rect 43804 45446 43806 45498
rect 43806 45446 43858 45498
rect 43858 45446 43860 45498
rect 43804 45444 43860 45446
rect 43908 45498 43964 45500
rect 43908 45446 43910 45498
rect 43910 45446 43962 45498
rect 43962 45446 43964 45498
rect 43908 45444 43964 45446
rect 44012 45498 44068 45500
rect 44012 45446 44014 45498
rect 44014 45446 44066 45498
rect 44066 45446 44068 45498
rect 44012 45444 44068 45446
rect 43820 44604 43876 44660
rect 43804 43930 43860 43932
rect 43804 43878 43806 43930
rect 43806 43878 43858 43930
rect 43858 43878 43860 43930
rect 43804 43876 43860 43878
rect 43908 43930 43964 43932
rect 43908 43878 43910 43930
rect 43910 43878 43962 43930
rect 43962 43878 43964 43930
rect 43908 43876 43964 43878
rect 44012 43930 44068 43932
rect 44012 43878 44014 43930
rect 44014 43878 44066 43930
rect 44066 43878 44068 43930
rect 44012 43876 44068 43878
rect 43708 43708 43764 43764
rect 43596 43260 43652 43316
rect 43372 42588 43428 42644
rect 43372 42364 43428 42420
rect 43484 42252 43540 42308
rect 43036 41858 43092 41860
rect 43036 41806 43038 41858
rect 43038 41806 43090 41858
rect 43090 41806 43092 41858
rect 43036 41804 43092 41806
rect 42924 41468 42980 41524
rect 42812 41356 42868 41412
rect 43372 41804 43428 41860
rect 43260 41692 43316 41748
rect 43148 41244 43204 41300
rect 42476 40796 42532 40852
rect 42252 39788 42308 39844
rect 42252 39452 42308 39508
rect 43372 40962 43428 40964
rect 43372 40910 43374 40962
rect 43374 40910 43426 40962
rect 43426 40910 43428 40962
rect 43372 40908 43428 40910
rect 42812 40514 42868 40516
rect 42812 40462 42814 40514
rect 42814 40462 42866 40514
rect 42866 40462 42868 40514
rect 42812 40460 42868 40462
rect 43372 40402 43428 40404
rect 43372 40350 43374 40402
rect 43374 40350 43426 40402
rect 43426 40350 43428 40402
rect 43372 40348 43428 40350
rect 43708 42924 43764 42980
rect 43932 43708 43988 43764
rect 44464 46282 44520 46284
rect 44464 46230 44466 46282
rect 44466 46230 44518 46282
rect 44518 46230 44520 46282
rect 44464 46228 44520 46230
rect 44568 46282 44624 46284
rect 44568 46230 44570 46282
rect 44570 46230 44622 46282
rect 44622 46230 44624 46282
rect 44568 46228 44624 46230
rect 44672 46282 44728 46284
rect 44672 46230 44674 46282
rect 44674 46230 44726 46282
rect 44726 46230 44728 46282
rect 44672 46228 44728 46230
rect 45052 45836 45108 45892
rect 44940 45666 44996 45668
rect 44940 45614 44942 45666
rect 44942 45614 44994 45666
rect 44994 45614 44996 45666
rect 44940 45612 44996 45614
rect 44828 45388 44884 45444
rect 44380 45276 44436 45332
rect 44464 44714 44520 44716
rect 44464 44662 44466 44714
rect 44466 44662 44518 44714
rect 44518 44662 44520 44714
rect 44464 44660 44520 44662
rect 44568 44714 44624 44716
rect 44568 44662 44570 44714
rect 44570 44662 44622 44714
rect 44622 44662 44624 44714
rect 44568 44660 44624 44662
rect 44672 44714 44728 44716
rect 44672 44662 44674 44714
rect 44674 44662 44726 44714
rect 44726 44662 44728 44714
rect 44672 44660 44728 44662
rect 45500 46956 45556 47012
rect 45164 45276 45220 45332
rect 45388 46396 45444 46452
rect 45052 44604 45108 44660
rect 44940 44380 44996 44436
rect 44268 43484 44324 43540
rect 44492 43538 44548 43540
rect 44492 43486 44494 43538
rect 44494 43486 44546 43538
rect 44546 43486 44548 43538
rect 44492 43484 44548 43486
rect 44156 43426 44212 43428
rect 44156 43374 44158 43426
rect 44158 43374 44210 43426
rect 44210 43374 44212 43426
rect 44156 43372 44212 43374
rect 44268 43148 44324 43204
rect 44464 43146 44520 43148
rect 44464 43094 44466 43146
rect 44466 43094 44518 43146
rect 44518 43094 44520 43146
rect 44464 43092 44520 43094
rect 44568 43146 44624 43148
rect 44568 43094 44570 43146
rect 44570 43094 44622 43146
rect 44622 43094 44624 43146
rect 44568 43092 44624 43094
rect 44672 43146 44728 43148
rect 44672 43094 44674 43146
rect 44674 43094 44726 43146
rect 44726 43094 44728 43146
rect 44672 43092 44728 43094
rect 43932 42700 43988 42756
rect 43804 42362 43860 42364
rect 43804 42310 43806 42362
rect 43806 42310 43858 42362
rect 43858 42310 43860 42362
rect 43804 42308 43860 42310
rect 43908 42362 43964 42364
rect 43908 42310 43910 42362
rect 43910 42310 43962 42362
rect 43962 42310 43964 42362
rect 43908 42308 43964 42310
rect 44012 42362 44068 42364
rect 44012 42310 44014 42362
rect 44014 42310 44066 42362
rect 44066 42310 44068 42362
rect 44012 42308 44068 42310
rect 43820 41410 43876 41412
rect 43820 41358 43822 41410
rect 43822 41358 43874 41410
rect 43874 41358 43876 41410
rect 43820 41356 43876 41358
rect 43804 40794 43860 40796
rect 43804 40742 43806 40794
rect 43806 40742 43858 40794
rect 43858 40742 43860 40794
rect 43804 40740 43860 40742
rect 43908 40794 43964 40796
rect 43908 40742 43910 40794
rect 43910 40742 43962 40794
rect 43962 40742 43964 40794
rect 43908 40740 43964 40742
rect 44012 40794 44068 40796
rect 44012 40742 44014 40794
rect 44014 40742 44066 40794
rect 44066 40742 44068 40794
rect 44012 40740 44068 40742
rect 44156 40796 44212 40852
rect 42476 39564 42532 39620
rect 42028 38780 42084 38836
rect 42588 39116 42644 39172
rect 41916 38668 41972 38724
rect 42476 38556 42532 38612
rect 42028 38220 42084 38276
rect 42476 37938 42532 37940
rect 42476 37886 42478 37938
rect 42478 37886 42530 37938
rect 42530 37886 42532 37938
rect 42476 37884 42532 37886
rect 41804 37324 41860 37380
rect 41132 36370 41188 36372
rect 41132 36318 41134 36370
rect 41134 36318 41186 36370
rect 41186 36318 41188 36370
rect 41132 36316 41188 36318
rect 41356 36204 41412 36260
rect 41804 36876 41860 36932
rect 41580 35868 41636 35924
rect 41692 36316 41748 36372
rect 41468 35420 41524 35476
rect 41356 34300 41412 34356
rect 41468 35084 41524 35140
rect 41244 33740 41300 33796
rect 41692 34748 41748 34804
rect 41580 34412 41636 34468
rect 42476 36876 42532 36932
rect 41916 35756 41972 35812
rect 42252 36652 42308 36708
rect 42028 35084 42084 35140
rect 42028 34524 42084 34580
rect 41468 33292 41524 33348
rect 41804 34188 41860 34244
rect 41132 32844 41188 32900
rect 41244 32956 41300 33012
rect 41020 31948 41076 32004
rect 41356 32338 41412 32340
rect 41356 32286 41358 32338
rect 41358 32286 41410 32338
rect 41410 32286 41412 32338
rect 41356 32284 41412 32286
rect 41580 32172 41636 32228
rect 41132 31724 41188 31780
rect 41132 30994 41188 30996
rect 41132 30942 41134 30994
rect 41134 30942 41186 30994
rect 41186 30942 41188 30994
rect 41132 30940 41188 30942
rect 42364 35532 42420 35588
rect 43260 38220 43316 38276
rect 42812 37324 42868 37380
rect 43260 37548 43316 37604
rect 42700 36988 42756 37044
rect 42924 35586 42980 35588
rect 42924 35534 42926 35586
rect 42926 35534 42978 35586
rect 42978 35534 42980 35586
rect 42924 35532 42980 35534
rect 43148 35532 43204 35588
rect 42700 35084 42756 35140
rect 42812 35196 42868 35252
rect 43036 33964 43092 34020
rect 42700 33292 42756 33348
rect 42476 32956 42532 33012
rect 45724 48860 45780 48916
rect 46508 52892 46564 52948
rect 46284 52444 46340 52500
rect 46060 50204 46116 50260
rect 46060 49756 46116 49812
rect 46620 52722 46676 52724
rect 46620 52670 46622 52722
rect 46622 52670 46674 52722
rect 46674 52670 46676 52722
rect 46620 52668 46676 52670
rect 46620 52220 46676 52276
rect 47292 54236 47348 54292
rect 47180 53676 47236 53732
rect 46956 53228 47012 53284
rect 46732 52108 46788 52164
rect 47516 53730 47572 53732
rect 47516 53678 47518 53730
rect 47518 53678 47570 53730
rect 47570 53678 47572 53730
rect 47516 53676 47572 53678
rect 46844 51996 46900 52052
rect 47516 51772 47572 51828
rect 46620 51212 46676 51268
rect 46396 50764 46452 50820
rect 46172 50428 46228 50484
rect 47068 50988 47124 51044
rect 46844 49810 46900 49812
rect 46844 49758 46846 49810
rect 46846 49758 46898 49810
rect 46898 49758 46900 49810
rect 46844 49756 46900 49758
rect 46396 49644 46452 49700
rect 45948 47180 46004 47236
rect 46396 48972 46452 49028
rect 46620 48860 46676 48916
rect 48636 56700 48692 56756
rect 49532 56812 49588 56868
rect 49084 56476 49140 56532
rect 49756 56476 49812 56532
rect 48188 56028 48244 56084
rect 49084 55970 49140 55972
rect 49084 55918 49086 55970
rect 49086 55918 49138 55970
rect 49138 55918 49140 55970
rect 49084 55916 49140 55918
rect 47852 55356 47908 55412
rect 48412 55858 48468 55860
rect 48412 55806 48414 55858
rect 48414 55806 48466 55858
rect 48466 55806 48468 55858
rect 48412 55804 48468 55806
rect 48748 55468 48804 55524
rect 48972 55692 49028 55748
rect 48076 55132 48132 55188
rect 48748 54684 48804 54740
rect 48636 54348 48692 54404
rect 48188 53730 48244 53732
rect 48188 53678 48190 53730
rect 48190 53678 48242 53730
rect 48242 53678 48244 53730
rect 48188 53676 48244 53678
rect 48412 52834 48468 52836
rect 48412 52782 48414 52834
rect 48414 52782 48466 52834
rect 48466 52782 48468 52834
rect 48412 52780 48468 52782
rect 48076 52108 48132 52164
rect 48300 52332 48356 52388
rect 48748 54124 48804 54180
rect 48972 54124 49028 54180
rect 49196 55692 49252 55748
rect 49420 55468 49476 55524
rect 49980 55468 50036 55524
rect 50540 57148 50596 57204
rect 50876 57036 50932 57092
rect 50876 55468 50932 55524
rect 51100 55580 51156 55636
rect 50428 55186 50484 55188
rect 50428 55134 50430 55186
rect 50430 55134 50482 55186
rect 50482 55134 50484 55186
rect 50428 55132 50484 55134
rect 50316 54908 50372 54964
rect 50652 54796 50708 54852
rect 49980 54684 50036 54740
rect 49420 54012 49476 54068
rect 49196 53788 49252 53844
rect 49084 53676 49140 53732
rect 48636 53228 48692 53284
rect 49868 53004 49924 53060
rect 48524 52332 48580 52388
rect 49196 52722 49252 52724
rect 49196 52670 49198 52722
rect 49198 52670 49250 52722
rect 49250 52670 49252 52722
rect 49196 52668 49252 52670
rect 48748 52220 48804 52276
rect 48860 52556 48916 52612
rect 48860 51996 48916 52052
rect 48300 51548 48356 51604
rect 48076 51100 48132 51156
rect 47628 50988 47684 51044
rect 47740 50876 47796 50932
rect 47180 50652 47236 50708
rect 47404 50706 47460 50708
rect 47404 50654 47406 50706
rect 47406 50654 47458 50706
rect 47458 50654 47460 50706
rect 47404 50652 47460 50654
rect 47516 50540 47572 50596
rect 47404 50204 47460 50260
rect 47068 48860 47124 48916
rect 46732 48748 46788 48804
rect 46844 47570 46900 47572
rect 46844 47518 46846 47570
rect 46846 47518 46898 47570
rect 46898 47518 46900 47570
rect 46844 47516 46900 47518
rect 46508 47404 46564 47460
rect 46732 46674 46788 46676
rect 46732 46622 46734 46674
rect 46734 46622 46786 46674
rect 46786 46622 46788 46674
rect 46732 46620 46788 46622
rect 47068 47740 47124 47796
rect 45612 45948 45668 46004
rect 45388 43484 45444 43540
rect 45388 42924 45444 42980
rect 45276 42812 45332 42868
rect 44940 41916 44996 41972
rect 45052 42700 45108 42756
rect 44828 41692 44884 41748
rect 44464 41578 44520 41580
rect 44464 41526 44466 41578
rect 44466 41526 44518 41578
rect 44518 41526 44520 41578
rect 44464 41524 44520 41526
rect 44568 41578 44624 41580
rect 44568 41526 44570 41578
rect 44570 41526 44622 41578
rect 44622 41526 44624 41578
rect 44568 41524 44624 41526
rect 44672 41578 44728 41580
rect 44672 41526 44674 41578
rect 44674 41526 44726 41578
rect 44726 41526 44728 41578
rect 44672 41524 44728 41526
rect 44940 41132 44996 41188
rect 45164 42588 45220 42644
rect 45388 41468 45444 41524
rect 45500 41692 45556 41748
rect 45500 40908 45556 40964
rect 44268 40460 44324 40516
rect 44492 40460 44548 40516
rect 44156 40012 44212 40068
rect 44828 40178 44884 40180
rect 44828 40126 44830 40178
rect 44830 40126 44882 40178
rect 44882 40126 44884 40178
rect 44828 40124 44884 40126
rect 43708 39452 43764 39508
rect 43804 39226 43860 39228
rect 43484 39116 43540 39172
rect 43804 39174 43806 39226
rect 43806 39174 43858 39226
rect 43858 39174 43860 39226
rect 43804 39172 43860 39174
rect 43908 39226 43964 39228
rect 43908 39174 43910 39226
rect 43910 39174 43962 39226
rect 43962 39174 43964 39226
rect 43908 39172 43964 39174
rect 44012 39226 44068 39228
rect 44012 39174 44014 39226
rect 44014 39174 44066 39226
rect 44066 39174 44068 39226
rect 44012 39172 44068 39174
rect 43932 38668 43988 38724
rect 44464 40010 44520 40012
rect 44464 39958 44466 40010
rect 44466 39958 44518 40010
rect 44518 39958 44520 40010
rect 44464 39956 44520 39958
rect 44568 40010 44624 40012
rect 44568 39958 44570 40010
rect 44570 39958 44622 40010
rect 44622 39958 44624 40010
rect 44568 39956 44624 39958
rect 44672 40010 44728 40012
rect 44672 39958 44674 40010
rect 44674 39958 44726 40010
rect 44726 39958 44728 40010
rect 44672 39956 44728 39958
rect 44716 39452 44772 39508
rect 44380 39116 44436 39172
rect 44380 38668 44436 38724
rect 44716 38722 44772 38724
rect 44716 38670 44718 38722
rect 44718 38670 44770 38722
rect 44770 38670 44772 38722
rect 44716 38668 44772 38670
rect 45276 40796 45332 40852
rect 45164 40684 45220 40740
rect 45052 39842 45108 39844
rect 45052 39790 45054 39842
rect 45054 39790 45106 39842
rect 45106 39790 45108 39842
rect 45052 39788 45108 39790
rect 45052 39340 45108 39396
rect 44268 38332 44324 38388
rect 44464 38442 44520 38444
rect 44464 38390 44466 38442
rect 44466 38390 44518 38442
rect 44518 38390 44520 38442
rect 44464 38388 44520 38390
rect 44568 38442 44624 38444
rect 44568 38390 44570 38442
rect 44570 38390 44622 38442
rect 44622 38390 44624 38442
rect 44568 38388 44624 38390
rect 44672 38442 44728 38444
rect 44672 38390 44674 38442
rect 44674 38390 44726 38442
rect 44726 38390 44728 38442
rect 44672 38388 44728 38390
rect 44492 37996 44548 38052
rect 43372 36652 43428 36708
rect 43804 37658 43860 37660
rect 43804 37606 43806 37658
rect 43806 37606 43858 37658
rect 43858 37606 43860 37658
rect 43804 37604 43860 37606
rect 43908 37658 43964 37660
rect 43908 37606 43910 37658
rect 43910 37606 43962 37658
rect 43962 37606 43964 37658
rect 43908 37604 43964 37606
rect 44012 37658 44068 37660
rect 44012 37606 44014 37658
rect 44014 37606 44066 37658
rect 44066 37606 44068 37658
rect 44156 37660 44212 37716
rect 44012 37604 44068 37606
rect 44492 37548 44548 37604
rect 43372 36428 43428 36484
rect 43596 37324 43652 37380
rect 43708 37212 43764 37268
rect 43484 36316 43540 36372
rect 44492 37212 44548 37268
rect 44156 37154 44212 37156
rect 44156 37102 44158 37154
rect 44158 37102 44210 37154
rect 44210 37102 44212 37154
rect 44156 37100 44212 37102
rect 44716 37154 44772 37156
rect 44716 37102 44718 37154
rect 44718 37102 44770 37154
rect 44770 37102 44772 37154
rect 44716 37100 44772 37102
rect 44464 36874 44520 36876
rect 44156 36764 44212 36820
rect 44464 36822 44466 36874
rect 44466 36822 44518 36874
rect 44518 36822 44520 36874
rect 44464 36820 44520 36822
rect 44568 36874 44624 36876
rect 44568 36822 44570 36874
rect 44570 36822 44622 36874
rect 44622 36822 44624 36874
rect 44568 36820 44624 36822
rect 44672 36874 44728 36876
rect 44672 36822 44674 36874
rect 44674 36822 44726 36874
rect 44726 36822 44728 36874
rect 44672 36820 44728 36822
rect 43708 36316 43764 36372
rect 43804 36090 43860 36092
rect 43804 36038 43806 36090
rect 43806 36038 43858 36090
rect 43858 36038 43860 36090
rect 43804 36036 43860 36038
rect 43908 36090 43964 36092
rect 43908 36038 43910 36090
rect 43910 36038 43962 36090
rect 43962 36038 43964 36090
rect 43908 36036 43964 36038
rect 44012 36090 44068 36092
rect 44012 36038 44014 36090
rect 44014 36038 44066 36090
rect 44066 36038 44068 36090
rect 44012 36036 44068 36038
rect 44380 35980 44436 36036
rect 44268 35922 44324 35924
rect 44268 35870 44270 35922
rect 44270 35870 44322 35922
rect 44322 35870 44324 35922
rect 44268 35868 44324 35870
rect 43484 35756 43540 35812
rect 43596 35644 43652 35700
rect 43372 35308 43428 35364
rect 43708 35586 43764 35588
rect 43708 35534 43710 35586
rect 43710 35534 43762 35586
rect 43762 35534 43764 35586
rect 43708 35532 43764 35534
rect 43596 35196 43652 35252
rect 44940 38274 44996 38276
rect 44940 38222 44942 38274
rect 44942 38222 44994 38274
rect 44994 38222 44996 38274
rect 44940 38220 44996 38222
rect 45052 38050 45108 38052
rect 45052 37998 45054 38050
rect 45054 37998 45106 38050
rect 45106 37998 45108 38050
rect 45052 37996 45108 37998
rect 44464 35306 44520 35308
rect 44464 35254 44466 35306
rect 44466 35254 44518 35306
rect 44518 35254 44520 35306
rect 44464 35252 44520 35254
rect 44568 35306 44624 35308
rect 44568 35254 44570 35306
rect 44570 35254 44622 35306
rect 44622 35254 44624 35306
rect 44568 35252 44624 35254
rect 44672 35306 44728 35308
rect 44672 35254 44674 35306
rect 44674 35254 44726 35306
rect 44726 35254 44728 35306
rect 44828 35308 44884 35364
rect 44940 37660 44996 37716
rect 45276 40124 45332 40180
rect 45500 39788 45556 39844
rect 45388 39116 45444 39172
rect 46284 45890 46340 45892
rect 46284 45838 46286 45890
rect 46286 45838 46338 45890
rect 46338 45838 46340 45890
rect 46284 45836 46340 45838
rect 45948 45330 46004 45332
rect 45948 45278 45950 45330
rect 45950 45278 46002 45330
rect 46002 45278 46004 45330
rect 45948 45276 46004 45278
rect 45836 44380 45892 44436
rect 45948 43484 46004 43540
rect 45724 43260 45780 43316
rect 45724 42866 45780 42868
rect 45724 42814 45726 42866
rect 45726 42814 45778 42866
rect 45778 42814 45780 42866
rect 45724 42812 45780 42814
rect 45724 42588 45780 42644
rect 46508 45218 46564 45220
rect 46508 45166 46510 45218
rect 46510 45166 46562 45218
rect 46562 45166 46564 45218
rect 46508 45164 46564 45166
rect 46396 45106 46452 45108
rect 46396 45054 46398 45106
rect 46398 45054 46450 45106
rect 46450 45054 46452 45106
rect 46396 45052 46452 45054
rect 46732 45666 46788 45668
rect 46732 45614 46734 45666
rect 46734 45614 46786 45666
rect 46786 45614 46788 45666
rect 46732 45612 46788 45614
rect 46620 44716 46676 44772
rect 46732 45388 46788 45444
rect 46284 43932 46340 43988
rect 46172 43148 46228 43204
rect 46060 42588 46116 42644
rect 45724 41580 45780 41636
rect 45724 39564 45780 39620
rect 45836 41468 45892 41524
rect 45612 39116 45668 39172
rect 45948 40908 46004 40964
rect 46284 42700 46340 42756
rect 46620 43314 46676 43316
rect 46620 43262 46622 43314
rect 46622 43262 46674 43314
rect 46674 43262 46676 43314
rect 46620 43260 46676 43262
rect 47404 46396 47460 46452
rect 47628 49868 47684 49924
rect 48076 50876 48132 50932
rect 47852 50316 47908 50372
rect 48748 51938 48804 51940
rect 48748 51886 48750 51938
rect 48750 51886 48802 51938
rect 48802 51886 48804 51938
rect 48748 51884 48804 51886
rect 48524 51490 48580 51492
rect 48524 51438 48526 51490
rect 48526 51438 48578 51490
rect 48578 51438 48580 51490
rect 48524 51436 48580 51438
rect 48748 51100 48804 51156
rect 48972 51884 49028 51940
rect 48860 50764 48916 50820
rect 48524 50594 48580 50596
rect 48524 50542 48526 50594
rect 48526 50542 48578 50594
rect 48578 50542 48580 50594
rect 48524 50540 48580 50542
rect 49308 51548 49364 51604
rect 49084 50706 49140 50708
rect 49084 50654 49086 50706
rect 49086 50654 49138 50706
rect 49138 50654 49140 50706
rect 49084 50652 49140 50654
rect 49196 50428 49252 50484
rect 48412 49868 48468 49924
rect 48860 49868 48916 49924
rect 47964 49698 48020 49700
rect 47964 49646 47966 49698
rect 47966 49646 48018 49698
rect 48018 49646 48020 49698
rect 47964 49644 48020 49646
rect 47740 47628 47796 47684
rect 48524 49644 48580 49700
rect 48300 49026 48356 49028
rect 48300 48974 48302 49026
rect 48302 48974 48354 49026
rect 48354 48974 48356 49026
rect 48300 48972 48356 48974
rect 48972 49810 49028 49812
rect 48972 49758 48974 49810
rect 48974 49758 49026 49810
rect 49026 49758 49028 49810
rect 48972 49756 49028 49758
rect 49084 49420 49140 49476
rect 47628 46450 47684 46452
rect 47628 46398 47630 46450
rect 47630 46398 47682 46450
rect 47682 46398 47684 46450
rect 47628 46396 47684 46398
rect 47404 46002 47460 46004
rect 47404 45950 47406 46002
rect 47406 45950 47458 46002
rect 47458 45950 47460 46002
rect 47404 45948 47460 45950
rect 47292 45778 47348 45780
rect 47292 45726 47294 45778
rect 47294 45726 47346 45778
rect 47346 45726 47348 45778
rect 47292 45724 47348 45726
rect 47180 45276 47236 45332
rect 46844 43484 46900 43540
rect 46956 44828 47012 44884
rect 46844 42924 46900 42980
rect 46060 38668 46116 38724
rect 46732 41916 46788 41972
rect 46620 40514 46676 40516
rect 46620 40462 46622 40514
rect 46622 40462 46674 40514
rect 46674 40462 46676 40514
rect 46620 40460 46676 40462
rect 46844 40796 46900 40852
rect 46396 38780 46452 38836
rect 46508 39340 46564 39396
rect 45164 37324 45220 37380
rect 44672 35252 44728 35254
rect 44828 35138 44884 35140
rect 44828 35086 44830 35138
rect 44830 35086 44882 35138
rect 44882 35086 44884 35138
rect 44828 35084 44884 35086
rect 43260 34636 43316 34692
rect 43372 34524 43428 34580
rect 43148 32956 43204 33012
rect 43260 34412 43316 34468
rect 43804 34522 43860 34524
rect 43804 34470 43806 34522
rect 43806 34470 43858 34522
rect 43858 34470 43860 34522
rect 43804 34468 43860 34470
rect 43908 34522 43964 34524
rect 43908 34470 43910 34522
rect 43910 34470 43962 34522
rect 43962 34470 43964 34522
rect 43908 34468 43964 34470
rect 44012 34522 44068 34524
rect 44012 34470 44014 34522
rect 44014 34470 44066 34522
rect 44066 34470 44068 34522
rect 44012 34468 44068 34470
rect 43372 33740 43428 33796
rect 43260 33628 43316 33684
rect 42252 32172 42308 32228
rect 42028 31778 42084 31780
rect 42028 31726 42030 31778
rect 42030 31726 42082 31778
rect 42082 31726 42084 31778
rect 42028 31724 42084 31726
rect 42252 31164 42308 31220
rect 42476 31724 42532 31780
rect 41132 30268 41188 30324
rect 41020 30210 41076 30212
rect 41020 30158 41022 30210
rect 41022 30158 41074 30210
rect 41074 30158 41076 30210
rect 41020 30156 41076 30158
rect 41244 30156 41300 30212
rect 40908 29260 40964 29316
rect 41020 28924 41076 28980
rect 42140 28924 42196 28980
rect 40908 28866 40964 28868
rect 40908 28814 40910 28866
rect 40910 28814 40962 28866
rect 40962 28814 40964 28866
rect 40908 28812 40964 28814
rect 40796 28140 40852 28196
rect 41916 28700 41972 28756
rect 40684 28028 40740 28084
rect 40684 27634 40740 27636
rect 40684 27582 40686 27634
rect 40686 27582 40738 27634
rect 40738 27582 40740 27634
rect 40684 27580 40740 27582
rect 40572 27132 40628 27188
rect 40460 26796 40516 26852
rect 40572 26684 40628 26740
rect 40684 27020 40740 27076
rect 41132 27074 41188 27076
rect 41132 27022 41134 27074
rect 41134 27022 41186 27074
rect 41186 27022 41188 27074
rect 41132 27020 41188 27022
rect 41804 27356 41860 27412
rect 41468 27132 41524 27188
rect 41692 27020 41748 27076
rect 40796 26460 40852 26516
rect 41468 26348 41524 26404
rect 40460 25788 40516 25844
rect 40684 25730 40740 25732
rect 40684 25678 40686 25730
rect 40686 25678 40738 25730
rect 40738 25678 40740 25730
rect 40684 25676 40740 25678
rect 40796 25618 40852 25620
rect 40796 25566 40798 25618
rect 40798 25566 40850 25618
rect 40850 25566 40852 25618
rect 40796 25564 40852 25566
rect 41244 26178 41300 26180
rect 41244 26126 41246 26178
rect 41246 26126 41298 26178
rect 41298 26126 41300 26178
rect 41244 26124 41300 26126
rect 41020 25618 41076 25620
rect 41020 25566 41022 25618
rect 41022 25566 41074 25618
rect 41074 25566 41076 25618
rect 41020 25564 41076 25566
rect 40460 25506 40516 25508
rect 40460 25454 40462 25506
rect 40462 25454 40514 25506
rect 40514 25454 40516 25506
rect 40460 25452 40516 25454
rect 41020 25340 41076 25396
rect 39340 21868 39396 21924
rect 39228 21586 39284 21588
rect 39228 21534 39230 21586
rect 39230 21534 39282 21586
rect 39282 21534 39284 21586
rect 39228 21532 39284 21534
rect 38892 20802 38948 20804
rect 38892 20750 38894 20802
rect 38894 20750 38946 20802
rect 38946 20750 38948 20802
rect 38892 20748 38948 20750
rect 38780 18396 38836 18452
rect 38892 19180 38948 19236
rect 38780 16882 38836 16884
rect 38780 16830 38782 16882
rect 38782 16830 38834 16882
rect 38834 16830 38836 16882
rect 38780 16828 38836 16830
rect 39228 21084 39284 21140
rect 39116 20972 39172 21028
rect 39116 20636 39172 20692
rect 39228 20524 39284 20580
rect 39564 21586 39620 21588
rect 39564 21534 39566 21586
rect 39566 21534 39618 21586
rect 39618 21534 39620 21586
rect 39564 21532 39620 21534
rect 39900 23436 39956 23492
rect 40012 21644 40068 21700
rect 39676 20802 39732 20804
rect 39676 20750 39678 20802
rect 39678 20750 39730 20802
rect 39730 20750 39732 20802
rect 39676 20748 39732 20750
rect 39340 20018 39396 20020
rect 39340 19966 39342 20018
rect 39342 19966 39394 20018
rect 39394 19966 39396 20018
rect 39340 19964 39396 19966
rect 39564 20636 39620 20692
rect 39788 19852 39844 19908
rect 39340 18732 39396 18788
rect 39676 18620 39732 18676
rect 39004 17500 39060 17556
rect 39228 16658 39284 16660
rect 39228 16606 39230 16658
rect 39230 16606 39282 16658
rect 39282 16606 39284 16658
rect 39228 16604 39284 16606
rect 39564 16492 39620 16548
rect 38892 16098 38948 16100
rect 38892 16046 38894 16098
rect 38894 16046 38946 16098
rect 38946 16046 38948 16098
rect 38892 16044 38948 16046
rect 38780 15148 38836 15204
rect 38780 14812 38836 14868
rect 38668 14028 38724 14084
rect 38892 13804 38948 13860
rect 39004 16380 39060 16436
rect 38332 11676 38388 11732
rect 38556 13580 38612 13636
rect 38892 12124 38948 12180
rect 39564 15148 39620 15204
rect 39340 14924 39396 14980
rect 39340 14364 39396 14420
rect 39004 12012 39060 12068
rect 39116 13356 39172 13412
rect 39004 11506 39060 11508
rect 39004 11454 39006 11506
rect 39006 11454 39058 11506
rect 39058 11454 39060 11506
rect 39004 11452 39060 11454
rect 39228 12796 39284 12852
rect 39452 12684 39508 12740
rect 39116 11340 39172 11396
rect 39340 12012 39396 12068
rect 38780 9324 38836 9380
rect 38444 8988 38500 9044
rect 38668 9042 38724 9044
rect 38668 8990 38670 9042
rect 38670 8990 38722 9042
rect 38722 8990 38724 9042
rect 38668 8988 38724 8990
rect 38332 8370 38388 8372
rect 38332 8318 38334 8370
rect 38334 8318 38386 8370
rect 38386 8318 38388 8370
rect 38332 8316 38388 8318
rect 38444 7420 38500 7476
rect 39004 10892 39060 10948
rect 37996 6300 38052 6356
rect 38108 5852 38164 5908
rect 37884 5068 37940 5124
rect 37996 5010 38052 5012
rect 37996 4958 37998 5010
rect 37998 4958 38050 5010
rect 38050 4958 38052 5010
rect 37996 4956 38052 4958
rect 38444 6802 38500 6804
rect 38444 6750 38446 6802
rect 38446 6750 38498 6802
rect 38498 6750 38500 6802
rect 38444 6748 38500 6750
rect 39340 10332 39396 10388
rect 39788 12684 39844 12740
rect 39676 12012 39732 12068
rect 39452 9548 39508 9604
rect 39452 9212 39508 9268
rect 39340 7474 39396 7476
rect 39340 7422 39342 7474
rect 39342 7422 39394 7474
rect 39394 7422 39396 7474
rect 39340 7420 39396 7422
rect 40236 23436 40292 23492
rect 40236 23154 40292 23156
rect 40236 23102 40238 23154
rect 40238 23102 40290 23154
rect 40290 23102 40292 23154
rect 40236 23100 40292 23102
rect 40460 22482 40516 22484
rect 40460 22430 40462 22482
rect 40462 22430 40514 22482
rect 40514 22430 40516 22482
rect 40460 22428 40516 22430
rect 41468 25788 41524 25844
rect 43932 33516 43988 33572
rect 43932 33292 43988 33348
rect 44380 34076 44436 34132
rect 44716 34748 44772 34804
rect 44828 34130 44884 34132
rect 44828 34078 44830 34130
rect 44830 34078 44882 34130
rect 44882 34078 44884 34130
rect 44828 34076 44884 34078
rect 45276 35644 45332 35700
rect 45388 36316 45444 36372
rect 45948 37938 46004 37940
rect 45948 37886 45950 37938
rect 45950 37886 46002 37938
rect 46002 37886 46004 37938
rect 45948 37884 46004 37886
rect 45500 35756 45556 35812
rect 45500 35420 45556 35476
rect 45052 35084 45108 35140
rect 44268 33740 44324 33796
rect 43260 32396 43316 32452
rect 43372 32844 43428 32900
rect 42588 30828 42644 30884
rect 42476 29820 42532 29876
rect 42364 28252 42420 28308
rect 42700 29148 42756 29204
rect 43260 31778 43316 31780
rect 43260 31726 43262 31778
rect 43262 31726 43314 31778
rect 43314 31726 43316 31778
rect 43260 31724 43316 31726
rect 43260 31388 43316 31444
rect 43148 28924 43204 28980
rect 43484 32562 43540 32564
rect 43484 32510 43486 32562
rect 43486 32510 43538 32562
rect 43538 32510 43540 32562
rect 43484 32508 43540 32510
rect 44464 33738 44520 33740
rect 44464 33686 44466 33738
rect 44466 33686 44518 33738
rect 44518 33686 44520 33738
rect 44464 33684 44520 33686
rect 44568 33738 44624 33740
rect 44568 33686 44570 33738
rect 44570 33686 44622 33738
rect 44622 33686 44624 33738
rect 44568 33684 44624 33686
rect 44672 33738 44728 33740
rect 44672 33686 44674 33738
rect 44674 33686 44726 33738
rect 44726 33686 44728 33738
rect 44672 33684 44728 33686
rect 44828 33628 44884 33684
rect 44380 33346 44436 33348
rect 44380 33294 44382 33346
rect 44382 33294 44434 33346
rect 44434 33294 44436 33346
rect 44380 33292 44436 33294
rect 43804 32954 43860 32956
rect 43804 32902 43806 32954
rect 43806 32902 43858 32954
rect 43858 32902 43860 32954
rect 43804 32900 43860 32902
rect 43908 32954 43964 32956
rect 43908 32902 43910 32954
rect 43910 32902 43962 32954
rect 43962 32902 43964 32954
rect 43908 32900 43964 32902
rect 44012 32954 44068 32956
rect 44012 32902 44014 32954
rect 44014 32902 44066 32954
rect 44066 32902 44068 32954
rect 44268 32956 44324 33012
rect 44012 32900 44068 32902
rect 43596 32060 43652 32116
rect 43596 31836 43652 31892
rect 44268 32508 44324 32564
rect 44492 32508 44548 32564
rect 45052 33740 45108 33796
rect 45052 33516 45108 33572
rect 44940 32508 44996 32564
rect 45052 32956 45108 33012
rect 44464 32170 44520 32172
rect 44464 32118 44466 32170
rect 44466 32118 44518 32170
rect 44518 32118 44520 32170
rect 44464 32116 44520 32118
rect 44568 32170 44624 32172
rect 44568 32118 44570 32170
rect 44570 32118 44622 32170
rect 44622 32118 44624 32170
rect 44568 32116 44624 32118
rect 44672 32170 44728 32172
rect 44672 32118 44674 32170
rect 44674 32118 44726 32170
rect 44726 32118 44728 32170
rect 44672 32116 44728 32118
rect 44492 31500 44548 31556
rect 43804 31386 43860 31388
rect 43804 31334 43806 31386
rect 43806 31334 43858 31386
rect 43858 31334 43860 31386
rect 43804 31332 43860 31334
rect 43908 31386 43964 31388
rect 43908 31334 43910 31386
rect 43910 31334 43962 31386
rect 43962 31334 43964 31386
rect 43908 31332 43964 31334
rect 44012 31386 44068 31388
rect 44012 31334 44014 31386
rect 44014 31334 44066 31386
rect 44066 31334 44068 31386
rect 44012 31332 44068 31334
rect 43484 31164 43540 31220
rect 44156 30828 44212 30884
rect 43596 30770 43652 30772
rect 43596 30718 43598 30770
rect 43598 30718 43650 30770
rect 43650 30718 43652 30770
rect 43596 30716 43652 30718
rect 43804 29818 43860 29820
rect 43804 29766 43806 29818
rect 43806 29766 43858 29818
rect 43858 29766 43860 29818
rect 43804 29764 43860 29766
rect 43908 29818 43964 29820
rect 43908 29766 43910 29818
rect 43910 29766 43962 29818
rect 43962 29766 43964 29818
rect 43908 29764 43964 29766
rect 44012 29818 44068 29820
rect 44012 29766 44014 29818
rect 44014 29766 44066 29818
rect 44066 29766 44068 29818
rect 44012 29764 44068 29766
rect 44156 29708 44212 29764
rect 44716 30882 44772 30884
rect 44716 30830 44718 30882
rect 44718 30830 44770 30882
rect 44770 30830 44772 30882
rect 44716 30828 44772 30830
rect 44464 30602 44520 30604
rect 44464 30550 44466 30602
rect 44466 30550 44518 30602
rect 44518 30550 44520 30602
rect 44464 30548 44520 30550
rect 44568 30602 44624 30604
rect 44568 30550 44570 30602
rect 44570 30550 44622 30602
rect 44622 30550 44624 30602
rect 44568 30548 44624 30550
rect 44672 30602 44728 30604
rect 44672 30550 44674 30602
rect 44674 30550 44726 30602
rect 44726 30550 44728 30602
rect 44672 30548 44728 30550
rect 44268 30156 44324 30212
rect 44492 30268 44548 30324
rect 44268 29372 44324 29428
rect 43372 28924 43428 28980
rect 43484 29036 43540 29092
rect 42588 28028 42644 28084
rect 42252 27186 42308 27188
rect 42252 27134 42254 27186
rect 42254 27134 42306 27186
rect 42306 27134 42308 27186
rect 42252 27132 42308 27134
rect 42028 27020 42084 27076
rect 41692 26124 41748 26180
rect 41804 25676 41860 25732
rect 42028 25730 42084 25732
rect 42028 25678 42030 25730
rect 42030 25678 42082 25730
rect 42082 25678 42084 25730
rect 42028 25676 42084 25678
rect 41580 25340 41636 25396
rect 41804 25228 41860 25284
rect 41580 25004 41636 25060
rect 41020 24108 41076 24164
rect 41356 24556 41412 24612
rect 40796 23548 40852 23604
rect 41468 24220 41524 24276
rect 41468 23884 41524 23940
rect 41356 23548 41412 23604
rect 41692 24444 41748 24500
rect 41580 22988 41636 23044
rect 41692 24220 41748 24276
rect 41916 24834 41972 24836
rect 41916 24782 41918 24834
rect 41918 24782 41970 24834
rect 41970 24782 41972 24834
rect 41916 24780 41972 24782
rect 42140 25004 42196 25060
rect 41804 23996 41860 24052
rect 41916 24108 41972 24164
rect 41580 22652 41636 22708
rect 40460 21868 40516 21924
rect 40348 21644 40404 21700
rect 40236 20636 40292 20692
rect 40908 21420 40964 21476
rect 40796 20972 40852 21028
rect 40684 20914 40740 20916
rect 40684 20862 40686 20914
rect 40686 20862 40738 20914
rect 40738 20862 40740 20914
rect 40684 20860 40740 20862
rect 40348 20748 40404 20804
rect 40796 20802 40852 20804
rect 40796 20750 40798 20802
rect 40798 20750 40850 20802
rect 40850 20750 40852 20802
rect 40796 20748 40852 20750
rect 40572 20636 40628 20692
rect 40908 20524 40964 20580
rect 41916 23436 41972 23492
rect 42028 23884 42084 23940
rect 41916 23100 41972 23156
rect 41916 22652 41972 22708
rect 41132 21420 41188 21476
rect 41020 20636 41076 20692
rect 40124 18060 40180 18116
rect 40460 19180 40516 19236
rect 40572 19122 40628 19124
rect 40572 19070 40574 19122
rect 40574 19070 40626 19122
rect 40626 19070 40628 19122
rect 40572 19068 40628 19070
rect 40572 18674 40628 18676
rect 40572 18622 40574 18674
rect 40574 18622 40626 18674
rect 40626 18622 40628 18674
rect 40572 18620 40628 18622
rect 41132 21084 41188 21140
rect 41356 21756 41412 21812
rect 42028 22428 42084 22484
rect 42140 21868 42196 21924
rect 41916 21756 41972 21812
rect 42476 25676 42532 25732
rect 42476 24780 42532 24836
rect 43708 28754 43764 28756
rect 43708 28702 43710 28754
rect 43710 28702 43762 28754
rect 43762 28702 43764 28754
rect 43708 28700 43764 28702
rect 44464 29034 44520 29036
rect 44464 28982 44466 29034
rect 44466 28982 44518 29034
rect 44518 28982 44520 29034
rect 44464 28980 44520 28982
rect 44568 29034 44624 29036
rect 44568 28982 44570 29034
rect 44570 28982 44622 29034
rect 44622 28982 44624 29034
rect 44568 28980 44624 28982
rect 44672 29034 44728 29036
rect 44672 28982 44674 29034
rect 44674 28982 44726 29034
rect 44726 28982 44728 29034
rect 44672 28980 44728 28982
rect 44604 28476 44660 28532
rect 43484 27468 43540 27524
rect 43596 28364 43652 28420
rect 43260 27186 43316 27188
rect 43260 27134 43262 27186
rect 43262 27134 43314 27186
rect 43314 27134 43316 27186
rect 43260 27132 43316 27134
rect 42812 27074 42868 27076
rect 42812 27022 42814 27074
rect 42814 27022 42866 27074
rect 42866 27022 42868 27074
rect 42812 27020 42868 27022
rect 43260 26908 43316 26964
rect 44268 28364 44324 28420
rect 43804 28250 43860 28252
rect 43804 28198 43806 28250
rect 43806 28198 43858 28250
rect 43858 28198 43860 28250
rect 43804 28196 43860 28198
rect 43908 28250 43964 28252
rect 43908 28198 43910 28250
rect 43910 28198 43962 28250
rect 43962 28198 43964 28250
rect 43908 28196 43964 28198
rect 44012 28250 44068 28252
rect 44012 28198 44014 28250
rect 44014 28198 44066 28250
rect 44066 28198 44068 28250
rect 44012 28196 44068 28198
rect 43596 26908 43652 26964
rect 44156 27468 44212 27524
rect 43148 26796 43204 26852
rect 43804 26682 43860 26684
rect 43804 26630 43806 26682
rect 43806 26630 43858 26682
rect 43858 26630 43860 26682
rect 43804 26628 43860 26630
rect 43908 26682 43964 26684
rect 43908 26630 43910 26682
rect 43910 26630 43962 26682
rect 43962 26630 43964 26682
rect 43908 26628 43964 26630
rect 44012 26682 44068 26684
rect 44012 26630 44014 26682
rect 44014 26630 44066 26682
rect 44066 26630 44068 26682
rect 44012 26628 44068 26630
rect 43596 26460 43652 26516
rect 43372 26178 43428 26180
rect 43372 26126 43374 26178
rect 43374 26126 43426 26178
rect 43426 26126 43428 26178
rect 43372 26124 43428 26126
rect 43260 26012 43316 26068
rect 43484 26012 43540 26068
rect 42700 25618 42756 25620
rect 42700 25566 42702 25618
rect 42702 25566 42754 25618
rect 42754 25566 42756 25618
rect 42700 25564 42756 25566
rect 42700 25394 42756 25396
rect 42700 25342 42702 25394
rect 42702 25342 42754 25394
rect 42754 25342 42756 25394
rect 42700 25340 42756 25342
rect 43036 25452 43092 25508
rect 42924 25340 42980 25396
rect 42700 23436 42756 23492
rect 42924 22988 42980 23044
rect 42364 21756 42420 21812
rect 41356 21420 41412 21476
rect 41468 21026 41524 21028
rect 41468 20974 41470 21026
rect 41470 20974 41522 21026
rect 41522 20974 41524 21026
rect 41468 20972 41524 20974
rect 41468 20748 41524 20804
rect 41132 20300 41188 20356
rect 41244 20524 41300 20580
rect 41132 19852 41188 19908
rect 41020 18732 41076 18788
rect 41132 19068 41188 19124
rect 41804 21084 41860 21140
rect 41356 20018 41412 20020
rect 41356 19966 41358 20018
rect 41358 19966 41410 20018
rect 41410 19966 41412 20018
rect 41356 19964 41412 19966
rect 42364 20802 42420 20804
rect 42364 20750 42366 20802
rect 42366 20750 42418 20802
rect 42418 20750 42420 20802
rect 42364 20748 42420 20750
rect 41580 19404 41636 19460
rect 41916 20300 41972 20356
rect 41244 18844 41300 18900
rect 41804 18956 41860 19012
rect 41580 18450 41636 18452
rect 41580 18398 41582 18450
rect 41582 18398 41634 18450
rect 41634 18398 41636 18450
rect 41580 18396 41636 18398
rect 40796 17948 40852 18004
rect 40236 15932 40292 15988
rect 40460 15986 40516 15988
rect 40460 15934 40462 15986
rect 40462 15934 40514 15986
rect 40514 15934 40516 15986
rect 40460 15932 40516 15934
rect 41020 17666 41076 17668
rect 41020 17614 41022 17666
rect 41022 17614 41074 17666
rect 41074 17614 41076 17666
rect 41020 17612 41076 17614
rect 41020 17164 41076 17220
rect 40908 16882 40964 16884
rect 40908 16830 40910 16882
rect 40910 16830 40962 16882
rect 40962 16830 40964 16882
rect 40908 16828 40964 16830
rect 40236 15596 40292 15652
rect 40236 12850 40292 12852
rect 40236 12798 40238 12850
rect 40238 12798 40290 12850
rect 40290 12798 40292 12850
rect 40236 12796 40292 12798
rect 40460 15260 40516 15316
rect 40684 15314 40740 15316
rect 40684 15262 40686 15314
rect 40686 15262 40738 15314
rect 40738 15262 40740 15314
rect 40684 15260 40740 15262
rect 40572 14140 40628 14196
rect 40348 11564 40404 11620
rect 40460 13468 40516 13524
rect 40236 11228 40292 11284
rect 40124 11116 40180 11172
rect 40460 10556 40516 10612
rect 39900 10444 39956 10500
rect 40124 10444 40180 10500
rect 39900 8988 39956 9044
rect 39900 8316 39956 8372
rect 39564 6690 39620 6692
rect 39564 6638 39566 6690
rect 39566 6638 39618 6690
rect 39618 6638 39620 6690
rect 39564 6636 39620 6638
rect 39676 6300 39732 6356
rect 38444 5628 38500 5684
rect 38108 4396 38164 4452
rect 38332 4450 38388 4452
rect 38332 4398 38334 4450
rect 38334 4398 38386 4450
rect 38386 4398 38388 4450
rect 38332 4396 38388 4398
rect 37996 3778 38052 3780
rect 37996 3726 37998 3778
rect 37998 3726 38050 3778
rect 38050 3726 38052 3778
rect 37996 3724 38052 3726
rect 37884 3442 37940 3444
rect 37884 3390 37886 3442
rect 37886 3390 37938 3442
rect 37938 3390 37940 3442
rect 37884 3388 37940 3390
rect 37996 2546 38052 2548
rect 37996 2494 37998 2546
rect 37998 2494 38050 2546
rect 38050 2494 38052 2546
rect 37996 2492 38052 2494
rect 37884 2268 37940 2324
rect 38220 2210 38276 2212
rect 38220 2158 38222 2210
rect 38222 2158 38274 2210
rect 38274 2158 38276 2210
rect 38220 2156 38276 2158
rect 37884 2098 37940 2100
rect 37884 2046 37886 2098
rect 37886 2046 37938 2098
rect 37938 2046 37940 2098
rect 37884 2044 37940 2046
rect 37660 1202 37716 1204
rect 37660 1150 37662 1202
rect 37662 1150 37714 1202
rect 37714 1150 37716 1202
rect 37660 1148 37716 1150
rect 37324 812 37380 868
rect 37436 924 37492 980
rect 37212 364 37268 420
rect 38556 5010 38612 5012
rect 38556 4958 38558 5010
rect 38558 4958 38610 5010
rect 38610 4958 38612 5010
rect 38556 4956 38612 4958
rect 38668 4844 38724 4900
rect 39340 5628 39396 5684
rect 39116 4898 39172 4900
rect 39116 4846 39118 4898
rect 39118 4846 39170 4898
rect 39170 4846 39172 4898
rect 39116 4844 39172 4846
rect 38780 4396 38836 4452
rect 39900 7474 39956 7476
rect 39900 7422 39902 7474
rect 39902 7422 39954 7474
rect 39954 7422 39956 7474
rect 39900 7420 39956 7422
rect 40348 9436 40404 9492
rect 40236 8652 40292 8708
rect 40460 7644 40516 7700
rect 41244 17388 41300 17444
rect 41468 17724 41524 17780
rect 41468 17164 41524 17220
rect 41468 16380 41524 16436
rect 41132 15484 41188 15540
rect 41580 15932 41636 15988
rect 41020 14812 41076 14868
rect 43260 25452 43316 25508
rect 43260 25004 43316 25060
rect 43148 24050 43204 24052
rect 43148 23998 43150 24050
rect 43150 23998 43202 24050
rect 43202 23998 43204 24050
rect 43148 23996 43204 23998
rect 43148 22764 43204 22820
rect 43036 22204 43092 22260
rect 43036 21868 43092 21924
rect 42924 21196 42980 21252
rect 43148 21420 43204 21476
rect 42812 20636 42868 20692
rect 42140 19458 42196 19460
rect 42140 19406 42142 19458
rect 42142 19406 42194 19458
rect 42194 19406 42196 19458
rect 42140 19404 42196 19406
rect 42028 19068 42084 19124
rect 42364 19404 42420 19460
rect 42252 18396 42308 18452
rect 42364 19068 42420 19124
rect 41916 18172 41972 18228
rect 42140 18060 42196 18116
rect 41916 17052 41972 17108
rect 41804 15372 41860 15428
rect 41916 16044 41972 16100
rect 41580 14476 41636 14532
rect 41804 14140 41860 14196
rect 40908 13692 40964 13748
rect 41580 13692 41636 13748
rect 41468 13580 41524 13636
rect 40908 13020 40964 13076
rect 40796 12178 40852 12180
rect 40796 12126 40798 12178
rect 40798 12126 40850 12178
rect 40850 12126 40852 12178
rect 40796 12124 40852 12126
rect 41020 12962 41076 12964
rect 41020 12910 41022 12962
rect 41022 12910 41074 12962
rect 41074 12910 41076 12962
rect 41020 12908 41076 12910
rect 41020 11676 41076 11732
rect 40908 11452 40964 11508
rect 41132 11452 41188 11508
rect 41020 10556 41076 10612
rect 41132 10220 41188 10276
rect 41020 9324 41076 9380
rect 41020 8652 41076 8708
rect 40908 8540 40964 8596
rect 40236 6578 40292 6580
rect 40236 6526 40238 6578
rect 40238 6526 40290 6578
rect 40290 6526 40292 6578
rect 40236 6524 40292 6526
rect 40124 5794 40180 5796
rect 40124 5742 40126 5794
rect 40126 5742 40178 5794
rect 40178 5742 40180 5794
rect 40124 5740 40180 5742
rect 40348 5180 40404 5236
rect 40796 7980 40852 8036
rect 41132 8540 41188 8596
rect 41020 8258 41076 8260
rect 41020 8206 41022 8258
rect 41022 8206 41074 8258
rect 41074 8206 41076 8258
rect 41020 8204 41076 8206
rect 41804 12460 41860 12516
rect 41468 10050 41524 10052
rect 41468 9998 41470 10050
rect 41470 9998 41522 10050
rect 41522 9998 41524 10050
rect 41468 9996 41524 9998
rect 41580 8316 41636 8372
rect 41356 8034 41412 8036
rect 41356 7982 41358 8034
rect 41358 7982 41410 8034
rect 41410 7982 41412 8034
rect 41356 7980 41412 7982
rect 41804 9884 41860 9940
rect 41692 7868 41748 7924
rect 41804 8316 41860 8372
rect 41244 7308 41300 7364
rect 41580 7308 41636 7364
rect 40572 6690 40628 6692
rect 40572 6638 40574 6690
rect 40574 6638 40626 6690
rect 40626 6638 40628 6690
rect 40572 6636 40628 6638
rect 40796 6636 40852 6692
rect 40460 5068 40516 5124
rect 38668 3724 38724 3780
rect 40012 3724 40068 3780
rect 38556 2770 38612 2772
rect 38556 2718 38558 2770
rect 38558 2718 38610 2770
rect 38610 2718 38612 2770
rect 38556 2716 38612 2718
rect 39228 3276 39284 3332
rect 39340 2770 39396 2772
rect 39340 2718 39342 2770
rect 39342 2718 39394 2770
rect 39394 2718 39396 2770
rect 39340 2716 39396 2718
rect 39564 2098 39620 2100
rect 39564 2046 39566 2098
rect 39566 2046 39618 2098
rect 39618 2046 39620 2098
rect 39564 2044 39620 2046
rect 39452 1484 39508 1540
rect 38780 1372 38836 1428
rect 37996 252 38052 308
rect 38332 700 38388 756
rect 39452 1202 39508 1204
rect 39452 1150 39454 1202
rect 39454 1150 39506 1202
rect 39506 1150 39508 1202
rect 39452 1148 39508 1150
rect 39116 476 39172 532
rect 39228 364 39284 420
rect 40572 3442 40628 3444
rect 40572 3390 40574 3442
rect 40574 3390 40626 3442
rect 40626 3390 40628 3442
rect 40572 3388 40628 3390
rect 40012 2994 40068 2996
rect 40012 2942 40014 2994
rect 40014 2942 40066 2994
rect 40066 2942 40068 2994
rect 40012 2940 40068 2942
rect 41020 6412 41076 6468
rect 41804 7084 41860 7140
rect 41580 6748 41636 6804
rect 42140 16716 42196 16772
rect 42028 11506 42084 11508
rect 42028 11454 42030 11506
rect 42030 11454 42082 11506
rect 42082 11454 42084 11506
rect 42028 11452 42084 11454
rect 42028 10498 42084 10500
rect 42028 10446 42030 10498
rect 42030 10446 42082 10498
rect 42082 10446 42084 10498
rect 42028 10444 42084 10446
rect 42364 16604 42420 16660
rect 42364 15260 42420 15316
rect 42700 20018 42756 20020
rect 42700 19966 42702 20018
rect 42702 19966 42754 20018
rect 42754 19966 42756 20018
rect 42700 19964 42756 19966
rect 42588 19234 42644 19236
rect 42588 19182 42590 19234
rect 42590 19182 42642 19234
rect 42642 19182 42644 19234
rect 42588 19180 42644 19182
rect 43036 20914 43092 20916
rect 43036 20862 43038 20914
rect 43038 20862 43090 20914
rect 43090 20862 43092 20914
rect 43036 20860 43092 20862
rect 42924 19740 42980 19796
rect 42700 19068 42756 19124
rect 42812 19458 42868 19460
rect 42812 19406 42814 19458
rect 42814 19406 42866 19458
rect 42866 19406 42868 19458
rect 42812 19404 42868 19406
rect 43036 19404 43092 19460
rect 42812 18620 42868 18676
rect 42588 17106 42644 17108
rect 42588 17054 42590 17106
rect 42590 17054 42642 17106
rect 42642 17054 42644 17106
rect 42588 17052 42644 17054
rect 43036 18508 43092 18564
rect 43708 26124 43764 26180
rect 43708 25900 43764 25956
rect 44044 25564 44100 25620
rect 44156 25452 44212 25508
rect 44492 28028 44548 28084
rect 44716 28140 44772 28196
rect 44716 27804 44772 27860
rect 44464 27466 44520 27468
rect 44464 27414 44466 27466
rect 44466 27414 44518 27466
rect 44518 27414 44520 27466
rect 44464 27412 44520 27414
rect 44568 27466 44624 27468
rect 44568 27414 44570 27466
rect 44570 27414 44622 27466
rect 44622 27414 44624 27466
rect 44568 27412 44624 27414
rect 44672 27466 44728 27468
rect 44672 27414 44674 27466
rect 44674 27414 44726 27466
rect 44726 27414 44728 27466
rect 44672 27412 44728 27414
rect 44380 26460 44436 26516
rect 44604 26236 44660 26292
rect 45052 32172 45108 32228
rect 45276 32732 45332 32788
rect 45500 34524 45556 34580
rect 45612 34354 45668 34356
rect 45612 34302 45614 34354
rect 45614 34302 45666 34354
rect 45666 34302 45668 34354
rect 45612 34300 45668 34302
rect 45612 33516 45668 33572
rect 45612 33068 45668 33124
rect 45388 31890 45444 31892
rect 45388 31838 45390 31890
rect 45390 31838 45442 31890
rect 45442 31838 45444 31890
rect 45388 31836 45444 31838
rect 44940 29932 44996 29988
rect 44940 29148 44996 29204
rect 45052 28364 45108 28420
rect 45164 30268 45220 30324
rect 45052 27858 45108 27860
rect 45052 27806 45054 27858
rect 45054 27806 45106 27858
rect 45106 27806 45108 27858
rect 45052 27804 45108 27806
rect 44940 26572 44996 26628
rect 45276 29932 45332 29988
rect 45612 30940 45668 30996
rect 45612 30492 45668 30548
rect 45612 30156 45668 30212
rect 45276 28700 45332 28756
rect 45500 28924 45556 28980
rect 44828 26236 44884 26292
rect 44940 26348 44996 26404
rect 44464 25898 44520 25900
rect 44464 25846 44466 25898
rect 44466 25846 44518 25898
rect 44518 25846 44520 25898
rect 44464 25844 44520 25846
rect 44568 25898 44624 25900
rect 44568 25846 44570 25898
rect 44570 25846 44622 25898
rect 44622 25846 44624 25898
rect 44568 25844 44624 25846
rect 44672 25898 44728 25900
rect 44672 25846 44674 25898
rect 44674 25846 44726 25898
rect 44726 25846 44728 25898
rect 44672 25844 44728 25846
rect 43804 25114 43860 25116
rect 43804 25062 43806 25114
rect 43806 25062 43858 25114
rect 43858 25062 43860 25114
rect 43804 25060 43860 25062
rect 43908 25114 43964 25116
rect 43908 25062 43910 25114
rect 43910 25062 43962 25114
rect 43962 25062 43964 25114
rect 43908 25060 43964 25062
rect 44012 25114 44068 25116
rect 44012 25062 44014 25114
rect 44014 25062 44066 25114
rect 44066 25062 44068 25114
rect 44012 25060 44068 25062
rect 44156 25004 44212 25060
rect 44156 24780 44212 24836
rect 43596 24668 43652 24724
rect 43596 24332 43652 24388
rect 44464 24330 44520 24332
rect 44464 24278 44466 24330
rect 44466 24278 44518 24330
rect 44518 24278 44520 24330
rect 44464 24276 44520 24278
rect 44568 24330 44624 24332
rect 44568 24278 44570 24330
rect 44570 24278 44622 24330
rect 44622 24278 44624 24330
rect 44568 24276 44624 24278
rect 44672 24330 44728 24332
rect 44672 24278 44674 24330
rect 44674 24278 44726 24330
rect 44726 24278 44728 24330
rect 44672 24276 44728 24278
rect 44380 23996 44436 24052
rect 43484 23548 43540 23604
rect 43804 23546 43860 23548
rect 43804 23494 43806 23546
rect 43806 23494 43858 23546
rect 43858 23494 43860 23546
rect 43804 23492 43860 23494
rect 43908 23546 43964 23548
rect 43908 23494 43910 23546
rect 43910 23494 43962 23546
rect 43962 23494 43964 23546
rect 43908 23492 43964 23494
rect 44012 23546 44068 23548
rect 44012 23494 44014 23546
rect 44014 23494 44066 23546
rect 44066 23494 44068 23546
rect 44012 23492 44068 23494
rect 43596 23100 43652 23156
rect 43484 22428 43540 22484
rect 43484 21868 43540 21924
rect 43372 19964 43428 20020
rect 43484 20748 43540 20804
rect 43148 17948 43204 18004
rect 43260 18396 43316 18452
rect 43260 17276 43316 17332
rect 44156 22540 44212 22596
rect 43804 21978 43860 21980
rect 43804 21926 43806 21978
rect 43806 21926 43858 21978
rect 43858 21926 43860 21978
rect 43804 21924 43860 21926
rect 43908 21978 43964 21980
rect 43908 21926 43910 21978
rect 43910 21926 43962 21978
rect 43962 21926 43964 21978
rect 43908 21924 43964 21926
rect 44012 21978 44068 21980
rect 44012 21926 44014 21978
rect 44014 21926 44066 21978
rect 44066 21926 44068 21978
rect 44012 21924 44068 21926
rect 44464 22762 44520 22764
rect 44464 22710 44466 22762
rect 44466 22710 44518 22762
rect 44518 22710 44520 22762
rect 44464 22708 44520 22710
rect 44568 22762 44624 22764
rect 44568 22710 44570 22762
rect 44570 22710 44622 22762
rect 44622 22710 44624 22762
rect 44568 22708 44624 22710
rect 44672 22762 44728 22764
rect 44672 22710 44674 22762
rect 44674 22710 44726 22762
rect 44726 22710 44728 22762
rect 44672 22708 44728 22710
rect 44380 22540 44436 22596
rect 44380 21756 44436 21812
rect 44828 21756 44884 21812
rect 44828 21308 44884 21364
rect 44464 21194 44520 21196
rect 44464 21142 44466 21194
rect 44466 21142 44518 21194
rect 44518 21142 44520 21194
rect 44464 21140 44520 21142
rect 44568 21194 44624 21196
rect 44568 21142 44570 21194
rect 44570 21142 44622 21194
rect 44622 21142 44624 21194
rect 44568 21140 44624 21142
rect 44672 21194 44728 21196
rect 44672 21142 44674 21194
rect 44674 21142 44726 21194
rect 44726 21142 44728 21194
rect 44672 21140 44728 21142
rect 43804 20410 43860 20412
rect 43804 20358 43806 20410
rect 43806 20358 43858 20410
rect 43858 20358 43860 20410
rect 43804 20356 43860 20358
rect 43908 20410 43964 20412
rect 43908 20358 43910 20410
rect 43910 20358 43962 20410
rect 43962 20358 43964 20410
rect 43908 20356 43964 20358
rect 44012 20410 44068 20412
rect 44012 20358 44014 20410
rect 44014 20358 44066 20410
rect 44066 20358 44068 20410
rect 44012 20356 44068 20358
rect 44268 19852 44324 19908
rect 43596 19404 43652 19460
rect 43708 19180 43764 19236
rect 44156 19628 44212 19684
rect 44268 19516 44324 19572
rect 44464 19626 44520 19628
rect 44464 19574 44466 19626
rect 44466 19574 44518 19626
rect 44518 19574 44520 19626
rect 44464 19572 44520 19574
rect 44568 19626 44624 19628
rect 44568 19574 44570 19626
rect 44570 19574 44622 19626
rect 44622 19574 44624 19626
rect 44568 19572 44624 19574
rect 44672 19626 44728 19628
rect 44672 19574 44674 19626
rect 44674 19574 44726 19626
rect 44726 19574 44728 19626
rect 44672 19572 44728 19574
rect 43804 18842 43860 18844
rect 43804 18790 43806 18842
rect 43806 18790 43858 18842
rect 43858 18790 43860 18842
rect 43804 18788 43860 18790
rect 43908 18842 43964 18844
rect 43908 18790 43910 18842
rect 43910 18790 43962 18842
rect 43962 18790 43964 18842
rect 43908 18788 43964 18790
rect 44012 18842 44068 18844
rect 44012 18790 44014 18842
rect 44014 18790 44066 18842
rect 44066 18790 44068 18842
rect 44156 18844 44212 18900
rect 44012 18788 44068 18790
rect 43932 18620 43988 18676
rect 43708 18508 43764 18564
rect 44828 18508 44884 18564
rect 45948 35644 46004 35700
rect 46060 36428 46116 36484
rect 45836 35084 45892 35140
rect 45948 35196 46004 35252
rect 45836 33740 45892 33796
rect 45836 33292 45892 33348
rect 46060 34130 46116 34132
rect 46060 34078 46062 34130
rect 46062 34078 46114 34130
rect 46114 34078 46116 34130
rect 46060 34076 46116 34078
rect 45948 32786 46004 32788
rect 45948 32734 45950 32786
rect 45950 32734 46002 32786
rect 46002 32734 46004 32786
rect 45948 32732 46004 32734
rect 45836 31276 45892 31332
rect 45948 31724 46004 31780
rect 45724 28812 45780 28868
rect 45612 27468 45668 27524
rect 45724 28642 45780 28644
rect 45724 28590 45726 28642
rect 45726 28590 45778 28642
rect 45778 28590 45780 28642
rect 45724 28588 45780 28590
rect 45500 27298 45556 27300
rect 45500 27246 45502 27298
rect 45502 27246 45554 27298
rect 45554 27246 45556 27298
rect 45500 27244 45556 27246
rect 45724 27244 45780 27300
rect 45388 26908 45444 26964
rect 45276 26572 45332 26628
rect 45500 27020 45556 27076
rect 45612 26290 45668 26292
rect 45612 26238 45614 26290
rect 45614 26238 45666 26290
rect 45666 26238 45668 26290
rect 45612 26236 45668 26238
rect 46284 37378 46340 37380
rect 46284 37326 46286 37378
rect 46286 37326 46338 37378
rect 46338 37326 46340 37378
rect 46284 37324 46340 37326
rect 46396 35308 46452 35364
rect 46284 35084 46340 35140
rect 46732 38108 46788 38164
rect 46844 38780 46900 38836
rect 46732 37938 46788 37940
rect 46732 37886 46734 37938
rect 46734 37886 46786 37938
rect 46786 37886 46788 37938
rect 46732 37884 46788 37886
rect 46620 35698 46676 35700
rect 46620 35646 46622 35698
rect 46622 35646 46674 35698
rect 46674 35646 46676 35698
rect 46620 35644 46676 35646
rect 46732 35756 46788 35812
rect 46508 35084 46564 35140
rect 46508 34748 46564 34804
rect 46620 34636 46676 34692
rect 46508 34188 46564 34244
rect 46284 34018 46340 34020
rect 46284 33966 46286 34018
rect 46286 33966 46338 34018
rect 46338 33966 46340 34018
rect 46284 33964 46340 33966
rect 46396 33516 46452 33572
rect 46620 33180 46676 33236
rect 46732 32956 46788 33012
rect 46508 32844 46564 32900
rect 46508 32396 46564 32452
rect 46732 32396 46788 32452
rect 46620 32172 46676 32228
rect 46620 31554 46676 31556
rect 46620 31502 46622 31554
rect 46622 31502 46674 31554
rect 46674 31502 46676 31554
rect 46620 31500 46676 31502
rect 46172 30604 46228 30660
rect 46284 30380 46340 30436
rect 46172 30210 46228 30212
rect 46172 30158 46174 30210
rect 46174 30158 46226 30210
rect 46226 30158 46228 30210
rect 46172 30156 46228 30158
rect 46060 29148 46116 29204
rect 45948 28700 46004 28756
rect 46172 28812 46228 28868
rect 46620 30156 46676 30212
rect 47516 44882 47572 44884
rect 47516 44830 47518 44882
rect 47518 44830 47570 44882
rect 47570 44830 47572 44882
rect 47516 44828 47572 44830
rect 47068 44380 47124 44436
rect 47404 43484 47460 43540
rect 47180 43260 47236 43316
rect 47068 42754 47124 42756
rect 47068 42702 47070 42754
rect 47070 42702 47122 42754
rect 47122 42702 47124 42754
rect 47068 42700 47124 42702
rect 47292 42812 47348 42868
rect 47852 46620 47908 46676
rect 48412 48748 48468 48804
rect 47740 45388 47796 45444
rect 47852 43426 47908 43428
rect 47852 43374 47854 43426
rect 47854 43374 47906 43426
rect 47906 43374 47908 43426
rect 47852 43372 47908 43374
rect 47852 42812 47908 42868
rect 47740 42476 47796 42532
rect 47404 41916 47460 41972
rect 47404 41692 47460 41748
rect 47740 40684 47796 40740
rect 47628 40124 47684 40180
rect 47068 39900 47124 39956
rect 47516 39900 47572 39956
rect 47404 39676 47460 39732
rect 47180 39004 47236 39060
rect 46956 38722 47012 38724
rect 46956 38670 46958 38722
rect 46958 38670 47010 38722
rect 47010 38670 47012 38722
rect 46956 38668 47012 38670
rect 47292 38162 47348 38164
rect 47292 38110 47294 38162
rect 47294 38110 47346 38162
rect 47346 38110 47348 38162
rect 47292 38108 47348 38110
rect 47292 37324 47348 37380
rect 47628 39564 47684 39620
rect 47740 39788 47796 39844
rect 47516 38780 47572 38836
rect 47516 38220 47572 38276
rect 47516 37660 47572 37716
rect 46956 36482 47012 36484
rect 46956 36430 46958 36482
rect 46958 36430 47010 36482
rect 47010 36430 47012 36482
rect 46956 36428 47012 36430
rect 46956 35756 47012 35812
rect 47516 35756 47572 35812
rect 47628 35980 47684 36036
rect 47516 35420 47572 35476
rect 47180 35138 47236 35140
rect 47180 35086 47182 35138
rect 47182 35086 47234 35138
rect 47234 35086 47236 35138
rect 47180 35084 47236 35086
rect 46956 34300 47012 34356
rect 47404 34636 47460 34692
rect 47628 34636 47684 34692
rect 47516 34300 47572 34356
rect 48076 47682 48132 47684
rect 48076 47630 48078 47682
rect 48078 47630 48130 47682
rect 48130 47630 48132 47682
rect 48076 47628 48132 47630
rect 48300 47458 48356 47460
rect 48300 47406 48302 47458
rect 48302 47406 48354 47458
rect 48354 47406 48356 47458
rect 48300 47404 48356 47406
rect 48188 47346 48244 47348
rect 48188 47294 48190 47346
rect 48190 47294 48242 47346
rect 48242 47294 48244 47346
rect 48188 47292 48244 47294
rect 48524 47404 48580 47460
rect 48412 45836 48468 45892
rect 48300 45724 48356 45780
rect 48188 44156 48244 44212
rect 48076 41692 48132 41748
rect 48860 49026 48916 49028
rect 48860 48974 48862 49026
rect 48862 48974 48914 49026
rect 48914 48974 48916 49026
rect 48860 48972 48916 48974
rect 48860 48748 48916 48804
rect 48636 45164 48692 45220
rect 48524 44380 48580 44436
rect 48412 43260 48468 43316
rect 48524 44210 48580 44212
rect 48524 44158 48526 44210
rect 48526 44158 48578 44210
rect 48578 44158 48580 44210
rect 48524 44156 48580 44158
rect 48748 44156 48804 44212
rect 49644 51602 49700 51604
rect 49644 51550 49646 51602
rect 49646 51550 49698 51602
rect 49698 51550 49700 51602
rect 49644 51548 49700 51550
rect 49644 50540 49700 50596
rect 50092 54236 50148 54292
rect 50540 53452 50596 53508
rect 49868 52162 49924 52164
rect 49868 52110 49870 52162
rect 49870 52110 49922 52162
rect 49922 52110 49924 52162
rect 49868 52108 49924 52110
rect 49868 51490 49924 51492
rect 49868 51438 49870 51490
rect 49870 51438 49922 51490
rect 49922 51438 49924 51490
rect 49868 51436 49924 51438
rect 50204 51548 50260 51604
rect 49868 51100 49924 51156
rect 49980 49980 50036 50036
rect 49532 49868 49588 49924
rect 50204 50764 50260 50820
rect 50092 49868 50148 49924
rect 49308 48972 49364 49028
rect 49420 48748 49476 48804
rect 49532 48412 49588 48468
rect 49196 47740 49252 47796
rect 48972 47404 49028 47460
rect 49196 47180 49252 47236
rect 48972 46508 49028 46564
rect 49532 47068 49588 47124
rect 49868 49420 49924 49476
rect 49644 46844 49700 46900
rect 49756 48972 49812 49028
rect 49868 48860 49924 48916
rect 49980 48412 50036 48468
rect 49868 47740 49924 47796
rect 50428 52108 50484 52164
rect 50764 53730 50820 53732
rect 50764 53678 50766 53730
rect 50766 53678 50818 53730
rect 50818 53678 50820 53730
rect 50764 53676 50820 53678
rect 51548 55858 51604 55860
rect 51548 55806 51550 55858
rect 51550 55806 51602 55858
rect 51602 55806 51604 55858
rect 51548 55804 51604 55806
rect 51324 55468 51380 55524
rect 51212 55356 51268 55412
rect 51324 54460 51380 54516
rect 51100 53004 51156 53060
rect 51212 52892 51268 52948
rect 50876 52722 50932 52724
rect 50876 52670 50878 52722
rect 50878 52670 50930 52722
rect 50930 52670 50932 52722
rect 50876 52668 50932 52670
rect 50652 52444 50708 52500
rect 51100 52444 51156 52500
rect 50540 50316 50596 50372
rect 50652 51436 50708 51492
rect 50540 49868 50596 49924
rect 50428 49756 50484 49812
rect 50316 49196 50372 49252
rect 50764 50706 50820 50708
rect 50764 50654 50766 50706
rect 50766 50654 50818 50706
rect 50818 50654 50820 50706
rect 50764 50652 50820 50654
rect 51212 52220 51268 52276
rect 52108 57148 52164 57204
rect 51996 56812 52052 56868
rect 51884 56252 51940 56308
rect 51996 55244 52052 55300
rect 52220 56476 52276 56532
rect 53116 56588 53172 56644
rect 53228 56700 53284 56756
rect 52668 56140 52724 56196
rect 52556 56028 52612 56084
rect 54012 57260 54068 57316
rect 55356 57260 55412 57316
rect 54908 56924 54964 56980
rect 54460 56364 54516 56420
rect 55020 56476 55076 56532
rect 51548 53730 51604 53732
rect 51548 53678 51550 53730
rect 51550 53678 51602 53730
rect 51602 53678 51604 53730
rect 51548 53676 51604 53678
rect 51436 51548 51492 51604
rect 51324 51378 51380 51380
rect 51324 51326 51326 51378
rect 51326 51326 51378 51378
rect 51378 51326 51380 51378
rect 51324 51324 51380 51326
rect 51212 51212 51268 51268
rect 50988 50540 51044 50596
rect 51548 50876 51604 50932
rect 50652 49420 50708 49476
rect 50540 48972 50596 49028
rect 50876 48524 50932 48580
rect 49980 47012 50036 47068
rect 50540 48412 50596 48468
rect 49868 46620 49924 46676
rect 50316 48130 50372 48132
rect 50316 48078 50318 48130
rect 50318 48078 50370 48130
rect 50370 48078 50372 48130
rect 50316 48076 50372 48078
rect 50204 47068 50260 47124
rect 50092 46508 50148 46564
rect 50316 46956 50372 47012
rect 50204 46450 50260 46452
rect 50204 46398 50206 46450
rect 50206 46398 50258 46450
rect 50258 46398 50260 46450
rect 50204 46396 50260 46398
rect 49084 46002 49140 46004
rect 49084 45950 49086 46002
rect 49086 45950 49138 46002
rect 49138 45950 49140 46002
rect 49084 45948 49140 45950
rect 50092 46284 50148 46340
rect 49980 45836 50036 45892
rect 50092 45724 50148 45780
rect 49532 45500 49588 45556
rect 48972 44434 49028 44436
rect 48972 44382 48974 44434
rect 48974 44382 49026 44434
rect 49026 44382 49028 44434
rect 48972 44380 49028 44382
rect 49196 44156 49252 44212
rect 49644 45388 49700 45444
rect 48636 43372 48692 43428
rect 48860 43314 48916 43316
rect 48860 43262 48862 43314
rect 48862 43262 48914 43314
rect 48914 43262 48916 43314
rect 48860 43260 48916 43262
rect 48524 41916 48580 41972
rect 48076 41298 48132 41300
rect 48076 41246 48078 41298
rect 48078 41246 48130 41298
rect 48130 41246 48132 41298
rect 48076 41244 48132 41246
rect 49196 43538 49252 43540
rect 49196 43486 49198 43538
rect 49198 43486 49250 43538
rect 49250 43486 49252 43538
rect 49196 43484 49252 43486
rect 48972 41356 49028 41412
rect 49084 43036 49140 43092
rect 48748 41244 48804 41300
rect 48300 41132 48356 41188
rect 48188 39730 48244 39732
rect 48188 39678 48190 39730
rect 48190 39678 48242 39730
rect 48242 39678 48244 39730
rect 48188 39676 48244 39678
rect 48412 40908 48468 40964
rect 48972 40962 49028 40964
rect 48972 40910 48974 40962
rect 48974 40910 49026 40962
rect 49026 40910 49028 40962
rect 48972 40908 49028 40910
rect 48748 40796 48804 40852
rect 48972 40684 49028 40740
rect 48524 39564 48580 39620
rect 48300 38668 48356 38724
rect 48188 38274 48244 38276
rect 48188 38222 48190 38274
rect 48190 38222 48242 38274
rect 48242 38222 48244 38274
rect 48188 38220 48244 38222
rect 48076 38162 48132 38164
rect 48076 38110 48078 38162
rect 48078 38110 48130 38162
rect 48130 38110 48132 38162
rect 48076 38108 48132 38110
rect 48188 37660 48244 37716
rect 47964 36428 48020 36484
rect 48188 35980 48244 36036
rect 47964 34188 48020 34244
rect 47852 34130 47908 34132
rect 47852 34078 47854 34130
rect 47854 34078 47906 34130
rect 47906 34078 47908 34130
rect 47852 34076 47908 34078
rect 46956 33740 47012 33796
rect 47292 34018 47348 34020
rect 47292 33966 47294 34018
rect 47294 33966 47346 34018
rect 47346 33966 47348 34018
rect 47292 33964 47348 33966
rect 47068 33292 47124 33348
rect 47180 32620 47236 32676
rect 46956 32450 47012 32452
rect 46956 32398 46958 32450
rect 46958 32398 47010 32450
rect 47010 32398 47012 32450
rect 46956 32396 47012 32398
rect 47068 30940 47124 30996
rect 47516 33572 47572 33628
rect 47628 33852 47684 33908
rect 47516 33458 47572 33460
rect 47516 33406 47518 33458
rect 47518 33406 47570 33458
rect 47570 33406 47572 33458
rect 47516 33404 47572 33406
rect 47516 31724 47572 31780
rect 47404 31500 47460 31556
rect 47516 31164 47572 31220
rect 47964 33740 48020 33796
rect 48076 34076 48132 34132
rect 47628 30940 47684 30996
rect 47852 33628 47908 33684
rect 47516 30882 47572 30884
rect 47516 30830 47518 30882
rect 47518 30830 47570 30882
rect 47570 30830 47572 30882
rect 47516 30828 47572 30830
rect 46956 30380 47012 30436
rect 47068 30268 47124 30324
rect 47180 30156 47236 30212
rect 47292 30268 47348 30324
rect 47404 30156 47460 30212
rect 46844 29538 46900 29540
rect 46844 29486 46846 29538
rect 46846 29486 46898 29538
rect 46898 29486 46900 29538
rect 46844 29484 46900 29486
rect 46956 29314 47012 29316
rect 46956 29262 46958 29314
rect 46958 29262 47010 29314
rect 47010 29262 47012 29314
rect 46956 29260 47012 29262
rect 47516 29426 47572 29428
rect 47516 29374 47518 29426
rect 47518 29374 47570 29426
rect 47570 29374 47572 29426
rect 47516 29372 47572 29374
rect 46284 27468 46340 27524
rect 46172 27244 46228 27300
rect 45388 25788 45444 25844
rect 45612 25452 45668 25508
rect 45276 25340 45332 25396
rect 45388 25116 45444 25172
rect 45276 24556 45332 24612
rect 45388 24498 45444 24500
rect 45388 24446 45390 24498
rect 45390 24446 45442 24498
rect 45442 24446 45444 24498
rect 45388 24444 45444 24446
rect 45052 23100 45108 23156
rect 45164 23212 45220 23268
rect 45164 22428 45220 22484
rect 45500 22316 45556 22372
rect 44828 18172 44884 18228
rect 44464 18058 44520 18060
rect 44464 18006 44466 18058
rect 44466 18006 44518 18058
rect 44518 18006 44520 18058
rect 44464 18004 44520 18006
rect 44568 18058 44624 18060
rect 44568 18006 44570 18058
rect 44570 18006 44622 18058
rect 44622 18006 44624 18058
rect 44568 18004 44624 18006
rect 44672 18058 44728 18060
rect 44672 18006 44674 18058
rect 44674 18006 44726 18058
rect 44726 18006 44728 18058
rect 44672 18004 44728 18006
rect 44044 17666 44100 17668
rect 44044 17614 44046 17666
rect 44046 17614 44098 17666
rect 44098 17614 44100 17666
rect 44044 17612 44100 17614
rect 43804 17274 43860 17276
rect 43804 17222 43806 17274
rect 43806 17222 43858 17274
rect 43858 17222 43860 17274
rect 43804 17220 43860 17222
rect 43908 17274 43964 17276
rect 43908 17222 43910 17274
rect 43910 17222 43962 17274
rect 43962 17222 43964 17274
rect 43908 17220 43964 17222
rect 44012 17274 44068 17276
rect 44012 17222 44014 17274
rect 44014 17222 44066 17274
rect 44066 17222 44068 17274
rect 44012 17220 44068 17222
rect 44156 17164 44212 17220
rect 43372 16604 43428 16660
rect 42812 16044 42868 16100
rect 43804 15706 43860 15708
rect 43804 15654 43806 15706
rect 43806 15654 43858 15706
rect 43858 15654 43860 15706
rect 43804 15652 43860 15654
rect 43908 15706 43964 15708
rect 43908 15654 43910 15706
rect 43910 15654 43962 15706
rect 43962 15654 43964 15706
rect 43908 15652 43964 15654
rect 44012 15706 44068 15708
rect 44012 15654 44014 15706
rect 44014 15654 44066 15706
rect 44066 15654 44068 15706
rect 44012 15652 44068 15654
rect 43708 15484 43764 15540
rect 43148 15372 43204 15428
rect 42476 14812 42532 14868
rect 42364 13468 42420 13524
rect 42252 12572 42308 12628
rect 42140 10108 42196 10164
rect 42252 11564 42308 11620
rect 42252 10556 42308 10612
rect 42476 11564 42532 11620
rect 43036 15148 43092 15204
rect 43036 14530 43092 14532
rect 43036 14478 43038 14530
rect 43038 14478 43090 14530
rect 43090 14478 43092 14530
rect 43036 14476 43092 14478
rect 43036 14140 43092 14196
rect 42924 13916 42980 13972
rect 43596 15372 43652 15428
rect 43148 13916 43204 13972
rect 43036 12572 43092 12628
rect 43148 13692 43204 13748
rect 42924 12124 42980 12180
rect 42812 11788 42868 11844
rect 43036 11618 43092 11620
rect 43036 11566 43038 11618
rect 43038 11566 43090 11618
rect 43090 11566 43092 11618
rect 43036 11564 43092 11566
rect 42812 11004 42868 11060
rect 44464 16490 44520 16492
rect 44464 16438 44466 16490
rect 44466 16438 44518 16490
rect 44518 16438 44520 16490
rect 44464 16436 44520 16438
rect 44568 16490 44624 16492
rect 44568 16438 44570 16490
rect 44570 16438 44622 16490
rect 44622 16438 44624 16490
rect 44568 16436 44624 16438
rect 44672 16490 44728 16492
rect 44672 16438 44674 16490
rect 44674 16438 44726 16490
rect 44726 16438 44728 16490
rect 44672 16436 44728 16438
rect 44380 15932 44436 15988
rect 44828 16098 44884 16100
rect 44828 16046 44830 16098
rect 44830 16046 44882 16098
rect 44882 16046 44884 16098
rect 44828 16044 44884 16046
rect 44268 15372 44324 15428
rect 44156 15260 44212 15316
rect 44044 15036 44100 15092
rect 44716 15036 44772 15092
rect 44464 14922 44520 14924
rect 44464 14870 44466 14922
rect 44466 14870 44518 14922
rect 44518 14870 44520 14922
rect 44464 14868 44520 14870
rect 44568 14922 44624 14924
rect 44568 14870 44570 14922
rect 44570 14870 44622 14922
rect 44622 14870 44624 14922
rect 44568 14868 44624 14870
rect 44672 14922 44728 14924
rect 44672 14870 44674 14922
rect 44674 14870 44726 14922
rect 44726 14870 44728 14922
rect 44672 14868 44728 14870
rect 44044 14700 44100 14756
rect 43932 14476 43988 14532
rect 45052 19906 45108 19908
rect 45052 19854 45054 19906
rect 45054 19854 45106 19906
rect 45106 19854 45108 19906
rect 45052 19852 45108 19854
rect 45948 25116 46004 25172
rect 45724 24332 45780 24388
rect 46060 23100 46116 23156
rect 46060 22482 46116 22484
rect 46060 22430 46062 22482
rect 46062 22430 46114 22482
rect 46114 22430 46116 22482
rect 46060 22428 46116 22430
rect 46060 22146 46116 22148
rect 46060 22094 46062 22146
rect 46062 22094 46114 22146
rect 46114 22094 46116 22146
rect 46060 22092 46116 22094
rect 45948 21868 46004 21924
rect 45948 21196 46004 21252
rect 45948 20860 46004 20916
rect 45836 20300 45892 20356
rect 45612 20076 45668 20132
rect 45836 19740 45892 19796
rect 46060 19794 46116 19796
rect 46060 19742 46062 19794
rect 46062 19742 46114 19794
rect 46114 19742 46116 19794
rect 46060 19740 46116 19742
rect 45500 19516 45556 19572
rect 45164 19404 45220 19460
rect 45052 19180 45108 19236
rect 45276 19346 45332 19348
rect 45276 19294 45278 19346
rect 45278 19294 45330 19346
rect 45330 19294 45332 19346
rect 45276 19292 45332 19294
rect 45612 19180 45668 19236
rect 45836 19234 45892 19236
rect 45836 19182 45838 19234
rect 45838 19182 45890 19234
rect 45890 19182 45892 19234
rect 45836 19180 45892 19182
rect 45612 18620 45668 18676
rect 45836 18620 45892 18676
rect 45388 18396 45444 18452
rect 45836 18172 45892 18228
rect 45052 16828 45108 16884
rect 45388 17724 45444 17780
rect 45500 17276 45556 17332
rect 45836 17164 45892 17220
rect 46620 26572 46676 26628
rect 46508 26460 46564 26516
rect 46396 25004 46452 25060
rect 46396 24332 46452 24388
rect 46508 23884 46564 23940
rect 46508 23714 46564 23716
rect 46508 23662 46510 23714
rect 46510 23662 46562 23714
rect 46562 23662 46564 23714
rect 46508 23660 46564 23662
rect 46508 23154 46564 23156
rect 46508 23102 46510 23154
rect 46510 23102 46562 23154
rect 46562 23102 46564 23154
rect 46508 23100 46564 23102
rect 46396 21980 46452 22036
rect 47628 28754 47684 28756
rect 47628 28702 47630 28754
rect 47630 28702 47682 28754
rect 47682 28702 47684 28754
rect 47628 28700 47684 28702
rect 47404 28364 47460 28420
rect 47292 28140 47348 28196
rect 47292 27468 47348 27524
rect 47180 26236 47236 26292
rect 47628 26460 47684 26516
rect 46844 24498 46900 24500
rect 46844 24446 46846 24498
rect 46846 24446 46898 24498
rect 46898 24446 46900 24498
rect 46844 24444 46900 24446
rect 46844 23548 46900 23604
rect 46844 22652 46900 22708
rect 47068 25228 47124 25284
rect 47404 24834 47460 24836
rect 47404 24782 47406 24834
rect 47406 24782 47458 24834
rect 47458 24782 47460 24834
rect 47404 24780 47460 24782
rect 47068 23548 47124 23604
rect 46956 21756 47012 21812
rect 48412 38220 48468 38276
rect 48300 34860 48356 34916
rect 48412 35644 48468 35700
rect 48300 34242 48356 34244
rect 48300 34190 48302 34242
rect 48302 34190 48354 34242
rect 48354 34190 48356 34242
rect 48300 34188 48356 34190
rect 48188 32732 48244 32788
rect 47852 31500 47908 31556
rect 48972 40236 49028 40292
rect 49420 41916 49476 41972
rect 49532 44380 49588 44436
rect 49420 41356 49476 41412
rect 49308 41186 49364 41188
rect 49308 41134 49310 41186
rect 49310 41134 49362 41186
rect 49362 41134 49364 41186
rect 49308 41132 49364 41134
rect 48860 39618 48916 39620
rect 48860 39566 48862 39618
rect 48862 39566 48914 39618
rect 48914 39566 48916 39618
rect 48860 39564 48916 39566
rect 48636 34018 48692 34020
rect 48636 33966 48638 34018
rect 48638 33966 48690 34018
rect 48690 33966 48692 34018
rect 48636 33964 48692 33966
rect 48860 37660 48916 37716
rect 48860 36204 48916 36260
rect 48860 34188 48916 34244
rect 48636 33516 48692 33572
rect 48748 33292 48804 33348
rect 48636 32732 48692 32788
rect 48412 31778 48468 31780
rect 48412 31726 48414 31778
rect 48414 31726 48466 31778
rect 48466 31726 48468 31778
rect 48412 31724 48468 31726
rect 48300 31500 48356 31556
rect 48524 31500 48580 31556
rect 48300 31164 48356 31220
rect 48524 31218 48580 31220
rect 48524 31166 48526 31218
rect 48526 31166 48578 31218
rect 48578 31166 48580 31218
rect 48524 31164 48580 31166
rect 48524 30940 48580 30996
rect 48076 30156 48132 30212
rect 48300 30268 48356 30324
rect 48412 30156 48468 30212
rect 48188 29484 48244 29540
rect 48412 29372 48468 29428
rect 48636 29986 48692 29988
rect 48636 29934 48638 29986
rect 48638 29934 48690 29986
rect 48690 29934 48692 29986
rect 48636 29932 48692 29934
rect 48524 29148 48580 29204
rect 48412 29036 48468 29092
rect 48188 28642 48244 28644
rect 48188 28590 48190 28642
rect 48190 28590 48242 28642
rect 48242 28590 48244 28642
rect 48188 28588 48244 28590
rect 47964 28476 48020 28532
rect 47852 24610 47908 24612
rect 47852 24558 47854 24610
rect 47854 24558 47906 24610
rect 47906 24558 47908 24610
rect 47852 24556 47908 24558
rect 47852 23996 47908 24052
rect 48188 26962 48244 26964
rect 48188 26910 48190 26962
rect 48190 26910 48242 26962
rect 48242 26910 48244 26962
rect 48188 26908 48244 26910
rect 48188 26460 48244 26516
rect 47852 23154 47908 23156
rect 47852 23102 47854 23154
rect 47854 23102 47906 23154
rect 47906 23102 47908 23154
rect 47852 23100 47908 23102
rect 47180 22876 47236 22932
rect 47404 22540 47460 22596
rect 47740 22540 47796 22596
rect 46844 21644 46900 21700
rect 46732 21532 46788 21588
rect 46620 20972 46676 21028
rect 46732 21308 46788 21364
rect 46508 20524 46564 20580
rect 46396 19964 46452 20020
rect 47180 21026 47236 21028
rect 47180 20974 47182 21026
rect 47182 20974 47234 21026
rect 47234 20974 47236 21026
rect 47180 20972 47236 20974
rect 46844 20914 46900 20916
rect 46844 20862 46846 20914
rect 46846 20862 46898 20914
rect 46898 20862 46900 20914
rect 46844 20860 46900 20862
rect 47180 20412 47236 20468
rect 46844 20300 46900 20356
rect 46508 19852 46564 19908
rect 46620 19180 46676 19236
rect 46732 18508 46788 18564
rect 46508 17164 46564 17220
rect 47068 20018 47124 20020
rect 47068 19966 47070 20018
rect 47070 19966 47122 20018
rect 47122 19966 47124 20018
rect 47068 19964 47124 19966
rect 47068 19740 47124 19796
rect 46956 18284 47012 18340
rect 47404 21980 47460 22036
rect 47516 21420 47572 21476
rect 47740 21420 47796 21476
rect 47852 22316 47908 22372
rect 47628 21362 47684 21364
rect 47628 21310 47630 21362
rect 47630 21310 47682 21362
rect 47682 21310 47684 21362
rect 47628 21308 47684 21310
rect 47852 21308 47908 21364
rect 47404 19964 47460 20020
rect 47292 18732 47348 18788
rect 47180 18284 47236 18340
rect 47068 17778 47124 17780
rect 47068 17726 47070 17778
rect 47070 17726 47122 17778
rect 47122 17726 47124 17778
rect 47068 17724 47124 17726
rect 45500 16492 45556 16548
rect 44940 15260 44996 15316
rect 45052 16156 45108 16212
rect 44940 14924 44996 14980
rect 43804 14138 43860 14140
rect 43804 14086 43806 14138
rect 43806 14086 43858 14138
rect 43858 14086 43860 14138
rect 43804 14084 43860 14086
rect 43908 14138 43964 14140
rect 43908 14086 43910 14138
rect 43910 14086 43962 14138
rect 43962 14086 43964 14138
rect 43908 14084 43964 14086
rect 44012 14138 44068 14140
rect 44012 14086 44014 14138
rect 44014 14086 44066 14138
rect 44066 14086 44068 14138
rect 44012 14084 44068 14086
rect 44156 14028 44212 14084
rect 43372 13580 43428 13636
rect 43708 13804 43764 13860
rect 44828 14140 44884 14196
rect 44492 13746 44548 13748
rect 44492 13694 44494 13746
rect 44494 13694 44546 13746
rect 44546 13694 44548 13746
rect 44492 13692 44548 13694
rect 44716 13692 44772 13748
rect 43596 13468 43652 13524
rect 44044 13468 44100 13524
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 43484 13132 43540 13188
rect 43260 12684 43316 12740
rect 43260 11788 43316 11844
rect 44604 13020 44660 13076
rect 43484 12908 43540 12964
rect 44380 12908 44436 12964
rect 44604 12684 44660 12740
rect 43804 12570 43860 12572
rect 43484 12460 43540 12516
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 43372 11340 43428 11396
rect 44940 13580 44996 13636
rect 44940 13244 44996 13300
rect 44940 13020 44996 13076
rect 44940 12572 44996 12628
rect 44828 11900 44884 11956
rect 44268 11788 44324 11844
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44044 11452 44100 11508
rect 44156 11394 44212 11396
rect 44156 11342 44158 11394
rect 44158 11342 44210 11394
rect 44210 11342 44212 11394
rect 44156 11340 44212 11342
rect 44044 11228 44100 11284
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 44268 11004 44324 11060
rect 44492 10892 44548 10948
rect 44492 10668 44548 10724
rect 45388 16210 45444 16212
rect 45388 16158 45390 16210
rect 45390 16158 45442 16210
rect 45442 16158 45444 16210
rect 45388 16156 45444 16158
rect 45388 15932 45444 15988
rect 45612 15932 45668 15988
rect 45388 15484 45444 15540
rect 45388 15260 45444 15316
rect 45164 14812 45220 14868
rect 46284 16882 46340 16884
rect 46284 16830 46286 16882
rect 46286 16830 46338 16882
rect 46338 16830 46340 16882
rect 46284 16828 46340 16830
rect 46956 16882 47012 16884
rect 46956 16830 46958 16882
rect 46958 16830 47010 16882
rect 47010 16830 47012 16882
rect 46956 16828 47012 16830
rect 45724 14530 45780 14532
rect 45724 14478 45726 14530
rect 45726 14478 45778 14530
rect 45778 14478 45780 14530
rect 45724 14476 45780 14478
rect 46620 16658 46676 16660
rect 46620 16606 46622 16658
rect 46622 16606 46674 16658
rect 46674 16606 46676 16658
rect 46620 16604 46676 16606
rect 45500 13916 45556 13972
rect 45164 13522 45220 13524
rect 45164 13470 45166 13522
rect 45166 13470 45218 13522
rect 45218 13470 45220 13522
rect 45164 13468 45220 13470
rect 45164 13020 45220 13076
rect 44716 10668 44772 10724
rect 44380 10498 44436 10500
rect 44380 10446 44382 10498
rect 44382 10446 44434 10498
rect 44434 10446 44436 10498
rect 44380 10444 44436 10446
rect 44604 10386 44660 10388
rect 44604 10334 44606 10386
rect 44606 10334 44658 10386
rect 44658 10334 44660 10386
rect 44604 10332 44660 10334
rect 43596 9996 43652 10052
rect 44268 10220 44324 10276
rect 44044 9884 44100 9940
rect 42700 9324 42756 9380
rect 42588 9042 42644 9044
rect 42588 8990 42590 9042
rect 42590 8990 42642 9042
rect 42642 8990 42644 9042
rect 42588 8988 42644 8990
rect 43036 8876 43092 8932
rect 42476 8370 42532 8372
rect 42476 8318 42478 8370
rect 42478 8318 42530 8370
rect 42530 8318 42532 8370
rect 42476 8316 42532 8318
rect 43036 8316 43092 8372
rect 42140 7362 42196 7364
rect 42140 7310 42142 7362
rect 42142 7310 42194 7362
rect 42194 7310 42196 7362
rect 42140 7308 42196 7310
rect 42252 6860 42308 6916
rect 41468 5740 41524 5796
rect 41356 5234 41412 5236
rect 41356 5182 41358 5234
rect 41358 5182 41410 5234
rect 41410 5182 41412 5234
rect 41356 5180 41412 5182
rect 41132 4844 41188 4900
rect 41244 5068 41300 5124
rect 40908 3666 40964 3668
rect 40908 3614 40910 3666
rect 40910 3614 40962 3666
rect 40962 3614 40964 3666
rect 40908 3612 40964 3614
rect 42140 6412 42196 6468
rect 42364 6748 42420 6804
rect 43148 8092 43204 8148
rect 42924 7084 42980 7140
rect 43932 9772 43988 9828
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 44268 9884 44324 9940
rect 44492 9996 44548 10052
rect 45388 12124 45444 12180
rect 45276 10556 45332 10612
rect 43804 9434 43860 9436
rect 43484 9324 43540 9380
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 44156 9324 44212 9380
rect 44604 9436 44660 9492
rect 44044 8876 44100 8932
rect 44828 8930 44884 8932
rect 44828 8878 44830 8930
rect 44830 8878 44882 8930
rect 44882 8878 44884 8930
rect 44828 8876 44884 8878
rect 44464 8650 44520 8652
rect 43820 8258 43876 8260
rect 43820 8206 43822 8258
rect 43822 8206 43874 8258
rect 43874 8206 43876 8258
rect 43820 8204 43876 8206
rect 43932 8146 43988 8148
rect 43932 8094 43934 8146
rect 43934 8094 43986 8146
rect 43986 8094 43988 8146
rect 43932 8092 43988 8094
rect 44268 8540 44324 8596
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 44940 8652 44996 8708
rect 45052 9436 45108 9492
rect 44044 7980 44100 8036
rect 43596 7868 43652 7924
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 44828 7756 44884 7812
rect 44268 7644 44324 7700
rect 44828 7362 44884 7364
rect 44828 7310 44830 7362
rect 44830 7310 44882 7362
rect 44882 7310 44884 7362
rect 44828 7308 44884 7310
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44380 6636 44436 6692
rect 44492 6412 44548 6468
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 45500 11676 45556 11732
rect 45388 9436 45444 9492
rect 45612 11452 45668 11508
rect 46620 15932 46676 15988
rect 46172 15148 46228 15204
rect 46172 14812 46228 14868
rect 46844 15484 46900 15540
rect 48188 25228 48244 25284
rect 48300 23660 48356 23716
rect 48188 22482 48244 22484
rect 48188 22430 48190 22482
rect 48190 22430 48242 22482
rect 48242 22430 48244 22482
rect 48188 22428 48244 22430
rect 47964 19964 48020 20020
rect 47628 17500 47684 17556
rect 47852 19180 47908 19236
rect 47404 16940 47460 16996
rect 47516 17276 47572 17332
rect 47292 16828 47348 16884
rect 47404 16658 47460 16660
rect 47404 16606 47406 16658
rect 47406 16606 47458 16658
rect 47458 16606 47460 16658
rect 47404 16604 47460 16606
rect 47180 16380 47236 16436
rect 46956 15372 47012 15428
rect 47180 15314 47236 15316
rect 47180 15262 47182 15314
rect 47182 15262 47234 15314
rect 47234 15262 47236 15314
rect 47180 15260 47236 15262
rect 47628 17164 47684 17220
rect 47516 16156 47572 16212
rect 46956 15202 47012 15204
rect 46956 15150 46958 15202
rect 46958 15150 47010 15202
rect 47010 15150 47012 15202
rect 46956 15148 47012 15150
rect 46620 14924 46676 14980
rect 46172 14476 46228 14532
rect 46060 14364 46116 14420
rect 46172 13804 46228 13860
rect 47516 15036 47572 15092
rect 47180 14812 47236 14868
rect 47740 15372 47796 15428
rect 48076 18956 48132 19012
rect 47852 14924 47908 14980
rect 47964 18620 48020 18676
rect 47628 14812 47684 14868
rect 47516 14700 47572 14756
rect 47404 14364 47460 14420
rect 48524 28418 48580 28420
rect 48524 28366 48526 28418
rect 48526 28366 48578 28418
rect 48578 28366 48580 28418
rect 48524 28364 48580 28366
rect 49084 38220 49140 38276
rect 49420 40348 49476 40404
rect 49308 40290 49364 40292
rect 49308 40238 49310 40290
rect 49310 40238 49362 40290
rect 49362 40238 49364 40290
rect 49308 40236 49364 40238
rect 49196 37884 49252 37940
rect 49308 38162 49364 38164
rect 49308 38110 49310 38162
rect 49310 38110 49362 38162
rect 49362 38110 49364 38162
rect 49308 38108 49364 38110
rect 49084 37660 49140 37716
rect 49084 36204 49140 36260
rect 49196 36092 49252 36148
rect 49756 44882 49812 44884
rect 49756 44830 49758 44882
rect 49758 44830 49810 44882
rect 49810 44830 49812 44882
rect 49756 44828 49812 44830
rect 49980 44828 50036 44884
rect 49756 43426 49812 43428
rect 49756 43374 49758 43426
rect 49758 43374 49810 43426
rect 49810 43374 49812 43426
rect 49756 43372 49812 43374
rect 50316 45890 50372 45892
rect 50316 45838 50318 45890
rect 50318 45838 50370 45890
rect 50370 45838 50372 45890
rect 50316 45836 50372 45838
rect 50204 45612 50260 45668
rect 50428 45612 50484 45668
rect 49756 42364 49812 42420
rect 49756 41020 49812 41076
rect 49868 41916 49924 41972
rect 49980 41468 50036 41524
rect 50876 48242 50932 48244
rect 50876 48190 50878 48242
rect 50878 48190 50930 48242
rect 50930 48190 50932 48242
rect 50876 48188 50932 48190
rect 51436 50316 51492 50372
rect 51212 49644 51268 49700
rect 51100 48412 51156 48468
rect 51100 48076 51156 48132
rect 51548 49308 51604 49364
rect 51884 53564 51940 53620
rect 51996 52444 52052 52500
rect 51884 52274 51940 52276
rect 51884 52222 51886 52274
rect 51886 52222 51938 52274
rect 51938 52222 51940 52274
rect 51884 52220 51940 52222
rect 51772 51436 51828 51492
rect 52892 55858 52948 55860
rect 52892 55806 52894 55858
rect 52894 55806 52946 55858
rect 52946 55806 52948 55858
rect 52892 55804 52948 55806
rect 52668 55468 52724 55524
rect 53564 55970 53620 55972
rect 53564 55918 53566 55970
rect 53566 55918 53618 55970
rect 53618 55918 53620 55970
rect 53564 55916 53620 55918
rect 53452 55020 53508 55076
rect 52556 53730 52612 53732
rect 52556 53678 52558 53730
rect 52558 53678 52610 53730
rect 52610 53678 52612 53730
rect 52556 53676 52612 53678
rect 52556 53452 52612 53508
rect 52332 52892 52388 52948
rect 52220 52668 52276 52724
rect 52220 52050 52276 52052
rect 52220 51998 52222 52050
rect 52222 51998 52274 52050
rect 52274 51998 52276 52050
rect 52220 51996 52276 51998
rect 52108 51378 52164 51380
rect 52108 51326 52110 51378
rect 52110 51326 52162 51378
rect 52162 51326 52164 51378
rect 52108 51324 52164 51326
rect 52108 51100 52164 51156
rect 52220 50652 52276 50708
rect 51884 49644 51940 49700
rect 52108 49868 52164 49924
rect 51996 49084 52052 49140
rect 51660 48748 51716 48804
rect 51772 48524 51828 48580
rect 51660 48188 51716 48244
rect 51548 47628 51604 47684
rect 51436 47404 51492 47460
rect 50764 46844 50820 46900
rect 50652 46620 50708 46676
rect 51436 47180 51492 47236
rect 50764 46284 50820 46340
rect 50764 45890 50820 45892
rect 50764 45838 50766 45890
rect 50766 45838 50818 45890
rect 50818 45838 50820 45890
rect 50764 45836 50820 45838
rect 51436 46396 51492 46452
rect 51436 46172 51492 46228
rect 50988 45890 51044 45892
rect 50988 45838 50990 45890
rect 50990 45838 51042 45890
rect 51042 45838 51044 45890
rect 50988 45836 51044 45838
rect 50652 44828 50708 44884
rect 51324 45388 51380 45444
rect 50764 44604 50820 44660
rect 50876 44940 50932 44996
rect 50316 44380 50372 44436
rect 49980 41074 50036 41076
rect 49980 41022 49982 41074
rect 49982 41022 50034 41074
rect 50034 41022 50036 41074
rect 49980 41020 50036 41022
rect 49868 40348 49924 40404
rect 50092 40348 50148 40404
rect 49756 40012 49812 40068
rect 49532 37042 49588 37044
rect 49532 36990 49534 37042
rect 49534 36990 49586 37042
rect 49586 36990 49588 37042
rect 49532 36988 49588 36990
rect 49420 35980 49476 36036
rect 49084 35420 49140 35476
rect 49532 35308 49588 35364
rect 49420 33516 49476 33572
rect 49532 34188 49588 34244
rect 49084 31612 49140 31668
rect 49420 31388 49476 31444
rect 49308 31164 49364 31220
rect 49756 37324 49812 37380
rect 50428 44156 50484 44212
rect 50988 44828 51044 44884
rect 50876 44044 50932 44100
rect 51212 44604 51268 44660
rect 51212 44044 51268 44100
rect 51548 44380 51604 44436
rect 51660 46620 51716 46676
rect 51660 45836 51716 45892
rect 51436 44322 51492 44324
rect 51436 44270 51438 44322
rect 51438 44270 51490 44322
rect 51490 44270 51492 44322
rect 51436 44268 51492 44270
rect 50540 43260 50596 43316
rect 50876 43596 50932 43652
rect 50764 43538 50820 43540
rect 50764 43486 50766 43538
rect 50766 43486 50818 43538
rect 50818 43486 50820 43538
rect 50764 43484 50820 43486
rect 50764 43260 50820 43316
rect 50428 41020 50484 41076
rect 50428 40178 50484 40180
rect 50428 40126 50430 40178
rect 50430 40126 50482 40178
rect 50482 40126 50484 40178
rect 50428 40124 50484 40126
rect 50316 39676 50372 39732
rect 50092 38892 50148 38948
rect 50204 39116 50260 39172
rect 49980 36876 50036 36932
rect 50092 37884 50148 37940
rect 50092 36652 50148 36708
rect 49868 35756 49924 35812
rect 50092 35420 50148 35476
rect 49868 33906 49924 33908
rect 49868 33854 49870 33906
rect 49870 33854 49922 33906
rect 49922 33854 49924 33906
rect 49868 33852 49924 33854
rect 49980 33628 50036 33684
rect 49868 33516 49924 33572
rect 49868 32620 49924 32676
rect 50428 38780 50484 38836
rect 50876 41692 50932 41748
rect 51436 44044 51492 44100
rect 50764 41356 50820 41412
rect 50876 41186 50932 41188
rect 50876 41134 50878 41186
rect 50878 41134 50930 41186
rect 50930 41134 50932 41186
rect 50876 41132 50932 41134
rect 51212 43484 51268 43540
rect 51324 43426 51380 43428
rect 51324 43374 51326 43426
rect 51326 43374 51378 43426
rect 51378 43374 51380 43426
rect 51324 43372 51380 43374
rect 52332 49868 52388 49924
rect 52220 49756 52276 49812
rect 52332 49586 52388 49588
rect 52332 49534 52334 49586
rect 52334 49534 52386 49586
rect 52386 49534 52388 49586
rect 52332 49532 52388 49534
rect 52332 49084 52388 49140
rect 52220 48748 52276 48804
rect 52332 48412 52388 48468
rect 51884 46956 51940 47012
rect 51884 45836 51940 45892
rect 51996 45778 52052 45780
rect 51996 45726 51998 45778
rect 51998 45726 52050 45778
rect 52050 45726 52052 45778
rect 51996 45724 52052 45726
rect 51884 45666 51940 45668
rect 51884 45614 51886 45666
rect 51886 45614 51938 45666
rect 51938 45614 51940 45666
rect 51884 45612 51940 45614
rect 52668 53228 52724 53284
rect 53340 52892 53396 52948
rect 52892 52444 52948 52500
rect 52780 52108 52836 52164
rect 52668 51996 52724 52052
rect 53116 51996 53172 52052
rect 52556 51548 52612 51604
rect 52444 46956 52500 47012
rect 52444 46674 52500 46676
rect 52444 46622 52446 46674
rect 52446 46622 52498 46674
rect 52498 46622 52500 46674
rect 52444 46620 52500 46622
rect 51660 44044 51716 44100
rect 51772 43708 51828 43764
rect 51660 43148 51716 43204
rect 51436 42140 51492 42196
rect 52108 44882 52164 44884
rect 52108 44830 52110 44882
rect 52110 44830 52162 44882
rect 52162 44830 52164 44882
rect 52108 44828 52164 44830
rect 52332 43708 52388 43764
rect 51996 43596 52052 43652
rect 54012 55298 54068 55300
rect 54012 55246 54014 55298
rect 54014 55246 54066 55298
rect 54066 55246 54068 55298
rect 54012 55244 54068 55246
rect 54348 55858 54404 55860
rect 54348 55806 54350 55858
rect 54350 55806 54402 55858
rect 54402 55806 54404 55858
rect 54348 55804 54404 55806
rect 53676 54684 53732 54740
rect 54236 55692 54292 55748
rect 53564 53900 53620 53956
rect 53564 53452 53620 53508
rect 53900 54236 53956 54292
rect 54684 55410 54740 55412
rect 54684 55358 54686 55410
rect 54686 55358 54738 55410
rect 54738 55358 54740 55410
rect 54684 55356 54740 55358
rect 54348 54290 54404 54292
rect 54348 54238 54350 54290
rect 54350 54238 54402 54290
rect 54402 54238 54404 54290
rect 54348 54236 54404 54238
rect 53900 53730 53956 53732
rect 53900 53678 53902 53730
rect 53902 53678 53954 53730
rect 53954 53678 53956 53730
rect 53900 53676 53956 53678
rect 55692 55858 55748 55860
rect 55692 55806 55694 55858
rect 55694 55806 55746 55858
rect 55746 55806 55748 55858
rect 55692 55804 55748 55806
rect 56252 56812 56308 56868
rect 55804 55468 55860 55524
rect 53788 53004 53844 53060
rect 53676 51660 53732 51716
rect 53564 51548 53620 51604
rect 53004 51100 53060 51156
rect 53452 50988 53508 51044
rect 52780 50482 52836 50484
rect 52780 50430 52782 50482
rect 52782 50430 52834 50482
rect 52834 50430 52836 50482
rect 52780 50428 52836 50430
rect 52668 48188 52724 48244
rect 52668 47628 52724 47684
rect 53004 49868 53060 49924
rect 53116 49756 53172 49812
rect 53004 49138 53060 49140
rect 53004 49086 53006 49138
rect 53006 49086 53058 49138
rect 53058 49086 53060 49138
rect 53004 49084 53060 49086
rect 52892 47628 52948 47684
rect 52892 46956 52948 47012
rect 53116 46620 53172 46676
rect 53004 46396 53060 46452
rect 52780 45388 52836 45444
rect 52892 44156 52948 44212
rect 52108 43538 52164 43540
rect 52108 43486 52110 43538
rect 52110 43486 52162 43538
rect 52162 43486 52164 43538
rect 52108 43484 52164 43486
rect 51996 43148 52052 43204
rect 52220 43372 52276 43428
rect 51212 41746 51268 41748
rect 51212 41694 51214 41746
rect 51214 41694 51266 41746
rect 51266 41694 51268 41746
rect 51212 41692 51268 41694
rect 51324 41298 51380 41300
rect 51324 41246 51326 41298
rect 51326 41246 51378 41298
rect 51378 41246 51380 41298
rect 51324 41244 51380 41246
rect 51100 41132 51156 41188
rect 51772 41132 51828 41188
rect 50988 40684 51044 40740
rect 50764 39228 50820 39284
rect 50988 39618 51044 39620
rect 50988 39566 50990 39618
rect 50990 39566 51042 39618
rect 51042 39566 51044 39618
rect 50988 39564 51044 39566
rect 51100 39340 51156 39396
rect 50876 39004 50932 39060
rect 51212 39116 51268 39172
rect 50764 38946 50820 38948
rect 50764 38894 50766 38946
rect 50766 38894 50818 38946
rect 50818 38894 50820 38946
rect 50764 38892 50820 38894
rect 51324 38444 51380 38500
rect 51996 40460 52052 40516
rect 51884 39004 51940 39060
rect 51996 40124 52052 40180
rect 51548 38332 51604 38388
rect 51100 37996 51156 38052
rect 51100 37772 51156 37828
rect 51436 37660 51492 37716
rect 51324 36428 51380 36484
rect 50988 35474 51044 35476
rect 50988 35422 50990 35474
rect 50990 35422 51042 35474
rect 51042 35422 51044 35474
rect 50988 35420 51044 35422
rect 50876 35196 50932 35252
rect 51212 35084 51268 35140
rect 51436 36092 51492 36148
rect 51548 35868 51604 35924
rect 51660 37996 51716 38052
rect 50876 34860 50932 34916
rect 50764 34524 50820 34580
rect 50764 34018 50820 34020
rect 50764 33966 50766 34018
rect 50766 33966 50818 34018
rect 50818 33966 50820 34018
rect 50764 33964 50820 33966
rect 50988 34018 51044 34020
rect 50988 33966 50990 34018
rect 50990 33966 51042 34018
rect 51042 33966 51044 34018
rect 50988 33964 51044 33966
rect 51100 33740 51156 33796
rect 50540 33628 50596 33684
rect 50540 33516 50596 33572
rect 50876 33572 50932 33628
rect 50204 33404 50260 33460
rect 50652 33404 50708 33460
rect 50092 32172 50148 32228
rect 49644 31612 49700 31668
rect 49084 31052 49140 31108
rect 48972 30322 49028 30324
rect 48972 30270 48974 30322
rect 48974 30270 49026 30322
rect 49026 30270 49028 30322
rect 48972 30268 49028 30270
rect 49084 29708 49140 29764
rect 49084 29202 49140 29204
rect 49084 29150 49086 29202
rect 49086 29150 49138 29202
rect 49138 29150 49140 29202
rect 49084 29148 49140 29150
rect 49084 27356 49140 27412
rect 48860 24050 48916 24052
rect 48860 23998 48862 24050
rect 48862 23998 48914 24050
rect 48914 23998 48916 24050
rect 48860 23996 48916 23998
rect 48748 23212 48804 23268
rect 48972 23100 49028 23156
rect 48748 23042 48804 23044
rect 48748 22990 48750 23042
rect 48750 22990 48802 23042
rect 48802 22990 48804 23042
rect 48748 22988 48804 22990
rect 48860 21756 48916 21812
rect 48748 21474 48804 21476
rect 48748 21422 48750 21474
rect 48750 21422 48802 21474
rect 48802 21422 48804 21474
rect 48748 21420 48804 21422
rect 48412 19964 48468 20020
rect 48300 18620 48356 18676
rect 48076 17500 48132 17556
rect 48300 17500 48356 17556
rect 48188 17276 48244 17332
rect 48300 16716 48356 16772
rect 48300 15538 48356 15540
rect 48300 15486 48302 15538
rect 48302 15486 48354 15538
rect 48354 15486 48356 15538
rect 48300 15484 48356 15486
rect 48188 15260 48244 15316
rect 48076 14700 48132 14756
rect 48748 20972 48804 21028
rect 48636 20690 48692 20692
rect 48636 20638 48638 20690
rect 48638 20638 48690 20690
rect 48690 20638 48692 20690
rect 48636 20636 48692 20638
rect 49308 28924 49364 28980
rect 49756 31276 49812 31332
rect 49644 30604 49700 30660
rect 49532 30210 49588 30212
rect 49532 30158 49534 30210
rect 49534 30158 49586 30210
rect 49586 30158 49588 30210
rect 49532 30156 49588 30158
rect 49532 29932 49588 29988
rect 49868 31164 49924 31220
rect 49868 30604 49924 30660
rect 49532 29426 49588 29428
rect 49532 29374 49534 29426
rect 49534 29374 49586 29426
rect 49586 29374 49588 29426
rect 49532 29372 49588 29374
rect 49868 29314 49924 29316
rect 49868 29262 49870 29314
rect 49870 29262 49922 29314
rect 49922 29262 49924 29314
rect 49868 29260 49924 29262
rect 49420 27356 49476 27412
rect 49756 29202 49812 29204
rect 49756 29150 49758 29202
rect 49758 29150 49810 29202
rect 49810 29150 49812 29202
rect 49756 29148 49812 29150
rect 49420 27020 49476 27076
rect 49644 28924 49700 28980
rect 49308 26460 49364 26516
rect 49084 22988 49140 23044
rect 49084 22316 49140 22372
rect 49308 25730 49364 25732
rect 49308 25678 49310 25730
rect 49310 25678 49362 25730
rect 49362 25678 49364 25730
rect 49308 25676 49364 25678
rect 49308 22594 49364 22596
rect 49308 22542 49310 22594
rect 49310 22542 49362 22594
rect 49362 22542 49364 22594
rect 49308 22540 49364 22542
rect 48860 19516 48916 19572
rect 48972 19234 49028 19236
rect 48972 19182 48974 19234
rect 48974 19182 49026 19234
rect 49026 19182 49028 19234
rect 48972 19180 49028 19182
rect 49196 21196 49252 21252
rect 49196 19458 49252 19460
rect 49196 19406 49198 19458
rect 49198 19406 49250 19458
rect 49250 19406 49252 19458
rect 49196 19404 49252 19406
rect 49084 18562 49140 18564
rect 49084 18510 49086 18562
rect 49086 18510 49138 18562
rect 49138 18510 49140 18562
rect 49084 18508 49140 18510
rect 49756 28642 49812 28644
rect 49756 28590 49758 28642
rect 49758 28590 49810 28642
rect 49810 28590 49812 28642
rect 49756 28588 49812 28590
rect 49868 27244 49924 27300
rect 49868 25676 49924 25732
rect 49756 25452 49812 25508
rect 49756 24780 49812 24836
rect 49644 23266 49700 23268
rect 49644 23214 49646 23266
rect 49646 23214 49698 23266
rect 49698 23214 49700 23266
rect 49644 23212 49700 23214
rect 49868 23772 49924 23828
rect 50876 33180 50932 33236
rect 50988 32956 51044 33012
rect 51772 37324 51828 37380
rect 51660 34636 51716 34692
rect 51772 36092 51828 36148
rect 51772 34300 51828 34356
rect 52556 43260 52612 43316
rect 52444 43036 52500 43092
rect 52444 42140 52500 42196
rect 52556 42252 52612 42308
rect 52332 42028 52388 42084
rect 52780 43372 52836 43428
rect 52780 43036 52836 43092
rect 52668 42140 52724 42196
rect 52332 41692 52388 41748
rect 52332 41132 52388 41188
rect 52220 41020 52276 41076
rect 52220 40684 52276 40740
rect 52892 41746 52948 41748
rect 52892 41694 52894 41746
rect 52894 41694 52946 41746
rect 52946 41694 52948 41746
rect 52892 41692 52948 41694
rect 52780 41580 52836 41636
rect 52892 41468 52948 41524
rect 52556 41074 52612 41076
rect 52556 41022 52558 41074
rect 52558 41022 52610 41074
rect 52610 41022 52612 41074
rect 52556 41020 52612 41022
rect 52444 40684 52500 40740
rect 52892 41132 52948 41188
rect 52668 39788 52724 39844
rect 52444 39228 52500 39284
rect 52556 39676 52612 39732
rect 52668 39394 52724 39396
rect 52668 39342 52670 39394
rect 52670 39342 52722 39394
rect 52722 39342 52724 39394
rect 52668 39340 52724 39342
rect 52556 39116 52612 39172
rect 52220 38946 52276 38948
rect 52220 38894 52222 38946
rect 52222 38894 52274 38946
rect 52274 38894 52276 38946
rect 52220 38892 52276 38894
rect 52444 38834 52500 38836
rect 52444 38782 52446 38834
rect 52446 38782 52498 38834
rect 52498 38782 52500 38834
rect 52444 38780 52500 38782
rect 52780 39116 52836 39172
rect 52444 37996 52500 38052
rect 52444 37660 52500 37716
rect 52556 36876 52612 36932
rect 52108 36428 52164 36484
rect 52444 36764 52500 36820
rect 51996 35868 52052 35924
rect 52108 35698 52164 35700
rect 52108 35646 52110 35698
rect 52110 35646 52162 35698
rect 52162 35646 52164 35698
rect 52108 35644 52164 35646
rect 51996 35420 52052 35476
rect 52332 35698 52388 35700
rect 52332 35646 52334 35698
rect 52334 35646 52386 35698
rect 52386 35646 52388 35698
rect 52332 35644 52388 35646
rect 52668 36652 52724 36708
rect 53116 45948 53172 46004
rect 53564 50652 53620 50708
rect 53676 50316 53732 50372
rect 53452 49868 53508 49924
rect 53564 49586 53620 49588
rect 53564 49534 53566 49586
rect 53566 49534 53618 49586
rect 53618 49534 53620 49586
rect 53564 49532 53620 49534
rect 54012 52162 54068 52164
rect 54012 52110 54014 52162
rect 54014 52110 54066 52162
rect 54066 52110 54068 52162
rect 54012 52108 54068 52110
rect 54236 53004 54292 53060
rect 54684 53676 54740 53732
rect 54572 52780 54628 52836
rect 54348 52444 54404 52500
rect 54124 51436 54180 51492
rect 54236 52332 54292 52388
rect 54348 51884 54404 51940
rect 55132 54124 55188 54180
rect 55132 53900 55188 53956
rect 56252 55580 56308 55636
rect 56028 54460 56084 54516
rect 55916 54348 55972 54404
rect 56028 54290 56084 54292
rect 56028 54238 56030 54290
rect 56030 54238 56082 54290
rect 56082 54238 56084 54290
rect 56028 54236 56084 54238
rect 55356 54124 55412 54180
rect 55244 53228 55300 53284
rect 55020 52892 55076 52948
rect 55356 52892 55412 52948
rect 54684 51660 54740 51716
rect 54796 51996 54852 52052
rect 54572 51436 54628 51492
rect 54124 51212 54180 51268
rect 54236 51154 54292 51156
rect 54236 51102 54238 51154
rect 54238 51102 54290 51154
rect 54290 51102 54292 51154
rect 54236 51100 54292 51102
rect 54124 50988 54180 51044
rect 54236 50482 54292 50484
rect 54236 50430 54238 50482
rect 54238 50430 54290 50482
rect 54290 50430 54292 50482
rect 54236 50428 54292 50430
rect 54572 51266 54628 51268
rect 54572 51214 54574 51266
rect 54574 51214 54626 51266
rect 54626 51214 54628 51266
rect 54572 51212 54628 51214
rect 54460 50988 54516 51044
rect 54684 50764 54740 50820
rect 54348 50204 54404 50260
rect 53900 50092 53956 50148
rect 53788 48188 53844 48244
rect 53900 48076 53956 48132
rect 53788 47740 53844 47796
rect 53788 47292 53844 47348
rect 53340 46674 53396 46676
rect 53340 46622 53342 46674
rect 53342 46622 53394 46674
rect 53394 46622 53396 46674
rect 53340 46620 53396 46622
rect 53228 45724 53284 45780
rect 53116 45612 53172 45668
rect 53228 42476 53284 42532
rect 53228 40460 53284 40516
rect 53116 40236 53172 40292
rect 53788 46674 53844 46676
rect 53788 46622 53790 46674
rect 53790 46622 53842 46674
rect 53842 46622 53844 46674
rect 53788 46620 53844 46622
rect 53676 46396 53732 46452
rect 53564 46172 53620 46228
rect 53788 46172 53844 46228
rect 53788 45612 53844 45668
rect 54236 48130 54292 48132
rect 54236 48078 54238 48130
rect 54238 48078 54290 48130
rect 54290 48078 54292 48130
rect 54236 48076 54292 48078
rect 54908 51324 54964 51380
rect 54908 50876 54964 50932
rect 55020 50764 55076 50820
rect 55356 51660 55412 51716
rect 55244 50988 55300 51044
rect 55020 50594 55076 50596
rect 55020 50542 55022 50594
rect 55022 50542 55074 50594
rect 55074 50542 55076 50594
rect 55020 50540 55076 50542
rect 54908 49420 54964 49476
rect 55020 48748 55076 48804
rect 54236 46620 54292 46676
rect 54684 48300 54740 48356
rect 54012 45612 54068 45668
rect 54796 47458 54852 47460
rect 54796 47406 54798 47458
rect 54798 47406 54850 47458
rect 54850 47406 54852 47458
rect 54796 47404 54852 47406
rect 54236 45388 54292 45444
rect 54796 46620 54852 46676
rect 55020 48130 55076 48132
rect 55020 48078 55022 48130
rect 55022 48078 55074 48130
rect 55074 48078 55076 48130
rect 55020 48076 55076 48078
rect 55692 50092 55748 50148
rect 55356 49250 55412 49252
rect 55356 49198 55358 49250
rect 55358 49198 55410 49250
rect 55410 49198 55412 49250
rect 55356 49196 55412 49198
rect 55020 46956 55076 47012
rect 54124 45276 54180 45332
rect 54012 44716 54068 44772
rect 54908 46450 54964 46452
rect 54908 46398 54910 46450
rect 54910 46398 54962 46450
rect 54962 46398 54964 46450
rect 54908 46396 54964 46398
rect 55244 46620 55300 46676
rect 55244 46396 55300 46452
rect 54684 45778 54740 45780
rect 54684 45726 54686 45778
rect 54686 45726 54738 45778
rect 54738 45726 54740 45778
rect 54684 45724 54740 45726
rect 54796 45276 54852 45332
rect 55132 45724 55188 45780
rect 54908 44882 54964 44884
rect 54908 44830 54910 44882
rect 54910 44830 54962 44882
rect 54962 44830 54964 44882
rect 54908 44828 54964 44830
rect 53676 43708 53732 43764
rect 54460 44380 54516 44436
rect 53564 43596 53620 43652
rect 53564 43314 53620 43316
rect 53564 43262 53566 43314
rect 53566 43262 53618 43314
rect 53618 43262 53620 43314
rect 53564 43260 53620 43262
rect 53676 42866 53732 42868
rect 53676 42814 53678 42866
rect 53678 42814 53730 42866
rect 53730 42814 53732 42866
rect 53676 42812 53732 42814
rect 53452 42588 53508 42644
rect 53452 42140 53508 42196
rect 54012 44044 54068 44100
rect 53900 43596 53956 43652
rect 53788 42140 53844 42196
rect 54572 43708 54628 43764
rect 54796 43708 54852 43764
rect 54124 43538 54180 43540
rect 54124 43486 54126 43538
rect 54126 43486 54178 43538
rect 54178 43486 54180 43538
rect 54124 43484 54180 43486
rect 54460 43596 54516 43652
rect 54348 43036 54404 43092
rect 54460 42642 54516 42644
rect 54460 42590 54462 42642
rect 54462 42590 54514 42642
rect 54514 42590 54516 42642
rect 54460 42588 54516 42590
rect 54572 42476 54628 42532
rect 54572 42194 54628 42196
rect 54572 42142 54574 42194
rect 54574 42142 54626 42194
rect 54626 42142 54628 42194
rect 54572 42140 54628 42142
rect 53564 41298 53620 41300
rect 53564 41246 53566 41298
rect 53566 41246 53618 41298
rect 53618 41246 53620 41298
rect 53564 41244 53620 41246
rect 54012 41244 54068 41300
rect 53452 41020 53508 41076
rect 53900 39564 53956 39620
rect 53116 39394 53172 39396
rect 53116 39342 53118 39394
rect 53118 39342 53170 39394
rect 53170 39342 53172 39394
rect 53116 39340 53172 39342
rect 53116 39116 53172 39172
rect 53340 39058 53396 39060
rect 53340 39006 53342 39058
rect 53342 39006 53394 39058
rect 53394 39006 53396 39058
rect 53340 39004 53396 39006
rect 53788 39340 53844 39396
rect 53452 38892 53508 38948
rect 53564 39228 53620 39284
rect 53564 38668 53620 38724
rect 52892 38556 52948 38612
rect 53676 38946 53732 38948
rect 53676 38894 53678 38946
rect 53678 38894 53730 38946
rect 53730 38894 53732 38946
rect 53676 38892 53732 38894
rect 53228 38556 53284 38612
rect 52892 37042 52948 37044
rect 52892 36990 52894 37042
rect 52894 36990 52946 37042
rect 52946 36990 52948 37042
rect 52892 36988 52948 36990
rect 52668 35980 52724 36036
rect 52780 36204 52836 36260
rect 52556 35810 52612 35812
rect 52556 35758 52558 35810
rect 52558 35758 52610 35810
rect 52610 35758 52612 35810
rect 52556 35756 52612 35758
rect 52892 35420 52948 35476
rect 52780 35084 52836 35140
rect 51436 33516 51492 33572
rect 51660 33516 51716 33572
rect 51212 33404 51268 33460
rect 50428 32508 50484 32564
rect 50428 31948 50484 32004
rect 50652 32060 50708 32116
rect 50428 31778 50484 31780
rect 50428 31726 50430 31778
rect 50430 31726 50482 31778
rect 50482 31726 50484 31778
rect 50428 31724 50484 31726
rect 50316 31612 50372 31668
rect 50204 31554 50260 31556
rect 50204 31502 50206 31554
rect 50206 31502 50258 31554
rect 50258 31502 50260 31554
rect 50204 31500 50260 31502
rect 50092 30434 50148 30436
rect 50092 30382 50094 30434
rect 50094 30382 50146 30434
rect 50146 30382 50148 30434
rect 50092 30380 50148 30382
rect 50204 30268 50260 30324
rect 50764 31276 50820 31332
rect 51436 32732 51492 32788
rect 51548 32620 51604 32676
rect 51436 32172 51492 32228
rect 51548 32284 51604 32340
rect 51548 31948 51604 32004
rect 51324 31666 51380 31668
rect 51324 31614 51326 31666
rect 51326 31614 51378 31666
rect 51378 31614 51380 31666
rect 51324 31612 51380 31614
rect 51324 31218 51380 31220
rect 51324 31166 51326 31218
rect 51326 31166 51378 31218
rect 51378 31166 51380 31218
rect 51324 31164 51380 31166
rect 51212 30994 51268 30996
rect 51212 30942 51214 30994
rect 51214 30942 51266 30994
rect 51266 30942 51268 30994
rect 51212 30940 51268 30942
rect 51324 30770 51380 30772
rect 51324 30718 51326 30770
rect 51326 30718 51378 30770
rect 51378 30718 51380 30770
rect 51324 30716 51380 30718
rect 51884 33516 51940 33572
rect 52556 34242 52612 34244
rect 52556 34190 52558 34242
rect 52558 34190 52610 34242
rect 52610 34190 52612 34242
rect 52556 34188 52612 34190
rect 52220 33516 52276 33572
rect 52668 33458 52724 33460
rect 52668 33406 52670 33458
rect 52670 33406 52722 33458
rect 52722 33406 52724 33458
rect 52668 33404 52724 33406
rect 51884 32508 51940 32564
rect 51660 30828 51716 30884
rect 51772 31890 51828 31892
rect 51772 31838 51774 31890
rect 51774 31838 51826 31890
rect 51826 31838 51828 31890
rect 51772 31836 51828 31838
rect 51548 30716 51604 30772
rect 51212 30322 51268 30324
rect 51212 30270 51214 30322
rect 51214 30270 51266 30322
rect 51266 30270 51268 30322
rect 51212 30268 51268 30270
rect 50764 30156 50820 30212
rect 50092 29596 50148 29652
rect 50204 29484 50260 29540
rect 50316 29426 50372 29428
rect 50316 29374 50318 29426
rect 50318 29374 50370 29426
rect 50370 29374 50372 29426
rect 50316 29372 50372 29374
rect 50764 29260 50820 29316
rect 50204 28028 50260 28084
rect 50316 29036 50372 29092
rect 51660 30210 51716 30212
rect 51660 30158 51662 30210
rect 51662 30158 51714 30210
rect 51714 30158 51716 30210
rect 51660 30156 51716 30158
rect 50988 28588 51044 28644
rect 51100 28924 51156 28980
rect 50876 27356 50932 27412
rect 51100 27020 51156 27076
rect 51884 31164 51940 31220
rect 50316 25676 50372 25732
rect 50204 25228 50260 25284
rect 50316 24892 50372 24948
rect 50092 22930 50148 22932
rect 50092 22878 50094 22930
rect 50094 22878 50146 22930
rect 50146 22878 50148 22930
rect 50092 22876 50148 22878
rect 50204 22764 50260 22820
rect 49644 22316 49700 22372
rect 49532 20748 49588 20804
rect 49644 22092 49700 22148
rect 49420 18396 49476 18452
rect 48860 18060 48916 18116
rect 48748 17836 48804 17892
rect 49196 16940 49252 16996
rect 48636 16770 48692 16772
rect 48636 16718 48638 16770
rect 48638 16718 48690 16770
rect 48690 16718 48692 16770
rect 48636 16716 48692 16718
rect 48860 16380 48916 16436
rect 48748 15986 48804 15988
rect 48748 15934 48750 15986
rect 48750 15934 48802 15986
rect 48802 15934 48804 15986
rect 48748 15932 48804 15934
rect 48636 15484 48692 15540
rect 48524 14700 48580 14756
rect 48636 14924 48692 14980
rect 48748 14812 48804 14868
rect 47964 14364 48020 14420
rect 48412 14418 48468 14420
rect 48412 14366 48414 14418
rect 48414 14366 48466 14418
rect 48466 14366 48468 14418
rect 48412 14364 48468 14366
rect 47404 14140 47460 14196
rect 47292 13580 47348 13636
rect 46172 13074 46228 13076
rect 46172 13022 46174 13074
rect 46174 13022 46226 13074
rect 46226 13022 46228 13074
rect 46172 13020 46228 13022
rect 46844 13020 46900 13076
rect 46508 12572 46564 12628
rect 46844 12460 46900 12516
rect 45836 7868 45892 7924
rect 45948 10444 46004 10500
rect 45612 7756 45668 7812
rect 45836 7644 45892 7700
rect 44940 6188 44996 6244
rect 44156 5740 44212 5796
rect 41692 3388 41748 3444
rect 40684 2940 40740 2996
rect 40572 2380 40628 2436
rect 40012 1596 40068 1652
rect 39788 978 39844 980
rect 39788 926 39790 978
rect 39790 926 39842 978
rect 39842 926 39844 978
rect 39788 924 39844 926
rect 40236 924 40292 980
rect 40460 700 40516 756
rect 40796 2210 40852 2212
rect 40796 2158 40798 2210
rect 40798 2158 40850 2210
rect 40850 2158 40852 2210
rect 40796 2156 40852 2158
rect 42140 5122 42196 5124
rect 42140 5070 42142 5122
rect 42142 5070 42194 5122
rect 42194 5070 42196 5122
rect 42140 5068 42196 5070
rect 42588 5180 42644 5236
rect 43596 5516 43652 5572
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 44828 5404 44884 5460
rect 42812 4956 42868 5012
rect 43484 5122 43540 5124
rect 43484 5070 43486 5122
rect 43486 5070 43538 5122
rect 43538 5070 43540 5122
rect 43484 5068 43540 5070
rect 44380 5122 44436 5124
rect 44380 5070 44382 5122
rect 44382 5070 44434 5122
rect 44434 5070 44436 5122
rect 44380 5068 44436 5070
rect 45612 6748 45668 6804
rect 45948 6860 46004 6916
rect 46060 10332 46116 10388
rect 46396 12124 46452 12180
rect 46284 11228 46340 11284
rect 46732 11788 46788 11844
rect 46396 10108 46452 10164
rect 46508 7756 46564 7812
rect 46732 11116 46788 11172
rect 46732 10444 46788 10500
rect 46956 12124 47012 12180
rect 47964 13916 48020 13972
rect 48524 13970 48580 13972
rect 48524 13918 48526 13970
rect 48526 13918 48578 13970
rect 48578 13918 48580 13970
rect 48524 13916 48580 13918
rect 49420 16716 49476 16772
rect 49420 15932 49476 15988
rect 48972 15708 49028 15764
rect 48972 15260 49028 15316
rect 49420 15260 49476 15316
rect 49756 20972 49812 21028
rect 49756 18844 49812 18900
rect 50204 21026 50260 21028
rect 50204 20974 50206 21026
rect 50206 20974 50258 21026
rect 50258 20974 50260 21026
rect 50204 20972 50260 20974
rect 50092 20076 50148 20132
rect 50204 18956 50260 19012
rect 50540 25676 50596 25732
rect 50540 25506 50596 25508
rect 50540 25454 50542 25506
rect 50542 25454 50594 25506
rect 50594 25454 50596 25506
rect 50540 25452 50596 25454
rect 50652 24892 50708 24948
rect 50652 24668 50708 24724
rect 50988 25452 51044 25508
rect 50428 23212 50484 23268
rect 50988 24892 51044 24948
rect 50540 22204 50596 22260
rect 50428 20188 50484 20244
rect 50316 18732 50372 18788
rect 50428 19516 50484 19572
rect 50540 19404 50596 19460
rect 50428 18844 50484 18900
rect 49644 18450 49700 18452
rect 49644 18398 49646 18450
rect 49646 18398 49698 18450
rect 49698 18398 49700 18450
rect 49644 18396 49700 18398
rect 50092 18172 50148 18228
rect 50092 17724 50148 17780
rect 50204 18396 50260 18452
rect 49980 16940 50036 16996
rect 50092 17276 50148 17332
rect 51100 24834 51156 24836
rect 51100 24782 51102 24834
rect 51102 24782 51154 24834
rect 51154 24782 51156 24834
rect 51100 24780 51156 24782
rect 50764 23212 50820 23268
rect 51324 25228 51380 25284
rect 51548 25116 51604 25172
rect 51660 29484 51716 29540
rect 52220 32956 52276 33012
rect 52332 31836 52388 31892
rect 52220 31612 52276 31668
rect 52220 30994 52276 30996
rect 52220 30942 52222 30994
rect 52222 30942 52274 30994
rect 52274 30942 52276 30994
rect 52220 30940 52276 30942
rect 52108 30322 52164 30324
rect 52108 30270 52110 30322
rect 52110 30270 52162 30322
rect 52162 30270 52164 30322
rect 52108 30268 52164 30270
rect 52332 29708 52388 29764
rect 52780 33292 52836 33348
rect 52892 34188 52948 34244
rect 53116 36988 53172 37044
rect 53116 36652 53172 36708
rect 53116 35532 53172 35588
rect 53004 33964 53060 34020
rect 53340 37212 53396 37268
rect 53564 38050 53620 38052
rect 53564 37998 53566 38050
rect 53566 37998 53618 38050
rect 53618 37998 53620 38050
rect 53564 37996 53620 37998
rect 53564 36988 53620 37044
rect 53788 37212 53844 37268
rect 55020 42028 55076 42084
rect 54908 41356 54964 41412
rect 54348 39618 54404 39620
rect 54348 39566 54350 39618
rect 54350 39566 54402 39618
rect 54402 39566 54404 39618
rect 54348 39564 54404 39566
rect 54236 39004 54292 39060
rect 53676 36652 53732 36708
rect 53900 36652 53956 36708
rect 54124 36988 54180 37044
rect 54460 38780 54516 38836
rect 54572 38892 54628 38948
rect 54348 38722 54404 38724
rect 54348 38670 54350 38722
rect 54350 38670 54402 38722
rect 54402 38670 54404 38722
rect 54348 38668 54404 38670
rect 54796 39676 54852 39732
rect 54348 36482 54404 36484
rect 54348 36430 54350 36482
rect 54350 36430 54402 36482
rect 54402 36430 54404 36482
rect 54348 36428 54404 36430
rect 54684 38610 54740 38612
rect 54684 38558 54686 38610
rect 54686 38558 54738 38610
rect 54738 38558 54740 38610
rect 54684 38556 54740 38558
rect 54796 38444 54852 38500
rect 54572 37996 54628 38052
rect 55356 45612 55412 45668
rect 56028 52386 56084 52388
rect 56028 52334 56030 52386
rect 56030 52334 56082 52386
rect 56082 52334 56084 52386
rect 56028 52332 56084 52334
rect 55916 51324 55972 51380
rect 55804 48076 55860 48132
rect 56028 49196 56084 49252
rect 56364 52892 56420 52948
rect 56364 52722 56420 52724
rect 56364 52670 56366 52722
rect 56366 52670 56418 52722
rect 56418 52670 56420 52722
rect 56364 52668 56420 52670
rect 56364 51548 56420 51604
rect 56364 51154 56420 51156
rect 56364 51102 56366 51154
rect 56366 51102 56418 51154
rect 56418 51102 56420 51154
rect 56364 51100 56420 51102
rect 56364 50706 56420 50708
rect 56364 50654 56366 50706
rect 56366 50654 56418 50706
rect 56418 50654 56420 50706
rect 56364 50652 56420 50654
rect 56252 49756 56308 49812
rect 56252 49586 56308 49588
rect 56252 49534 56254 49586
rect 56254 49534 56306 49586
rect 56306 49534 56308 49586
rect 56252 49532 56308 49534
rect 55916 47852 55972 47908
rect 56028 49026 56084 49028
rect 56028 48974 56030 49026
rect 56030 48974 56082 49026
rect 56082 48974 56084 49026
rect 56028 48972 56084 48974
rect 56028 47740 56084 47796
rect 55692 47628 55748 47684
rect 55580 47516 55636 47572
rect 55468 43260 55524 43316
rect 55244 42978 55300 42980
rect 55244 42926 55246 42978
rect 55246 42926 55298 42978
rect 55298 42926 55300 42978
rect 55244 42924 55300 42926
rect 55244 42700 55300 42756
rect 55244 42476 55300 42532
rect 55468 41804 55524 41860
rect 55356 41186 55412 41188
rect 55356 41134 55358 41186
rect 55358 41134 55410 41186
rect 55410 41134 55412 41186
rect 55356 41132 55412 41134
rect 55244 39116 55300 39172
rect 55356 40236 55412 40292
rect 55244 38556 55300 38612
rect 55132 37548 55188 37604
rect 55132 37042 55188 37044
rect 55132 36990 55134 37042
rect 55134 36990 55186 37042
rect 55186 36990 55188 37042
rect 55132 36988 55188 36990
rect 53452 35196 53508 35252
rect 53676 35308 53732 35364
rect 53340 35084 53396 35140
rect 53228 34076 53284 34132
rect 53564 34972 53620 35028
rect 53564 34076 53620 34132
rect 53116 33628 53172 33684
rect 53788 35196 53844 35252
rect 54684 36428 54740 36484
rect 54124 35698 54180 35700
rect 54124 35646 54126 35698
rect 54126 35646 54178 35698
rect 54178 35646 54180 35698
rect 54124 35644 54180 35646
rect 54124 35420 54180 35476
rect 53900 34748 53956 34804
rect 54908 36428 54964 36484
rect 54796 35980 54852 36036
rect 54684 35196 54740 35252
rect 54684 35026 54740 35028
rect 54684 34974 54686 35026
rect 54686 34974 54738 35026
rect 54738 34974 54740 35026
rect 54684 34972 54740 34974
rect 54348 34802 54404 34804
rect 54348 34750 54350 34802
rect 54350 34750 54402 34802
rect 54402 34750 54404 34802
rect 54348 34748 54404 34750
rect 56028 46450 56084 46452
rect 56028 46398 56030 46450
rect 56030 46398 56082 46450
rect 56082 46398 56084 46450
rect 56028 46396 56084 46398
rect 55804 45276 55860 45332
rect 55804 43426 55860 43428
rect 55804 43374 55806 43426
rect 55806 43374 55858 43426
rect 55858 43374 55860 43426
rect 55804 43372 55860 43374
rect 55692 42924 55748 42980
rect 55804 42364 55860 42420
rect 55692 41746 55748 41748
rect 55692 41694 55694 41746
rect 55694 41694 55746 41746
rect 55746 41694 55748 41746
rect 55692 41692 55748 41694
rect 56028 45164 56084 45220
rect 56252 48188 56308 48244
rect 56812 55580 56868 55636
rect 56812 48972 56868 49028
rect 57036 53004 57092 53060
rect 56588 48636 56644 48692
rect 56476 47740 56532 47796
rect 56364 47570 56420 47572
rect 56364 47518 56366 47570
rect 56366 47518 56418 47570
rect 56418 47518 56420 47570
rect 56364 47516 56420 47518
rect 56252 46732 56308 46788
rect 56252 45388 56308 45444
rect 56364 45276 56420 45332
rect 56476 45164 56532 45220
rect 56252 44716 56308 44772
rect 56364 44434 56420 44436
rect 56364 44382 56366 44434
rect 56366 44382 56418 44434
rect 56418 44382 56420 44434
rect 56364 44380 56420 44382
rect 56476 43932 56532 43988
rect 56364 43426 56420 43428
rect 56364 43374 56366 43426
rect 56366 43374 56418 43426
rect 56418 43374 56420 43426
rect 56364 43372 56420 43374
rect 55916 41356 55972 41412
rect 55916 41186 55972 41188
rect 55916 41134 55918 41186
rect 55918 41134 55970 41186
rect 55970 41134 55972 41186
rect 55916 41132 55972 41134
rect 55804 40908 55860 40964
rect 55916 40514 55972 40516
rect 55916 40462 55918 40514
rect 55918 40462 55970 40514
rect 55970 40462 55972 40514
rect 55916 40460 55972 40462
rect 56252 42700 56308 42756
rect 56140 42082 56196 42084
rect 56140 42030 56142 42082
rect 56142 42030 56194 42082
rect 56194 42030 56196 42082
rect 56140 42028 56196 42030
rect 56364 41356 56420 41412
rect 56028 39618 56084 39620
rect 56028 39566 56030 39618
rect 56030 39566 56082 39618
rect 56082 39566 56084 39618
rect 56028 39564 56084 39566
rect 55580 39452 55636 39508
rect 55804 39004 55860 39060
rect 55692 38946 55748 38948
rect 55692 38894 55694 38946
rect 55694 38894 55746 38946
rect 55746 38894 55748 38946
rect 55692 38892 55748 38894
rect 55580 38834 55636 38836
rect 55580 38782 55582 38834
rect 55582 38782 55634 38834
rect 55634 38782 55636 38834
rect 55580 38780 55636 38782
rect 55468 37100 55524 37156
rect 55580 38556 55636 38612
rect 55356 36370 55412 36372
rect 55356 36318 55358 36370
rect 55358 36318 55410 36370
rect 55410 36318 55412 36370
rect 55356 36316 55412 36318
rect 55468 35980 55524 36036
rect 55132 35532 55188 35588
rect 55244 35644 55300 35700
rect 55020 34748 55076 34804
rect 53788 33852 53844 33908
rect 54012 33964 54068 34020
rect 53116 33292 53172 33348
rect 52892 32620 52948 32676
rect 52556 31948 52612 32004
rect 53564 32508 53620 32564
rect 53116 31948 53172 32004
rect 53340 32172 53396 32228
rect 53004 31276 53060 31332
rect 52668 30882 52724 30884
rect 52668 30830 52670 30882
rect 52670 30830 52722 30882
rect 52722 30830 52724 30882
rect 52668 30828 52724 30830
rect 52668 30044 52724 30100
rect 52332 29036 52388 29092
rect 52556 29202 52612 29204
rect 52556 29150 52558 29202
rect 52558 29150 52610 29202
rect 52610 29150 52612 29202
rect 52556 29148 52612 29150
rect 52780 29426 52836 29428
rect 52780 29374 52782 29426
rect 52782 29374 52834 29426
rect 52834 29374 52836 29426
rect 52780 29372 52836 29374
rect 53228 30044 53284 30100
rect 53340 29820 53396 29876
rect 53340 29484 53396 29540
rect 52108 28812 52164 28868
rect 52556 28812 52612 28868
rect 51996 28700 52052 28756
rect 52220 28418 52276 28420
rect 52220 28366 52222 28418
rect 52222 28366 52274 28418
rect 52274 28366 52276 28418
rect 52220 28364 52276 28366
rect 52108 28140 52164 28196
rect 51884 27692 51940 27748
rect 52220 26572 52276 26628
rect 52220 26012 52276 26068
rect 53340 29036 53396 29092
rect 52892 28700 52948 28756
rect 52556 27858 52612 27860
rect 52556 27806 52558 27858
rect 52558 27806 52610 27858
rect 52610 27806 52612 27858
rect 52556 27804 52612 27806
rect 52780 27468 52836 27524
rect 52668 27186 52724 27188
rect 52668 27134 52670 27186
rect 52670 27134 52722 27186
rect 52722 27134 52724 27186
rect 52668 27132 52724 27134
rect 53788 33404 53844 33460
rect 54012 33068 54068 33124
rect 53900 32844 53956 32900
rect 54012 32172 54068 32228
rect 53788 31948 53844 32004
rect 53676 30940 53732 30996
rect 53676 30716 53732 30772
rect 53900 29820 53956 29876
rect 53900 29260 53956 29316
rect 53564 28252 53620 28308
rect 53676 29148 53732 29204
rect 53340 28082 53396 28084
rect 53340 28030 53342 28082
rect 53342 28030 53394 28082
rect 53394 28030 53396 28082
rect 53340 28028 53396 28030
rect 53340 27746 53396 27748
rect 53340 27694 53342 27746
rect 53342 27694 53394 27746
rect 53394 27694 53396 27746
rect 53340 27692 53396 27694
rect 53228 27244 53284 27300
rect 53116 27132 53172 27188
rect 53452 26908 53508 26964
rect 53564 27132 53620 27188
rect 52444 26572 52500 26628
rect 52556 26402 52612 26404
rect 52556 26350 52558 26402
rect 52558 26350 52610 26402
rect 52610 26350 52612 26402
rect 52556 26348 52612 26350
rect 52668 26290 52724 26292
rect 52668 26238 52670 26290
rect 52670 26238 52722 26290
rect 52722 26238 52724 26290
rect 52668 26236 52724 26238
rect 52556 26124 52612 26180
rect 52892 26572 52948 26628
rect 51660 24556 51716 24612
rect 51324 24332 51380 24388
rect 50876 22988 50932 23044
rect 50876 22540 50932 22596
rect 50764 21474 50820 21476
rect 50764 21422 50766 21474
rect 50766 21422 50818 21474
rect 50818 21422 50820 21474
rect 50764 21420 50820 21422
rect 50988 22316 51044 22372
rect 51100 22876 51156 22932
rect 50652 17836 50708 17892
rect 50428 17276 50484 17332
rect 50876 19852 50932 19908
rect 51548 23772 51604 23828
rect 51212 21868 51268 21924
rect 51772 25340 51828 25396
rect 52108 25340 52164 25396
rect 52108 25004 52164 25060
rect 52444 24946 52500 24948
rect 52444 24894 52446 24946
rect 52446 24894 52498 24946
rect 52498 24894 52500 24946
rect 52444 24892 52500 24894
rect 52556 24332 52612 24388
rect 52108 23996 52164 24052
rect 51772 22540 51828 22596
rect 51660 20748 51716 20804
rect 51324 20242 51380 20244
rect 51324 20190 51326 20242
rect 51326 20190 51378 20242
rect 51378 20190 51380 20242
rect 51324 20188 51380 20190
rect 51996 20578 52052 20580
rect 51996 20526 51998 20578
rect 51998 20526 52050 20578
rect 52050 20526 52052 20578
rect 51996 20524 52052 20526
rect 51884 20188 51940 20244
rect 52220 23266 52276 23268
rect 52220 23214 52222 23266
rect 52222 23214 52274 23266
rect 52274 23214 52276 23266
rect 52220 23212 52276 23214
rect 52668 23042 52724 23044
rect 52668 22990 52670 23042
rect 52670 22990 52722 23042
rect 52722 22990 52724 23042
rect 52668 22988 52724 22990
rect 52332 21084 52388 21140
rect 52108 19906 52164 19908
rect 52108 19854 52110 19906
rect 52110 19854 52162 19906
rect 52162 19854 52164 19906
rect 52108 19852 52164 19854
rect 51884 19516 51940 19572
rect 51324 18620 51380 18676
rect 50876 18508 50932 18564
rect 51212 18562 51268 18564
rect 51212 18510 51214 18562
rect 51214 18510 51266 18562
rect 51266 18510 51268 18562
rect 51212 18508 51268 18510
rect 51324 18450 51380 18452
rect 51324 18398 51326 18450
rect 51326 18398 51378 18450
rect 51378 18398 51380 18450
rect 51324 18396 51380 18398
rect 50876 18338 50932 18340
rect 50876 18286 50878 18338
rect 50878 18286 50930 18338
rect 50930 18286 50932 18338
rect 50876 18284 50932 18286
rect 51100 17612 51156 17668
rect 50316 16380 50372 16436
rect 49644 15484 49700 15540
rect 49644 15260 49700 15316
rect 50764 16604 50820 16660
rect 50204 16156 50260 16212
rect 50092 15986 50148 15988
rect 50092 15934 50094 15986
rect 50094 15934 50146 15986
rect 50146 15934 50148 15986
rect 50092 15932 50148 15934
rect 50204 15148 50260 15204
rect 49532 14924 49588 14980
rect 50988 16882 51044 16884
rect 50988 16830 50990 16882
rect 50990 16830 51042 16882
rect 51042 16830 51044 16882
rect 50988 16828 51044 16830
rect 50876 16156 50932 16212
rect 49868 15036 49924 15092
rect 49532 14642 49588 14644
rect 49532 14590 49534 14642
rect 49534 14590 49586 14642
rect 49586 14590 49588 14642
rect 49532 14588 49588 14590
rect 48860 13916 48916 13972
rect 48972 14364 49028 14420
rect 50428 15820 50484 15876
rect 50540 15484 50596 15540
rect 50652 15932 50708 15988
rect 50876 15874 50932 15876
rect 50876 15822 50878 15874
rect 50878 15822 50930 15874
rect 50930 15822 50932 15874
rect 50876 15820 50932 15822
rect 50764 15708 50820 15764
rect 51324 17106 51380 17108
rect 51324 17054 51326 17106
rect 51326 17054 51378 17106
rect 51378 17054 51380 17106
rect 51324 17052 51380 17054
rect 51884 19292 51940 19348
rect 51660 18732 51716 18788
rect 51548 17276 51604 17332
rect 51212 16156 51268 16212
rect 50092 14364 50148 14420
rect 48972 13244 49028 13300
rect 49196 14140 49252 14196
rect 48076 13132 48132 13188
rect 48636 13132 48692 13188
rect 48860 13186 48916 13188
rect 48860 13134 48862 13186
rect 48862 13134 48914 13186
rect 48914 13134 48916 13186
rect 48860 13132 48916 13134
rect 47852 12460 47908 12516
rect 46956 11004 47012 11060
rect 47068 11900 47124 11956
rect 46620 7084 46676 7140
rect 46844 8764 46900 8820
rect 46956 7868 47012 7924
rect 47292 11788 47348 11844
rect 47852 11900 47908 11956
rect 47404 11506 47460 11508
rect 47404 11454 47406 11506
rect 47406 11454 47458 11506
rect 47458 11454 47460 11506
rect 47404 11452 47460 11454
rect 47852 11340 47908 11396
rect 48300 12460 48356 12516
rect 48300 12012 48356 12068
rect 48524 12012 48580 12068
rect 48300 11788 48356 11844
rect 48972 12460 49028 12516
rect 48748 11900 48804 11956
rect 48636 11788 48692 11844
rect 47628 11004 47684 11060
rect 47404 10108 47460 10164
rect 47404 9660 47460 9716
rect 47180 9602 47236 9604
rect 47180 9550 47182 9602
rect 47182 9550 47234 9602
rect 47234 9550 47236 9602
rect 47180 9548 47236 9550
rect 47740 10610 47796 10612
rect 47740 10558 47742 10610
rect 47742 10558 47794 10610
rect 47794 10558 47796 10610
rect 47740 10556 47796 10558
rect 47964 10498 48020 10500
rect 47964 10446 47966 10498
rect 47966 10446 48018 10498
rect 48018 10446 48020 10498
rect 47964 10444 48020 10446
rect 48076 10108 48132 10164
rect 48524 11394 48580 11396
rect 48524 11342 48526 11394
rect 48526 11342 48578 11394
rect 48578 11342 48580 11394
rect 48524 11340 48580 11342
rect 48524 11004 48580 11060
rect 48412 10610 48468 10612
rect 48412 10558 48414 10610
rect 48414 10558 48466 10610
rect 48466 10558 48468 10610
rect 48412 10556 48468 10558
rect 48524 10108 48580 10164
rect 47852 9772 47908 9828
rect 47180 8930 47236 8932
rect 47180 8878 47182 8930
rect 47182 8878 47234 8930
rect 47234 8878 47236 8930
rect 47180 8876 47236 8878
rect 47516 8316 47572 8372
rect 47180 7868 47236 7924
rect 47180 7420 47236 7476
rect 46620 6860 46676 6916
rect 46284 6802 46340 6804
rect 46284 6750 46286 6802
rect 46286 6750 46338 6802
rect 46338 6750 46340 6802
rect 46284 6748 46340 6750
rect 45836 6300 45892 6356
rect 44604 5068 44660 5124
rect 44156 4844 44212 4900
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 44604 4396 44660 4452
rect 44492 4338 44548 4340
rect 44492 4286 44494 4338
rect 44494 4286 44546 4338
rect 44546 4286 44548 4338
rect 44492 4284 44548 4286
rect 42140 2770 42196 2772
rect 42140 2718 42142 2770
rect 42142 2718 42194 2770
rect 42194 2718 42196 2770
rect 42140 2716 42196 2718
rect 41132 2658 41188 2660
rect 41132 2606 41134 2658
rect 41134 2606 41186 2658
rect 41186 2606 41188 2658
rect 41132 2604 41188 2606
rect 41468 2492 41524 2548
rect 41132 1372 41188 1428
rect 41916 1708 41972 1764
rect 41468 1036 41524 1092
rect 41020 476 41076 532
rect 44044 4172 44100 4228
rect 44940 4844 44996 4900
rect 44828 4508 44884 4564
rect 44464 3946 44520 3948
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 44156 3666 44212 3668
rect 44156 3614 44158 3666
rect 44158 3614 44210 3666
rect 44210 3614 44212 3666
rect 44156 3612 44212 3614
rect 44492 3612 44548 3668
rect 44044 3388 44100 3444
rect 43804 3162 43860 3164
rect 43484 3052 43540 3108
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 43596 2770 43652 2772
rect 43596 2718 43598 2770
rect 43598 2718 43650 2770
rect 43650 2718 43652 2770
rect 43596 2716 43652 2718
rect 44828 3276 44884 3332
rect 43372 2604 43428 2660
rect 44156 2658 44212 2660
rect 44156 2606 44158 2658
rect 44158 2606 44210 2658
rect 44210 2606 44212 2658
rect 44156 2604 44212 2606
rect 43148 2546 43204 2548
rect 43148 2494 43150 2546
rect 43150 2494 43202 2546
rect 43202 2494 43204 2546
rect 43148 2492 43204 2494
rect 43932 2492 43988 2548
rect 42476 1932 42532 1988
rect 42364 812 42420 868
rect 42924 2210 42980 2212
rect 42924 2158 42926 2210
rect 42926 2158 42978 2210
rect 42978 2158 42980 2210
rect 42924 2156 42980 2158
rect 44268 2492 44324 2548
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 43484 2044 43540 2100
rect 43260 1148 43316 1204
rect 43372 1820 43428 1876
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 44604 1596 44660 1652
rect 45164 3500 45220 3556
rect 46172 3836 46228 3892
rect 45724 2940 45780 2996
rect 45500 2770 45556 2772
rect 45500 2718 45502 2770
rect 45502 2718 45554 2770
rect 45554 2718 45556 2770
rect 45500 2716 45556 2718
rect 45724 2716 45780 2772
rect 45388 2604 45444 2660
rect 45164 2268 45220 2324
rect 45164 1484 45220 1540
rect 45276 1372 45332 1428
rect 43596 1036 43652 1092
rect 44044 1036 44100 1092
rect 43148 364 43204 420
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 45612 2210 45668 2212
rect 45612 2158 45614 2210
rect 45614 2158 45666 2210
rect 45666 2158 45668 2210
rect 45612 2156 45668 2158
rect 46508 4284 46564 4340
rect 46620 5068 46676 5124
rect 46844 4956 46900 5012
rect 46508 3836 46564 3892
rect 46284 2828 46340 2884
rect 46396 3612 46452 3668
rect 45836 2546 45892 2548
rect 45836 2494 45838 2546
rect 45838 2494 45890 2546
rect 45890 2494 45892 2546
rect 45836 2492 45892 2494
rect 45948 2380 46004 2436
rect 45836 1986 45892 1988
rect 45836 1934 45838 1986
rect 45838 1934 45890 1986
rect 45890 1934 45892 1986
rect 45836 1932 45892 1934
rect 45052 978 45108 980
rect 45052 926 45054 978
rect 45054 926 45106 978
rect 45106 926 45108 978
rect 45052 924 45108 926
rect 44044 588 44100 644
rect 44156 364 44212 420
rect 43820 252 43876 308
rect 46284 2210 46340 2212
rect 46284 2158 46286 2210
rect 46286 2158 46338 2210
rect 46338 2158 46340 2210
rect 46284 2156 46340 2158
rect 46732 3500 46788 3556
rect 46620 1932 46676 1988
rect 47180 6524 47236 6580
rect 47068 6076 47124 6132
rect 47068 3836 47124 3892
rect 47068 3666 47124 3668
rect 47068 3614 47070 3666
rect 47070 3614 47122 3666
rect 47122 3614 47124 3666
rect 47068 3612 47124 3614
rect 47404 3554 47460 3556
rect 47404 3502 47406 3554
rect 47406 3502 47458 3554
rect 47458 3502 47460 3554
rect 47404 3500 47460 3502
rect 47740 7980 47796 8036
rect 48076 8876 48132 8932
rect 48188 9660 48244 9716
rect 48188 8988 48244 9044
rect 47964 8258 48020 8260
rect 47964 8206 47966 8258
rect 47966 8206 48018 8258
rect 48018 8206 48020 8258
rect 47964 8204 48020 8206
rect 48412 9772 48468 9828
rect 49084 11564 49140 11620
rect 48748 11506 48804 11508
rect 48748 11454 48750 11506
rect 48750 11454 48802 11506
rect 48802 11454 48804 11506
rect 48748 11452 48804 11454
rect 48860 10220 48916 10276
rect 48188 7980 48244 8036
rect 48300 7756 48356 7812
rect 48300 7420 48356 7476
rect 47852 3612 47908 3668
rect 48412 6188 48468 6244
rect 47516 3164 47572 3220
rect 46956 3052 47012 3108
rect 48412 2940 48468 2996
rect 47852 2546 47908 2548
rect 47852 2494 47854 2546
rect 47854 2494 47906 2546
rect 47906 2494 47908 2546
rect 47852 2492 47908 2494
rect 48188 2546 48244 2548
rect 48188 2494 48190 2546
rect 48190 2494 48242 2546
rect 48242 2494 48244 2546
rect 48188 2492 48244 2494
rect 47516 2380 47572 2436
rect 48412 2380 48468 2436
rect 47180 2156 47236 2212
rect 47292 2268 47348 2324
rect 48076 2210 48132 2212
rect 48076 2158 48078 2210
rect 48078 2158 48130 2210
rect 48130 2158 48132 2210
rect 48076 2156 48132 2158
rect 46956 1820 47012 1876
rect 46732 1372 46788 1428
rect 47404 1708 47460 1764
rect 46956 1202 47012 1204
rect 46956 1150 46958 1202
rect 46958 1150 47010 1202
rect 47010 1150 47012 1202
rect 46956 1148 47012 1150
rect 47292 1036 47348 1092
rect 46732 476 46788 532
rect 46844 924 46900 980
rect 47628 1596 47684 1652
rect 48412 2210 48468 2212
rect 48412 2158 48414 2210
rect 48414 2158 48466 2210
rect 48466 2158 48468 2210
rect 48412 2156 48468 2158
rect 48188 1820 48244 1876
rect 47740 700 47796 756
rect 48636 8540 48692 8596
rect 48972 9884 49028 9940
rect 49532 13916 49588 13972
rect 49308 13692 49364 13748
rect 49420 12348 49476 12404
rect 49420 10668 49476 10724
rect 49756 13692 49812 13748
rect 49644 13522 49700 13524
rect 49644 13470 49646 13522
rect 49646 13470 49698 13522
rect 49698 13470 49700 13522
rect 49644 13468 49700 13470
rect 50204 14812 50260 14868
rect 50428 14418 50484 14420
rect 50428 14366 50430 14418
rect 50430 14366 50482 14418
rect 50482 14366 50484 14418
rect 50428 14364 50484 14366
rect 50428 12908 50484 12964
rect 49308 10610 49364 10612
rect 49308 10558 49310 10610
rect 49310 10558 49362 10610
rect 49362 10558 49364 10610
rect 49308 10556 49364 10558
rect 49308 10108 49364 10164
rect 49644 10108 49700 10164
rect 49420 9884 49476 9940
rect 49308 9826 49364 9828
rect 49308 9774 49310 9826
rect 49310 9774 49362 9826
rect 49362 9774 49364 9826
rect 49308 9772 49364 9774
rect 49196 9660 49252 9716
rect 49308 9212 49364 9268
rect 48972 8540 49028 8596
rect 48860 7308 48916 7364
rect 48748 5852 48804 5908
rect 48636 5628 48692 5684
rect 48748 4508 48804 4564
rect 48972 5740 49028 5796
rect 48636 2828 48692 2884
rect 48748 3500 48804 3556
rect 48860 2716 48916 2772
rect 49084 3388 49140 3444
rect 49756 9884 49812 9940
rect 50316 12066 50372 12068
rect 50316 12014 50318 12066
rect 50318 12014 50370 12066
rect 50370 12014 50372 12066
rect 50316 12012 50372 12014
rect 50204 11788 50260 11844
rect 49532 8764 49588 8820
rect 49420 5180 49476 5236
rect 50204 9996 50260 10052
rect 49980 9212 50036 9268
rect 50876 14754 50932 14756
rect 50876 14702 50878 14754
rect 50878 14702 50930 14754
rect 50930 14702 50932 14754
rect 50876 14700 50932 14702
rect 50764 13580 50820 13636
rect 50652 12348 50708 12404
rect 50876 13356 50932 13412
rect 50988 12684 51044 12740
rect 51100 12348 51156 12404
rect 50764 11618 50820 11620
rect 50764 11566 50766 11618
rect 50766 11566 50818 11618
rect 50818 11566 50820 11618
rect 50764 11564 50820 11566
rect 50316 8764 50372 8820
rect 49868 7980 49924 8036
rect 49980 8652 50036 8708
rect 49868 7644 49924 7700
rect 49532 3276 49588 3332
rect 49756 5068 49812 5124
rect 49308 2604 49364 2660
rect 49196 2156 49252 2212
rect 48636 1484 48692 1540
rect 48300 588 48356 644
rect 48972 252 49028 308
rect 49196 1932 49252 1988
rect 49420 1036 49476 1092
rect 49868 1372 49924 1428
rect 50316 7980 50372 8036
rect 50204 3948 50260 4004
rect 50092 700 50148 756
rect 49644 364 49700 420
rect 49980 588 50036 644
rect 50316 252 50372 308
rect 49980 140 50036 196
rect 50540 9266 50596 9268
rect 50540 9214 50542 9266
rect 50542 9214 50594 9266
rect 50594 9214 50596 9266
rect 50540 9212 50596 9214
rect 50764 9826 50820 9828
rect 50764 9774 50766 9826
rect 50766 9774 50818 9826
rect 50818 9774 50820 9826
rect 50764 9772 50820 9774
rect 50764 8988 50820 9044
rect 50652 8092 50708 8148
rect 50540 6636 50596 6692
rect 50764 6300 50820 6356
rect 50764 3724 50820 3780
rect 51548 16380 51604 16436
rect 51436 16098 51492 16100
rect 51436 16046 51438 16098
rect 51438 16046 51490 16098
rect 51490 16046 51492 16098
rect 51436 16044 51492 16046
rect 52108 18562 52164 18564
rect 52108 18510 52110 18562
rect 52110 18510 52162 18562
rect 52162 18510 52164 18562
rect 52108 18508 52164 18510
rect 52108 18284 52164 18340
rect 51996 17890 52052 17892
rect 51996 17838 51998 17890
rect 51998 17838 52050 17890
rect 52050 17838 52052 17890
rect 51996 17836 52052 17838
rect 52108 17612 52164 17668
rect 52108 16380 52164 16436
rect 52108 15538 52164 15540
rect 52108 15486 52110 15538
rect 52110 15486 52162 15538
rect 52162 15486 52164 15538
rect 52108 15484 52164 15486
rect 51996 14700 52052 14756
rect 51884 13916 51940 13972
rect 51996 13804 52052 13860
rect 51772 12796 51828 12852
rect 51436 12738 51492 12740
rect 51436 12686 51438 12738
rect 51438 12686 51490 12738
rect 51490 12686 51492 12738
rect 51436 12684 51492 12686
rect 51324 11788 51380 11844
rect 50988 8316 51044 8372
rect 51436 9996 51492 10052
rect 51660 10108 51716 10164
rect 52556 21362 52612 21364
rect 52556 21310 52558 21362
rect 52558 21310 52610 21362
rect 52610 21310 52612 21362
rect 52556 21308 52612 21310
rect 54236 32284 54292 32340
rect 54348 34076 54404 34132
rect 54124 31890 54180 31892
rect 54124 31838 54126 31890
rect 54126 31838 54178 31890
rect 54178 31838 54180 31890
rect 54124 31836 54180 31838
rect 54348 31612 54404 31668
rect 54460 33964 54516 34020
rect 54460 31388 54516 31444
rect 54236 31276 54292 31332
rect 54348 30994 54404 30996
rect 54348 30942 54350 30994
rect 54350 30942 54402 30994
rect 54402 30942 54404 30994
rect 54348 30940 54404 30942
rect 54236 29932 54292 29988
rect 55692 36876 55748 36932
rect 56028 38050 56084 38052
rect 56028 37998 56030 38050
rect 56030 37998 56082 38050
rect 56082 37998 56084 38050
rect 56028 37996 56084 37998
rect 56588 41020 56644 41076
rect 56476 39452 56532 39508
rect 56588 38556 56644 38612
rect 57260 52892 57316 52948
rect 57036 47740 57092 47796
rect 57148 47852 57204 47908
rect 57036 47516 57092 47572
rect 56812 42028 56868 42084
rect 56924 44380 56980 44436
rect 56812 41580 56868 41636
rect 56812 38668 56868 38724
rect 56700 38444 56756 38500
rect 56588 38332 56644 38388
rect 56364 38162 56420 38164
rect 56364 38110 56366 38162
rect 56366 38110 56418 38162
rect 56418 38110 56420 38162
rect 56364 38108 56420 38110
rect 56476 37324 56532 37380
rect 55916 36594 55972 36596
rect 55916 36542 55918 36594
rect 55918 36542 55970 36594
rect 55970 36542 55972 36594
rect 55916 36540 55972 36542
rect 55804 36316 55860 36372
rect 55804 35868 55860 35924
rect 55916 34860 55972 34916
rect 55916 34690 55972 34692
rect 55916 34638 55918 34690
rect 55918 34638 55970 34690
rect 55970 34638 55972 34690
rect 55916 34636 55972 34638
rect 56252 36428 56308 36484
rect 56140 36316 56196 36372
rect 56252 36258 56308 36260
rect 56252 36206 56254 36258
rect 56254 36206 56306 36258
rect 56306 36206 56308 36258
rect 56252 36204 56308 36206
rect 56140 35474 56196 35476
rect 56140 35422 56142 35474
rect 56142 35422 56194 35474
rect 56194 35422 56196 35474
rect 56140 35420 56196 35422
rect 56140 35026 56196 35028
rect 56140 34974 56142 35026
rect 56142 34974 56194 35026
rect 56194 34974 56196 35026
rect 56140 34972 56196 34974
rect 56140 34802 56196 34804
rect 56140 34750 56142 34802
rect 56142 34750 56194 34802
rect 56194 34750 56196 34802
rect 56140 34748 56196 34750
rect 55692 34242 55748 34244
rect 55692 34190 55694 34242
rect 55694 34190 55746 34242
rect 55746 34190 55748 34242
rect 55692 34188 55748 34190
rect 55244 34076 55300 34132
rect 54796 31164 54852 31220
rect 55132 32338 55188 32340
rect 55132 32286 55134 32338
rect 55134 32286 55186 32338
rect 55186 32286 55188 32338
rect 55132 32284 55188 32286
rect 55244 32172 55300 32228
rect 55356 32060 55412 32116
rect 54908 30492 54964 30548
rect 55020 29708 55076 29764
rect 56476 36092 56532 36148
rect 56364 33852 56420 33908
rect 56812 38108 56868 38164
rect 56588 33628 56644 33684
rect 56700 37996 56756 38052
rect 55692 32450 55748 32452
rect 55692 32398 55694 32450
rect 55694 32398 55746 32450
rect 55746 32398 55748 32450
rect 55692 32396 55748 32398
rect 56028 31500 56084 31556
rect 55580 30604 55636 30660
rect 54348 29260 54404 29316
rect 55132 29036 55188 29092
rect 54012 28530 54068 28532
rect 54012 28478 54014 28530
rect 54014 28478 54066 28530
rect 54066 28478 54068 28530
rect 54012 28476 54068 28478
rect 54124 28140 54180 28196
rect 53900 28082 53956 28084
rect 53900 28030 53902 28082
rect 53902 28030 53954 28082
rect 53954 28030 53956 28082
rect 53900 28028 53956 28030
rect 53676 26684 53732 26740
rect 53788 27356 53844 27412
rect 53788 26460 53844 26516
rect 55020 28866 55076 28868
rect 55020 28814 55022 28866
rect 55022 28814 55074 28866
rect 55074 28814 55076 28866
rect 55020 28812 55076 28814
rect 54348 28700 54404 28756
rect 54796 28588 54852 28644
rect 54236 27132 54292 27188
rect 53900 26236 53956 26292
rect 54012 26796 54068 26852
rect 53564 26124 53620 26180
rect 54908 28252 54964 28308
rect 55020 27746 55076 27748
rect 55020 27694 55022 27746
rect 55022 27694 55074 27746
rect 55074 27694 55076 27746
rect 55020 27692 55076 27694
rect 55020 27298 55076 27300
rect 55020 27246 55022 27298
rect 55022 27246 55074 27298
rect 55074 27246 55076 27298
rect 55020 27244 55076 27246
rect 56140 30434 56196 30436
rect 56140 30382 56142 30434
rect 56142 30382 56194 30434
rect 56194 30382 56196 30434
rect 56140 30380 56196 30382
rect 55580 28588 55636 28644
rect 55804 30156 55860 30212
rect 54460 26684 54516 26740
rect 55244 27020 55300 27076
rect 54236 26124 54292 26180
rect 53564 25676 53620 25732
rect 53004 23996 53060 24052
rect 52892 23212 52948 23268
rect 54348 26012 54404 26068
rect 53900 25618 53956 25620
rect 53900 25566 53902 25618
rect 53902 25566 53954 25618
rect 53954 25566 53956 25618
rect 53900 25564 53956 25566
rect 54012 25116 54068 25172
rect 53340 24332 53396 24388
rect 53116 22876 53172 22932
rect 53228 23884 53284 23940
rect 53004 22146 53060 22148
rect 53004 22094 53006 22146
rect 53006 22094 53058 22146
rect 53058 22094 53060 22146
rect 53004 22092 53060 22094
rect 52892 21756 52948 21812
rect 52780 21196 52836 21252
rect 52892 21084 52948 21140
rect 52556 20802 52612 20804
rect 52556 20750 52558 20802
rect 52558 20750 52610 20802
rect 52610 20750 52612 20802
rect 52556 20748 52612 20750
rect 53004 20636 53060 20692
rect 52444 20300 52500 20356
rect 52668 19906 52724 19908
rect 52668 19854 52670 19906
rect 52670 19854 52722 19906
rect 52722 19854 52724 19906
rect 52668 19852 52724 19854
rect 52780 19516 52836 19572
rect 52444 18396 52500 18452
rect 52332 18338 52388 18340
rect 52332 18286 52334 18338
rect 52334 18286 52386 18338
rect 52386 18286 52388 18338
rect 52332 18284 52388 18286
rect 52668 18396 52724 18452
rect 52444 17948 52500 18004
rect 52332 17724 52388 17780
rect 52668 17948 52724 18004
rect 53228 19852 53284 19908
rect 53228 19292 53284 19348
rect 53116 19068 53172 19124
rect 53004 18674 53060 18676
rect 53004 18622 53006 18674
rect 53006 18622 53058 18674
rect 53058 18622 53060 18674
rect 53004 18620 53060 18622
rect 53116 18508 53172 18564
rect 53564 23212 53620 23268
rect 53788 23266 53844 23268
rect 53788 23214 53790 23266
rect 53790 23214 53842 23266
rect 53842 23214 53844 23266
rect 53788 23212 53844 23214
rect 53564 21756 53620 21812
rect 53452 19852 53508 19908
rect 53788 21532 53844 21588
rect 54236 24610 54292 24612
rect 54236 24558 54238 24610
rect 54238 24558 54290 24610
rect 54290 24558 54292 24610
rect 54236 24556 54292 24558
rect 54012 23938 54068 23940
rect 54012 23886 54014 23938
rect 54014 23886 54066 23938
rect 54066 23886 54068 23938
rect 54012 23884 54068 23886
rect 54236 23772 54292 23828
rect 55468 28028 55524 28084
rect 55356 26908 55412 26964
rect 55244 26684 55300 26740
rect 54796 26348 54852 26404
rect 54572 24780 54628 24836
rect 55580 26572 55636 26628
rect 55580 26236 55636 26292
rect 56476 32284 56532 32340
rect 56028 29372 56084 29428
rect 56476 30380 56532 30436
rect 56588 29820 56644 29876
rect 57148 41580 57204 41636
rect 57260 45276 57316 45332
rect 57036 41132 57092 41188
rect 57036 38444 57092 38500
rect 57036 32508 57092 32564
rect 57260 39676 57316 39732
rect 57260 37212 57316 37268
rect 57260 36988 57316 37044
rect 57260 36764 57316 36820
rect 57260 32060 57316 32116
rect 57372 33628 57428 33684
rect 57148 31612 57204 31668
rect 56924 31164 56980 31220
rect 57260 30716 57316 30772
rect 56812 30268 56868 30324
rect 56364 29372 56420 29428
rect 55916 29202 55972 29204
rect 55916 29150 55918 29202
rect 55918 29150 55970 29202
rect 55970 29150 55972 29202
rect 55916 29148 55972 29150
rect 55916 28866 55972 28868
rect 55916 28814 55918 28866
rect 55918 28814 55970 28866
rect 55970 28814 55972 28866
rect 55916 28812 55972 28814
rect 56364 28924 56420 28980
rect 55916 28588 55972 28644
rect 56140 28476 56196 28532
rect 56028 27634 56084 27636
rect 56028 27582 56030 27634
rect 56030 27582 56082 27634
rect 56082 27582 56084 27634
rect 56028 27580 56084 27582
rect 56476 28476 56532 28532
rect 55916 26962 55972 26964
rect 55916 26910 55918 26962
rect 55918 26910 55970 26962
rect 55970 26910 55972 26962
rect 55916 26908 55972 26910
rect 56140 27020 56196 27076
rect 56140 26290 56196 26292
rect 56140 26238 56142 26290
rect 56142 26238 56194 26290
rect 56194 26238 56196 26290
rect 56140 26236 56196 26238
rect 55692 25788 55748 25844
rect 55468 25228 55524 25284
rect 55020 24444 55076 24500
rect 54460 23212 54516 23268
rect 55244 24780 55300 24836
rect 54908 22876 54964 22932
rect 54684 22764 54740 22820
rect 54124 22594 54180 22596
rect 54124 22542 54126 22594
rect 54126 22542 54178 22594
rect 54178 22542 54180 22594
rect 54124 22540 54180 22542
rect 53676 19852 53732 19908
rect 54012 22092 54068 22148
rect 54012 21532 54068 21588
rect 53564 19346 53620 19348
rect 53564 19294 53566 19346
rect 53566 19294 53618 19346
rect 53618 19294 53620 19346
rect 53564 19292 53620 19294
rect 52892 18172 52948 18228
rect 53452 19180 53508 19236
rect 52444 17164 52500 17220
rect 52332 16098 52388 16100
rect 52332 16046 52334 16098
rect 52334 16046 52386 16098
rect 52386 16046 52388 16098
rect 52332 16044 52388 16046
rect 52556 14812 52612 14868
rect 53004 17164 53060 17220
rect 52780 14924 52836 14980
rect 52892 16492 52948 16548
rect 53116 16770 53172 16772
rect 53116 16718 53118 16770
rect 53118 16718 53170 16770
rect 53170 16718 53172 16770
rect 53116 16716 53172 16718
rect 53004 15484 53060 15540
rect 53676 18620 53732 18676
rect 53564 18508 53620 18564
rect 53452 17948 53508 18004
rect 53676 18060 53732 18116
rect 53564 17106 53620 17108
rect 53564 17054 53566 17106
rect 53566 17054 53618 17106
rect 53618 17054 53620 17106
rect 53564 17052 53620 17054
rect 53340 16380 53396 16436
rect 53452 16322 53508 16324
rect 53452 16270 53454 16322
rect 53454 16270 53506 16322
rect 53506 16270 53508 16322
rect 53452 16268 53508 16270
rect 53340 15260 53396 15316
rect 52668 14476 52724 14532
rect 53004 14924 53060 14980
rect 52556 13634 52612 13636
rect 52556 13582 52558 13634
rect 52558 13582 52610 13634
rect 52610 13582 52612 13634
rect 52556 13580 52612 13582
rect 52220 13356 52276 13412
rect 51996 12348 52052 12404
rect 52332 12962 52388 12964
rect 52332 12910 52334 12962
rect 52334 12910 52386 12962
rect 52386 12910 52388 12962
rect 52332 12908 52388 12910
rect 52556 12348 52612 12404
rect 52108 11788 52164 11844
rect 51884 11618 51940 11620
rect 51884 11566 51886 11618
rect 51886 11566 51938 11618
rect 51938 11566 51940 11618
rect 51884 11564 51940 11566
rect 51996 10610 52052 10612
rect 51996 10558 51998 10610
rect 51998 10558 52050 10610
rect 52050 10558 52052 10610
rect 51996 10556 52052 10558
rect 51772 9548 51828 9604
rect 51884 10108 51940 10164
rect 51996 9996 52052 10052
rect 51100 7868 51156 7924
rect 51436 7644 51492 7700
rect 51548 7420 51604 7476
rect 51212 6188 51268 6244
rect 51324 7084 51380 7140
rect 51100 3388 51156 3444
rect 50876 1260 50932 1316
rect 50876 1036 50932 1092
rect 50540 978 50596 980
rect 50540 926 50542 978
rect 50542 926 50594 978
rect 50594 926 50596 978
rect 50540 924 50596 926
rect 51772 6076 51828 6132
rect 51548 4732 51604 4788
rect 51996 8092 52052 8148
rect 52892 14530 52948 14532
rect 52892 14478 52894 14530
rect 52894 14478 52946 14530
rect 52946 14478 52948 14530
rect 52892 14476 52948 14478
rect 53340 14754 53396 14756
rect 53340 14702 53342 14754
rect 53342 14702 53394 14754
rect 53394 14702 53396 14754
rect 53340 14700 53396 14702
rect 53116 14028 53172 14084
rect 53676 16492 53732 16548
rect 53900 19852 53956 19908
rect 54124 21756 54180 21812
rect 54460 20748 54516 20804
rect 54124 20636 54180 20692
rect 54460 20188 54516 20244
rect 54348 19794 54404 19796
rect 54348 19742 54350 19794
rect 54350 19742 54402 19794
rect 54402 19742 54404 19794
rect 54348 19740 54404 19742
rect 54572 19740 54628 19796
rect 54236 19346 54292 19348
rect 54236 19294 54238 19346
rect 54238 19294 54290 19346
rect 54290 19294 54292 19346
rect 54236 19292 54292 19294
rect 54012 18172 54068 18228
rect 54124 17276 54180 17332
rect 54460 19234 54516 19236
rect 54460 19182 54462 19234
rect 54462 19182 54514 19234
rect 54514 19182 54516 19234
rect 54460 19180 54516 19182
rect 54460 18172 54516 18228
rect 54012 17052 54068 17108
rect 54236 16716 54292 16772
rect 54348 15820 54404 15876
rect 53676 15484 53732 15540
rect 53564 15148 53620 15204
rect 53788 14364 53844 14420
rect 53676 14028 53732 14084
rect 53116 13804 53172 13860
rect 53004 13634 53060 13636
rect 53004 13582 53006 13634
rect 53006 13582 53058 13634
rect 53058 13582 53060 13634
rect 53004 13580 53060 13582
rect 53452 13522 53508 13524
rect 53452 13470 53454 13522
rect 53454 13470 53506 13522
rect 53506 13470 53508 13522
rect 53452 13468 53508 13470
rect 53340 12796 53396 12852
rect 52332 11564 52388 11620
rect 52444 11788 52500 11844
rect 53004 11788 53060 11844
rect 52556 11564 52612 11620
rect 52220 10386 52276 10388
rect 52220 10334 52222 10386
rect 52222 10334 52274 10386
rect 52274 10334 52276 10386
rect 52220 10332 52276 10334
rect 53116 11228 53172 11284
rect 53004 11004 53060 11060
rect 52892 10556 52948 10612
rect 52220 9772 52276 9828
rect 52668 10444 52724 10500
rect 52332 9100 52388 9156
rect 52220 8764 52276 8820
rect 52332 8092 52388 8148
rect 52220 7868 52276 7924
rect 52108 6188 52164 6244
rect 51884 1372 51940 1428
rect 52108 2940 52164 2996
rect 51772 700 51828 756
rect 52108 700 52164 756
rect 52556 9548 52612 9604
rect 52668 9042 52724 9044
rect 52668 8990 52670 9042
rect 52670 8990 52722 9042
rect 52722 8990 52724 9042
rect 52668 8988 52724 8990
rect 52668 8764 52724 8820
rect 52892 9324 52948 9380
rect 52780 8428 52836 8484
rect 52892 8204 52948 8260
rect 52556 7362 52612 7364
rect 52556 7310 52558 7362
rect 52558 7310 52610 7362
rect 52610 7310 52612 7362
rect 52556 7308 52612 7310
rect 52444 6130 52500 6132
rect 52444 6078 52446 6130
rect 52446 6078 52498 6130
rect 52498 6078 52500 6130
rect 52444 6076 52500 6078
rect 52668 6076 52724 6132
rect 52556 5180 52612 5236
rect 52332 4060 52388 4116
rect 52556 4732 52612 4788
rect 52668 4508 52724 4564
rect 52668 1036 52724 1092
rect 53004 7644 53060 7700
rect 53452 12124 53508 12180
rect 53564 12012 53620 12068
rect 53564 11564 53620 11620
rect 53452 9996 53508 10052
rect 53564 10892 53620 10948
rect 53340 8988 53396 9044
rect 53452 9100 53508 9156
rect 54124 13244 54180 13300
rect 54012 12178 54068 12180
rect 54012 12126 54014 12178
rect 54014 12126 54066 12178
rect 54066 12126 54068 12178
rect 54012 12124 54068 12126
rect 53788 10892 53844 10948
rect 53676 10556 53732 10612
rect 53788 10668 53844 10724
rect 53676 9996 53732 10052
rect 54012 9938 54068 9940
rect 54012 9886 54014 9938
rect 54014 9886 54066 9938
rect 54066 9886 54068 9938
rect 54012 9884 54068 9886
rect 53228 8764 53284 8820
rect 53340 7868 53396 7924
rect 53340 7644 53396 7700
rect 53228 7196 53284 7252
rect 53340 6524 53396 6580
rect 53564 8930 53620 8932
rect 53564 8878 53566 8930
rect 53566 8878 53618 8930
rect 53618 8878 53620 8930
rect 53564 8876 53620 8878
rect 54124 9212 54180 9268
rect 53788 8764 53844 8820
rect 53676 7868 53732 7924
rect 53900 8428 53956 8484
rect 53564 7532 53620 7588
rect 53788 7250 53844 7252
rect 53788 7198 53790 7250
rect 53790 7198 53842 7250
rect 53842 7198 53844 7250
rect 53788 7196 53844 7198
rect 53564 6636 53620 6692
rect 53676 6578 53732 6580
rect 53676 6526 53678 6578
rect 53678 6526 53730 6578
rect 53730 6526 53732 6578
rect 53676 6524 53732 6526
rect 53564 5964 53620 6020
rect 53116 5068 53172 5124
rect 54124 8370 54180 8372
rect 54124 8318 54126 8370
rect 54126 8318 54178 8370
rect 54178 8318 54180 8370
rect 54124 8316 54180 8318
rect 54124 6914 54180 6916
rect 54124 6862 54126 6914
rect 54126 6862 54178 6914
rect 54178 6862 54180 6914
rect 54124 6860 54180 6862
rect 54684 19404 54740 19460
rect 54684 18396 54740 18452
rect 54796 18284 54852 18340
rect 54684 17500 54740 17556
rect 55244 22146 55300 22148
rect 55244 22094 55246 22146
rect 55246 22094 55298 22146
rect 55298 22094 55300 22146
rect 55244 22092 55300 22094
rect 55468 24498 55524 24500
rect 55468 24446 55470 24498
rect 55470 24446 55522 24498
rect 55522 24446 55524 24498
rect 55468 24444 55524 24446
rect 55356 21980 55412 22036
rect 55020 20188 55076 20244
rect 55916 25340 55972 25396
rect 55916 23436 55972 23492
rect 57148 27580 57204 27636
rect 57036 27132 57092 27188
rect 56588 26684 56644 26740
rect 56924 26236 56980 26292
rect 56812 24892 56868 24948
rect 56252 23212 56308 23268
rect 55692 21868 55748 21924
rect 56588 23884 56644 23940
rect 55692 21698 55748 21700
rect 55692 21646 55694 21698
rect 55694 21646 55746 21698
rect 55746 21646 55748 21698
rect 55692 21644 55748 21646
rect 55580 20972 55636 21028
rect 55692 21196 55748 21252
rect 55356 20188 55412 20244
rect 55468 19794 55524 19796
rect 55468 19742 55470 19794
rect 55470 19742 55522 19794
rect 55522 19742 55524 19794
rect 55468 19740 55524 19742
rect 55356 19068 55412 19124
rect 55244 18172 55300 18228
rect 54908 17778 54964 17780
rect 54908 17726 54910 17778
rect 54910 17726 54962 17778
rect 54962 17726 54964 17778
rect 54908 17724 54964 17726
rect 55020 17666 55076 17668
rect 55020 17614 55022 17666
rect 55022 17614 55074 17666
rect 55074 17614 55076 17666
rect 55020 17612 55076 17614
rect 54684 16940 54740 16996
rect 54908 16716 54964 16772
rect 54684 16098 54740 16100
rect 54684 16046 54686 16098
rect 54686 16046 54738 16098
rect 54738 16046 54740 16098
rect 54684 16044 54740 16046
rect 55132 17164 55188 17220
rect 55020 16268 55076 16324
rect 55132 16604 55188 16660
rect 54572 15820 54628 15876
rect 54572 15484 54628 15540
rect 54460 14642 54516 14644
rect 54460 14590 54462 14642
rect 54462 14590 54514 14642
rect 54514 14590 54516 14642
rect 54460 14588 54516 14590
rect 54908 15202 54964 15204
rect 54908 15150 54910 15202
rect 54910 15150 54962 15202
rect 54962 15150 54964 15202
rect 54908 15148 54964 15150
rect 54348 13580 54404 13636
rect 54572 14140 54628 14196
rect 54908 13244 54964 13300
rect 54684 13186 54740 13188
rect 54684 13134 54686 13186
rect 54686 13134 54738 13186
rect 54738 13134 54740 13186
rect 54684 13132 54740 13134
rect 54460 12066 54516 12068
rect 54460 12014 54462 12066
rect 54462 12014 54514 12066
rect 54514 12014 54516 12066
rect 54460 12012 54516 12014
rect 54460 10332 54516 10388
rect 54348 8764 54404 8820
rect 54460 6412 54516 6468
rect 54348 6300 54404 6356
rect 53564 4284 53620 4340
rect 53564 4060 53620 4116
rect 52780 812 52836 868
rect 53116 3052 53172 3108
rect 54012 3724 54068 3780
rect 56812 23884 56868 23940
rect 56700 23772 56756 23828
rect 56028 22092 56084 22148
rect 56028 21362 56084 21364
rect 56028 21310 56030 21362
rect 56030 21310 56082 21362
rect 56082 21310 56084 21362
rect 56028 21308 56084 21310
rect 56140 20188 56196 20244
rect 56364 21026 56420 21028
rect 56364 20974 56366 21026
rect 56366 20974 56418 21026
rect 56418 20974 56420 21026
rect 56364 20972 56420 20974
rect 55916 19628 55972 19684
rect 56028 19458 56084 19460
rect 56028 19406 56030 19458
rect 56030 19406 56082 19458
rect 56082 19406 56084 19458
rect 56028 19404 56084 19406
rect 56364 19458 56420 19460
rect 56364 19406 56366 19458
rect 56366 19406 56418 19458
rect 56418 19406 56420 19458
rect 56364 19404 56420 19406
rect 56252 19180 56308 19236
rect 55356 17836 55412 17892
rect 55468 18172 55524 18228
rect 55132 13468 55188 13524
rect 55244 15708 55300 15764
rect 55132 12124 55188 12180
rect 55132 11900 55188 11956
rect 55020 11676 55076 11732
rect 55020 10386 55076 10388
rect 55020 10334 55022 10386
rect 55022 10334 55074 10386
rect 55074 10334 55076 10386
rect 55020 10332 55076 10334
rect 55356 15484 55412 15540
rect 55356 10556 55412 10612
rect 54796 7980 54852 8036
rect 54908 5794 54964 5796
rect 54908 5742 54910 5794
rect 54910 5742 54962 5794
rect 54962 5742 54964 5794
rect 54908 5740 54964 5742
rect 55692 17948 55748 18004
rect 55804 17724 55860 17780
rect 55804 17276 55860 17332
rect 55580 14812 55636 14868
rect 55692 13916 55748 13972
rect 55692 12348 55748 12404
rect 55580 11954 55636 11956
rect 55580 11902 55582 11954
rect 55582 11902 55634 11954
rect 55634 11902 55636 11954
rect 55580 11900 55636 11902
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 55468 8540 55524 8596
rect 55020 4620 55076 4676
rect 55468 6524 55524 6580
rect 55468 5292 55524 5348
rect 55356 3778 55412 3780
rect 55356 3726 55358 3778
rect 55358 3726 55410 3778
rect 55410 3726 55412 3778
rect 55356 3724 55412 3726
rect 54348 1484 54404 1540
rect 54908 3612 54964 3668
rect 54236 140 54292 196
rect 54460 1372 54516 1428
rect 56364 18338 56420 18340
rect 56364 18286 56366 18338
rect 56366 18286 56418 18338
rect 56418 18286 56420 18338
rect 56364 18284 56420 18286
rect 56364 17890 56420 17892
rect 56364 17838 56366 17890
rect 56366 17838 56418 17890
rect 56418 17838 56420 17890
rect 56364 17836 56420 17838
rect 56028 16322 56084 16324
rect 56028 16270 56030 16322
rect 56030 16270 56082 16322
rect 56082 16270 56084 16322
rect 56028 16268 56084 16270
rect 56028 16044 56084 16100
rect 56364 16322 56420 16324
rect 56364 16270 56366 16322
rect 56366 16270 56418 16322
rect 56418 16270 56420 16322
rect 56364 16268 56420 16270
rect 56252 16156 56308 16212
rect 56140 15538 56196 15540
rect 56140 15486 56142 15538
rect 56142 15486 56194 15538
rect 56194 15486 56196 15538
rect 56140 15484 56196 15486
rect 56028 14754 56084 14756
rect 56028 14702 56030 14754
rect 56030 14702 56082 14754
rect 56082 14702 56084 14754
rect 56028 14700 56084 14702
rect 56140 14252 56196 14308
rect 56140 13468 56196 13524
rect 55916 12236 55972 12292
rect 56028 11116 56084 11172
rect 56028 10610 56084 10612
rect 56028 10558 56030 10610
rect 56030 10558 56082 10610
rect 56082 10558 56084 10610
rect 56028 10556 56084 10558
rect 56364 14364 56420 14420
rect 56812 23212 56868 23268
rect 56700 19180 56756 19236
rect 56700 16268 56756 16324
rect 56588 14476 56644 14532
rect 56924 19292 56980 19348
rect 56812 14252 56868 14308
rect 56924 19068 56980 19124
rect 56588 13020 56644 13076
rect 56140 10332 56196 10388
rect 56252 11900 56308 11956
rect 55916 9660 55972 9716
rect 56028 9100 56084 9156
rect 56364 11618 56420 11620
rect 56364 11566 56366 11618
rect 56366 11566 56418 11618
rect 56418 11566 56420 11618
rect 56364 11564 56420 11566
rect 56364 10498 56420 10500
rect 56364 10446 56366 10498
rect 56366 10446 56418 10498
rect 56418 10446 56420 10498
rect 56364 10444 56420 10446
rect 56364 10050 56420 10052
rect 56364 9998 56366 10050
rect 56366 9998 56418 10050
rect 56418 9998 56420 10050
rect 56364 9996 56420 9998
rect 56364 8988 56420 9044
rect 56028 7756 56084 7812
rect 55916 6636 55972 6692
rect 55916 4956 55972 5012
rect 57260 25340 57316 25396
rect 57260 23772 57316 23828
rect 57260 22652 57316 22708
rect 57148 19404 57204 19460
rect 57036 17836 57092 17892
rect 57148 17724 57204 17780
rect 57036 14588 57092 14644
rect 56252 7084 56308 7140
rect 56364 8204 56420 8260
rect 57148 8204 57204 8260
rect 56252 6412 56308 6468
rect 56140 5740 56196 5796
rect 56252 5122 56308 5124
rect 56252 5070 56254 5122
rect 56254 5070 56306 5122
rect 56306 5070 56308 5122
rect 56252 5068 56308 5070
rect 55916 4172 55972 4228
rect 57260 14140 57316 14196
rect 56588 7644 56644 7700
rect 57372 8988 57428 9044
rect 55804 3164 55860 3220
rect 55244 2658 55300 2660
rect 55244 2606 55246 2658
rect 55246 2606 55298 2658
rect 55298 2606 55300 2658
rect 55244 2604 55300 2606
rect 55916 2828 55972 2884
rect 56252 3052 56308 3108
rect 56924 3052 56980 3108
rect 57036 5068 57092 5124
rect 55804 1484 55860 1540
rect 55356 1260 55412 1316
rect 24276 28 24332 84
<< metal3 >>
rect 41692 57372 46844 57428
rect 46900 57372 46910 57428
rect 48514 57372 48524 57428
rect 48580 57372 55412 57428
rect 41692 57316 41748 57372
rect 55356 57316 55412 57372
rect 2156 57260 10108 57316
rect 10164 57260 10174 57316
rect 41682 57260 41692 57316
rect 41748 57260 41758 57316
rect 43698 57260 43708 57316
rect 43764 57260 45276 57316
rect 45332 57260 45342 57316
rect 46162 57260 46172 57316
rect 46228 57260 54012 57316
rect 54068 57260 54078 57316
rect 55346 57260 55356 57316
rect 55412 57260 55422 57316
rect 0 57204 112 57232
rect 2156 57204 2212 57260
rect 57344 57204 57456 57232
rect 0 57148 924 57204
rect 980 57148 990 57204
rect 2146 57148 2156 57204
rect 2212 57148 2222 57204
rect 2370 57148 2380 57204
rect 2436 57148 4284 57204
rect 4340 57148 4350 57204
rect 4620 57148 6188 57204
rect 6244 57148 6254 57204
rect 22754 57148 22764 57204
rect 22820 57148 32060 57204
rect 32116 57148 32126 57204
rect 34514 57148 34524 57204
rect 34580 57148 50540 57204
rect 50596 57148 50606 57204
rect 52098 57148 52108 57204
rect 52164 57148 57456 57204
rect 0 57120 112 57148
rect 4620 57092 4676 57148
rect 57344 57120 57456 57148
rect 1586 57036 1596 57092
rect 1652 57036 4676 57092
rect 5730 57036 5740 57092
rect 5796 57036 14140 57092
rect 14196 57036 14206 57092
rect 21298 57036 21308 57092
rect 21364 57036 26908 57092
rect 30594 57036 30604 57092
rect 30660 57036 38444 57092
rect 38500 57036 38510 57092
rect 40786 57036 40796 57092
rect 40852 57036 46620 57092
rect 46676 57036 46686 57092
rect 46834 57036 46844 57092
rect 46900 57036 50876 57092
rect 50932 57036 50942 57092
rect 26852 56980 26908 57036
rect 1698 56924 1708 56980
rect 1764 56924 9212 56980
rect 9268 56924 9278 56980
rect 16482 56924 16492 56980
rect 16548 56924 25340 56980
rect 25396 56924 25406 56980
rect 26852 56924 41020 56980
rect 41076 56924 41086 56980
rect 43474 56924 43484 56980
rect 43540 56924 54908 56980
rect 54964 56924 54974 56980
rect 578 56812 588 56868
rect 644 56812 2380 56868
rect 2436 56812 2446 56868
rect 3042 56812 3052 56868
rect 3108 56812 11452 56868
rect 11508 56812 11518 56868
rect 11890 56812 11900 56868
rect 11956 56812 24892 56868
rect 24948 56812 24958 56868
rect 26674 56812 26684 56868
rect 26740 56812 27804 56868
rect 27860 56812 27870 56868
rect 31378 56812 31388 56868
rect 31444 56812 37324 56868
rect 37380 56812 37390 56868
rect 44258 56812 44268 56868
rect 44324 56812 45052 56868
rect 45108 56812 45118 56868
rect 45266 56812 45276 56868
rect 45332 56812 49532 56868
rect 49588 56812 49598 56868
rect 51986 56812 51996 56868
rect 52052 56812 56252 56868
rect 56308 56812 56318 56868
rect 0 56756 112 56784
rect 57344 56756 57456 56784
rect 0 56700 476 56756
rect 532 56700 542 56756
rect 690 56700 700 56756
rect 756 56700 3388 56756
rect 3602 56700 3612 56756
rect 3668 56700 13244 56756
rect 13300 56700 13310 56756
rect 13458 56700 13468 56756
rect 13524 56700 18620 56756
rect 18676 56700 18686 56756
rect 18834 56700 18844 56756
rect 18900 56700 22204 56756
rect 22260 56700 22270 56756
rect 31714 56700 31724 56756
rect 31780 56700 45164 56756
rect 45220 56700 45230 56756
rect 48626 56700 48636 56756
rect 48692 56700 53228 56756
rect 53284 56700 53294 56756
rect 55794 56700 55804 56756
rect 55860 56700 57456 56756
rect 0 56672 112 56700
rect 3332 56644 3388 56700
rect 57344 56672 57456 56700
rect 3332 56588 11676 56644
rect 11732 56588 11742 56644
rect 11890 56588 11900 56644
rect 11956 56588 18172 56644
rect 18228 56588 18238 56644
rect 28242 56588 28252 56644
rect 28308 56588 38668 56644
rect 42130 56588 42140 56644
rect 42196 56588 44212 56644
rect 44370 56588 44380 56644
rect 44436 56588 44828 56644
rect 44884 56588 44894 56644
rect 47058 56588 47068 56644
rect 47124 56588 53116 56644
rect 53172 56588 53182 56644
rect 38612 56532 38668 56588
rect 44156 56532 44212 56588
rect 4274 56476 4284 56532
rect 4340 56476 5068 56532
rect 5124 56476 5134 56532
rect 10770 56476 10780 56532
rect 10836 56476 17724 56532
rect 17780 56476 17790 56532
rect 18610 56476 18620 56532
rect 18676 56476 20412 56532
rect 20468 56476 20478 56532
rect 24434 56476 24444 56532
rect 24500 56476 30380 56532
rect 30436 56476 30446 56532
rect 31826 56476 31836 56532
rect 31892 56476 36820 56532
rect 38612 56476 38780 56532
rect 38836 56476 38846 56532
rect 41010 56476 41020 56532
rect 41076 56476 43596 56532
rect 43652 56476 43662 56532
rect 44156 56476 46284 56532
rect 46340 56476 46350 56532
rect 48626 56476 48636 56532
rect 48692 56476 49084 56532
rect 49140 56476 49150 56532
rect 49746 56476 49756 56532
rect 49812 56476 52220 56532
rect 52276 56476 52286 56532
rect 52434 56476 52444 56532
rect 52500 56476 55020 56532
rect 55076 56476 55086 56532
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 36764 56420 36820 56476
rect 43794 56420 43804 56476
rect 43860 56420 43908 56476
rect 43964 56420 44012 56476
rect 44068 56420 44078 56476
rect 3378 56364 3388 56420
rect 3444 56364 3482 56420
rect 4162 56364 4172 56420
rect 4228 56364 7420 56420
rect 7476 56364 7486 56420
rect 7858 56364 7868 56420
rect 7924 56364 9324 56420
rect 9380 56364 9390 56420
rect 10098 56364 10108 56420
rect 10164 56364 16828 56420
rect 16884 56364 16894 56420
rect 17602 56364 17612 56420
rect 17668 56364 21644 56420
rect 21700 56364 21710 56420
rect 24332 56364 25116 56420
rect 25172 56364 25182 56420
rect 27580 56364 34972 56420
rect 35028 56364 35038 56420
rect 35522 56364 35532 56420
rect 35588 56364 36540 56420
rect 36596 56364 36606 56420
rect 36764 56364 38668 56420
rect 42802 56364 42812 56420
rect 42868 56364 43260 56420
rect 43316 56364 43326 56420
rect 44146 56364 44156 56420
rect 44212 56364 54460 56420
rect 54516 56364 54526 56420
rect 0 56308 112 56336
rect 24332 56308 24388 56364
rect 27580 56308 27636 56364
rect 38612 56308 38668 56364
rect 57344 56308 57456 56336
rect 0 56252 252 56308
rect 308 56252 318 56308
rect 2370 56252 2380 56308
rect 2436 56252 4732 56308
rect 4788 56252 4798 56308
rect 5058 56252 5068 56308
rect 5124 56252 6076 56308
rect 6132 56252 6142 56308
rect 8204 56252 12348 56308
rect 12404 56252 12414 56308
rect 13234 56252 13244 56308
rect 13300 56252 18732 56308
rect 18788 56252 18798 56308
rect 19068 56252 24388 56308
rect 24546 56252 24556 56308
rect 24612 56252 27636 56308
rect 27794 56252 27804 56308
rect 27860 56252 31612 56308
rect 31668 56252 31678 56308
rect 33170 56252 33180 56308
rect 33236 56252 37716 56308
rect 38612 56252 43820 56308
rect 43876 56252 43886 56308
rect 44146 56252 44156 56308
rect 44212 56252 44548 56308
rect 44706 56252 44716 56308
rect 44772 56252 51884 56308
rect 51940 56252 51950 56308
rect 53900 56252 57456 56308
rect 0 56224 112 56252
rect 8204 56196 8260 56252
rect 19068 56196 19124 56252
rect 37660 56196 37716 56252
rect 44492 56196 44548 56252
rect 2258 56140 2268 56196
rect 2324 56140 8260 56196
rect 9426 56140 9436 56196
rect 9492 56140 19124 56196
rect 19282 56140 19292 56196
rect 19348 56140 28140 56196
rect 28196 56140 28206 56196
rect 29474 56140 29484 56196
rect 29540 56140 30492 56196
rect 30548 56140 31500 56196
rect 31556 56140 31566 56196
rect 36866 56140 36876 56196
rect 36932 56140 37436 56196
rect 37492 56140 37502 56196
rect 37660 56140 44268 56196
rect 44324 56140 44334 56196
rect 44492 56140 45276 56196
rect 45332 56140 45342 56196
rect 45490 56140 45500 56196
rect 45556 56140 46284 56196
rect 46340 56140 46350 56196
rect 47730 56140 47740 56196
rect 47796 56140 52668 56196
rect 52724 56140 52734 56196
rect 2902 56028 2940 56084
rect 2996 56028 3006 56084
rect 3332 56028 5628 56084
rect 5684 56028 5694 56084
rect 6290 56028 6300 56084
rect 6356 56028 14588 56084
rect 14644 56028 14654 56084
rect 18162 56028 18172 56084
rect 18228 56028 20860 56084
rect 20916 56028 20926 56084
rect 27094 56028 27132 56084
rect 27188 56028 27198 56084
rect 30258 56028 30268 56084
rect 30324 56028 31724 56084
rect 31780 56028 31790 56084
rect 32470 56028 32508 56084
rect 32564 56028 32574 56084
rect 33366 56028 33404 56084
rect 33460 56028 33470 56084
rect 34710 56028 34748 56084
rect 34804 56028 34814 56084
rect 36418 56028 36428 56084
rect 36484 56028 36988 56084
rect 37044 56028 37054 56084
rect 42326 56028 42364 56084
rect 42420 56028 42430 56084
rect 42588 56028 45836 56084
rect 45892 56028 45902 56084
rect 48178 56028 48188 56084
rect 48244 56028 52556 56084
rect 52612 56028 52622 56084
rect 0 55860 112 55888
rect 0 55804 812 55860
rect 868 55804 878 55860
rect 0 55776 112 55804
rect 690 55692 700 55748
rect 756 55692 1148 55748
rect 1204 55692 1214 55748
rect 3332 55524 3388 56028
rect 42588 55972 42644 56028
rect 3938 55916 3948 55972
rect 4004 55916 11004 55972
rect 11060 55916 11070 55972
rect 11228 55916 15036 55972
rect 15092 55916 15102 55972
rect 16818 55916 16828 55972
rect 16884 55916 19068 55972
rect 19124 55916 19134 55972
rect 19954 55916 19964 55972
rect 20020 55916 20412 55972
rect 20468 55916 20478 55972
rect 21942 55916 21980 55972
rect 22036 55916 22046 55972
rect 22642 55916 22652 55972
rect 22708 55916 23100 55972
rect 23156 55916 23166 55972
rect 25778 55916 25788 55972
rect 25844 55916 25900 55972
rect 25956 55916 25966 55972
rect 26898 55916 26908 55972
rect 26964 55916 29932 55972
rect 29988 55916 29998 55972
rect 32722 55916 32732 55972
rect 32788 55916 42644 55972
rect 43026 55916 43036 55972
rect 43092 55916 45948 55972
rect 46004 55916 46014 55972
rect 49074 55916 49084 55972
rect 49140 55916 53564 55972
rect 53620 55916 53630 55972
rect 11228 55860 11284 55916
rect 3490 55804 3500 55860
rect 3556 55804 6804 55860
rect 6962 55804 6972 55860
rect 7028 55804 11284 55860
rect 11554 55804 11564 55860
rect 11620 55804 17164 55860
rect 17220 55804 17230 55860
rect 19506 55804 19516 55860
rect 19572 55804 22540 55860
rect 22596 55804 22606 55860
rect 22978 55804 22988 55860
rect 23044 55804 25340 55860
rect 25396 55804 25406 55860
rect 26422 55804 26460 55860
rect 26516 55804 26526 55860
rect 27458 55804 27468 55860
rect 27524 55804 27916 55860
rect 27972 55804 27982 55860
rect 29558 55804 29596 55860
rect 29652 55804 29662 55860
rect 30034 55804 30044 55860
rect 30100 55804 30268 55860
rect 30324 55804 30334 55860
rect 31714 55804 31724 55860
rect 31780 55804 32284 55860
rect 32340 55804 32350 55860
rect 33730 55804 33740 55860
rect 33796 55804 34300 55860
rect 34356 55804 34366 55860
rect 35746 55804 35756 55860
rect 35812 55804 36092 55860
rect 36148 55804 36158 55860
rect 37090 55804 37100 55860
rect 37156 55804 37324 55860
rect 37380 55804 37390 55860
rect 38098 55804 38108 55860
rect 38164 55804 38556 55860
rect 38612 55804 38622 55860
rect 39078 55804 39116 55860
rect 39172 55804 39182 55860
rect 41122 55804 41132 55860
rect 41188 55804 44492 55860
rect 44548 55804 44558 55860
rect 44818 55804 44828 55860
rect 44884 55804 44940 55860
rect 44996 55804 45006 55860
rect 47366 55804 47404 55860
rect 47460 55804 47470 55860
rect 48402 55804 48412 55860
rect 48468 55804 51548 55860
rect 51604 55804 51614 55860
rect 52098 55804 52108 55860
rect 52164 55804 52892 55860
rect 52948 55804 52958 55860
rect 6748 55748 6804 55804
rect 53900 55748 53956 56252
rect 57344 56224 57456 56252
rect 57344 55860 57456 55888
rect 54310 55804 54348 55860
rect 54404 55804 54414 55860
rect 55570 55804 55580 55860
rect 55636 55804 55692 55860
rect 55748 55804 55758 55860
rect 55916 55804 57456 55860
rect 55916 55748 55972 55804
rect 57344 55776 57456 55804
rect 6748 55692 10668 55748
rect 10724 55692 10734 55748
rect 11778 55692 11788 55748
rect 11844 55692 13356 55748
rect 13412 55692 13422 55748
rect 28802 55692 28812 55748
rect 28868 55692 29820 55748
rect 29876 55692 29886 55748
rect 30930 55692 30940 55748
rect 30996 55692 33516 55748
rect 33572 55692 33582 55748
rect 33842 55692 33852 55748
rect 33908 55692 35196 55748
rect 35252 55692 35262 55748
rect 38658 55692 38668 55748
rect 38724 55692 44156 55748
rect 44212 55692 44222 55748
rect 45276 55692 48972 55748
rect 49028 55692 49038 55748
rect 49186 55692 49196 55748
rect 49252 55692 53956 55748
rect 54226 55692 54236 55748
rect 54292 55692 55972 55748
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 44454 55636 44464 55692
rect 44520 55636 44568 55692
rect 44624 55636 44672 55692
rect 44728 55636 44738 55692
rect 4918 55580 4956 55636
rect 5012 55580 5022 55636
rect 6738 55580 6748 55636
rect 6804 55580 7308 55636
rect 7364 55580 7374 55636
rect 7634 55580 7644 55636
rect 7700 55580 14812 55636
rect 14868 55580 14878 55636
rect 19170 55580 19180 55636
rect 19236 55580 21756 55636
rect 21812 55580 21822 55636
rect 26114 55580 26124 55636
rect 26180 55580 27692 55636
rect 27748 55580 27758 55636
rect 29250 55580 29260 55636
rect 29316 55580 35308 55636
rect 35364 55580 35374 55636
rect 41430 55580 41468 55636
rect 41524 55580 41534 55636
rect 42802 55580 42812 55636
rect 42868 55580 43260 55636
rect 43316 55580 43326 55636
rect 43586 55580 43596 55636
rect 43652 55580 44268 55636
rect 44324 55580 44334 55636
rect 44930 55580 44940 55636
rect 44996 55580 45052 55636
rect 45108 55580 45118 55636
rect 45276 55524 45332 55692
rect 45490 55580 45500 55636
rect 45556 55580 45948 55636
rect 46004 55580 46014 55636
rect 46722 55580 46732 55636
rect 46788 55580 47628 55636
rect 47684 55580 47694 55636
rect 51090 55580 51100 55636
rect 51156 55580 53732 55636
rect 56242 55580 56252 55636
rect 56308 55580 56812 55636
rect 56868 55580 56878 55636
rect 53676 55524 53732 55580
rect 2258 55468 2268 55524
rect 2324 55468 3388 55524
rect 4498 55468 4508 55524
rect 4564 55468 5964 55524
rect 6020 55468 6030 55524
rect 6514 55468 6524 55524
rect 6580 55468 8148 55524
rect 8754 55468 8764 55524
rect 8820 55468 9436 55524
rect 9492 55468 9502 55524
rect 9622 55468 9660 55524
rect 9716 55468 9726 55524
rect 10434 55468 10444 55524
rect 10500 55468 15148 55524
rect 17938 55468 17948 55524
rect 18004 55468 19796 55524
rect 23202 55468 23212 55524
rect 23268 55468 25284 55524
rect 25778 55468 25788 55524
rect 25844 55468 26236 55524
rect 26292 55468 26302 55524
rect 27542 55468 27580 55524
rect 27636 55468 27646 55524
rect 27990 55468 28028 55524
rect 28084 55468 28094 55524
rect 29334 55468 29372 55524
rect 29428 55468 29438 55524
rect 30678 55468 30716 55524
rect 30772 55468 30782 55524
rect 34290 55468 34300 55524
rect 34356 55468 34524 55524
rect 34580 55468 34590 55524
rect 35410 55468 35420 55524
rect 35476 55468 35756 55524
rect 35812 55468 35822 55524
rect 37762 55468 37772 55524
rect 37828 55468 38332 55524
rect 38388 55468 38398 55524
rect 40226 55468 40236 55524
rect 40292 55468 41916 55524
rect 41972 55468 41982 55524
rect 43474 55468 43484 55524
rect 43540 55468 45332 55524
rect 46050 55468 46060 55524
rect 46116 55468 46396 55524
rect 46452 55468 46462 55524
rect 46806 55468 46844 55524
rect 46900 55468 46910 55524
rect 47254 55468 47292 55524
rect 47348 55468 47358 55524
rect 48738 55468 48748 55524
rect 48804 55468 48972 55524
rect 49028 55468 49038 55524
rect 49382 55468 49420 55524
rect 49476 55468 49486 55524
rect 49942 55468 49980 55524
rect 50036 55468 50046 55524
rect 50838 55468 50876 55524
rect 50932 55468 50942 55524
rect 51314 55468 51324 55524
rect 51380 55468 52668 55524
rect 52724 55468 52734 55524
rect 53676 55468 55804 55524
rect 55860 55468 55870 55524
rect 0 55412 112 55440
rect 8092 55412 8148 55468
rect 15092 55412 15148 55468
rect 19740 55412 19796 55468
rect 25228 55412 25284 55468
rect 57344 55412 57456 55440
rect 0 55356 1092 55412
rect 1250 55356 1260 55412
rect 1316 55356 1708 55412
rect 1764 55356 1774 55412
rect 3490 55356 3500 55412
rect 3556 55356 4956 55412
rect 5012 55356 5022 55412
rect 6850 55356 6860 55412
rect 6916 55356 6972 55412
rect 7028 55356 7038 55412
rect 8092 55356 9548 55412
rect 9604 55356 9614 55412
rect 9874 55356 9884 55412
rect 9940 55356 14476 55412
rect 14532 55356 14542 55412
rect 15092 55356 15820 55412
rect 15876 55356 15886 55412
rect 17490 55356 17500 55412
rect 17556 55356 19516 55412
rect 19572 55356 19582 55412
rect 19740 55356 20860 55412
rect 20916 55356 20926 55412
rect 21084 55356 23548 55412
rect 23604 55356 23614 55412
rect 25228 55356 29484 55412
rect 29540 55356 29550 55412
rect 29810 55356 29820 55412
rect 29876 55356 30156 55412
rect 30212 55356 30222 55412
rect 30454 55356 30492 55412
rect 30548 55356 30558 55412
rect 30818 55356 30828 55412
rect 30884 55356 32396 55412
rect 32452 55356 32462 55412
rect 33814 55356 33852 55412
rect 33908 55356 33918 55412
rect 34178 55356 34188 55412
rect 34244 55356 34524 55412
rect 34580 55356 34590 55412
rect 36278 55356 36316 55412
rect 36372 55356 36382 55412
rect 37538 55356 37548 55412
rect 37604 55356 37884 55412
rect 37940 55356 37950 55412
rect 38882 55356 38892 55412
rect 38948 55356 39452 55412
rect 39508 55356 39518 55412
rect 40562 55356 40572 55412
rect 40628 55356 40684 55412
rect 40740 55356 40750 55412
rect 41122 55356 41132 55412
rect 41188 55356 44492 55412
rect 44548 55356 44558 55412
rect 46172 55356 46508 55412
rect 46564 55356 46574 55412
rect 47842 55356 47852 55412
rect 47908 55356 51212 55412
rect 51268 55356 51278 55412
rect 52434 55356 52444 55412
rect 52500 55356 54684 55412
rect 54740 55356 54750 55412
rect 54908 55356 57456 55412
rect 0 55328 112 55356
rect 1036 55300 1092 55356
rect 21084 55300 21140 55356
rect 46172 55300 46228 55356
rect 1036 55244 3052 55300
rect 3108 55244 3118 55300
rect 3266 55244 3276 55300
rect 3332 55244 4508 55300
rect 4564 55244 4574 55300
rect 6066 55244 6076 55300
rect 6132 55244 6524 55300
rect 6580 55244 6590 55300
rect 8082 55244 8092 55300
rect 8148 55244 8204 55300
rect 8260 55244 8270 55300
rect 8530 55244 8540 55300
rect 8596 55244 9100 55300
rect 9156 55244 9166 55300
rect 10406 55244 10444 55300
rect 10500 55244 10510 55300
rect 11890 55244 11900 55300
rect 11956 55244 13804 55300
rect 13860 55244 13870 55300
rect 14802 55244 14812 55300
rect 14868 55244 15372 55300
rect 15428 55244 15438 55300
rect 15586 55244 15596 55300
rect 15652 55244 17612 55300
rect 17668 55244 17678 55300
rect 17826 55244 17836 55300
rect 17892 55244 19404 55300
rect 19460 55244 19470 55300
rect 19730 55244 19740 55300
rect 19796 55244 21140 55300
rect 21634 55244 21644 55300
rect 21700 55244 21756 55300
rect 21812 55244 21822 55300
rect 22502 55244 22540 55300
rect 22596 55244 22606 55300
rect 26898 55244 26908 55300
rect 26964 55244 27002 55300
rect 29586 55244 29596 55300
rect 29652 55244 30828 55300
rect 30884 55244 30894 55300
rect 31154 55244 31164 55300
rect 31220 55244 32172 55300
rect 32228 55244 32238 55300
rect 32498 55244 32508 55300
rect 32564 55244 32732 55300
rect 32788 55244 32798 55300
rect 33618 55244 33628 55300
rect 33684 55244 35196 55300
rect 35252 55244 35262 55300
rect 40002 55244 40012 55300
rect 40068 55244 43820 55300
rect 43876 55244 43886 55300
rect 44118 55244 44156 55300
rect 44212 55244 44222 55300
rect 44370 55244 44380 55300
rect 44436 55244 46228 55300
rect 46358 55244 46396 55300
rect 46452 55244 46462 55300
rect 46610 55244 46620 55300
rect 46676 55244 51996 55300
rect 52052 55244 52062 55300
rect 53974 55244 54012 55300
rect 54068 55244 54078 55300
rect 54908 55188 54964 55356
rect 57344 55328 57456 55356
rect 3266 55132 3276 55188
rect 3332 55132 4060 55188
rect 4116 55132 4126 55188
rect 5058 55132 5068 55188
rect 5124 55132 6972 55188
rect 7028 55132 7038 55188
rect 8306 55132 8316 55188
rect 8372 55132 24780 55188
rect 24836 55132 24846 55188
rect 28802 55132 28812 55188
rect 28868 55132 33180 55188
rect 33236 55132 33246 55188
rect 33394 55132 33404 55188
rect 33460 55132 38668 55188
rect 38724 55132 38734 55188
rect 42578 55132 42588 55188
rect 42644 55132 46060 55188
rect 46116 55132 46126 55188
rect 48066 55132 48076 55188
rect 48132 55132 50428 55188
rect 50484 55132 50494 55188
rect 51426 55132 51436 55188
rect 51492 55132 54964 55188
rect 3378 55020 3388 55076
rect 3444 55020 4284 55076
rect 4340 55020 4844 55076
rect 4900 55020 4910 55076
rect 5282 55020 5292 55076
rect 5348 55020 12460 55076
rect 12516 55020 12526 55076
rect 12786 55020 12796 55076
rect 12852 55020 13132 55076
rect 13188 55020 13198 55076
rect 13458 55020 13468 55076
rect 13524 55020 15372 55076
rect 15428 55020 15438 55076
rect 15586 55020 15596 55076
rect 15652 55020 16716 55076
rect 16772 55020 16782 55076
rect 17154 55020 17164 55076
rect 17220 55020 17388 55076
rect 17444 55020 18284 55076
rect 18340 55020 18350 55076
rect 18498 55020 18508 55076
rect 18564 55020 22876 55076
rect 22932 55020 22942 55076
rect 26852 55020 41356 55076
rect 41412 55020 41422 55076
rect 43250 55020 43260 55076
rect 43316 55020 46732 55076
rect 46788 55020 46798 55076
rect 47964 55020 53452 55076
rect 53508 55020 53518 55076
rect 0 54964 112 54992
rect 0 54908 140 54964
rect 196 54908 206 54964
rect 6402 54908 6412 54964
rect 6468 54908 10220 54964
rect 10276 54908 10286 54964
rect 12114 54908 12124 54964
rect 12180 54908 16380 54964
rect 16436 54908 16446 54964
rect 16818 54908 16828 54964
rect 16884 54908 20076 54964
rect 20132 54908 20142 54964
rect 0 54880 112 54908
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 3378 54796 3388 54852
rect 3444 54796 3482 54852
rect 4274 54796 4284 54852
rect 4340 54796 13692 54852
rect 13748 54796 13758 54852
rect 16482 54796 16492 54852
rect 16548 54796 19740 54852
rect 19796 54796 19806 54852
rect 20290 54796 20300 54852
rect 20356 54796 20636 54852
rect 20692 54796 20702 54852
rect 26852 54740 26908 55020
rect 47964 54964 48020 55020
rect 57344 54964 57456 54992
rect 29138 54908 29148 54964
rect 29204 54908 33292 54964
rect 33348 54908 33358 54964
rect 33506 54908 33516 54964
rect 33572 54908 41804 54964
rect 41860 54908 41870 54964
rect 42354 54908 42364 54964
rect 42420 54908 43596 54964
rect 43652 54908 43662 54964
rect 44146 54908 44156 54964
rect 44212 54908 45724 54964
rect 45780 54908 45790 54964
rect 45938 54908 45948 54964
rect 46004 54908 48020 54964
rect 48178 54908 48188 54964
rect 48244 54908 50316 54964
rect 50372 54908 50382 54964
rect 53900 54908 57456 54964
rect 43794 54852 43804 54908
rect 43860 54852 43908 54908
rect 43964 54852 44012 54908
rect 44068 54852 44078 54908
rect 27122 54796 27132 54852
rect 27188 54796 30380 54852
rect 30436 54796 30446 54852
rect 32386 54796 32396 54852
rect 32452 54796 37772 54852
rect 37828 54796 37838 54852
rect 38098 54796 38108 54852
rect 38164 54796 41580 54852
rect 41636 54796 41646 54852
rect 42018 54796 42028 54852
rect 42084 54796 43484 54852
rect 43540 54796 43550 54852
rect 44258 54796 44268 54852
rect 44324 54796 45220 54852
rect 45350 54796 45388 54852
rect 45444 54796 45454 54852
rect 45836 54796 50652 54852
rect 50708 54796 50718 54852
rect 45164 54740 45220 54796
rect 45836 54740 45892 54796
rect 1922 54684 1932 54740
rect 1988 54684 10332 54740
rect 10388 54684 10398 54740
rect 11442 54684 11452 54740
rect 11508 54684 12796 54740
rect 12852 54684 12862 54740
rect 13010 54684 13020 54740
rect 13076 54684 21756 54740
rect 21812 54684 21822 54740
rect 23762 54684 23772 54740
rect 23828 54684 26908 54740
rect 28578 54684 28588 54740
rect 28644 54684 29148 54740
rect 29204 54684 29214 54740
rect 30258 54684 30268 54740
rect 30324 54684 37548 54740
rect 37604 54684 37614 54740
rect 37762 54684 37772 54740
rect 37828 54684 38668 54740
rect 38724 54684 38734 54740
rect 41234 54684 41244 54740
rect 41300 54684 44940 54740
rect 44996 54684 45006 54740
rect 45164 54684 45892 54740
rect 46050 54684 46060 54740
rect 46116 54684 48524 54740
rect 48580 54684 48590 54740
rect 48738 54684 48748 54740
rect 48804 54684 49980 54740
rect 50036 54684 50046 54740
rect 51986 54684 51996 54740
rect 52052 54684 53676 54740
rect 53732 54684 53742 54740
rect 53900 54628 53956 54908
rect 57344 54880 57456 54908
rect 2594 54572 2604 54628
rect 2660 54572 8988 54628
rect 9044 54572 9054 54628
rect 10658 54572 10668 54628
rect 10724 54572 11004 54628
rect 11060 54572 11070 54628
rect 11890 54572 11900 54628
rect 11956 54572 13132 54628
rect 13188 54572 13198 54628
rect 13346 54572 13356 54628
rect 13412 54572 14924 54628
rect 14980 54572 14990 54628
rect 15474 54572 15484 54628
rect 15540 54572 16044 54628
rect 16100 54572 16110 54628
rect 16370 54572 16380 54628
rect 16436 54572 17276 54628
rect 17332 54572 17342 54628
rect 17500 54572 24556 54628
rect 24612 54572 24622 54628
rect 28690 54572 28700 54628
rect 28756 54572 29372 54628
rect 29428 54572 29438 54628
rect 31266 54572 31276 54628
rect 31332 54572 32844 54628
rect 32900 54572 32910 54628
rect 33170 54572 33180 54628
rect 33236 54572 36540 54628
rect 36596 54572 36606 54628
rect 38770 54572 38780 54628
rect 38836 54572 39564 54628
rect 39620 54572 39630 54628
rect 39890 54572 39900 54628
rect 39956 54572 40460 54628
rect 40516 54572 40526 54628
rect 42130 54572 42140 54628
rect 42196 54572 53956 54628
rect 54460 54572 56308 54628
rect 0 54516 112 54544
rect 17500 54516 17556 54572
rect 54460 54516 54516 54572
rect 56252 54516 56308 54572
rect 57344 54516 57456 54544
rect 0 54460 1372 54516
rect 1428 54460 1438 54516
rect 2706 54460 2716 54516
rect 2772 54460 3276 54516
rect 3332 54460 3342 54516
rect 4274 54460 4284 54516
rect 4340 54460 6692 54516
rect 7074 54460 7084 54516
rect 7140 54460 9772 54516
rect 9828 54460 9838 54516
rect 10882 54460 10892 54516
rect 10948 54460 17556 54516
rect 18274 54460 18284 54516
rect 18340 54460 21196 54516
rect 21252 54460 21262 54516
rect 25666 54460 25676 54516
rect 25732 54460 26572 54516
rect 26628 54460 26638 54516
rect 27570 54460 27580 54516
rect 27636 54460 27646 54516
rect 28914 54460 28924 54516
rect 28980 54460 39844 54516
rect 0 54432 112 54460
rect 6636 54404 6692 54460
rect 27580 54404 27636 54460
rect 39788 54404 39844 54460
rect 40684 54460 40908 54516
rect 40964 54460 42700 54516
rect 42756 54460 42766 54516
rect 44482 54460 44492 54516
rect 44548 54460 46004 54516
rect 46134 54460 46172 54516
rect 46228 54460 46238 54516
rect 46498 54460 46508 54516
rect 46564 54460 50092 54516
rect 50148 54460 50158 54516
rect 51314 54460 51324 54516
rect 51380 54460 54516 54516
rect 54674 54460 54684 54516
rect 54740 54460 56028 54516
rect 56084 54460 56094 54516
rect 56252 54460 57456 54516
rect 40684 54404 40740 54460
rect 45948 54404 46004 54460
rect 57344 54432 57456 54460
rect 914 54348 924 54404
rect 980 54348 2492 54404
rect 2548 54348 2558 54404
rect 2930 54348 2940 54404
rect 2996 54348 3164 54404
rect 3220 54348 3230 54404
rect 3332 54348 4452 54404
rect 5926 54348 5964 54404
rect 6020 54348 6030 54404
rect 6636 54348 7532 54404
rect 7588 54348 7598 54404
rect 8978 54348 8988 54404
rect 9044 54348 11900 54404
rect 11956 54348 11966 54404
rect 12124 54348 14756 54404
rect 14914 54348 14924 54404
rect 14980 54348 18340 54404
rect 18498 54348 18508 54404
rect 18564 54348 18620 54404
rect 18676 54348 18686 54404
rect 18946 54348 18956 54404
rect 19012 54348 22428 54404
rect 22484 54348 22494 54404
rect 26114 54348 26124 54404
rect 26180 54348 26460 54404
rect 26516 54348 26526 54404
rect 26674 54348 26684 54404
rect 26740 54348 27524 54404
rect 27580 54348 34916 54404
rect 35074 54348 35084 54404
rect 35140 54348 39564 54404
rect 39620 54348 39630 54404
rect 39788 54348 40740 54404
rect 41906 54348 41916 54404
rect 41972 54348 45388 54404
rect 45444 54348 45454 54404
rect 45948 54348 48636 54404
rect 48692 54348 48702 54404
rect 48860 54348 55916 54404
rect 55972 54348 55982 54404
rect 3332 54292 3388 54348
rect 1810 54236 1820 54292
rect 1876 54236 3388 54292
rect 4396 54292 4452 54348
rect 12124 54292 12180 54348
rect 4396 54236 7644 54292
rect 7700 54236 7710 54292
rect 9734 54236 9772 54292
rect 9828 54236 9838 54292
rect 10546 54236 10556 54292
rect 10612 54236 12180 54292
rect 14130 54236 14140 54292
rect 14196 54236 14476 54292
rect 14532 54236 14542 54292
rect 14700 54180 14756 54348
rect 18284 54292 18340 54348
rect 27468 54292 27524 54348
rect 34860 54292 34916 54348
rect 48860 54292 48916 54348
rect 15138 54236 15148 54292
rect 15204 54236 15242 54292
rect 15362 54236 15372 54292
rect 15428 54236 15820 54292
rect 15876 54236 16268 54292
rect 16324 54236 16334 54292
rect 18284 54236 23100 54292
rect 23156 54236 23166 54292
rect 23398 54236 23436 54292
rect 23492 54236 23502 54292
rect 23874 54236 23884 54292
rect 23940 54236 26908 54292
rect 27206 54236 27244 54292
rect 27300 54236 27310 54292
rect 27458 54236 27468 54292
rect 27524 54236 27534 54292
rect 27878 54236 27916 54292
rect 27972 54236 27982 54292
rect 28140 54236 32396 54292
rect 32452 54236 32462 54292
rect 32834 54236 32844 54292
rect 32900 54236 33068 54292
rect 33124 54236 33134 54292
rect 34860 54236 36876 54292
rect 36932 54236 36942 54292
rect 40422 54236 40460 54292
rect 40516 54236 40526 54292
rect 41794 54236 41804 54292
rect 41860 54236 44716 54292
rect 44772 54236 44782 54292
rect 47282 54236 47292 54292
rect 47348 54236 48916 54292
rect 50082 54236 50092 54292
rect 50148 54236 53900 54292
rect 53956 54236 53966 54292
rect 54338 54236 54348 54292
rect 54404 54236 55468 54292
rect 55524 54236 55534 54292
rect 55682 54236 55692 54292
rect 55748 54236 56028 54292
rect 56084 54236 56094 54292
rect 26852 54180 26908 54236
rect 28140 54180 28196 54236
rect 690 54124 700 54180
rect 756 54124 4340 54180
rect 4844 54124 5292 54180
rect 5348 54124 5358 54180
rect 6626 54124 6636 54180
rect 6692 54124 7644 54180
rect 7700 54124 7710 54180
rect 7858 54124 7868 54180
rect 7924 54124 12684 54180
rect 12740 54124 12750 54180
rect 14018 54124 14028 54180
rect 14084 54124 14476 54180
rect 14532 54124 14542 54180
rect 14700 54124 18396 54180
rect 18452 54124 18462 54180
rect 18722 54124 18732 54180
rect 18788 54124 19292 54180
rect 19348 54124 19358 54180
rect 20822 54124 20860 54180
rect 20916 54124 20926 54180
rect 25330 54124 25340 54180
rect 25396 54124 25564 54180
rect 25620 54124 25630 54180
rect 26852 54124 28196 54180
rect 28466 54124 28476 54180
rect 28532 54124 42812 54180
rect 42868 54124 43036 54180
rect 43092 54124 43102 54180
rect 45154 54124 45164 54180
rect 45220 54124 48748 54180
rect 48804 54124 48814 54180
rect 48962 54124 48972 54180
rect 49028 54124 50428 54180
rect 55122 54124 55132 54180
rect 55188 54124 55356 54180
rect 55412 54124 55422 54180
rect 0 54068 112 54096
rect 0 54012 1260 54068
rect 1316 54012 1326 54068
rect 3602 54012 3612 54068
rect 3668 54012 3724 54068
rect 3780 54012 3790 54068
rect 0 53984 112 54012
rect 4284 53956 4340 54124
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 4844 53956 4900 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 44454 54068 44464 54124
rect 44520 54068 44568 54124
rect 44624 54068 44672 54124
rect 44728 54068 44738 54124
rect 50372 54068 50428 54124
rect 57344 54068 57456 54096
rect 5394 54012 5404 54068
rect 5460 54012 18564 54068
rect 18722 54012 18732 54068
rect 18788 54012 19516 54068
rect 19572 54012 19582 54068
rect 19926 54012 19964 54068
rect 20020 54012 20030 54068
rect 20178 54012 20188 54068
rect 20244 54012 22092 54068
rect 22148 54012 22158 54068
rect 24892 54012 27804 54068
rect 27860 54012 27870 54068
rect 32386 54012 32396 54068
rect 32452 54012 32844 54068
rect 32900 54012 32910 54068
rect 35634 54012 35644 54068
rect 35700 54012 36652 54068
rect 36708 54012 36718 54068
rect 36866 54012 36876 54068
rect 36932 54012 40908 54068
rect 40964 54012 40974 54068
rect 43362 54012 43372 54068
rect 43428 54012 43988 54068
rect 46274 54012 46284 54068
rect 46340 54012 48524 54068
rect 48580 54012 48590 54068
rect 48850 54012 48860 54068
rect 48916 54012 49420 54068
rect 49476 54012 49486 54068
rect 50372 54012 57456 54068
rect 18508 53956 18564 54012
rect 24892 53956 24948 54012
rect 43932 53956 43988 54012
rect 57344 53984 57456 54012
rect 1138 53900 1148 53956
rect 1204 53900 4060 53956
rect 4116 53900 4126 53956
rect 4284 53900 4900 53956
rect 5058 53900 5068 53956
rect 5124 53900 6412 53956
rect 6468 53900 6478 53956
rect 7970 53900 7980 53956
rect 8036 53900 8428 53956
rect 8484 53900 8494 53956
rect 9874 53900 9884 53956
rect 9940 53900 13244 53956
rect 13300 53900 13310 53956
rect 15092 53900 15932 53956
rect 15988 53900 15998 53956
rect 18508 53900 20524 53956
rect 20580 53900 20590 53956
rect 23090 53900 23100 53956
rect 23156 53900 24948 53956
rect 26338 53900 26348 53956
rect 26404 53900 28476 53956
rect 28532 53900 28542 53956
rect 31938 53900 31948 53956
rect 32004 53900 32508 53956
rect 32564 53900 32574 53956
rect 34178 53900 34188 53956
rect 34244 53900 35084 53956
rect 35140 53900 35150 53956
rect 35298 53900 35308 53956
rect 35364 53900 38668 53956
rect 43474 53900 43484 53956
rect 43540 53900 43876 53956
rect 43932 53900 53564 53956
rect 53620 53900 53630 53956
rect 53778 53900 53788 53956
rect 53844 53900 55132 53956
rect 55188 53900 55198 53956
rect 15092 53844 15148 53900
rect 38612 53844 38668 53900
rect 43820 53844 43876 53900
rect 3154 53788 3164 53844
rect 3220 53788 3388 53844
rect 3444 53788 3454 53844
rect 3602 53788 3612 53844
rect 3668 53788 5180 53844
rect 5236 53788 5246 53844
rect 7270 53788 7308 53844
rect 7364 53788 7374 53844
rect 8316 53788 15148 53844
rect 18386 53788 18396 53844
rect 18452 53788 18462 53844
rect 18610 53788 18620 53844
rect 18676 53788 21980 53844
rect 22036 53788 22046 53844
rect 24098 53788 24108 53844
rect 24164 53788 25564 53844
rect 25620 53788 25630 53844
rect 25778 53788 25788 53844
rect 25844 53788 26628 53844
rect 26786 53788 26796 53844
rect 26852 53788 27132 53844
rect 27188 53788 27198 53844
rect 27458 53788 27468 53844
rect 27524 53788 31108 53844
rect 31266 53788 31276 53844
rect 31332 53788 35196 53844
rect 35252 53788 35262 53844
rect 35522 53788 35532 53844
rect 35588 53788 35756 53844
rect 35812 53788 35822 53844
rect 36754 53788 36764 53844
rect 36820 53788 36876 53844
rect 36932 53788 36942 53844
rect 38612 53788 39452 53844
rect 39508 53788 39518 53844
rect 43138 53788 43148 53844
rect 43204 53788 43596 53844
rect 43652 53788 43764 53844
rect 43820 53788 49196 53844
rect 49252 53788 49262 53844
rect 53676 53788 54180 53844
rect 8316 53732 8372 53788
rect 18396 53732 18452 53788
rect 1922 53676 1932 53732
rect 1988 53676 8372 53732
rect 9986 53676 9996 53732
rect 10052 53676 12012 53732
rect 12068 53676 12078 53732
rect 12422 53676 12460 53732
rect 12516 53676 12526 53732
rect 12674 53676 12684 53732
rect 12740 53676 13804 53732
rect 13860 53676 14252 53732
rect 14308 53676 14318 53732
rect 15026 53676 15036 53732
rect 15092 53676 15708 53732
rect 15764 53676 15774 53732
rect 18396 53676 21924 53732
rect 22054 53676 22092 53732
rect 22148 53676 22158 53732
rect 22950 53676 22988 53732
rect 23044 53676 23054 53732
rect 24658 53676 24668 53732
rect 24724 53676 25452 53732
rect 25508 53676 25518 53732
rect 25666 53676 25676 53732
rect 25732 53676 26348 53732
rect 26404 53676 26414 53732
rect 0 53620 112 53648
rect 21868 53620 21924 53676
rect 0 53564 924 53620
rect 980 53564 990 53620
rect 1250 53564 1260 53620
rect 1316 53564 5628 53620
rect 5684 53564 6636 53620
rect 6692 53564 6702 53620
rect 7410 53564 7420 53620
rect 7476 53564 9660 53620
rect 9716 53564 9726 53620
rect 10994 53564 11004 53620
rect 11060 53564 11340 53620
rect 11396 53564 11564 53620
rect 11620 53564 11630 53620
rect 13682 53564 13692 53620
rect 13748 53564 20188 53620
rect 20244 53564 20254 53620
rect 21074 53564 21084 53620
rect 21140 53564 21196 53620
rect 21252 53564 21532 53620
rect 21588 53564 21598 53620
rect 21868 53564 23324 53620
rect 23380 53564 23390 53620
rect 23548 53564 24220 53620
rect 24276 53564 24286 53620
rect 25218 53564 25228 53620
rect 25284 53564 25788 53620
rect 25844 53564 25854 53620
rect 0 53536 112 53564
rect 3378 53452 3388 53508
rect 3444 53452 3482 53508
rect 3612 53452 6972 53508
rect 7028 53452 7038 53508
rect 7186 53452 7196 53508
rect 7252 53452 8876 53508
rect 8932 53452 9772 53508
rect 9828 53452 9838 53508
rect 10322 53452 10332 53508
rect 10388 53452 10668 53508
rect 10724 53452 11676 53508
rect 11732 53452 11742 53508
rect 12908 53452 15820 53508
rect 15876 53452 15886 53508
rect 16930 53452 16940 53508
rect 16996 53452 18844 53508
rect 18900 53452 18910 53508
rect 19068 53452 22092 53508
rect 22148 53452 22158 53508
rect 22418 53452 22428 53508
rect 22484 53452 22764 53508
rect 22820 53452 23324 53508
rect 23380 53452 23390 53508
rect 3612 53396 3668 53452
rect 12908 53396 12964 53452
rect 16940 53396 16996 53452
rect 19068 53396 19124 53452
rect 23548 53396 23604 53564
rect 26572 53508 26628 53788
rect 27794 53676 27804 53732
rect 27860 53676 29260 53732
rect 29316 53676 29326 53732
rect 31052 53620 31108 53788
rect 43708 53732 43764 53788
rect 31462 53676 31500 53732
rect 31556 53676 31566 53732
rect 31714 53676 31724 53732
rect 31780 53676 32396 53732
rect 32452 53676 32462 53732
rect 32722 53676 32732 53732
rect 32788 53676 34860 53732
rect 34916 53676 34926 53732
rect 42130 53676 42140 53732
rect 42196 53676 43372 53732
rect 43428 53676 43438 53732
rect 43708 53676 44604 53732
rect 44660 53676 44670 53732
rect 45266 53676 45276 53732
rect 45332 53676 47180 53732
rect 47236 53676 47246 53732
rect 47478 53676 47516 53732
rect 47572 53676 47582 53732
rect 48178 53676 48188 53732
rect 48244 53676 49084 53732
rect 49140 53676 49150 53732
rect 50726 53676 50764 53732
rect 50820 53676 50830 53732
rect 51510 53676 51548 53732
rect 51604 53676 51614 53732
rect 52518 53676 52556 53732
rect 52612 53676 52622 53732
rect 53676 53620 53732 53788
rect 54124 53732 54180 53788
rect 53862 53676 53900 53732
rect 53956 53676 53966 53732
rect 54124 53676 54684 53732
rect 54740 53676 54750 53732
rect 57344 53620 57456 53648
rect 27682 53564 27692 53620
rect 27748 53564 30828 53620
rect 30884 53564 30894 53620
rect 31052 53564 31556 53620
rect 32162 53564 32172 53620
rect 32228 53564 34972 53620
rect 35028 53564 35038 53620
rect 35252 53564 35420 53620
rect 35476 53564 36540 53620
rect 36596 53564 37772 53620
rect 37828 53564 37838 53620
rect 43250 53564 43260 53620
rect 43316 53564 46508 53620
rect 46564 53564 46574 53620
rect 48514 53564 48524 53620
rect 48580 53564 51884 53620
rect 51940 53564 51950 53620
rect 52108 53564 53732 53620
rect 53788 53564 57456 53620
rect 31500 53508 31556 53564
rect 35252 53508 35308 53564
rect 52108 53508 52164 53564
rect 3490 53340 3500 53396
rect 3556 53340 3668 53396
rect 5730 53340 5740 53396
rect 5796 53340 7420 53396
rect 7476 53340 7486 53396
rect 7634 53340 7644 53396
rect 7700 53340 9996 53396
rect 10052 53340 10062 53396
rect 10770 53340 10780 53396
rect 10836 53340 12964 53396
rect 14018 53340 14028 53396
rect 14084 53340 16996 53396
rect 17378 53340 17388 53396
rect 17444 53340 19124 53396
rect 20290 53340 20300 53396
rect 20356 53340 23604 53396
rect 23660 53452 26796 53508
rect 26852 53452 26862 53508
rect 27346 53452 27356 53508
rect 27412 53452 30604 53508
rect 30660 53452 30670 53508
rect 31126 53452 31164 53508
rect 31220 53452 31230 53508
rect 31490 53452 31500 53508
rect 31556 53452 31566 53508
rect 32834 53452 32844 53508
rect 32900 53452 34076 53508
rect 34132 53452 34636 53508
rect 34692 53452 35308 53508
rect 40450 53452 40460 53508
rect 40516 53452 42700 53508
rect 42756 53452 44212 53508
rect 44482 53452 44492 53508
rect 44548 53452 45164 53508
rect 45220 53452 45230 53508
rect 45938 53452 45948 53508
rect 46004 53452 50540 53508
rect 50596 53452 50606 53508
rect 51090 53452 51100 53508
rect 51156 53452 52164 53508
rect 52546 53452 52556 53508
rect 52612 53452 53564 53508
rect 53620 53452 53630 53508
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 14028 53284 14084 53340
rect 17388 53284 17444 53340
rect 23660 53284 23716 53452
rect 24210 53340 24220 53396
rect 24276 53340 25116 53396
rect 25172 53340 26796 53396
rect 26852 53340 26862 53396
rect 28690 53340 28700 53396
rect 28756 53340 41132 53396
rect 41188 53340 41198 53396
rect 41570 53340 41580 53396
rect 41636 53340 43652 53396
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 4162 53228 4172 53284
rect 4228 53228 6076 53284
rect 6132 53228 6142 53284
rect 6850 53228 6860 53284
rect 6916 53228 8652 53284
rect 8708 53228 8718 53284
rect 9314 53228 9324 53284
rect 9380 53228 10444 53284
rect 10500 53228 10510 53284
rect 10658 53228 10668 53284
rect 10724 53228 14084 53284
rect 14242 53228 14252 53284
rect 14308 53228 17444 53284
rect 19954 53228 19964 53284
rect 20020 53228 23100 53284
rect 23156 53228 23716 53284
rect 24210 53228 24220 53284
rect 24276 53228 26236 53284
rect 26292 53228 27916 53284
rect 27972 53228 27982 53284
rect 28466 53228 28476 53284
rect 28532 53228 43372 53284
rect 43428 53228 43438 53284
rect 0 53172 112 53200
rect 43596 53172 43652 53340
rect 43794 53284 43804 53340
rect 43860 53284 43908 53340
rect 43964 53284 44012 53340
rect 44068 53284 44078 53340
rect 44156 53284 44212 53452
rect 53788 53396 53844 53564
rect 57344 53536 57456 53564
rect 44370 53340 44380 53396
rect 44436 53340 45276 53396
rect 45332 53340 45342 53396
rect 45490 53340 45500 53396
rect 45556 53340 53844 53396
rect 44156 53228 46956 53284
rect 47012 53228 47022 53284
rect 48626 53228 48636 53284
rect 48692 53228 52668 53284
rect 52724 53228 52734 53284
rect 53442 53228 53452 53284
rect 53508 53228 55244 53284
rect 55300 53228 55310 53284
rect 57344 53172 57456 53200
rect 0 53116 812 53172
rect 868 53116 878 53172
rect 2818 53116 2828 53172
rect 2884 53116 3276 53172
rect 3332 53116 7980 53172
rect 8036 53116 8046 53172
rect 8418 53116 8428 53172
rect 8484 53116 13244 53172
rect 13300 53116 13310 53172
rect 13906 53116 13916 53172
rect 13972 53116 15596 53172
rect 15652 53116 16492 53172
rect 16548 53116 16558 53172
rect 17714 53116 17724 53172
rect 17780 53116 19852 53172
rect 19908 53116 19918 53172
rect 20066 53116 20076 53172
rect 20132 53116 24108 53172
rect 24164 53116 24780 53172
rect 24836 53116 24846 53172
rect 26114 53116 26124 53172
rect 26180 53116 26572 53172
rect 26628 53116 26638 53172
rect 26796 53116 30100 53172
rect 31798 53116 31836 53172
rect 31892 53116 31902 53172
rect 32050 53116 32060 53172
rect 32116 53116 33068 53172
rect 33124 53116 33134 53172
rect 33954 53116 33964 53172
rect 34020 53116 43204 53172
rect 43596 53116 43820 53172
rect 43876 53116 43886 53172
rect 44818 53116 44828 53172
rect 44884 53116 45164 53172
rect 45220 53116 45230 53172
rect 46162 53116 46172 53172
rect 46228 53116 57456 53172
rect 0 53088 112 53116
rect 26796 53060 26852 53116
rect 3154 53004 3164 53060
rect 3220 53004 6188 53060
rect 6244 53004 6254 53060
rect 7298 53004 7308 53060
rect 7364 53004 11788 53060
rect 11844 53004 11854 53060
rect 12124 53004 13356 53060
rect 13412 53004 13422 53060
rect 13570 53004 13580 53060
rect 13636 53004 15148 53060
rect 15204 53004 15214 53060
rect 15698 53004 15708 53060
rect 15764 53004 24892 53060
rect 24948 53004 26852 53060
rect 27346 53004 27356 53060
rect 27412 53004 28588 53060
rect 28644 53004 28654 53060
rect 12124 52948 12180 53004
rect 30044 52948 30100 53116
rect 43148 53060 43204 53116
rect 57344 53088 57456 53116
rect 33618 53004 33628 53060
rect 33684 53004 42700 53060
rect 42756 53004 42924 53060
rect 42980 53004 42990 53060
rect 43148 53004 44324 53060
rect 45042 53004 45052 53060
rect 45108 53004 45724 53060
rect 45780 53004 45790 53060
rect 45938 53004 45948 53060
rect 46004 53004 49868 53060
rect 49924 53004 49934 53060
rect 50082 53004 50092 53060
rect 50148 53004 51100 53060
rect 51156 53004 51166 53060
rect 51314 53004 51324 53060
rect 51380 53004 53788 53060
rect 53844 53004 53854 53060
rect 54226 53004 54236 53060
rect 54292 53004 57036 53060
rect 57092 53004 57102 53060
rect 44268 52948 44324 53004
rect 1922 52892 1932 52948
rect 1988 52892 2828 52948
rect 2884 52892 2940 52948
rect 2996 52892 4172 52948
rect 4228 52892 4238 52948
rect 4946 52892 4956 52948
rect 5012 52892 6524 52948
rect 6580 52892 6748 52948
rect 6804 52892 6814 52948
rect 6962 52892 6972 52948
rect 7028 52892 12180 52948
rect 12338 52892 12348 52948
rect 12404 52892 16044 52948
rect 16100 52892 16110 52948
rect 16258 52892 16268 52948
rect 16324 52892 17724 52948
rect 17780 52892 17790 52948
rect 17938 52892 17948 52948
rect 18004 52892 20188 52948
rect 20244 52892 20254 52948
rect 21634 52892 21644 52948
rect 21700 52892 22652 52948
rect 22708 52892 22718 52948
rect 23650 52892 23660 52948
rect 23716 52892 24220 52948
rect 24276 52892 24286 52948
rect 24994 52892 25004 52948
rect 25060 52892 25900 52948
rect 25956 52892 25966 52948
rect 26898 52892 26908 52948
rect 26964 52892 28252 52948
rect 28308 52892 28318 52948
rect 29362 52892 29372 52948
rect 29428 52892 29820 52948
rect 29876 52892 29886 52948
rect 30044 52892 32620 52948
rect 32676 52892 32686 52948
rect 33058 52892 33068 52948
rect 33124 52892 35868 52948
rect 35924 52892 35934 52948
rect 41794 52892 41804 52948
rect 41860 52892 43932 52948
rect 43988 52892 43998 52948
rect 44268 52892 45332 52948
rect 46498 52892 46508 52948
rect 46564 52892 51212 52948
rect 51268 52892 51278 52948
rect 52322 52892 52332 52948
rect 52388 52892 53340 52948
rect 53396 52892 53406 52948
rect 55010 52892 55020 52948
rect 55076 52892 55086 52948
rect 55234 52892 55244 52948
rect 55300 52892 55356 52948
rect 55412 52892 55422 52948
rect 56354 52892 56364 52948
rect 56420 52892 57260 52948
rect 57316 52892 57326 52948
rect 1026 52780 1036 52836
rect 1092 52780 1596 52836
rect 1652 52780 1662 52836
rect 2594 52780 2604 52836
rect 2660 52780 3276 52836
rect 3332 52780 3342 52836
rect 4162 52780 4172 52836
rect 4228 52780 5292 52836
rect 5348 52780 5358 52836
rect 6738 52780 6748 52836
rect 6804 52780 9324 52836
rect 9380 52780 9390 52836
rect 10994 52780 11004 52836
rect 11060 52780 11676 52836
rect 11732 52780 15708 52836
rect 15764 52780 15774 52836
rect 15922 52780 15932 52836
rect 15988 52780 21980 52836
rect 22036 52780 22046 52836
rect 22418 52780 22428 52836
rect 22484 52780 24668 52836
rect 24724 52780 26348 52836
rect 26404 52780 26414 52836
rect 27570 52780 27580 52836
rect 27636 52780 30940 52836
rect 30996 52780 31006 52836
rect 31154 52780 31164 52836
rect 31220 52780 35924 52836
rect 36530 52780 36540 52836
rect 36596 52780 45052 52836
rect 45108 52780 45118 52836
rect 0 52724 112 52752
rect 31164 52724 31220 52780
rect 35868 52724 35924 52780
rect 0 52668 476 52724
rect 532 52668 2940 52724
rect 2996 52668 3006 52724
rect 3378 52668 3388 52724
rect 3444 52668 4228 52724
rect 4386 52668 4396 52724
rect 4452 52668 5852 52724
rect 5908 52668 5918 52724
rect 6066 52668 6076 52724
rect 6132 52668 7084 52724
rect 7140 52668 7868 52724
rect 7924 52668 7934 52724
rect 10546 52668 10556 52724
rect 10612 52668 13580 52724
rect 13636 52668 14140 52724
rect 14196 52668 14206 52724
rect 15250 52668 15260 52724
rect 15316 52668 17948 52724
rect 18004 52668 18014 52724
rect 19282 52668 19292 52724
rect 19348 52668 19516 52724
rect 19572 52668 19628 52724
rect 19684 52668 19694 52724
rect 19842 52668 19852 52724
rect 19908 52668 20244 52724
rect 22278 52668 22316 52724
rect 22372 52668 22382 52724
rect 25330 52668 25340 52724
rect 25396 52668 27020 52724
rect 27076 52668 27086 52724
rect 28998 52668 29036 52724
rect 29092 52668 31220 52724
rect 31490 52668 31500 52724
rect 31556 52668 33068 52724
rect 33124 52668 33134 52724
rect 33404 52668 35644 52724
rect 35700 52668 35710 52724
rect 35868 52668 36876 52724
rect 36932 52668 37436 52724
rect 37492 52668 37502 52724
rect 38098 52668 38108 52724
rect 38164 52668 39004 52724
rect 39060 52668 39070 52724
rect 41766 52668 41804 52724
rect 41860 52668 41870 52724
rect 43334 52668 43372 52724
rect 43428 52668 43438 52724
rect 44268 52668 44884 52724
rect 0 52640 112 52668
rect 1474 52556 1484 52612
rect 1540 52556 3500 52612
rect 3556 52556 3566 52612
rect 3266 52444 3276 52500
rect 3332 52444 3612 52500
rect 3668 52444 3678 52500
rect 4172 52388 4228 52668
rect 20188 52612 20244 52668
rect 33404 52612 33460 52668
rect 44268 52612 44324 52668
rect 5506 52556 5516 52612
rect 5572 52556 7644 52612
rect 7700 52556 7710 52612
rect 10098 52556 10108 52612
rect 10164 52556 14364 52612
rect 14420 52556 14430 52612
rect 15138 52556 15148 52612
rect 15204 52556 15484 52612
rect 15540 52556 16380 52612
rect 16436 52556 16446 52612
rect 18162 52556 18172 52612
rect 18228 52556 18732 52612
rect 18788 52556 19404 52612
rect 19460 52556 19470 52612
rect 19730 52556 19740 52612
rect 19796 52556 19964 52612
rect 20020 52556 20030 52612
rect 20188 52556 24220 52612
rect 24276 52556 24286 52612
rect 26114 52556 26124 52612
rect 26180 52556 26908 52612
rect 26964 52556 26974 52612
rect 27346 52556 27356 52612
rect 27412 52556 33460 52612
rect 33842 52556 33852 52612
rect 33908 52556 39900 52612
rect 39956 52556 39966 52612
rect 41132 52556 44324 52612
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 41132 52500 41188 52556
rect 44454 52500 44464 52556
rect 44520 52500 44568 52556
rect 44624 52500 44672 52556
rect 44728 52500 44738 52556
rect 44828 52500 44884 52668
rect 45276 52612 45332 52892
rect 48402 52780 48412 52836
rect 48468 52780 49476 52836
rect 50978 52780 50988 52836
rect 51044 52780 54572 52836
rect 54628 52780 54638 52836
rect 49420 52724 49476 52780
rect 55020 52724 55076 52892
rect 57344 52724 57456 52752
rect 46610 52668 46620 52724
rect 46676 52668 48300 52724
rect 48356 52668 48366 52724
rect 49158 52668 49196 52724
rect 49252 52668 49262 52724
rect 49420 52668 50876 52724
rect 50932 52668 50942 52724
rect 52210 52668 52220 52724
rect 52276 52668 55076 52724
rect 56354 52668 56364 52724
rect 56420 52668 56924 52724
rect 56980 52668 56990 52724
rect 57148 52668 57456 52724
rect 57148 52612 57204 52668
rect 57344 52640 57456 52668
rect 45276 52556 48636 52612
rect 48692 52556 48702 52612
rect 48850 52556 48860 52612
rect 48916 52556 57204 52612
rect 5394 52444 5404 52500
rect 5460 52444 8428 52500
rect 8484 52444 8494 52500
rect 8642 52444 8652 52500
rect 8708 52444 23548 52500
rect 23604 52444 23614 52500
rect 25666 52444 25676 52500
rect 25732 52444 27804 52500
rect 27860 52444 27870 52500
rect 29474 52444 29484 52500
rect 29540 52444 30156 52500
rect 30212 52444 30222 52500
rect 30594 52444 30604 52500
rect 30660 52444 33068 52500
rect 33124 52444 33134 52500
rect 33282 52444 33292 52500
rect 33348 52444 34916 52500
rect 35074 52444 35084 52500
rect 35140 52444 41188 52500
rect 41346 52444 41356 52500
rect 41412 52444 44156 52500
rect 44212 52444 44222 52500
rect 44828 52444 46284 52500
rect 46340 52444 48412 52500
rect 48468 52444 48860 52500
rect 48916 52444 48926 52500
rect 50642 52444 50652 52500
rect 50708 52444 51100 52500
rect 51156 52444 51166 52500
rect 51986 52444 51996 52500
rect 52052 52444 52892 52500
rect 52948 52444 52958 52500
rect 53106 52444 53116 52500
rect 53172 52444 54348 52500
rect 54404 52444 54414 52500
rect 34860 52388 34916 52444
rect 1138 52332 1148 52388
rect 1204 52332 3500 52388
rect 3556 52332 3566 52388
rect 4172 52332 8092 52388
rect 8148 52332 8158 52388
rect 8950 52332 8988 52388
rect 9044 52332 9054 52388
rect 9314 52332 9324 52388
rect 9380 52332 12124 52388
rect 12180 52332 12190 52388
rect 13122 52332 13132 52388
rect 13188 52332 16716 52388
rect 16772 52332 16782 52388
rect 16930 52332 16940 52388
rect 16996 52332 20636 52388
rect 20692 52332 20702 52388
rect 22082 52332 22092 52388
rect 22148 52332 22764 52388
rect 22820 52332 25004 52388
rect 25060 52332 25070 52388
rect 25862 52332 25900 52388
rect 25956 52332 25966 52388
rect 26562 52332 26572 52388
rect 26628 52332 26908 52388
rect 26964 52332 26974 52388
rect 28690 52332 28700 52388
rect 28756 52332 29708 52388
rect 29764 52332 29774 52388
rect 29922 52332 29932 52388
rect 29988 52332 34636 52388
rect 34692 52332 34702 52388
rect 34860 52332 36596 52388
rect 36754 52332 36764 52388
rect 36820 52332 43036 52388
rect 43092 52332 43102 52388
rect 43586 52332 43596 52388
rect 43652 52332 48300 52388
rect 48356 52332 48366 52388
rect 48514 52332 48524 52388
rect 48580 52332 53956 52388
rect 54226 52332 54236 52388
rect 54292 52332 56028 52388
rect 56084 52332 56094 52388
rect 0 52276 112 52304
rect 36540 52276 36596 52332
rect 53900 52276 53956 52332
rect 57344 52276 57456 52304
rect 0 52220 1876 52276
rect 2034 52220 2044 52276
rect 2100 52220 2716 52276
rect 2772 52220 2782 52276
rect 2930 52220 2940 52276
rect 2996 52220 4732 52276
rect 4788 52220 4798 52276
rect 6598 52220 6636 52276
rect 6692 52220 6702 52276
rect 9090 52220 9100 52276
rect 9156 52220 10668 52276
rect 10724 52220 10734 52276
rect 11788 52220 13244 52276
rect 13300 52220 13310 52276
rect 14466 52220 14476 52276
rect 14532 52220 16828 52276
rect 16884 52220 16894 52276
rect 17042 52220 17052 52276
rect 17108 52220 18508 52276
rect 18564 52220 18574 52276
rect 18946 52220 18956 52276
rect 19012 52220 20860 52276
rect 20916 52220 20926 52276
rect 21308 52220 23660 52276
rect 23716 52220 23726 52276
rect 23874 52220 23884 52276
rect 23940 52220 25228 52276
rect 25284 52220 26292 52276
rect 0 52192 112 52220
rect 1820 52164 1876 52220
rect 11788 52164 11844 52220
rect 21308 52164 21364 52220
rect 26236 52164 26292 52220
rect 26852 52220 31500 52276
rect 31556 52220 31566 52276
rect 32610 52220 32620 52276
rect 32676 52220 33740 52276
rect 33796 52220 33806 52276
rect 34626 52220 34636 52276
rect 34692 52220 34748 52276
rect 34804 52220 34814 52276
rect 35830 52220 35868 52276
rect 35924 52220 35934 52276
rect 36540 52220 37156 52276
rect 37426 52220 37436 52276
rect 37492 52220 40348 52276
rect 40404 52220 40414 52276
rect 40562 52220 40572 52276
rect 40628 52220 40908 52276
rect 40964 52220 40974 52276
rect 41234 52220 41244 52276
rect 41300 52220 41580 52276
rect 41636 52220 41646 52276
rect 43026 52220 43036 52276
rect 43092 52220 46620 52276
rect 46676 52220 46686 52276
rect 48738 52220 48748 52276
rect 48804 52220 50988 52276
rect 51044 52220 51054 52276
rect 51202 52220 51212 52276
rect 51268 52220 51884 52276
rect 51940 52220 51950 52276
rect 53900 52220 57456 52276
rect 1820 52108 2604 52164
rect 2660 52108 2670 52164
rect 2818 52108 2828 52164
rect 2884 52108 6244 52164
rect 6738 52108 6748 52164
rect 6804 52108 7980 52164
rect 8036 52108 8046 52164
rect 8194 52108 8204 52164
rect 8260 52108 11788 52164
rect 11844 52108 11854 52164
rect 12450 52108 12460 52164
rect 12516 52108 12908 52164
rect 12964 52108 13412 52164
rect 14242 52108 14252 52164
rect 14308 52108 14924 52164
rect 14980 52108 14990 52164
rect 15138 52108 15148 52164
rect 15204 52108 15932 52164
rect 15988 52108 17276 52164
rect 17332 52108 17342 52164
rect 19142 52108 19180 52164
rect 19236 52108 19246 52164
rect 19394 52108 19404 52164
rect 19460 52108 21364 52164
rect 21494 52108 21532 52164
rect 21588 52108 21598 52164
rect 24210 52108 24220 52164
rect 24276 52108 25900 52164
rect 25956 52108 25966 52164
rect 26226 52108 26236 52164
rect 26292 52108 26302 52164
rect 6188 52052 6244 52108
rect 13356 52052 13412 52108
rect 2594 51996 2604 52052
rect 2660 51996 4172 52052
rect 4228 51996 4238 52052
rect 4386 51996 4396 52052
rect 4452 51996 5964 52052
rect 6020 51996 6030 52052
rect 6188 51996 7308 52052
rect 7364 51996 7374 52052
rect 9986 51996 9996 52052
rect 10052 51996 11116 52052
rect 11172 51996 11182 52052
rect 11666 51996 11676 52052
rect 11732 51996 12012 52052
rect 12068 51996 13020 52052
rect 13076 51996 13086 52052
rect 13356 51996 16940 52052
rect 16996 51996 17006 52052
rect 17164 51940 17220 52108
rect 26852 52052 26908 52220
rect 33740 52164 33796 52220
rect 37100 52164 37156 52220
rect 57344 52192 57456 52220
rect 28578 52108 28588 52164
rect 28644 52108 29372 52164
rect 29428 52108 29438 52164
rect 29698 52108 29708 52164
rect 29764 52108 30268 52164
rect 30324 52108 30828 52164
rect 30884 52108 30894 52164
rect 31042 52108 31052 52164
rect 31108 52108 32508 52164
rect 32564 52108 32574 52164
rect 32946 52108 32956 52164
rect 33012 52108 33180 52164
rect 33236 52108 33246 52164
rect 33740 52108 34412 52164
rect 34468 52108 34478 52164
rect 36418 52108 36428 52164
rect 36484 52108 37044 52164
rect 37100 52108 40236 52164
rect 40292 52108 40302 52164
rect 43586 52108 43596 52164
rect 43652 52108 45388 52164
rect 45444 52108 45454 52164
rect 45602 52108 45612 52164
rect 45668 52108 46732 52164
rect 46788 52108 46798 52164
rect 48066 52108 48076 52164
rect 48132 52108 49868 52164
rect 49924 52108 49934 52164
rect 50418 52108 50428 52164
rect 50484 52108 52780 52164
rect 52836 52108 52846 52164
rect 54002 52108 54012 52164
rect 54068 52108 54124 52164
rect 54180 52108 54190 52164
rect 36988 52052 37044 52108
rect 18386 51996 18396 52052
rect 18452 51996 19516 52052
rect 19572 51996 19582 52052
rect 20626 51996 20636 52052
rect 20692 51996 20972 52052
rect 21028 51996 21038 52052
rect 21410 51996 21420 52052
rect 21476 51996 26908 52052
rect 29446 51996 29484 52052
rect 29540 51996 33628 52052
rect 33684 51996 33694 52052
rect 34066 51996 34076 52052
rect 34132 51996 35420 52052
rect 35476 51996 35486 52052
rect 36988 51996 38108 52052
rect 38164 51996 38174 52052
rect 40674 51996 40684 52052
rect 40740 51996 40796 52052
rect 40852 51996 40862 52052
rect 41234 51996 41244 52052
rect 41300 51996 43260 52052
rect 43316 51996 43326 52052
rect 43474 51996 43484 52052
rect 43540 51996 45164 52052
rect 45220 51996 45230 52052
rect 46834 51996 46844 52052
rect 46900 51996 48860 52052
rect 48916 51996 48926 52052
rect 49634 51996 49644 52052
rect 49700 51996 52220 52052
rect 52276 51996 52286 52052
rect 52630 51996 52668 52052
rect 52724 51996 52734 52052
rect 53106 51996 53116 52052
rect 53172 51996 54796 52052
rect 54852 51996 54862 52052
rect 1922 51884 1932 51940
rect 1988 51884 3164 51940
rect 3220 51884 3230 51940
rect 3378 51884 3388 51940
rect 3444 51884 4284 51940
rect 4340 51884 4350 51940
rect 6626 51884 6636 51940
rect 6692 51884 9548 51940
rect 9604 51884 10108 51940
rect 10164 51884 10174 51940
rect 13234 51884 13244 51940
rect 13300 51884 14252 51940
rect 14308 51884 14318 51940
rect 17164 51884 20524 51940
rect 20580 51884 20590 51940
rect 27234 51884 27244 51940
rect 27300 51884 44212 51940
rect 44370 51884 44380 51940
rect 44436 51884 48748 51940
rect 48804 51884 48814 51940
rect 48962 51884 48972 51940
rect 49028 51884 54348 51940
rect 54404 51884 54414 51940
rect 0 51828 112 51856
rect 0 51772 1932 51828
rect 1988 51772 1998 51828
rect 2146 51772 2156 51828
rect 2212 51772 3388 51828
rect 6290 51772 6300 51828
rect 6356 51772 8876 51828
rect 8932 51772 8942 51828
rect 9762 51772 9772 51828
rect 9828 51772 14252 51828
rect 14308 51772 14318 51828
rect 14914 51772 14924 51828
rect 14980 51772 18620 51828
rect 18676 51772 18686 51828
rect 19506 51772 19516 51828
rect 19572 51772 19964 51828
rect 20020 51772 21532 51828
rect 21588 51772 21598 51828
rect 26852 51772 32172 51828
rect 32228 51772 33180 51828
rect 33236 51772 33246 51828
rect 34962 51772 34972 51828
rect 35028 51772 35196 51828
rect 35252 51772 35262 51828
rect 35634 51772 35644 51828
rect 35700 51772 36932 51828
rect 0 51744 112 51772
rect 3332 51604 3388 51772
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 4162 51660 4172 51716
rect 4228 51660 8036 51716
rect 8418 51660 8428 51716
rect 8484 51660 12516 51716
rect 12674 51660 12684 51716
rect 12740 51660 13580 51716
rect 13636 51660 13646 51716
rect 14690 51660 14700 51716
rect 14756 51660 18172 51716
rect 18228 51660 19740 51716
rect 19796 51660 23100 51716
rect 23156 51660 23166 51716
rect 26450 51660 26460 51716
rect 26516 51660 26796 51716
rect 26852 51660 26908 51772
rect 36876 51716 36932 51772
rect 43794 51716 43804 51772
rect 43860 51716 43908 51772
rect 43964 51716 44012 51772
rect 44068 51716 44078 51772
rect 44156 51716 44212 51884
rect 57344 51828 57456 51856
rect 44482 51772 44492 51828
rect 44548 51772 44940 51828
rect 44996 51772 45006 51828
rect 47506 51772 47516 51828
rect 47572 51772 57456 51828
rect 57344 51744 57456 51772
rect 29026 51660 29036 51716
rect 29092 51660 36820 51716
rect 36876 51660 39340 51716
rect 39396 51660 39406 51716
rect 44156 51660 53676 51716
rect 53732 51660 53742 51716
rect 54226 51660 54236 51716
rect 54292 51660 54684 51716
rect 54740 51660 54750 51716
rect 55122 51660 55132 51716
rect 55188 51660 55356 51716
rect 55412 51660 55422 51716
rect 7980 51604 8036 51660
rect 12460 51604 12516 51660
rect 36764 51604 36820 51660
rect 1586 51548 1596 51604
rect 1652 51548 1708 51604
rect 1764 51548 1774 51604
rect 3332 51548 6636 51604
rect 6692 51548 6702 51604
rect 6850 51548 6860 51604
rect 6916 51548 7756 51604
rect 7812 51548 7822 51604
rect 7980 51548 8764 51604
rect 8820 51548 8830 51604
rect 9538 51548 9548 51604
rect 9604 51548 10556 51604
rect 10612 51548 10622 51604
rect 12114 51548 12124 51604
rect 12180 51548 12404 51604
rect 12460 51548 21756 51604
rect 21812 51548 21822 51604
rect 22540 51548 23772 51604
rect 23828 51548 23838 51604
rect 23986 51548 23996 51604
rect 24052 51548 25004 51604
rect 25060 51548 25070 51604
rect 28690 51548 28700 51604
rect 28756 51548 36540 51604
rect 36596 51548 36606 51604
rect 36764 51548 42700 51604
rect 42756 51548 42766 51604
rect 43250 51548 43260 51604
rect 43316 51548 44604 51604
rect 44660 51548 44670 51604
rect 48290 51548 48300 51604
rect 48356 51548 49308 51604
rect 49364 51548 49374 51604
rect 49634 51548 49644 51604
rect 49700 51548 49868 51604
rect 49924 51548 49934 51604
rect 50082 51548 50092 51604
rect 50148 51548 50204 51604
rect 50260 51548 51436 51604
rect 51492 51548 51502 51604
rect 52546 51548 52556 51604
rect 52612 51548 52622 51604
rect 53554 51548 53564 51604
rect 53620 51548 55356 51604
rect 55412 51548 55422 51604
rect 56354 51548 56364 51604
rect 56420 51548 57260 51604
rect 57316 51548 57326 51604
rect 12348 51492 12404 51548
rect 1372 51436 3388 51492
rect 3444 51436 3454 51492
rect 4172 51436 7196 51492
rect 7252 51436 7262 51492
rect 7410 51436 7420 51492
rect 7476 51436 11284 51492
rect 11442 51436 11452 51492
rect 11508 51436 12124 51492
rect 12180 51436 12190 51492
rect 12348 51436 15708 51492
rect 15764 51436 15774 51492
rect 16146 51436 16156 51492
rect 16212 51436 17164 51492
rect 17220 51436 18284 51492
rect 18340 51436 18350 51492
rect 18498 51436 18508 51492
rect 18564 51436 21868 51492
rect 21924 51436 22316 51492
rect 22372 51436 22382 51492
rect 0 51380 112 51408
rect 0 51324 140 51380
rect 196 51324 1092 51380
rect 0 51296 112 51324
rect 1036 51044 1092 51324
rect 1372 51156 1428 51436
rect 4172 51380 4228 51436
rect 1250 51100 1260 51156
rect 1316 51100 1428 51156
rect 1596 51324 3612 51380
rect 3668 51324 3678 51380
rect 4162 51324 4172 51380
rect 4228 51324 4238 51380
rect 6188 51324 8260 51380
rect 8390 51324 8428 51380
rect 8484 51324 8494 51380
rect 1596 51044 1652 51324
rect 6188 51268 6244 51324
rect 8204 51268 8260 51324
rect 11228 51268 11284 51436
rect 22540 51380 22596 51548
rect 12338 51324 12348 51380
rect 12404 51324 13804 51380
rect 13860 51324 13870 51380
rect 15026 51324 15036 51380
rect 15092 51324 15484 51380
rect 15540 51324 15550 51380
rect 16034 51324 16044 51380
rect 16100 51324 20636 51380
rect 20692 51324 20702 51380
rect 21746 51324 21756 51380
rect 21812 51324 22596 51380
rect 22652 51436 27692 51492
rect 27748 51436 27758 51492
rect 28578 51436 28588 51492
rect 28644 51436 42140 51492
rect 42196 51436 42206 51492
rect 43138 51436 43148 51492
rect 43204 51436 45164 51492
rect 45220 51436 45230 51492
rect 48514 51436 48524 51492
rect 48580 51436 49868 51492
rect 49924 51436 49934 51492
rect 50092 51436 50204 51492
rect 50260 51436 50270 51492
rect 50642 51436 50652 51492
rect 50708 51436 51772 51492
rect 51828 51436 51838 51492
rect 22652 51268 22708 51436
rect 50092 51380 50148 51436
rect 23090 51324 23100 51380
rect 23156 51324 24668 51380
rect 24724 51324 24734 51380
rect 24994 51324 25004 51380
rect 25060 51324 26348 51380
rect 26404 51324 26414 51380
rect 27356 51324 30044 51380
rect 30100 51324 30110 51380
rect 30258 51324 30268 51380
rect 30324 51324 30996 51380
rect 31126 51324 31164 51380
rect 31220 51324 31230 51380
rect 32722 51324 32732 51380
rect 32788 51324 33964 51380
rect 34020 51324 36540 51380
rect 36596 51324 36764 51380
rect 36820 51324 37436 51380
rect 37492 51324 37772 51380
rect 37828 51324 37838 51380
rect 38444 51324 38892 51380
rect 38948 51324 39228 51380
rect 39284 51324 39294 51380
rect 39452 51324 40460 51380
rect 40516 51324 41916 51380
rect 41972 51324 41982 51380
rect 42466 51324 42476 51380
rect 42532 51324 44492 51380
rect 44548 51324 44558 51380
rect 44930 51324 44940 51380
rect 44996 51324 45724 51380
rect 45780 51324 45790 51380
rect 45938 51324 45948 51380
rect 46004 51324 50148 51380
rect 50306 51324 50316 51380
rect 50372 51324 51324 51380
rect 51380 51324 51390 51380
rect 51650 51324 51660 51380
rect 51716 51324 52108 51380
rect 52164 51324 52174 51380
rect 1810 51212 1820 51268
rect 1876 51212 6244 51268
rect 6402 51212 6412 51268
rect 6468 51212 7308 51268
rect 7364 51212 7374 51268
rect 8204 51212 9548 51268
rect 9604 51212 9614 51268
rect 10630 51212 10668 51268
rect 10724 51212 10734 51268
rect 11228 51212 12460 51268
rect 12516 51212 12526 51268
rect 12674 51212 12684 51268
rect 12740 51212 12796 51268
rect 12852 51212 12862 51268
rect 13570 51212 13580 51268
rect 13636 51212 15036 51268
rect 15092 51212 15102 51268
rect 16930 51212 16940 51268
rect 16996 51212 17612 51268
rect 17668 51212 17678 51268
rect 17826 51212 17836 51268
rect 17892 51212 19628 51268
rect 19684 51212 19694 51268
rect 20738 51212 20748 51268
rect 20804 51212 22708 51268
rect 24322 51212 24332 51268
rect 24388 51212 25564 51268
rect 25620 51212 25630 51268
rect 17612 51156 17668 51212
rect 27356 51156 27412 51324
rect 30940 51268 30996 51324
rect 29138 51212 29148 51268
rect 29204 51212 29820 51268
rect 29876 51212 29886 51268
rect 30940 51212 32620 51268
rect 32676 51212 32686 51268
rect 38098 51212 38108 51268
rect 38164 51212 38220 51268
rect 38276 51212 38286 51268
rect 38444 51156 38500 51324
rect 39452 51268 39508 51324
rect 52556 51268 52612 51548
rect 52770 51436 52780 51492
rect 52836 51436 54124 51492
rect 54180 51436 54190 51492
rect 54562 51436 54572 51492
rect 54628 51436 56196 51492
rect 56140 51380 56196 51436
rect 57344 51380 57456 51408
rect 54450 51324 54460 51380
rect 54516 51324 54628 51380
rect 54898 51324 54908 51380
rect 54964 51324 55916 51380
rect 55972 51324 55982 51380
rect 56140 51324 57456 51380
rect 54572 51268 54628 51324
rect 57344 51296 57456 51324
rect 39106 51212 39116 51268
rect 39172 51212 39508 51268
rect 40338 51212 40348 51268
rect 40404 51212 41132 51268
rect 41188 51212 41916 51268
rect 41972 51212 41982 51268
rect 44258 51212 44268 51268
rect 44324 51212 45276 51268
rect 45332 51212 45342 51268
rect 46610 51212 46620 51268
rect 46676 51212 51212 51268
rect 51268 51212 51278 51268
rect 51884 51212 52612 51268
rect 53004 51212 54124 51268
rect 54180 51212 54190 51268
rect 54562 51212 54572 51268
rect 54628 51212 54638 51268
rect 51884 51156 51940 51212
rect 53004 51156 53060 51212
rect 2370 51100 2380 51156
rect 2436 51100 2940 51156
rect 2996 51100 3006 51156
rect 3350 51100 3388 51156
rect 3444 51100 3454 51156
rect 5618 51100 5628 51156
rect 5684 51100 6524 51156
rect 6580 51100 6590 51156
rect 12226 51100 12236 51156
rect 12292 51100 13468 51156
rect 13524 51100 13534 51156
rect 15138 51100 15148 51156
rect 15204 51100 16828 51156
rect 16884 51100 16894 51156
rect 17612 51100 18620 51156
rect 18676 51100 22764 51156
rect 22820 51100 22830 51156
rect 23202 51100 23212 51156
rect 23268 51100 27412 51156
rect 27682 51100 27692 51156
rect 27748 51100 29484 51156
rect 29540 51100 29550 51156
rect 30034 51100 30044 51156
rect 30100 51100 31948 51156
rect 32004 51100 32014 51156
rect 32162 51100 32172 51156
rect 32228 51100 32620 51156
rect 32676 51100 32686 51156
rect 33478 51100 33516 51156
rect 33572 51100 33582 51156
rect 34850 51100 34860 51156
rect 34916 51100 35196 51156
rect 35252 51100 35262 51156
rect 35410 51100 35420 51156
rect 35476 51100 38500 51156
rect 38658 51100 38668 51156
rect 38724 51100 39228 51156
rect 39284 51100 39294 51156
rect 40086 51100 40124 51156
rect 40180 51100 40190 51156
rect 40674 51100 40684 51156
rect 40740 51100 41244 51156
rect 41300 51100 43372 51156
rect 43428 51100 43438 51156
rect 44370 51100 44380 51156
rect 44436 51100 45164 51156
rect 45220 51100 45230 51156
rect 45826 51100 45836 51156
rect 45892 51100 48076 51156
rect 48132 51100 48142 51156
rect 48738 51100 48748 51156
rect 48804 51100 49868 51156
rect 49924 51100 49934 51156
rect 50194 51100 50204 51156
rect 50260 51100 51940 51156
rect 52098 51100 52108 51156
rect 52164 51100 53004 51156
rect 53060 51100 53070 51156
rect 53666 51100 53676 51156
rect 53732 51100 54236 51156
rect 54292 51100 54302 51156
rect 56354 51100 56364 51156
rect 56420 51100 57148 51156
rect 57204 51100 57214 51156
rect 16828 51044 16884 51100
rect 1036 50988 1652 51044
rect 7046 50988 7084 51044
rect 7140 50988 7150 51044
rect 8082 50988 8092 51044
rect 8148 50988 12684 51044
rect 12740 50988 12750 51044
rect 16828 50988 19124 51044
rect 19954 50988 19964 51044
rect 20020 50988 21084 51044
rect 21140 50988 21150 51044
rect 21522 50988 21532 51044
rect 21588 50988 23100 51044
rect 23156 50988 23166 51044
rect 23426 50988 23436 51044
rect 23492 50988 23660 51044
rect 23716 50988 24108 51044
rect 24164 50988 24174 51044
rect 27794 50988 27804 51044
rect 27860 50988 28588 51044
rect 28644 50988 28654 51044
rect 29250 50988 29260 51044
rect 29316 50988 38668 51044
rect 41542 50988 41580 51044
rect 41636 50988 41646 51044
rect 43474 50988 43484 51044
rect 43540 50988 44268 51044
rect 44324 50988 44334 51044
rect 45490 50988 45500 51044
rect 45556 50988 47068 51044
rect 47124 50988 47134 51044
rect 47618 50988 47628 51044
rect 47684 50988 53452 51044
rect 53508 50988 53518 51044
rect 54114 50988 54124 51044
rect 54180 50988 54460 51044
rect 54516 50988 54526 51044
rect 54908 50988 55244 51044
rect 55300 50988 55310 51044
rect 0 50932 112 50960
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 19068 50932 19124 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 38612 50932 38668 50988
rect 44454 50932 44464 50988
rect 44520 50932 44568 50988
rect 44624 50932 44672 50988
rect 44728 50932 44738 50988
rect 54908 50932 54964 50988
rect 57344 50932 57456 50960
rect 0 50876 700 50932
rect 756 50876 766 50932
rect 2706 50876 2716 50932
rect 2772 50876 2828 50932
rect 2884 50876 2894 50932
rect 3462 50876 3500 50932
rect 3556 50876 3566 50932
rect 5180 50876 11676 50932
rect 11732 50876 11742 50932
rect 12450 50876 12460 50932
rect 12516 50876 12628 50932
rect 0 50848 112 50876
rect 5180 50820 5236 50876
rect 12572 50820 12628 50876
rect 16940 50876 17500 50932
rect 17556 50876 17566 50932
rect 17714 50876 17724 50932
rect 17780 50876 18844 50932
rect 18900 50876 18910 50932
rect 19068 50876 21756 50932
rect 21812 50876 21822 50932
rect 22754 50876 22764 50932
rect 22820 50876 23548 50932
rect 23604 50876 23614 50932
rect 23772 50876 24388 50932
rect 25890 50876 25900 50932
rect 25956 50876 27580 50932
rect 27636 50876 29372 50932
rect 29428 50876 29438 50932
rect 30370 50876 30380 50932
rect 30436 50876 33292 50932
rect 33348 50876 33358 50932
rect 36194 50876 36204 50932
rect 36260 50876 37884 50932
rect 37940 50876 37950 50932
rect 38612 50876 44268 50932
rect 44324 50876 44334 50932
rect 44930 50876 44940 50932
rect 44996 50876 47740 50932
rect 47796 50876 47806 50932
rect 48066 50876 48076 50932
rect 48132 50876 50092 50932
rect 50148 50876 50158 50932
rect 50418 50876 50428 50932
rect 50484 50876 51212 50932
rect 51268 50876 51278 50932
rect 51538 50876 51548 50932
rect 51604 50876 52444 50932
rect 52500 50876 52510 50932
rect 52658 50876 52668 50932
rect 52724 50876 54068 50932
rect 54898 50876 54908 50932
rect 54964 50876 54974 50932
rect 55346 50876 55356 50932
rect 55412 50876 57456 50932
rect 16940 50820 16996 50876
rect 23772 50820 23828 50876
rect 24332 50820 24388 50876
rect 1474 50764 1484 50820
rect 1540 50764 1550 50820
rect 1810 50764 1820 50820
rect 1876 50764 5236 50820
rect 5394 50764 5404 50820
rect 5460 50764 6300 50820
rect 6356 50764 6366 50820
rect 6962 50764 6972 50820
rect 7028 50764 8092 50820
rect 8148 50764 8158 50820
rect 9874 50764 9884 50820
rect 9940 50764 12348 50820
rect 12404 50764 12414 50820
rect 12572 50764 16996 50820
rect 17154 50764 17164 50820
rect 17220 50764 22316 50820
rect 22372 50764 23828 50820
rect 24098 50764 24108 50820
rect 24164 50764 24174 50820
rect 24332 50764 30268 50820
rect 30324 50764 30334 50820
rect 30482 50764 30492 50820
rect 30548 50764 32732 50820
rect 32788 50764 32798 50820
rect 35970 50764 35980 50820
rect 36036 50764 37212 50820
rect 37268 50764 37278 50820
rect 40226 50764 40236 50820
rect 40292 50764 42812 50820
rect 42868 50764 42878 50820
rect 43932 50764 45500 50820
rect 45556 50764 45566 50820
rect 46386 50764 46396 50820
rect 46452 50764 48860 50820
rect 48916 50764 48926 50820
rect 50166 50764 50204 50820
rect 50260 50764 50270 50820
rect 50530 50764 50540 50820
rect 50596 50764 53564 50820
rect 53620 50764 53630 50820
rect 1484 50708 1540 50764
rect 24108 50708 24164 50764
rect 43932 50708 43988 50764
rect 1484 50652 5292 50708
rect 5348 50652 5358 50708
rect 5618 50652 5628 50708
rect 5684 50652 6860 50708
rect 6916 50652 6926 50708
rect 7186 50652 7196 50708
rect 7252 50652 12012 50708
rect 12068 50652 12078 50708
rect 12338 50652 12348 50708
rect 12404 50652 13804 50708
rect 13860 50652 14588 50708
rect 14644 50652 14654 50708
rect 15026 50652 15036 50708
rect 15092 50652 16268 50708
rect 16324 50652 17836 50708
rect 17892 50652 17902 50708
rect 19282 50652 19292 50708
rect 19348 50652 21756 50708
rect 21812 50652 21822 50708
rect 24108 50652 25004 50708
rect 25060 50652 25070 50708
rect 25302 50652 25340 50708
rect 25396 50652 27468 50708
rect 27524 50652 27534 50708
rect 29810 50652 29820 50708
rect 29876 50652 30940 50708
rect 30996 50652 31006 50708
rect 31602 50652 31612 50708
rect 31668 50652 36204 50708
rect 36260 50652 36270 50708
rect 36418 50652 36428 50708
rect 36484 50652 36988 50708
rect 37044 50652 37054 50708
rect 37650 50652 37660 50708
rect 37716 50652 43932 50708
rect 43988 50652 43998 50708
rect 45042 50652 45052 50708
rect 45108 50652 47180 50708
rect 47236 50652 47246 50708
rect 47394 50652 47404 50708
rect 47460 50652 49084 50708
rect 49140 50652 49150 50708
rect 50726 50652 50764 50708
rect 50820 50652 50830 50708
rect 52210 50652 52220 50708
rect 52276 50652 53564 50708
rect 53620 50652 53630 50708
rect 54012 50596 54068 50876
rect 57344 50848 57456 50876
rect 54674 50764 54684 50820
rect 54740 50764 54796 50820
rect 54852 50764 54862 50820
rect 54982 50764 55020 50820
rect 55076 50764 55086 50820
rect 54226 50652 54236 50708
rect 54292 50652 56364 50708
rect 56420 50652 56430 50708
rect 578 50540 588 50596
rect 644 50540 1484 50596
rect 1540 50540 1550 50596
rect 7522 50540 7532 50596
rect 7588 50540 7868 50596
rect 7924 50540 7934 50596
rect 8306 50540 8316 50596
rect 8372 50540 11172 50596
rect 11330 50540 11340 50596
rect 11396 50540 12460 50596
rect 12516 50540 12526 50596
rect 14130 50540 14140 50596
rect 14196 50540 14476 50596
rect 14532 50540 14542 50596
rect 15222 50540 15260 50596
rect 15316 50540 15326 50596
rect 15698 50540 15708 50596
rect 15764 50540 17220 50596
rect 17490 50540 17500 50596
rect 17556 50540 18172 50596
rect 18228 50540 19516 50596
rect 19572 50540 19582 50596
rect 21074 50540 21084 50596
rect 21140 50540 24220 50596
rect 24276 50540 24286 50596
rect 24994 50540 25004 50596
rect 25060 50540 26124 50596
rect 26180 50540 26190 50596
rect 29250 50540 29260 50596
rect 29316 50540 30044 50596
rect 30100 50540 30110 50596
rect 30258 50540 30268 50596
rect 30324 50540 30604 50596
rect 30660 50540 30670 50596
rect 30818 50540 30828 50596
rect 30884 50540 32396 50596
rect 32452 50540 32462 50596
rect 35634 50540 35644 50596
rect 35700 50540 37436 50596
rect 37492 50540 37502 50596
rect 37874 50540 37884 50596
rect 37940 50540 38556 50596
rect 38612 50540 39116 50596
rect 39172 50540 39182 50596
rect 39554 50540 39564 50596
rect 39620 50540 40348 50596
rect 40404 50540 40414 50596
rect 41458 50540 41468 50596
rect 41524 50540 43260 50596
rect 43316 50540 43326 50596
rect 43586 50540 43596 50596
rect 43652 50540 44268 50596
rect 44324 50540 44334 50596
rect 45266 50540 45276 50596
rect 45332 50540 47516 50596
rect 47572 50540 47582 50596
rect 48486 50540 48524 50596
rect 48580 50540 48590 50596
rect 49634 50540 49644 50596
rect 49700 50540 50988 50596
rect 51044 50540 51054 50596
rect 51202 50540 51212 50596
rect 51268 50540 52332 50596
rect 52388 50540 52398 50596
rect 54012 50540 54628 50596
rect 54786 50540 54796 50596
rect 54852 50540 55020 50596
rect 55076 50540 55086 50596
rect 0 50484 112 50512
rect 11116 50484 11172 50540
rect 0 50428 1820 50484
rect 1876 50428 1886 50484
rect 2818 50428 2828 50484
rect 2884 50428 3276 50484
rect 3332 50428 3342 50484
rect 4498 50428 4508 50484
rect 4564 50428 6468 50484
rect 8754 50428 8764 50484
rect 8820 50428 10164 50484
rect 11116 50428 12348 50484
rect 12404 50428 12414 50484
rect 12674 50428 12684 50484
rect 12740 50428 16940 50484
rect 16996 50428 17006 50484
rect 0 50400 112 50428
rect 6412 50372 6468 50428
rect 1138 50316 1148 50372
rect 1204 50316 6076 50372
rect 6132 50316 6142 50372
rect 6412 50316 8764 50372
rect 8820 50316 8830 50372
rect 10108 50260 10164 50428
rect 17164 50372 17220 50540
rect 54572 50484 54628 50540
rect 57344 50484 57456 50512
rect 17826 50428 17836 50484
rect 17892 50428 22932 50484
rect 24322 50428 24332 50484
rect 24388 50428 24556 50484
rect 24612 50428 24622 50484
rect 24780 50428 25900 50484
rect 25956 50428 25966 50484
rect 26450 50428 26460 50484
rect 26516 50428 29932 50484
rect 29988 50428 29998 50484
rect 31826 50428 31836 50484
rect 31892 50428 35364 50484
rect 35858 50428 35868 50484
rect 35924 50428 36876 50484
rect 36932 50428 36942 50484
rect 37314 50428 37324 50484
rect 37380 50428 38892 50484
rect 38948 50428 38958 50484
rect 43362 50428 43372 50484
rect 43428 50428 44380 50484
rect 44436 50428 45948 50484
rect 46004 50428 46014 50484
rect 46162 50428 46172 50484
rect 46228 50428 49196 50484
rect 49252 50428 49262 50484
rect 49522 50428 49532 50484
rect 49588 50428 51996 50484
rect 52052 50428 52062 50484
rect 52742 50428 52780 50484
rect 52836 50428 52846 50484
rect 52994 50428 53004 50484
rect 53060 50428 54236 50484
rect 54292 50428 54302 50484
rect 54572 50428 57456 50484
rect 11330 50316 11340 50372
rect 11396 50316 12460 50372
rect 12516 50316 12526 50372
rect 15810 50316 15820 50372
rect 15876 50316 16492 50372
rect 16548 50316 17108 50372
rect 17164 50316 20076 50372
rect 20132 50316 20142 50372
rect 17052 50260 17108 50316
rect 22876 50260 22932 50428
rect 23492 50372 23604 50428
rect 24780 50372 24836 50428
rect 35308 50372 35364 50428
rect 57344 50400 57456 50428
rect 23090 50316 23100 50372
rect 23156 50316 24836 50372
rect 26786 50316 26796 50372
rect 26852 50316 29484 50372
rect 29540 50316 29550 50372
rect 29810 50316 29820 50372
rect 29876 50316 32508 50372
rect 32564 50316 32574 50372
rect 32722 50316 32732 50372
rect 32788 50316 33068 50372
rect 33124 50316 33964 50372
rect 34020 50316 34030 50372
rect 35308 50316 37548 50372
rect 37604 50316 37614 50372
rect 37762 50316 37772 50372
rect 37828 50316 43148 50372
rect 43204 50316 43214 50372
rect 43362 50316 43372 50372
rect 43428 50316 47852 50372
rect 47908 50316 47918 50372
rect 48076 50316 49644 50372
rect 49700 50316 49710 50372
rect 50530 50316 50540 50372
rect 50596 50316 50652 50372
rect 50708 50316 50718 50372
rect 51398 50316 51436 50372
rect 51492 50316 51502 50372
rect 52210 50316 52220 50372
rect 52276 50316 53676 50372
rect 53732 50316 53742 50372
rect 45836 50260 45892 50316
rect 48076 50260 48132 50316
rect 4722 50204 4732 50260
rect 4788 50204 6860 50260
rect 6916 50204 6926 50260
rect 7522 50204 7532 50260
rect 7588 50204 9324 50260
rect 9380 50204 9390 50260
rect 10108 50204 16828 50260
rect 16884 50204 16894 50260
rect 17042 50204 17052 50260
rect 17108 50204 17118 50260
rect 20178 50204 20188 50260
rect 20244 50204 20524 50260
rect 20580 50204 20590 50260
rect 20850 50204 20860 50260
rect 20916 50204 22652 50260
rect 22708 50204 22718 50260
rect 22876 50204 23436 50260
rect 23492 50204 23502 50260
rect 23622 50204 23660 50260
rect 23716 50204 23726 50260
rect 24780 50204 25564 50260
rect 25620 50204 25630 50260
rect 28690 50204 28700 50260
rect 28756 50204 41804 50260
rect 41860 50204 41870 50260
rect 44146 50204 44156 50260
rect 44212 50204 45164 50260
rect 45220 50204 45230 50260
rect 45826 50204 45836 50260
rect 45892 50204 45902 50260
rect 46050 50204 46060 50260
rect 46116 50204 47404 50260
rect 47460 50204 48132 50260
rect 48738 50204 48748 50260
rect 48804 50204 52556 50260
rect 52612 50204 52622 50260
rect 52882 50204 52892 50260
rect 52948 50204 54348 50260
rect 54404 50204 54414 50260
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 24780 50148 24836 50204
rect 43794 50148 43804 50204
rect 43860 50148 43908 50204
rect 43964 50148 44012 50204
rect 44068 50148 44078 50204
rect 4844 50092 6300 50148
rect 6356 50092 6366 50148
rect 6626 50092 6636 50148
rect 6692 50092 19740 50148
rect 19796 50092 19806 50148
rect 19954 50092 19964 50148
rect 20020 50092 23716 50148
rect 24210 50092 24220 50148
rect 24276 50092 24836 50148
rect 24994 50092 25004 50148
rect 25060 50092 28140 50148
rect 28196 50092 28206 50148
rect 30034 50092 30044 50148
rect 30100 50092 31276 50148
rect 31332 50092 31342 50148
rect 31602 50092 31612 50148
rect 31668 50092 31724 50148
rect 31780 50092 31790 50148
rect 32274 50092 32284 50148
rect 32340 50092 35308 50148
rect 36530 50092 36540 50148
rect 36596 50092 42924 50148
rect 42980 50092 42990 50148
rect 44482 50092 44492 50148
rect 44548 50092 45052 50148
rect 45108 50092 45118 50148
rect 45490 50092 45500 50148
rect 45556 50092 53900 50148
rect 53956 50092 53966 50148
rect 54450 50092 54460 50148
rect 54516 50092 55692 50148
rect 55748 50092 55758 50148
rect 0 50036 112 50064
rect 4844 50036 4900 50092
rect 23660 50036 23716 50092
rect 0 49980 700 50036
rect 756 49980 766 50036
rect 3042 49980 3052 50036
rect 3108 49980 4900 50036
rect 5058 49980 5068 50036
rect 5124 49980 8204 50036
rect 8260 49980 8270 50036
rect 9314 49980 9324 50036
rect 9380 49980 12012 50036
rect 12068 49980 12078 50036
rect 12226 49980 12236 50036
rect 12292 49980 15708 50036
rect 15764 49980 15774 50036
rect 16930 49980 16940 50036
rect 16996 49980 23436 50036
rect 23492 49980 23502 50036
rect 23660 49980 23996 50036
rect 24052 49980 24062 50036
rect 24210 49980 24220 50036
rect 24276 49980 28924 50036
rect 28980 49980 31388 50036
rect 31444 49980 31454 50036
rect 31612 49980 32396 50036
rect 32452 49980 32462 50036
rect 34962 49980 34972 50036
rect 35028 49980 35084 50036
rect 35140 49980 35150 50036
rect 0 49952 112 49980
rect 31612 49924 31668 49980
rect 35252 49924 35308 50092
rect 57344 50036 57456 50064
rect 36418 49980 36428 50036
rect 36484 49980 37212 50036
rect 37268 49980 37278 50036
rect 38098 49980 38108 50036
rect 38164 49980 39228 50036
rect 39284 49980 39294 50036
rect 43362 49980 43372 50036
rect 43428 49980 45612 50036
rect 45668 49980 45678 50036
rect 45836 49980 49812 50036
rect 49970 49980 49980 50036
rect 50036 49980 57456 50036
rect 45836 49924 45892 49980
rect 49756 49924 49812 49980
rect 57344 49952 57456 49980
rect 1586 49868 1596 49924
rect 1652 49868 2044 49924
rect 2100 49868 6972 49924
rect 7028 49868 7038 49924
rect 7186 49868 7196 49924
rect 7252 49868 7532 49924
rect 7588 49868 7598 49924
rect 8306 49868 8316 49924
rect 8372 49868 10892 49924
rect 10948 49868 14140 49924
rect 14196 49868 14206 49924
rect 14802 49868 14812 49924
rect 14868 49868 15036 49924
rect 15092 49868 16828 49924
rect 16884 49868 16894 49924
rect 18722 49868 18732 49924
rect 18788 49868 21084 49924
rect 21140 49868 21150 49924
rect 21308 49868 26460 49924
rect 26516 49868 26526 49924
rect 29698 49868 29708 49924
rect 29764 49868 30380 49924
rect 30436 49868 30446 49924
rect 30930 49868 30940 49924
rect 30996 49868 31668 49924
rect 32274 49868 32284 49924
rect 32340 49868 32732 49924
rect 32788 49868 32798 49924
rect 35252 49868 37324 49924
rect 37380 49868 37390 49924
rect 37538 49868 37548 49924
rect 37604 49868 44828 49924
rect 44884 49868 44894 49924
rect 45042 49868 45052 49924
rect 45108 49868 45892 49924
rect 47618 49868 47628 49924
rect 47684 49868 48412 49924
rect 48468 49868 48478 49924
rect 48850 49868 48860 49924
rect 48916 49868 49532 49924
rect 49588 49868 49598 49924
rect 49756 49868 50092 49924
rect 50148 49868 50158 49924
rect 50530 49868 50540 49924
rect 50596 49868 52108 49924
rect 52164 49868 52332 49924
rect 52388 49868 53004 49924
rect 53060 49868 53452 49924
rect 53508 49868 53518 49924
rect 21308 49812 21364 49868
rect 1922 49756 1932 49812
rect 1988 49756 2268 49812
rect 2324 49756 2334 49812
rect 4386 49756 4396 49812
rect 4452 49756 7868 49812
rect 7924 49756 7934 49812
rect 8418 49756 8428 49812
rect 8484 49756 9100 49812
rect 9156 49756 9166 49812
rect 9762 49756 9772 49812
rect 9828 49756 10220 49812
rect 10276 49756 10286 49812
rect 10658 49756 10668 49812
rect 10724 49756 11788 49812
rect 11844 49756 11854 49812
rect 12002 49756 12012 49812
rect 12068 49756 13524 49812
rect 14690 49756 14700 49812
rect 14756 49756 15484 49812
rect 15540 49756 15550 49812
rect 15698 49756 15708 49812
rect 15764 49756 15932 49812
rect 15988 49756 16940 49812
rect 16996 49756 17006 49812
rect 18834 49756 18844 49812
rect 18900 49756 19180 49812
rect 19236 49756 19246 49812
rect 20066 49756 20076 49812
rect 20132 49756 21364 49812
rect 21522 49756 21532 49812
rect 21588 49756 23660 49812
rect 23716 49756 29036 49812
rect 29092 49756 29102 49812
rect 30258 49756 30268 49812
rect 30324 49756 32956 49812
rect 33012 49756 33022 49812
rect 34402 49756 34412 49812
rect 34468 49756 35644 49812
rect 35700 49756 35710 49812
rect 37090 49756 37100 49812
rect 37156 49756 38108 49812
rect 38164 49756 38174 49812
rect 38434 49756 38444 49812
rect 38500 49756 41356 49812
rect 41412 49756 41422 49812
rect 42354 49756 42364 49812
rect 42420 49756 44716 49812
rect 44772 49756 44782 49812
rect 45266 49756 45276 49812
rect 45332 49756 46060 49812
rect 46116 49756 46126 49812
rect 46834 49756 46844 49812
rect 46900 49756 48972 49812
rect 49028 49756 49038 49812
rect 50418 49756 50428 49812
rect 50484 49756 52220 49812
rect 52276 49756 52286 49812
rect 53106 49756 53116 49812
rect 53172 49756 56252 49812
rect 56308 49756 56318 49812
rect 13468 49700 13524 49756
rect 34412 49700 34468 49756
rect 1558 49644 1596 49700
rect 1652 49644 1662 49700
rect 3490 49644 3500 49700
rect 3556 49644 4956 49700
rect 5012 49644 5022 49700
rect 6066 49644 6076 49700
rect 6132 49644 11004 49700
rect 11060 49644 12236 49700
rect 12292 49644 12302 49700
rect 13458 49644 13468 49700
rect 13524 49644 15148 49700
rect 15204 49644 15214 49700
rect 16454 49644 16492 49700
rect 16548 49644 16558 49700
rect 17042 49644 17052 49700
rect 17108 49644 19068 49700
rect 19124 49644 19740 49700
rect 19796 49644 19806 49700
rect 19954 49644 19964 49700
rect 20020 49644 25228 49700
rect 25284 49644 25294 49700
rect 29586 49644 29596 49700
rect 29652 49644 31612 49700
rect 31668 49644 31948 49700
rect 32004 49644 34468 49700
rect 34598 49644 34636 49700
rect 34692 49644 34702 49700
rect 39330 49644 39340 49700
rect 39396 49644 41804 49700
rect 41860 49644 41870 49700
rect 42102 49644 42140 49700
rect 42196 49644 42206 49700
rect 43138 49644 43148 49700
rect 43204 49644 46396 49700
rect 46452 49644 46462 49700
rect 47954 49644 47964 49700
rect 48020 49644 48524 49700
rect 48580 49644 48590 49700
rect 51174 49644 51212 49700
rect 51268 49644 51884 49700
rect 51940 49644 51950 49700
rect 52108 49644 55804 49700
rect 55860 49644 55870 49700
rect 0 49588 112 49616
rect 52108 49588 52164 49644
rect 57344 49588 57456 49616
rect 0 49532 252 49588
rect 308 49532 318 49588
rect 3154 49532 3164 49588
rect 3220 49532 3388 49588
rect 3444 49532 3454 49588
rect 4162 49532 4172 49588
rect 4228 49532 8428 49588
rect 8484 49532 8494 49588
rect 8754 49532 8764 49588
rect 8820 49532 11340 49588
rect 11396 49532 11406 49588
rect 12002 49532 12012 49588
rect 12068 49532 13580 49588
rect 13636 49532 13646 49588
rect 13804 49532 18172 49588
rect 18228 49532 18238 49588
rect 18946 49532 18956 49588
rect 19012 49532 22428 49588
rect 22484 49532 23212 49588
rect 23268 49532 23278 49588
rect 23426 49532 23436 49588
rect 23492 49532 24220 49588
rect 24276 49532 24286 49588
rect 26450 49532 26460 49588
rect 26516 49532 27860 49588
rect 28018 49532 28028 49588
rect 28084 49532 29708 49588
rect 29764 49532 29774 49588
rect 30594 49532 30604 49588
rect 30660 49532 37100 49588
rect 37156 49532 37166 49588
rect 38882 49532 38892 49588
rect 38948 49532 39676 49588
rect 39732 49532 39742 49588
rect 40450 49532 40460 49588
rect 40516 49532 52164 49588
rect 52294 49532 52332 49588
rect 52388 49532 52398 49588
rect 52546 49532 52556 49588
rect 52612 49532 53564 49588
rect 53620 49532 53630 49588
rect 56242 49532 56252 49588
rect 56308 49532 56588 49588
rect 56644 49532 56654 49588
rect 56812 49532 57456 49588
rect 0 49504 112 49532
rect 13804 49476 13860 49532
rect 2370 49420 2380 49476
rect 2436 49420 3948 49476
rect 4004 49420 4014 49476
rect 5394 49420 5404 49476
rect 5460 49420 7980 49476
rect 8036 49420 9212 49476
rect 9268 49420 13860 49476
rect 15138 49420 15148 49476
rect 15204 49420 17948 49476
rect 18004 49420 18014 49476
rect 18498 49420 18508 49476
rect 18564 49420 21420 49476
rect 21476 49420 21486 49476
rect 23538 49420 23548 49476
rect 23604 49420 24220 49476
rect 24276 49420 24286 49476
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 1586 49308 1596 49364
rect 1652 49308 2716 49364
rect 2772 49308 2940 49364
rect 2996 49308 3006 49364
rect 3602 49308 3612 49364
rect 3668 49308 4060 49364
rect 4116 49308 4126 49364
rect 6178 49308 6188 49364
rect 6244 49308 21644 49364
rect 21700 49308 21710 49364
rect 24892 49308 26684 49364
rect 26740 49308 26750 49364
rect 24892 49252 24948 49308
rect 27804 49252 27860 49532
rect 56812 49476 56868 49532
rect 57344 49504 57456 49532
rect 28242 49420 28252 49476
rect 28308 49420 37716 49476
rect 38210 49420 38220 49476
rect 38276 49420 38444 49476
rect 38500 49420 40908 49476
rect 40964 49420 40974 49476
rect 42018 49420 42028 49476
rect 42084 49420 44268 49476
rect 44324 49420 44334 49476
rect 44930 49420 44940 49476
rect 44996 49420 49084 49476
rect 49140 49420 49150 49476
rect 49858 49420 49868 49476
rect 49924 49420 50652 49476
rect 50708 49420 50718 49476
rect 51762 49420 51772 49476
rect 51828 49420 54908 49476
rect 54964 49420 54974 49476
rect 56018 49420 56028 49476
rect 56084 49420 56868 49476
rect 37660 49364 37716 49420
rect 44454 49364 44464 49420
rect 44520 49364 44568 49420
rect 44624 49364 44672 49420
rect 44728 49364 44738 49420
rect 28130 49308 28140 49364
rect 28196 49308 30940 49364
rect 30996 49308 31006 49364
rect 31378 49308 31388 49364
rect 31444 49308 32172 49364
rect 32228 49308 34076 49364
rect 34132 49308 34142 49364
rect 34290 49308 34300 49364
rect 34356 49308 37436 49364
rect 37492 49308 37502 49364
rect 37660 49308 44156 49364
rect 44212 49308 44222 49364
rect 44818 49308 44828 49364
rect 44884 49308 51548 49364
rect 51604 49308 51614 49364
rect 1138 49196 1148 49252
rect 1204 49196 2492 49252
rect 2548 49196 2558 49252
rect 2818 49196 2828 49252
rect 2884 49196 3388 49252
rect 3444 49196 5404 49252
rect 5460 49196 5470 49252
rect 6066 49196 6076 49252
rect 6132 49196 9772 49252
rect 9828 49196 9838 49252
rect 10098 49196 10108 49252
rect 10164 49196 11340 49252
rect 11396 49196 11406 49252
rect 14578 49196 14588 49252
rect 14644 49196 17164 49252
rect 17220 49196 17230 49252
rect 17938 49196 17948 49252
rect 18004 49196 18396 49252
rect 18452 49196 18462 49252
rect 19618 49196 19628 49252
rect 19684 49196 19852 49252
rect 19908 49196 19918 49252
rect 20178 49196 20188 49252
rect 20244 49196 23212 49252
rect 23268 49196 23278 49252
rect 23436 49196 24948 49252
rect 25106 49196 25116 49252
rect 25172 49196 26796 49252
rect 26852 49196 26862 49252
rect 27804 49196 30604 49252
rect 30660 49196 30670 49252
rect 30818 49196 30828 49252
rect 30884 49196 34188 49252
rect 34244 49196 34254 49252
rect 34514 49196 34524 49252
rect 34580 49196 36316 49252
rect 36372 49196 36382 49252
rect 37538 49196 37548 49252
rect 37604 49196 38332 49252
rect 38388 49196 38398 49252
rect 39666 49196 39676 49252
rect 39732 49196 40572 49252
rect 40628 49196 40638 49252
rect 41794 49196 41804 49252
rect 41860 49196 45500 49252
rect 45556 49196 45566 49252
rect 45714 49196 45724 49252
rect 45780 49196 49980 49252
rect 50036 49196 50046 49252
rect 50306 49196 50316 49252
rect 50372 49196 55188 49252
rect 55346 49196 55356 49252
rect 55412 49196 56028 49252
rect 56084 49196 56094 49252
rect 0 49140 112 49168
rect 14588 49140 14644 49196
rect 23436 49140 23492 49196
rect 55132 49140 55188 49196
rect 57344 49140 57456 49168
rect 0 49084 1596 49140
rect 1652 49084 1932 49140
rect 1988 49084 1998 49140
rect 2706 49084 2716 49140
rect 2772 49084 5068 49140
rect 5124 49084 5134 49140
rect 6710 49084 6748 49140
rect 6804 49084 6814 49140
rect 8306 49084 8316 49140
rect 8372 49084 10332 49140
rect 10388 49084 10398 49140
rect 10658 49084 10668 49140
rect 10724 49084 14644 49140
rect 15474 49084 15484 49140
rect 15540 49084 17052 49140
rect 17108 49084 17118 49140
rect 19170 49084 19180 49140
rect 19236 49084 22204 49140
rect 22260 49084 22270 49140
rect 22754 49084 22764 49140
rect 22820 49084 23436 49140
rect 23492 49084 23502 49140
rect 23650 49084 23660 49140
rect 23716 49084 25004 49140
rect 25060 49084 25070 49140
rect 26226 49084 26236 49140
rect 26292 49084 27692 49140
rect 27748 49084 27758 49140
rect 30370 49084 30380 49140
rect 30436 49084 34636 49140
rect 34692 49084 34702 49140
rect 35298 49084 35308 49140
rect 35364 49084 51996 49140
rect 52052 49084 52062 49140
rect 52322 49084 52332 49140
rect 52388 49084 53004 49140
rect 53060 49084 53070 49140
rect 55132 49084 57456 49140
rect 0 49056 112 49084
rect 57344 49056 57456 49084
rect 2230 48972 2268 49028
rect 2324 48972 2334 49028
rect 3462 48972 3500 49028
rect 3556 48972 3566 49028
rect 3938 48972 3948 49028
rect 4004 48972 5628 49028
rect 5684 48972 5694 49028
rect 8194 48972 8204 49028
rect 8260 48972 9436 49028
rect 9492 48972 9772 49028
rect 9828 48972 10556 49028
rect 10612 48972 10622 49028
rect 12450 48972 12460 49028
rect 12516 48972 15036 49028
rect 15092 48972 15102 49028
rect 16006 48972 16044 49028
rect 16100 48972 16110 49028
rect 17266 48972 17276 49028
rect 17332 48972 18844 49028
rect 18900 48972 18910 49028
rect 21858 48972 21868 49028
rect 21924 48972 25676 49028
rect 25732 48972 25742 49028
rect 25890 48972 25900 49028
rect 25956 48972 27356 49028
rect 27412 48972 27422 49028
rect 28466 48972 28476 49028
rect 28532 48972 30492 49028
rect 30548 48972 31500 49028
rect 31556 48972 31566 49028
rect 33506 48972 33516 49028
rect 33572 48972 35980 49028
rect 36036 48972 36820 49028
rect 37986 48972 37996 49028
rect 38052 48972 40348 49028
rect 40404 48972 41692 49028
rect 41748 48972 41758 49028
rect 43250 48972 43260 49028
rect 43316 48972 45052 49028
rect 45108 48972 45118 49028
rect 45378 48972 45388 49028
rect 45444 48972 45612 49028
rect 45668 48972 45678 49028
rect 46386 48972 46396 49028
rect 46452 48972 48300 49028
rect 48356 48972 48366 49028
rect 48850 48972 48860 49028
rect 48916 48972 49308 49028
rect 49364 48972 49374 49028
rect 49746 48972 49756 49028
rect 49812 48972 50540 49028
rect 50596 48972 50606 49028
rect 56018 48972 56028 49028
rect 56084 48972 56812 49028
rect 56868 48972 56878 49028
rect 36764 48916 36820 48972
rect 2482 48860 2492 48916
rect 2548 48860 4284 48916
rect 4340 48860 5012 48916
rect 5170 48860 5180 48916
rect 5236 48860 5516 48916
rect 5572 48860 5582 48916
rect 6188 48860 9100 48916
rect 9156 48860 13076 48916
rect 14914 48860 14924 48916
rect 14980 48860 17052 48916
rect 17108 48860 17118 48916
rect 19170 48860 19180 48916
rect 19236 48860 20748 48916
rect 20804 48860 20814 48916
rect 20962 48860 20972 48916
rect 21028 48860 21980 48916
rect 22036 48860 22046 48916
rect 22194 48860 22204 48916
rect 22260 48860 26796 48916
rect 26852 48860 26862 48916
rect 27570 48860 27580 48916
rect 27636 48860 29036 48916
rect 29092 48860 29102 48916
rect 31266 48860 31276 48916
rect 31332 48860 36540 48916
rect 36596 48860 36606 48916
rect 36764 48860 40908 48916
rect 40964 48860 41356 48916
rect 41412 48860 41422 48916
rect 41570 48860 41580 48916
rect 41636 48860 41674 48916
rect 43026 48860 43036 48916
rect 43092 48860 44156 48916
rect 44212 48860 44222 48916
rect 44594 48860 44604 48916
rect 44660 48860 45724 48916
rect 45780 48860 45836 48916
rect 45892 48860 45902 48916
rect 46582 48860 46620 48916
rect 46676 48860 46686 48916
rect 47058 48860 47068 48916
rect 47124 48860 48636 48916
rect 48692 48860 49868 48916
rect 49924 48860 49934 48916
rect 51090 48860 51100 48916
rect 51156 48860 53676 48916
rect 53732 48860 53742 48916
rect 4956 48804 5012 48860
rect 578 48748 588 48804
rect 644 48748 812 48804
rect 868 48748 878 48804
rect 2930 48748 2940 48804
rect 2996 48748 3164 48804
rect 3220 48748 3230 48804
rect 3612 48748 3836 48804
rect 3892 48748 3902 48804
rect 4956 48748 5348 48804
rect 5506 48748 5516 48804
rect 5572 48748 5964 48804
rect 6020 48748 6030 48804
rect 0 48692 112 48720
rect 0 48636 1036 48692
rect 1092 48636 1484 48692
rect 1540 48636 1550 48692
rect 1810 48636 1820 48692
rect 1876 48636 3388 48692
rect 3444 48636 3454 48692
rect 0 48608 112 48636
rect 3612 48580 3668 48748
rect 5292 48692 5348 48748
rect 6188 48692 6244 48860
rect 13020 48804 13076 48860
rect 8866 48748 8876 48804
rect 8932 48748 12796 48804
rect 12852 48748 12862 48804
rect 13020 48748 15764 48804
rect 15922 48748 15932 48804
rect 15988 48748 19740 48804
rect 19796 48748 19806 48804
rect 20290 48748 20300 48804
rect 20356 48748 21084 48804
rect 21140 48748 21150 48804
rect 22642 48748 22652 48804
rect 22708 48748 23772 48804
rect 23828 48748 23838 48804
rect 25442 48748 25452 48804
rect 25508 48748 27692 48804
rect 27748 48748 27758 48804
rect 29362 48748 29372 48804
rect 29428 48748 31500 48804
rect 31556 48748 31566 48804
rect 31826 48748 31836 48804
rect 31892 48748 32508 48804
rect 32564 48748 32574 48804
rect 33282 48748 33292 48804
rect 33348 48748 33964 48804
rect 34020 48748 34188 48804
rect 34244 48748 34524 48804
rect 34580 48748 34590 48804
rect 34738 48748 34748 48804
rect 34804 48748 35084 48804
rect 35140 48748 35150 48804
rect 36306 48748 36316 48804
rect 36372 48748 37996 48804
rect 38052 48748 38062 48804
rect 40236 48748 42812 48804
rect 42868 48748 43932 48804
rect 43988 48748 43998 48804
rect 44146 48748 44156 48804
rect 44212 48748 45724 48804
rect 45780 48748 45790 48804
rect 46722 48748 46732 48804
rect 46788 48748 48412 48804
rect 48468 48748 48478 48804
rect 48850 48748 48860 48804
rect 48916 48748 49420 48804
rect 49476 48748 49486 48804
rect 50372 48748 51660 48804
rect 51716 48748 51726 48804
rect 52210 48748 52220 48804
rect 52276 48748 55020 48804
rect 55076 48748 55086 48804
rect 15708 48692 15764 48748
rect 40236 48692 40292 48748
rect 50372 48692 50428 48748
rect 57344 48692 57456 48720
rect 5292 48636 6244 48692
rect 7186 48636 7196 48692
rect 7252 48636 10108 48692
rect 10164 48636 10332 48692
rect 10388 48636 10398 48692
rect 10994 48636 11004 48692
rect 11060 48636 11116 48692
rect 11172 48636 11182 48692
rect 12786 48636 12796 48692
rect 12852 48636 15484 48692
rect 15540 48636 15550 48692
rect 15708 48636 16492 48692
rect 16548 48636 16558 48692
rect 18162 48636 18172 48692
rect 18228 48636 20636 48692
rect 20692 48636 20702 48692
rect 24210 48636 24220 48692
rect 24276 48636 26572 48692
rect 26628 48636 26684 48692
rect 26740 48636 26750 48692
rect 27682 48636 27692 48692
rect 27748 48636 29708 48692
rect 29764 48636 29774 48692
rect 30706 48636 30716 48692
rect 30772 48636 33516 48692
rect 33572 48636 33582 48692
rect 34066 48636 34076 48692
rect 34132 48636 40292 48692
rect 40450 48636 40460 48692
rect 40516 48636 40796 48692
rect 40852 48636 40862 48692
rect 45042 48636 45052 48692
rect 45108 48636 50428 48692
rect 50652 48636 56588 48692
rect 56644 48636 56654 48692
rect 56812 48636 57456 48692
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 43794 48580 43804 48636
rect 43860 48580 43908 48636
rect 43964 48580 44012 48636
rect 44068 48580 44078 48636
rect 50652 48580 50708 48636
rect 56812 48580 56868 48636
rect 57344 48608 57456 48636
rect 2146 48524 2156 48580
rect 2212 48524 3668 48580
rect 4162 48524 4172 48580
rect 4228 48524 6748 48580
rect 6804 48524 6814 48580
rect 7196 48524 9884 48580
rect 9940 48524 9950 48580
rect 11218 48524 11228 48580
rect 11284 48524 11564 48580
rect 11620 48524 12964 48580
rect 14466 48524 14476 48580
rect 14532 48524 17500 48580
rect 17556 48524 17566 48580
rect 17714 48524 17724 48580
rect 17780 48524 20972 48580
rect 21028 48524 21038 48580
rect 24210 48524 24220 48580
rect 24276 48524 28364 48580
rect 28420 48524 28430 48580
rect 30594 48524 30604 48580
rect 30660 48524 31500 48580
rect 31556 48524 31566 48580
rect 33954 48524 33964 48580
rect 34020 48524 34412 48580
rect 34468 48524 34478 48580
rect 34962 48524 34972 48580
rect 35028 48524 38332 48580
rect 38388 48524 38398 48580
rect 41906 48524 41916 48580
rect 41972 48524 42812 48580
rect 42868 48524 42878 48580
rect 43026 48524 43036 48580
rect 43092 48524 43596 48580
rect 43652 48524 43662 48580
rect 44146 48524 44156 48580
rect 44212 48524 50708 48580
rect 50866 48524 50876 48580
rect 50932 48524 51772 48580
rect 51828 48524 51838 48580
rect 53330 48524 53340 48580
rect 53396 48524 56868 48580
rect 1698 48412 1708 48468
rect 1764 48412 2044 48468
rect 2100 48412 2110 48468
rect 3154 48412 3164 48468
rect 3220 48412 4508 48468
rect 4564 48412 4574 48468
rect 4946 48412 4956 48468
rect 5012 48412 5068 48468
rect 5124 48412 5134 48468
rect 5618 48412 5628 48468
rect 5684 48412 6412 48468
rect 6468 48412 6478 48468
rect 7196 48356 7252 48524
rect 7410 48412 7420 48468
rect 7476 48412 9772 48468
rect 9828 48412 12684 48468
rect 12740 48412 12750 48468
rect 12908 48356 12964 48524
rect 16034 48412 16044 48468
rect 16100 48412 18508 48468
rect 18564 48412 18574 48468
rect 19842 48412 19852 48468
rect 19908 48412 19964 48468
rect 20020 48412 20030 48468
rect 21970 48412 21980 48468
rect 22036 48412 23324 48468
rect 23380 48412 23390 48468
rect 23538 48412 23548 48468
rect 23604 48412 25340 48468
rect 25396 48412 25406 48468
rect 25554 48412 25564 48468
rect 25620 48412 30044 48468
rect 30100 48412 30110 48468
rect 32274 48412 32284 48468
rect 32340 48412 35308 48468
rect 35364 48412 35374 48468
rect 38994 48412 39004 48468
rect 39060 48412 49196 48468
rect 49252 48412 49262 48468
rect 49522 48412 49532 48468
rect 49588 48412 49980 48468
rect 50036 48412 50046 48468
rect 50530 48412 50540 48468
rect 50596 48412 51100 48468
rect 51156 48412 51166 48468
rect 52322 48412 52332 48468
rect 52388 48412 52398 48468
rect 52332 48356 52388 48412
rect 1138 48300 1148 48356
rect 1204 48300 2940 48356
rect 2996 48300 3006 48356
rect 3378 48300 3388 48356
rect 3444 48300 7252 48356
rect 7942 48300 7980 48356
rect 8036 48300 8046 48356
rect 8642 48300 8652 48356
rect 8708 48300 12348 48356
rect 12404 48300 12414 48356
rect 12908 48300 15260 48356
rect 15316 48300 15326 48356
rect 15810 48300 15820 48356
rect 15876 48300 16380 48356
rect 16436 48300 16446 48356
rect 16604 48300 21980 48356
rect 22036 48300 22046 48356
rect 22530 48300 22540 48356
rect 22596 48300 26460 48356
rect 26516 48300 26526 48356
rect 30146 48300 30156 48356
rect 30212 48300 34860 48356
rect 34916 48300 35084 48356
rect 35140 48300 35150 48356
rect 35298 48300 35308 48356
rect 35364 48300 39732 48356
rect 39890 48300 39900 48356
rect 39956 48300 48748 48356
rect 48804 48300 48814 48356
rect 49420 48300 52388 48356
rect 52444 48300 53116 48356
rect 53172 48300 53182 48356
rect 54674 48300 54684 48356
rect 54740 48300 54908 48356
rect 54964 48300 54974 48356
rect 0 48244 112 48272
rect 0 48188 364 48244
rect 420 48188 430 48244
rect 2370 48188 2380 48244
rect 2436 48188 2716 48244
rect 2772 48188 2782 48244
rect 3042 48188 3052 48244
rect 3108 48188 5292 48244
rect 5348 48188 5358 48244
rect 6514 48188 6524 48244
rect 6580 48188 10108 48244
rect 10164 48188 10174 48244
rect 10882 48188 10892 48244
rect 10948 48188 11004 48244
rect 11060 48188 11070 48244
rect 11218 48188 11228 48244
rect 11284 48188 11452 48244
rect 11508 48188 13692 48244
rect 13748 48188 13758 48244
rect 0 48160 112 48188
rect 16604 48132 16660 48300
rect 39676 48244 39732 48300
rect 49420 48244 49476 48300
rect 17266 48188 17276 48244
rect 17332 48188 17612 48244
rect 17668 48188 17678 48244
rect 20962 48188 20972 48244
rect 21028 48188 27972 48244
rect 29474 48188 29484 48244
rect 29540 48188 31388 48244
rect 31444 48188 31454 48244
rect 31602 48188 31612 48244
rect 31668 48188 35532 48244
rect 35588 48188 35598 48244
rect 39676 48188 41244 48244
rect 41300 48188 41310 48244
rect 41906 48188 41916 48244
rect 41972 48188 45276 48244
rect 45332 48188 45342 48244
rect 48290 48188 48300 48244
rect 48356 48188 49308 48244
rect 49364 48188 49476 48244
rect 50866 48188 50876 48244
rect 50932 48188 51212 48244
rect 51268 48188 51660 48244
rect 51716 48188 51726 48244
rect 1596 48076 5796 48132
rect 5954 48076 5964 48132
rect 6020 48076 16660 48132
rect 16818 48076 16828 48132
rect 16884 48076 22092 48132
rect 22148 48076 24332 48132
rect 24388 48076 24398 48132
rect 25666 48076 25676 48132
rect 25732 48076 26124 48132
rect 26180 48076 26572 48132
rect 26628 48076 26638 48132
rect 1596 48020 1652 48076
rect 5740 48020 5796 48076
rect 27916 48020 27972 48188
rect 28130 48076 28140 48132
rect 28196 48076 35308 48132
rect 35364 48076 35374 48132
rect 37202 48076 37212 48132
rect 37268 48076 39676 48132
rect 39732 48076 39742 48132
rect 41010 48076 41020 48132
rect 41076 48076 44660 48132
rect 44818 48076 44828 48132
rect 44884 48076 50316 48132
rect 50372 48076 51100 48132
rect 51156 48076 51166 48132
rect 44604 48020 44660 48076
rect 52444 48020 52500 48300
rect 57344 48244 57456 48272
rect 52658 48188 52668 48244
rect 52724 48188 52734 48244
rect 53750 48188 53788 48244
rect 53844 48188 53854 48244
rect 56242 48188 56252 48244
rect 56308 48188 57456 48244
rect 1586 47964 1596 48020
rect 1652 47964 1662 48020
rect 3154 47964 3164 48020
rect 3220 47964 5068 48020
rect 5124 47964 5134 48020
rect 5740 47964 7756 48020
rect 7812 47964 7822 48020
rect 9660 47964 10332 48020
rect 10388 47964 10398 48020
rect 10658 47964 10668 48020
rect 10724 47964 13468 48020
rect 13524 47964 13534 48020
rect 13682 47964 13692 48020
rect 13748 47964 13786 48020
rect 14242 47964 14252 48020
rect 14308 47964 16828 48020
rect 16884 47964 16894 48020
rect 19142 47964 19180 48020
rect 19236 47964 19246 48020
rect 19842 47964 19852 48020
rect 19908 47964 20076 48020
rect 20132 47964 20142 48020
rect 20300 47964 21420 48020
rect 21476 47964 24948 48020
rect 25554 47964 25564 48020
rect 25620 47964 27244 48020
rect 27300 47964 27310 48020
rect 27916 47964 30380 48020
rect 30436 47964 30446 48020
rect 31266 47964 31276 48020
rect 31332 47964 33516 48020
rect 33572 47964 33582 48020
rect 35186 47964 35196 48020
rect 35252 47964 38668 48020
rect 38724 47964 38734 48020
rect 42242 47964 42252 48020
rect 42308 47964 43484 48020
rect 43540 47964 43550 48020
rect 43698 47964 43708 48020
rect 43764 47964 43774 48020
rect 44594 47964 44604 48020
rect 44660 47964 44670 48020
rect 44930 47964 44940 48020
rect 44996 47964 52500 48020
rect 9660 47908 9716 47964
rect 20300 47908 20356 47964
rect 3378 47852 3388 47908
rect 3444 47852 4172 47908
rect 4228 47852 4238 47908
rect 4946 47852 4956 47908
rect 5012 47852 9716 47908
rect 9874 47852 9884 47908
rect 9940 47852 13468 47908
rect 13524 47852 13534 47908
rect 14018 47852 14028 47908
rect 14084 47852 14812 47908
rect 14868 47852 14878 47908
rect 15698 47852 15708 47908
rect 15764 47852 15932 47908
rect 15988 47852 15998 47908
rect 16258 47852 16268 47908
rect 16324 47852 16716 47908
rect 16772 47852 16782 47908
rect 19058 47852 19068 47908
rect 19124 47852 20356 47908
rect 0 47796 112 47824
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 24892 47796 24948 47964
rect 43708 47908 43764 47964
rect 52668 47908 52724 48188
rect 57344 48160 57456 48188
rect 53890 48076 53900 48132
rect 53956 48076 54236 48132
rect 54292 48076 54302 48132
rect 55010 48076 55020 48132
rect 55076 48076 55804 48132
rect 55860 48076 55870 48132
rect 26852 47852 30716 47908
rect 30772 47852 30782 47908
rect 30940 47852 38220 47908
rect 38276 47852 38286 47908
rect 43138 47852 43148 47908
rect 43204 47852 43372 47908
rect 43428 47852 43438 47908
rect 43586 47852 43596 47908
rect 43652 47852 43764 47908
rect 44818 47852 44828 47908
rect 44884 47852 52724 47908
rect 55906 47852 55916 47908
rect 55972 47852 57148 47908
rect 57204 47852 57214 47908
rect 26852 47796 26908 47852
rect 30940 47796 30996 47852
rect 44454 47796 44464 47852
rect 44520 47796 44568 47852
rect 44624 47796 44672 47852
rect 44728 47796 44738 47852
rect 57344 47796 57456 47824
rect 0 47740 1708 47796
rect 1764 47740 1774 47796
rect 3602 47740 3612 47796
rect 3668 47740 4284 47796
rect 4340 47740 4350 47796
rect 5730 47740 5740 47796
rect 5796 47740 5964 47796
rect 6020 47740 6030 47796
rect 6178 47740 6188 47796
rect 6244 47740 7420 47796
rect 7476 47740 11116 47796
rect 11172 47740 11182 47796
rect 11732 47740 13468 47796
rect 13524 47740 13916 47796
rect 13972 47740 13982 47796
rect 15026 47740 15036 47796
rect 15092 47740 24220 47796
rect 24276 47740 24286 47796
rect 24892 47740 26908 47796
rect 29586 47740 29596 47796
rect 29652 47740 30996 47796
rect 31052 47740 32396 47796
rect 32452 47740 32462 47796
rect 32834 47740 32844 47796
rect 32900 47740 44100 47796
rect 45042 47740 45052 47796
rect 45108 47740 47068 47796
rect 47124 47740 47134 47796
rect 49186 47740 49196 47796
rect 49252 47740 49868 47796
rect 49924 47740 49934 47796
rect 50082 47740 50092 47796
rect 50148 47740 51324 47796
rect 51380 47740 51390 47796
rect 53778 47740 53788 47796
rect 53844 47740 55020 47796
rect 55076 47740 55086 47796
rect 56018 47740 56028 47796
rect 56084 47740 56476 47796
rect 56532 47740 56542 47796
rect 57026 47740 57036 47796
rect 57092 47740 57456 47796
rect 0 47712 112 47740
rect 11732 47684 11788 47740
rect 31052 47684 31108 47740
rect 2818 47628 2828 47684
rect 2884 47628 4172 47684
rect 4228 47628 4620 47684
rect 4676 47628 4686 47684
rect 4844 47628 6076 47684
rect 6132 47628 6142 47684
rect 8978 47628 8988 47684
rect 9044 47628 9212 47684
rect 9268 47628 11228 47684
rect 11284 47628 11294 47684
rect 11442 47628 11452 47684
rect 11508 47628 11788 47684
rect 13020 47628 18060 47684
rect 18116 47628 18126 47684
rect 18386 47628 18396 47684
rect 18452 47628 22764 47684
rect 22820 47628 22830 47684
rect 23314 47628 23324 47684
rect 23380 47628 28140 47684
rect 28196 47628 28206 47684
rect 28354 47628 28364 47684
rect 28420 47628 31108 47684
rect 31378 47628 31388 47684
rect 31444 47628 32396 47684
rect 32452 47628 32462 47684
rect 34066 47628 34076 47684
rect 34132 47628 37772 47684
rect 37828 47628 37838 47684
rect 39442 47628 39452 47684
rect 39508 47628 40124 47684
rect 40180 47628 40190 47684
rect 41346 47628 41356 47684
rect 41412 47628 43596 47684
rect 43652 47628 43662 47684
rect 4844 47572 4900 47628
rect 476 47516 4900 47572
rect 5058 47516 5068 47572
rect 5124 47516 7196 47572
rect 7252 47516 7262 47572
rect 7746 47516 7756 47572
rect 7812 47516 8540 47572
rect 8596 47516 8606 47572
rect 10098 47516 10108 47572
rect 10164 47516 12684 47572
rect 12740 47516 12750 47572
rect 0 47348 112 47376
rect 476 47348 532 47516
rect 13020 47460 13076 47628
rect 13346 47516 13356 47572
rect 13412 47516 17164 47572
rect 17220 47516 17230 47572
rect 19842 47516 19852 47572
rect 19908 47516 20300 47572
rect 20356 47516 25340 47572
rect 25396 47516 25406 47572
rect 27794 47516 27804 47572
rect 27860 47516 28252 47572
rect 28308 47516 28318 47572
rect 29810 47516 29820 47572
rect 29876 47516 30380 47572
rect 30436 47516 30446 47572
rect 30706 47516 30716 47572
rect 30772 47516 31108 47572
rect 33730 47516 33740 47572
rect 33796 47516 34524 47572
rect 34580 47516 34590 47572
rect 35634 47516 35644 47572
rect 35700 47516 38444 47572
rect 38500 47516 38510 47572
rect 31052 47460 31108 47516
rect 44044 47460 44100 47740
rect 57344 47712 57456 47740
rect 44258 47628 44268 47684
rect 44324 47628 44334 47684
rect 47730 47628 47740 47684
rect 47796 47628 48076 47684
rect 48132 47628 48142 47684
rect 51538 47628 51548 47684
rect 51604 47628 52668 47684
rect 52724 47628 52734 47684
rect 52882 47628 52892 47684
rect 52948 47628 53004 47684
rect 53060 47628 53676 47684
rect 53732 47628 53742 47684
rect 55682 47628 55692 47684
rect 55748 47628 55860 47684
rect 44268 47572 44324 47628
rect 44258 47516 44268 47572
rect 44324 47516 44772 47572
rect 44716 47460 44772 47516
rect 46284 47516 46844 47572
rect 46900 47516 46910 47572
rect 49970 47516 49980 47572
rect 50036 47516 55580 47572
rect 55636 47516 55646 47572
rect 46284 47460 46340 47516
rect 55804 47460 55860 47628
rect 56354 47516 56364 47572
rect 56420 47516 57036 47572
rect 57092 47516 57102 47572
rect 3042 47404 3052 47460
rect 3108 47404 4396 47460
rect 4452 47404 4462 47460
rect 5170 47404 5180 47460
rect 5236 47404 6412 47460
rect 6468 47404 7084 47460
rect 7140 47404 7150 47460
rect 7970 47404 7980 47460
rect 8036 47404 8988 47460
rect 9044 47404 9054 47460
rect 9650 47404 9660 47460
rect 9716 47404 12012 47460
rect 12068 47404 12078 47460
rect 13010 47404 13020 47460
rect 13076 47404 13086 47460
rect 14690 47404 14700 47460
rect 14756 47404 16604 47460
rect 16660 47404 16670 47460
rect 17266 47404 17276 47460
rect 17332 47404 17836 47460
rect 17892 47404 19404 47460
rect 19460 47404 19470 47460
rect 19954 47404 19964 47460
rect 20020 47404 20636 47460
rect 20692 47404 20702 47460
rect 21858 47404 21868 47460
rect 21924 47404 25004 47460
rect 25060 47404 25070 47460
rect 26450 47404 26460 47460
rect 26516 47404 27356 47460
rect 27412 47404 27422 47460
rect 27570 47404 27580 47460
rect 27636 47404 28476 47460
rect 28532 47404 28542 47460
rect 29250 47404 29260 47460
rect 29316 47404 29484 47460
rect 29540 47404 29550 47460
rect 29698 47404 29708 47460
rect 29764 47404 30828 47460
rect 30884 47404 30894 47460
rect 31052 47404 31276 47460
rect 31332 47404 31342 47460
rect 33170 47404 33180 47460
rect 33236 47404 35252 47460
rect 36754 47404 36764 47460
rect 36820 47404 38556 47460
rect 38612 47404 38622 47460
rect 39554 47404 39564 47460
rect 39620 47404 40236 47460
rect 40292 47404 40302 47460
rect 40786 47404 40796 47460
rect 40852 47404 43596 47460
rect 43652 47404 43662 47460
rect 44044 47404 44492 47460
rect 44548 47404 44558 47460
rect 44716 47404 46340 47460
rect 46498 47404 46508 47460
rect 46564 47404 48300 47460
rect 48356 47404 48524 47460
rect 48580 47404 48590 47460
rect 48962 47404 48972 47460
rect 49028 47404 51436 47460
rect 51492 47404 51502 47460
rect 52434 47404 52444 47460
rect 52500 47404 54796 47460
rect 54852 47404 54862 47460
rect 55020 47404 55860 47460
rect 13020 47348 13076 47404
rect 27356 47348 27412 47404
rect 0 47292 532 47348
rect 3378 47292 3388 47348
rect 3444 47292 5180 47348
rect 5236 47292 12124 47348
rect 12180 47292 13076 47348
rect 13458 47292 13468 47348
rect 13524 47292 14364 47348
rect 14420 47292 15260 47348
rect 15316 47292 15326 47348
rect 16146 47292 16156 47348
rect 16212 47292 16492 47348
rect 16548 47292 16558 47348
rect 18274 47292 18284 47348
rect 18340 47292 20524 47348
rect 20580 47292 20590 47348
rect 21634 47292 21644 47348
rect 21700 47292 26684 47348
rect 26740 47292 26750 47348
rect 27356 47292 28700 47348
rect 28756 47292 28766 47348
rect 30258 47292 30268 47348
rect 30324 47292 32732 47348
rect 32788 47292 32798 47348
rect 33170 47292 33180 47348
rect 33236 47292 34860 47348
rect 34916 47292 34926 47348
rect 0 47264 112 47292
rect 35196 47236 35252 47404
rect 36306 47292 36316 47348
rect 36372 47292 36988 47348
rect 37044 47292 37054 47348
rect 37314 47292 37324 47348
rect 37380 47292 39284 47348
rect 40338 47292 40348 47348
rect 40404 47292 42924 47348
rect 42980 47292 42990 47348
rect 43148 47292 47964 47348
rect 48020 47292 48030 47348
rect 48150 47292 48188 47348
rect 48244 47292 48254 47348
rect 51426 47292 51436 47348
rect 51492 47292 53788 47348
rect 53844 47292 53854 47348
rect 39228 47236 39284 47292
rect 43148 47236 43204 47292
rect 55020 47236 55076 47404
rect 57344 47348 57456 47376
rect 3714 47180 3724 47236
rect 3780 47180 5628 47236
rect 5684 47180 5694 47236
rect 5954 47180 5964 47236
rect 6020 47180 7476 47236
rect 7746 47180 7756 47236
rect 7812 47180 7980 47236
rect 8036 47180 8046 47236
rect 9202 47180 9212 47236
rect 9268 47180 18508 47236
rect 18564 47180 18574 47236
rect 19730 47180 19740 47236
rect 19796 47180 20076 47236
rect 20132 47180 20142 47236
rect 20738 47180 20748 47236
rect 20804 47180 22316 47236
rect 22372 47180 24276 47236
rect 24434 47180 24444 47236
rect 24500 47180 29596 47236
rect 29652 47180 29662 47236
rect 30706 47180 30716 47236
rect 30772 47180 34860 47236
rect 34916 47180 34926 47236
rect 35196 47180 36708 47236
rect 38434 47180 38444 47236
rect 38500 47180 39004 47236
rect 39060 47180 39070 47236
rect 39228 47180 43204 47236
rect 43698 47180 43708 47236
rect 43764 47180 44660 47236
rect 44818 47180 44828 47236
rect 44884 47180 45164 47236
rect 45220 47180 45948 47236
rect 46004 47180 49196 47236
rect 49252 47180 49262 47236
rect 51426 47180 51436 47236
rect 51492 47180 55076 47236
rect 55468 47292 57456 47348
rect 7420 47124 7476 47180
rect 24220 47124 24276 47180
rect 36652 47124 36708 47180
rect 44604 47124 44660 47180
rect 1922 47068 1932 47124
rect 1988 47068 3052 47124
rect 3108 47068 3118 47124
rect 4162 47068 4172 47124
rect 4228 47068 4956 47124
rect 5012 47068 5022 47124
rect 5170 47068 5180 47124
rect 5236 47068 6748 47124
rect 6804 47068 6814 47124
rect 7410 47068 7420 47124
rect 7476 47068 7868 47124
rect 7924 47068 7934 47124
rect 8194 47068 8204 47124
rect 8260 47068 9884 47124
rect 9940 47068 9950 47124
rect 10322 47068 10332 47124
rect 10388 47068 13020 47124
rect 13076 47068 13086 47124
rect 13682 47068 13692 47124
rect 13748 47068 14588 47124
rect 14644 47068 14654 47124
rect 15922 47068 15932 47124
rect 15988 47068 16492 47124
rect 16548 47068 16558 47124
rect 16930 47068 16940 47124
rect 16996 47068 19068 47124
rect 19124 47068 19134 47124
rect 19394 47068 19404 47124
rect 19460 47068 21420 47124
rect 21476 47068 21486 47124
rect 21644 47068 22764 47124
rect 22820 47068 22830 47124
rect 24220 47068 26460 47124
rect 26516 47068 26526 47124
rect 26674 47068 26684 47124
rect 26740 47068 30044 47124
rect 30100 47068 30110 47124
rect 31154 47068 31164 47124
rect 31220 47068 31612 47124
rect 31668 47068 31678 47124
rect 32274 47068 32284 47124
rect 32340 47068 32844 47124
rect 32900 47068 32910 47124
rect 33058 47068 33068 47124
rect 33124 47068 36428 47124
rect 36484 47068 36494 47124
rect 36652 47068 42140 47124
rect 42196 47068 42206 47124
rect 44604 47068 49084 47124
rect 49140 47068 49150 47124
rect 49522 47068 49532 47124
rect 49588 47068 49598 47124
rect 50166 47068 50204 47124
rect 50260 47068 50270 47124
rect 50372 47068 52668 47124
rect 52724 47068 52734 47124
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 4956 47012 5012 47068
rect 21644 47012 21700 47068
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 43794 47012 43804 47068
rect 43860 47012 43908 47068
rect 43964 47012 44012 47068
rect 44068 47012 44078 47068
rect 49308 47012 49588 47068
rect 49970 47012 49980 47068
rect 50036 47012 50046 47068
rect 1922 46956 1932 47012
rect 1988 46956 3612 47012
rect 3668 46956 3678 47012
rect 4956 46956 5964 47012
rect 6020 46956 6030 47012
rect 6178 46956 6188 47012
rect 6244 46956 6748 47012
rect 6804 46956 6814 47012
rect 7522 46956 7532 47012
rect 7588 46956 9324 47012
rect 9380 46956 9390 47012
rect 10322 46956 10332 47012
rect 10388 46956 14252 47012
rect 14308 46956 14318 47012
rect 14802 46956 14812 47012
rect 14868 46956 18956 47012
rect 19012 46956 19022 47012
rect 19180 46956 21700 47012
rect 24210 46956 24220 47012
rect 24276 46956 26236 47012
rect 26292 46956 26302 47012
rect 27458 46956 27468 47012
rect 27524 46956 27636 47012
rect 28242 46956 28252 47012
rect 28308 46956 29036 47012
rect 29092 46956 29102 47012
rect 30482 46956 30492 47012
rect 30548 46956 30660 47012
rect 33394 46956 33404 47012
rect 33460 46956 34972 47012
rect 35028 46956 35038 47012
rect 35298 46956 35308 47012
rect 35364 46956 36876 47012
rect 36932 46956 36942 47012
rect 37090 46956 37100 47012
rect 37156 46956 40012 47012
rect 40068 46956 40078 47012
rect 41010 46956 41020 47012
rect 41076 46956 42252 47012
rect 42308 46956 42318 47012
rect 42690 46956 42700 47012
rect 42756 46956 43372 47012
rect 43428 46956 43438 47012
rect 44146 46956 44156 47012
rect 44212 46956 45500 47012
rect 45556 46956 45566 47012
rect 48290 46956 48300 47012
rect 48356 46956 49364 47012
rect 0 46900 112 46928
rect 19180 46900 19236 46956
rect 27580 46900 27636 46956
rect 30604 46900 30660 46956
rect 0 46844 16940 46900
rect 16996 46844 17006 46900
rect 17266 46844 17276 46900
rect 17332 46844 19236 46900
rect 20066 46844 20076 46900
rect 20132 46844 20748 46900
rect 20804 46844 20814 46900
rect 22726 46844 22764 46900
rect 22820 46844 22830 46900
rect 23314 46844 23324 46900
rect 23380 46844 26796 46900
rect 26852 46844 26862 46900
rect 27580 46844 28140 46900
rect 28196 46844 28206 46900
rect 0 46816 112 46844
rect 17276 46788 17332 46844
rect 1138 46732 1148 46788
rect 1204 46732 3388 46788
rect 3444 46732 3454 46788
rect 3602 46732 3612 46788
rect 3668 46732 5740 46788
rect 5796 46732 5806 46788
rect 5954 46732 5964 46788
rect 6020 46732 7756 46788
rect 7812 46732 7822 46788
rect 7970 46732 7980 46788
rect 8036 46732 13804 46788
rect 13860 46732 13870 46788
rect 14550 46732 14588 46788
rect 14644 46732 14654 46788
rect 14998 46732 15036 46788
rect 15092 46732 15102 46788
rect 15260 46732 17332 46788
rect 20290 46732 20300 46788
rect 20356 46732 27020 46788
rect 27076 46732 27086 46788
rect 15260 46676 15316 46732
rect 2482 46620 2492 46676
rect 2548 46620 3164 46676
rect 3220 46620 5068 46676
rect 5124 46620 5134 46676
rect 7746 46620 7756 46676
rect 7812 46620 7868 46676
rect 7924 46620 7934 46676
rect 10210 46620 10220 46676
rect 10276 46620 12908 46676
rect 12964 46620 12974 46676
rect 14242 46620 14252 46676
rect 14308 46620 15260 46676
rect 15316 46620 15326 46676
rect 15474 46620 15484 46676
rect 15540 46620 15708 46676
rect 15764 46620 15774 46676
rect 16706 46620 16716 46676
rect 16772 46620 20860 46676
rect 20916 46620 20926 46676
rect 24434 46620 24444 46676
rect 24500 46620 25116 46676
rect 25172 46620 27860 46676
rect 354 46508 364 46564
rect 420 46508 924 46564
rect 980 46508 1596 46564
rect 1652 46508 1662 46564
rect 3164 46508 3388 46564
rect 3444 46508 3454 46564
rect 3938 46508 3948 46564
rect 4004 46508 6692 46564
rect 6850 46508 6860 46564
rect 6916 46508 8652 46564
rect 8708 46508 8718 46564
rect 10546 46508 10556 46564
rect 10612 46508 12908 46564
rect 12964 46508 12974 46564
rect 13570 46508 13580 46564
rect 13636 46508 13804 46564
rect 13860 46508 13870 46564
rect 14914 46508 14924 46564
rect 14980 46508 15764 46564
rect 16034 46508 16044 46564
rect 16100 46508 20748 46564
rect 20804 46508 20814 46564
rect 21970 46508 21980 46564
rect 22036 46508 22092 46564
rect 22148 46508 22540 46564
rect 22596 46508 22606 46564
rect 23538 46508 23548 46564
rect 23604 46508 25004 46564
rect 25060 46508 25070 46564
rect 0 46452 112 46480
rect 3164 46452 3220 46508
rect 6636 46452 6692 46508
rect 15708 46452 15764 46508
rect 27804 46452 27860 46620
rect 28364 46564 28420 46900
rect 28476 46844 28486 46900
rect 30604 46844 31612 46900
rect 31668 46844 33628 46900
rect 33684 46844 33694 46900
rect 34626 46844 34636 46900
rect 34692 46844 49196 46900
rect 49252 46844 49262 46900
rect 49634 46844 49644 46900
rect 49700 46844 49738 46900
rect 49980 46788 50036 47012
rect 50306 46956 50316 47012
rect 50372 46956 50428 47068
rect 50642 46956 50652 47012
rect 50708 46956 51884 47012
rect 51940 46956 51950 47012
rect 52434 46956 52444 47012
rect 52500 46956 52892 47012
rect 52948 46956 52958 47012
rect 54982 46956 55020 47012
rect 55076 46956 55086 47012
rect 55468 46900 55524 47292
rect 57344 47264 57456 47292
rect 57344 46900 57456 46928
rect 50754 46844 50764 46900
rect 50820 46844 55524 46900
rect 55794 46844 55804 46900
rect 55860 46844 57456 46900
rect 57344 46816 57456 46844
rect 29026 46732 29036 46788
rect 29092 46732 29764 46788
rect 30146 46732 30156 46788
rect 30212 46732 31948 46788
rect 32004 46732 32014 46788
rect 32946 46732 32956 46788
rect 33012 46732 36764 46788
rect 36820 46732 36830 46788
rect 37426 46732 37436 46788
rect 37492 46732 41804 46788
rect 41860 46732 41870 46788
rect 42028 46732 42700 46788
rect 42756 46732 42766 46788
rect 43026 46732 43036 46788
rect 43092 46732 49420 46788
rect 49476 46732 49486 46788
rect 49980 46732 50316 46788
rect 50372 46732 50382 46788
rect 52994 46732 53004 46788
rect 53060 46732 56252 46788
rect 56308 46732 56318 46788
rect 29708 46676 29764 46732
rect 42028 46676 42084 46732
rect 29708 46620 30604 46676
rect 30660 46620 30670 46676
rect 30818 46620 30828 46676
rect 30884 46620 32844 46676
rect 32900 46620 32910 46676
rect 34738 46620 34748 46676
rect 34804 46620 35420 46676
rect 35476 46620 35486 46676
rect 36754 46620 36764 46676
rect 36820 46620 40404 46676
rect 41794 46620 41804 46676
rect 41860 46620 42084 46676
rect 42802 46620 42812 46676
rect 42868 46620 45444 46676
rect 46722 46620 46732 46676
rect 46788 46620 47852 46676
rect 47908 46620 47918 46676
rect 49858 46620 49868 46676
rect 49924 46620 50652 46676
rect 50708 46620 50718 46676
rect 51650 46620 51660 46676
rect 51716 46620 52444 46676
rect 52500 46620 52510 46676
rect 53078 46620 53116 46676
rect 53172 46620 53182 46676
rect 53330 46620 53340 46676
rect 53396 46620 53788 46676
rect 53844 46620 53854 46676
rect 54226 46620 54236 46676
rect 54292 46620 54796 46676
rect 54852 46620 54862 46676
rect 55234 46620 55244 46676
rect 55300 46620 56252 46676
rect 56308 46620 56318 46676
rect 28130 46508 28140 46564
rect 28196 46508 28420 46564
rect 28578 46508 28588 46564
rect 28644 46508 28812 46564
rect 28868 46508 28878 46564
rect 29138 46508 29148 46564
rect 29204 46508 40124 46564
rect 40180 46508 40190 46564
rect 40348 46452 40404 46620
rect 45388 46564 45444 46620
rect 40562 46508 40572 46564
rect 40628 46508 42756 46564
rect 43810 46508 43820 46564
rect 43876 46508 45164 46564
rect 45220 46508 45230 46564
rect 45388 46508 48972 46564
rect 49028 46508 49038 46564
rect 49196 46508 50092 46564
rect 50148 46508 50158 46564
rect 0 46396 364 46452
rect 420 46396 430 46452
rect 3154 46396 3164 46452
rect 3220 46396 3230 46452
rect 3378 46396 3388 46452
rect 3444 46396 4284 46452
rect 4340 46396 4350 46452
rect 5702 46396 5740 46452
rect 5796 46396 5806 46452
rect 6636 46396 10668 46452
rect 10724 46396 10734 46452
rect 10882 46396 10892 46452
rect 10948 46396 11004 46452
rect 11060 46396 11070 46452
rect 11778 46396 11788 46452
rect 11844 46396 12460 46452
rect 12516 46396 14588 46452
rect 14644 46396 14654 46452
rect 15708 46396 15932 46452
rect 15988 46396 16716 46452
rect 16772 46396 16782 46452
rect 17266 46396 17276 46452
rect 17332 46396 18172 46452
rect 18228 46396 18238 46452
rect 20066 46396 20076 46452
rect 20132 46396 24668 46452
rect 24724 46396 24734 46452
rect 27804 46396 28420 46452
rect 28914 46396 28924 46452
rect 28980 46396 29708 46452
rect 29764 46396 30604 46452
rect 30660 46396 30670 46452
rect 32722 46396 32732 46452
rect 32788 46396 35644 46452
rect 35700 46396 35710 46452
rect 36082 46396 36092 46452
rect 36148 46396 37548 46452
rect 37604 46396 37614 46452
rect 37762 46396 37772 46452
rect 37828 46396 38556 46452
rect 38612 46396 38622 46452
rect 38770 46396 38780 46452
rect 38836 46396 39340 46452
rect 39396 46396 39406 46452
rect 40348 46396 41132 46452
rect 41188 46396 41692 46452
rect 41748 46396 41758 46452
rect 42242 46396 42252 46452
rect 42308 46396 42476 46452
rect 42532 46396 42542 46452
rect 0 46368 112 46396
rect 28364 46340 28420 46396
rect 42700 46340 42756 46508
rect 49196 46452 49252 46508
rect 57344 46452 57456 46480
rect 42914 46396 42924 46452
rect 42980 46396 45388 46452
rect 45444 46396 45454 46452
rect 46946 46396 46956 46452
rect 47012 46396 47404 46452
rect 47460 46396 47470 46452
rect 47618 46396 47628 46452
rect 47684 46396 48300 46452
rect 48356 46396 48366 46452
rect 48524 46396 49252 46452
rect 49634 46396 49644 46452
rect 49700 46396 50204 46452
rect 50260 46396 50270 46452
rect 51426 46396 51436 46452
rect 51492 46396 53004 46452
rect 53060 46396 53676 46452
rect 53732 46396 53742 46452
rect 54898 46396 54908 46452
rect 54964 46396 54974 46452
rect 55234 46396 55244 46452
rect 55300 46396 56028 46452
rect 56084 46396 56094 46452
rect 57036 46396 57456 46452
rect 48524 46340 48580 46396
rect 54908 46340 54964 46396
rect 2034 46284 2044 46340
rect 2100 46284 4060 46340
rect 4116 46284 4126 46340
rect 5170 46284 5180 46340
rect 5236 46284 8764 46340
rect 8820 46284 8830 46340
rect 11330 46284 11340 46340
rect 11396 46284 12124 46340
rect 12180 46284 12190 46340
rect 13794 46284 13804 46340
rect 13860 46284 16828 46340
rect 16884 46284 16894 46340
rect 18274 46284 18284 46340
rect 18340 46284 23884 46340
rect 23940 46284 23950 46340
rect 24994 46284 25004 46340
rect 25060 46284 25676 46340
rect 25732 46284 25742 46340
rect 26226 46284 26236 46340
rect 26292 46284 28308 46340
rect 28364 46284 29036 46340
rect 29092 46284 29102 46340
rect 29922 46284 29932 46340
rect 29988 46284 31052 46340
rect 31108 46284 31118 46340
rect 31378 46284 31388 46340
rect 31444 46284 36764 46340
rect 36820 46284 36830 46340
rect 36978 46284 36988 46340
rect 37044 46284 37996 46340
rect 38052 46284 40348 46340
rect 40404 46284 40414 46340
rect 41570 46284 41580 46340
rect 41636 46284 41692 46340
rect 41748 46284 41758 46340
rect 42700 46284 44156 46340
rect 44212 46284 44222 46340
rect 47170 46284 47180 46340
rect 47236 46284 48580 46340
rect 48738 46284 48748 46340
rect 48804 46284 49868 46340
rect 49924 46284 49934 46340
rect 50082 46284 50092 46340
rect 50148 46284 50764 46340
rect 50820 46284 50830 46340
rect 51202 46284 51212 46340
rect 51268 46284 54964 46340
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 12124 46228 12180 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 28252 46228 28308 46284
rect 44454 46228 44464 46284
rect 44520 46228 44568 46284
rect 44624 46228 44672 46284
rect 44728 46228 44738 46284
rect 57036 46228 57092 46396
rect 57344 46368 57456 46396
rect 3042 46172 3052 46228
rect 3108 46172 3836 46228
rect 3892 46172 3902 46228
rect 12124 46172 17500 46228
rect 17556 46172 19404 46228
rect 19460 46172 19470 46228
rect 19628 46172 23660 46228
rect 23716 46172 23726 46228
rect 25330 46172 25340 46228
rect 25396 46172 28028 46228
rect 28084 46172 28094 46228
rect 28252 46172 34860 46228
rect 34916 46172 34926 46228
rect 35308 46172 36652 46228
rect 36708 46172 37436 46228
rect 37492 46172 37502 46228
rect 39228 46172 43372 46228
rect 43428 46172 43438 46228
rect 49074 46172 49084 46228
rect 49140 46172 51436 46228
rect 51492 46172 51502 46228
rect 51874 46172 51884 46228
rect 51940 46172 53564 46228
rect 53620 46172 53630 46228
rect 53778 46172 53788 46228
rect 53844 46172 57092 46228
rect 19628 46116 19684 46172
rect 35308 46116 35364 46172
rect 39228 46116 39284 46172
rect 1362 46060 1372 46116
rect 1428 46060 9212 46116
rect 9268 46060 9278 46116
rect 9986 46060 9996 46116
rect 10052 46060 12236 46116
rect 12292 46060 12302 46116
rect 12898 46060 12908 46116
rect 12964 46060 14252 46116
rect 14308 46060 14812 46116
rect 14868 46060 14878 46116
rect 15372 46060 16940 46116
rect 16996 46060 17006 46116
rect 17938 46060 17948 46116
rect 18004 46060 18508 46116
rect 18564 46060 18574 46116
rect 18946 46060 18956 46116
rect 19012 46060 19684 46116
rect 19954 46060 19964 46116
rect 20020 46060 21756 46116
rect 21812 46060 21822 46116
rect 21970 46060 21980 46116
rect 22036 46060 23212 46116
rect 23268 46060 26348 46116
rect 26404 46060 26414 46116
rect 27458 46060 27468 46116
rect 27524 46060 27692 46116
rect 27748 46060 27758 46116
rect 27906 46060 27916 46116
rect 27972 46060 28924 46116
rect 28980 46060 28990 46116
rect 30818 46060 30828 46116
rect 30884 46060 30894 46116
rect 31266 46060 31276 46116
rect 31332 46060 32620 46116
rect 32676 46060 32686 46116
rect 32834 46060 32844 46116
rect 32900 46060 34636 46116
rect 34692 46060 35364 46116
rect 35522 46060 35532 46116
rect 35588 46060 35980 46116
rect 36036 46060 36046 46116
rect 38994 46060 39004 46116
rect 39060 46060 39228 46116
rect 39284 46060 39294 46116
rect 41234 46060 41244 46116
rect 41300 46060 55804 46116
rect 55860 46060 55870 46116
rect 0 46004 112 46032
rect 0 45948 1148 46004
rect 1204 45948 1214 46004
rect 2006 45948 2044 46004
rect 2100 45948 2110 46004
rect 3490 45948 3500 46004
rect 3556 45948 4060 46004
rect 4116 45948 4126 46004
rect 5618 45948 5628 46004
rect 5684 45948 6076 46004
rect 6132 45948 6142 46004
rect 7410 45948 7420 46004
rect 7476 45948 14924 46004
rect 14980 45948 14990 46004
rect 0 45920 112 45948
rect 15372 45892 15428 46060
rect 30828 46004 30884 46060
rect 57344 46004 57456 46032
rect 17052 45948 21196 46004
rect 21252 45948 21262 46004
rect 21522 45948 21532 46004
rect 21588 45948 28364 46004
rect 28420 45948 28430 46004
rect 28578 45948 28588 46004
rect 28644 45948 30884 46004
rect 32050 45948 32060 46004
rect 32116 45948 35084 46004
rect 35140 45948 35150 46004
rect 35298 45948 35308 46004
rect 35364 45948 35532 46004
rect 35588 45948 35598 46004
rect 35858 45948 35868 46004
rect 35924 45948 37772 46004
rect 37828 45948 37838 46004
rect 41794 45948 41804 46004
rect 41860 45948 42476 46004
rect 42532 45948 42542 46004
rect 43362 45948 43372 46004
rect 43428 45948 45612 46004
rect 45668 45948 47404 46004
rect 47460 45948 47470 46004
rect 49046 45948 49084 46004
rect 49140 45948 49532 46004
rect 49588 45948 49598 46004
rect 49858 45948 49868 46004
rect 49924 45948 50540 46004
rect 50596 45948 50606 46004
rect 53106 45948 53116 46004
rect 53172 45948 54908 46004
rect 54964 45948 54974 46004
rect 55356 45948 57456 46004
rect 17052 45892 17108 45948
rect 55356 45892 55412 45948
rect 57344 45920 57456 45948
rect 2818 45836 2828 45892
rect 2884 45836 3388 45892
rect 3444 45836 3454 45892
rect 3612 45836 9212 45892
rect 9268 45836 9278 45892
rect 9762 45836 9772 45892
rect 9828 45836 9884 45892
rect 9940 45836 11004 45892
rect 11060 45836 11070 45892
rect 11778 45836 11788 45892
rect 11844 45836 12460 45892
rect 12516 45836 12526 45892
rect 13122 45836 13132 45892
rect 13188 45836 14028 45892
rect 14084 45836 15428 45892
rect 15708 45836 17052 45892
rect 17108 45836 17118 45892
rect 19730 45836 19740 45892
rect 19796 45836 22092 45892
rect 22148 45836 22158 45892
rect 22754 45836 22764 45892
rect 22820 45836 23100 45892
rect 23156 45836 23166 45892
rect 23874 45836 23884 45892
rect 23940 45836 24892 45892
rect 24948 45836 24958 45892
rect 27458 45836 27468 45892
rect 27524 45836 28364 45892
rect 28420 45836 28430 45892
rect 29026 45836 29036 45892
rect 29092 45836 30492 45892
rect 30548 45836 30558 45892
rect 30790 45836 30828 45892
rect 30884 45836 30894 45892
rect 31378 45836 31388 45892
rect 31444 45836 32396 45892
rect 32452 45836 32462 45892
rect 33618 45836 33628 45892
rect 33684 45836 37660 45892
rect 37716 45836 38668 45892
rect 39526 45836 39564 45892
rect 39620 45836 39630 45892
rect 39778 45836 39788 45892
rect 39844 45836 41692 45892
rect 41748 45836 41758 45892
rect 41906 45836 41916 45892
rect 41972 45836 45052 45892
rect 45108 45836 45118 45892
rect 46274 45836 46284 45892
rect 46340 45836 48412 45892
rect 48468 45836 48478 45892
rect 49186 45836 49196 45892
rect 49252 45836 49980 45892
rect 50036 45836 50046 45892
rect 50306 45836 50316 45892
rect 50372 45836 50764 45892
rect 50820 45836 50830 45892
rect 50978 45836 50988 45892
rect 51044 45836 51660 45892
rect 51716 45836 51726 45892
rect 51874 45836 51884 45892
rect 51940 45836 55412 45892
rect 3612 45780 3668 45836
rect 2706 45724 2716 45780
rect 2772 45724 3668 45780
rect 3724 45724 15484 45780
rect 15540 45724 15550 45780
rect 3724 45668 3780 45724
rect 15708 45668 15764 45836
rect 38612 45780 38668 45836
rect 16930 45724 16940 45780
rect 16996 45724 18172 45780
rect 18228 45724 18238 45780
rect 20514 45724 20524 45780
rect 20580 45724 25340 45780
rect 25396 45724 25406 45780
rect 25554 45724 25564 45780
rect 25620 45724 32788 45780
rect 33282 45724 33292 45780
rect 33348 45724 34076 45780
rect 34132 45724 36316 45780
rect 36372 45724 37436 45780
rect 37492 45724 38220 45780
rect 38276 45724 38286 45780
rect 38612 45724 43820 45780
rect 43876 45724 43886 45780
rect 47282 45724 47292 45780
rect 47348 45724 48300 45780
rect 48356 45724 48366 45780
rect 50082 45724 50092 45780
rect 50148 45724 51996 45780
rect 52052 45724 52062 45780
rect 53218 45724 53228 45780
rect 53284 45724 54684 45780
rect 54740 45724 54750 45780
rect 54898 45724 54908 45780
rect 54964 45724 55132 45780
rect 55188 45724 55198 45780
rect 32732 45668 32788 45724
rect 3266 45612 3276 45668
rect 3332 45612 3388 45668
rect 3444 45612 3454 45668
rect 3612 45612 3780 45668
rect 3938 45612 3948 45668
rect 4004 45612 7532 45668
rect 7588 45612 7598 45668
rect 8950 45612 8988 45668
rect 9044 45612 9054 45668
rect 9874 45612 9884 45668
rect 9940 45612 10668 45668
rect 10724 45612 10734 45668
rect 11442 45612 11452 45668
rect 11508 45612 13132 45668
rect 13188 45612 15764 45668
rect 15820 45612 19068 45668
rect 19124 45612 19134 45668
rect 19292 45612 20580 45668
rect 21186 45612 21196 45668
rect 21252 45612 21644 45668
rect 21700 45612 21710 45668
rect 21970 45612 21980 45668
rect 22036 45612 22764 45668
rect 22820 45612 29820 45668
rect 29876 45612 29886 45668
rect 30146 45612 30156 45668
rect 30212 45612 30604 45668
rect 30660 45612 31612 45668
rect 31668 45612 31678 45668
rect 31826 45612 31836 45668
rect 31892 45612 32508 45668
rect 32564 45612 32574 45668
rect 32732 45612 44324 45668
rect 44930 45612 44940 45668
rect 44996 45612 46732 45668
rect 46788 45612 46798 45668
rect 48850 45612 48860 45668
rect 48916 45612 50204 45668
rect 50260 45612 50270 45668
rect 50418 45612 50428 45668
rect 50484 45612 51884 45668
rect 51940 45612 51950 45668
rect 53078 45612 53116 45668
rect 53172 45612 53182 45668
rect 53564 45612 53788 45668
rect 53844 45612 53854 45668
rect 54002 45612 54012 45668
rect 54068 45612 55356 45668
rect 55412 45612 55422 45668
rect 0 45556 112 45584
rect 3612 45556 3668 45612
rect 15820 45556 15876 45612
rect 19292 45556 19348 45612
rect 0 45500 3668 45556
rect 4946 45500 4956 45556
rect 5012 45500 5068 45556
rect 5124 45500 5134 45556
rect 5282 45500 5292 45556
rect 5348 45500 6524 45556
rect 6580 45500 6972 45556
rect 7028 45500 7532 45556
rect 7588 45500 7598 45556
rect 8194 45500 8204 45556
rect 8260 45500 10892 45556
rect 10948 45500 10958 45556
rect 11106 45500 11116 45556
rect 11172 45500 15876 45556
rect 15932 45500 19348 45556
rect 20524 45556 20580 45612
rect 44268 45556 44324 45612
rect 20524 45500 23660 45556
rect 23716 45500 23726 45556
rect 25218 45500 25228 45556
rect 25284 45500 33964 45556
rect 34020 45500 34030 45556
rect 35634 45500 35644 45556
rect 35700 45500 37324 45556
rect 37380 45500 37390 45556
rect 39666 45500 39676 45556
rect 39732 45500 39788 45556
rect 39844 45500 39854 45556
rect 40674 45500 40684 45556
rect 40740 45500 43428 45556
rect 44268 45500 48748 45556
rect 48804 45500 48814 45556
rect 49522 45500 49532 45556
rect 49588 45500 49756 45556
rect 49812 45500 49822 45556
rect 0 45472 112 45500
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 15932 45444 15988 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 43372 45444 43428 45500
rect 43794 45444 43804 45500
rect 43860 45444 43908 45500
rect 43964 45444 44012 45500
rect 44068 45444 44078 45500
rect 2258 45388 2268 45444
rect 2324 45388 2716 45444
rect 2772 45388 2782 45444
rect 3154 45388 3164 45444
rect 3220 45388 3556 45444
rect 4162 45388 4172 45444
rect 4228 45388 5180 45444
rect 5236 45388 5246 45444
rect 6626 45388 6636 45444
rect 6692 45388 7420 45444
rect 7476 45388 7486 45444
rect 9202 45388 9212 45444
rect 9268 45388 15988 45444
rect 16146 45388 16156 45444
rect 16212 45388 16940 45444
rect 16996 45388 17006 45444
rect 17490 45388 17500 45444
rect 17556 45388 22652 45444
rect 22708 45388 22718 45444
rect 23492 45388 23716 45444
rect 24322 45388 24332 45444
rect 24388 45388 25452 45444
rect 25508 45388 25518 45444
rect 27906 45388 27916 45444
rect 27972 45388 30044 45444
rect 30100 45388 30110 45444
rect 30706 45388 30716 45444
rect 30772 45388 31332 45444
rect 31938 45388 31948 45444
rect 32004 45388 33740 45444
rect 33796 45388 33852 45444
rect 33908 45388 33918 45444
rect 34850 45388 34860 45444
rect 34916 45388 35532 45444
rect 35588 45388 35598 45444
rect 36530 45388 36540 45444
rect 36596 45388 38668 45444
rect 39330 45388 39340 45444
rect 39396 45388 42252 45444
rect 42308 45388 42318 45444
rect 43362 45388 43372 45444
rect 43428 45388 43652 45444
rect 44818 45388 44828 45444
rect 44884 45388 45612 45444
rect 45668 45388 45678 45444
rect 46722 45388 46732 45444
rect 46788 45388 47740 45444
rect 47796 45388 47806 45444
rect 49634 45388 49644 45444
rect 49700 45388 51324 45444
rect 51380 45388 51390 45444
rect 51986 45388 51996 45444
rect 52052 45388 52780 45444
rect 52836 45388 52846 45444
rect 3500 45332 3556 45388
rect 23492 45332 23548 45388
rect 2594 45276 2604 45332
rect 2660 45276 3388 45332
rect 3490 45276 3500 45332
rect 3556 45276 3566 45332
rect 4274 45276 4284 45332
rect 4340 45276 4396 45332
rect 4452 45276 4462 45332
rect 4610 45276 4620 45332
rect 4676 45276 5628 45332
rect 5684 45276 5694 45332
rect 6178 45276 6188 45332
rect 6244 45276 6300 45332
rect 6356 45276 6366 45332
rect 8754 45276 8764 45332
rect 8820 45276 9996 45332
rect 10052 45276 10062 45332
rect 10210 45276 10220 45332
rect 10276 45276 14028 45332
rect 14084 45276 23548 45332
rect 23660 45332 23716 45388
rect 31276 45332 31332 45388
rect 38612 45332 38668 45388
rect 43596 45332 43652 45388
rect 53564 45332 53620 45612
rect 57344 45556 57456 45584
rect 53778 45500 53788 45556
rect 53844 45500 57456 45556
rect 57344 45472 57456 45500
rect 54226 45388 54236 45444
rect 54292 45388 55356 45444
rect 55412 45388 55422 45444
rect 56140 45388 56252 45444
rect 56308 45388 56318 45444
rect 56140 45332 56196 45388
rect 23660 45276 28532 45332
rect 28690 45276 28700 45332
rect 28756 45276 29036 45332
rect 29092 45276 29102 45332
rect 30930 45276 30940 45332
rect 30996 45276 31052 45332
rect 31108 45276 31118 45332
rect 31276 45276 38220 45332
rect 38276 45276 38286 45332
rect 38612 45276 38780 45332
rect 38836 45276 38846 45332
rect 39890 45276 39900 45332
rect 39956 45276 41020 45332
rect 41076 45276 41086 45332
rect 42578 45276 42588 45332
rect 42644 45276 43036 45332
rect 43092 45276 43102 45332
rect 43596 45276 44380 45332
rect 44436 45276 45164 45332
rect 45220 45276 45230 45332
rect 45938 45276 45948 45332
rect 46004 45276 47180 45332
rect 47236 45276 47246 45332
rect 47618 45276 47628 45332
rect 47684 45276 50428 45332
rect 50484 45276 50494 45332
rect 53106 45276 53116 45332
rect 53172 45276 53620 45332
rect 54114 45276 54124 45332
rect 54180 45276 54796 45332
rect 54852 45276 54862 45332
rect 55794 45276 55804 45332
rect 55860 45276 56140 45332
rect 56196 45276 56206 45332
rect 56354 45276 56364 45332
rect 56420 45276 57260 45332
rect 57316 45276 57326 45332
rect 3332 45220 3388 45276
rect 28476 45220 28532 45276
rect 3332 45164 3612 45220
rect 3668 45164 3678 45220
rect 4162 45164 4172 45220
rect 4228 45164 4844 45220
rect 4900 45164 5292 45220
rect 5348 45164 5358 45220
rect 6178 45164 6188 45220
rect 6244 45164 8316 45220
rect 8372 45164 11676 45220
rect 11732 45164 11742 45220
rect 11890 45164 11900 45220
rect 11956 45164 13916 45220
rect 13972 45164 13982 45220
rect 14466 45164 14476 45220
rect 14532 45164 14700 45220
rect 14756 45164 14766 45220
rect 17602 45164 17612 45220
rect 17668 45164 21980 45220
rect 22036 45164 22046 45220
rect 22530 45164 22540 45220
rect 22596 45164 23548 45220
rect 23604 45164 23614 45220
rect 23762 45164 23772 45220
rect 23828 45164 25452 45220
rect 25508 45164 25518 45220
rect 28476 45164 34188 45220
rect 34244 45164 34254 45220
rect 34412 45164 38668 45220
rect 38724 45164 38734 45220
rect 38882 45164 38892 45220
rect 38948 45164 39564 45220
rect 39620 45164 39630 45220
rect 40002 45164 40012 45220
rect 40068 45164 46508 45220
rect 46564 45164 46574 45220
rect 48626 45164 48636 45220
rect 48692 45164 56028 45220
rect 56084 45164 56094 45220
rect 56438 45164 56476 45220
rect 56532 45164 56542 45220
rect 0 45108 112 45136
rect 34412 45108 34468 45164
rect 57344 45108 57456 45136
rect 0 45052 2268 45108
rect 2324 45052 2334 45108
rect 3266 45052 3276 45108
rect 3332 45052 3388 45108
rect 3444 45052 3948 45108
rect 4004 45052 6188 45108
rect 6244 45052 6254 45108
rect 7746 45052 7756 45108
rect 7812 45052 8092 45108
rect 8148 45052 8158 45108
rect 8642 45052 8652 45108
rect 8708 45052 13244 45108
rect 13300 45052 13310 45108
rect 14690 45052 14700 45108
rect 14756 45052 14812 45108
rect 14868 45052 14878 45108
rect 16006 45052 16044 45108
rect 16100 45052 21196 45108
rect 21252 45052 21262 45108
rect 21634 45052 21644 45108
rect 21700 45052 24668 45108
rect 24724 45052 24734 45108
rect 27010 45052 27020 45108
rect 27076 45052 27636 45108
rect 28690 45052 28700 45108
rect 28756 45052 30156 45108
rect 30212 45052 30222 45108
rect 30370 45052 30380 45108
rect 30436 45052 30940 45108
rect 30996 45052 33180 45108
rect 33236 45052 33246 45108
rect 33618 45052 33628 45108
rect 33684 45052 34468 45108
rect 37202 45052 37212 45108
rect 37268 45052 39788 45108
rect 39844 45052 39854 45108
rect 40114 45052 40124 45108
rect 40180 45052 41356 45108
rect 41412 45052 41422 45108
rect 41794 45052 41804 45108
rect 41860 45052 41916 45108
rect 41972 45052 41982 45108
rect 42214 45052 42252 45108
rect 42308 45052 42318 45108
rect 42914 45052 42924 45108
rect 42980 45052 43372 45108
rect 43428 45052 46396 45108
rect 46452 45052 46462 45108
rect 46620 45052 57456 45108
rect 0 45024 112 45052
rect 27580 44996 27636 45052
rect 46620 44996 46676 45052
rect 57344 45024 57456 45052
rect 1026 44940 1036 44996
rect 1092 44940 1260 44996
rect 1316 44940 1326 44996
rect 1810 44940 1820 44996
rect 1876 44940 2604 44996
rect 2660 44940 3164 44996
rect 3220 44940 3230 44996
rect 3378 44940 3388 44996
rect 3444 44940 4956 44996
rect 5012 44940 5022 44996
rect 5618 44940 5628 44996
rect 5684 44940 9716 44996
rect 9874 44940 9884 44996
rect 9940 44940 11564 44996
rect 11620 44940 11630 44996
rect 12114 44940 12124 44996
rect 12180 44940 14252 44996
rect 14308 44940 14318 44996
rect 16258 44940 16268 44996
rect 16324 44940 18620 44996
rect 18676 44940 20916 44996
rect 22502 44940 22540 44996
rect 22596 44940 22606 44996
rect 23492 44940 23940 44996
rect 24434 44940 24444 44996
rect 24500 44940 27356 44996
rect 27412 44940 27422 44996
rect 27580 44940 30156 44996
rect 30212 44940 30222 44996
rect 32050 44940 32060 44996
rect 32116 44940 37884 44996
rect 37940 44940 39844 44996
rect 40002 44940 40012 44996
rect 40068 44940 46676 44996
rect 46732 44940 48524 44996
rect 48580 44940 48590 44996
rect 49186 44940 49196 44996
rect 49252 44940 50316 44996
rect 50372 44940 50382 44996
rect 50866 44940 50876 44996
rect 50932 44940 51436 44996
rect 51492 44940 51502 44996
rect 53340 44940 55412 44996
rect 3042 44828 3052 44884
rect 3108 44828 3500 44884
rect 3556 44828 3566 44884
rect 4834 44828 4844 44884
rect 4900 44828 5068 44884
rect 5124 44828 5134 44884
rect 9660 44772 9716 44940
rect 20860 44884 20916 44940
rect 23492 44884 23548 44940
rect 10322 44828 10332 44884
rect 10388 44828 10780 44884
rect 10836 44828 10846 44884
rect 12348 44828 15036 44884
rect 15092 44828 15102 44884
rect 16828 44828 20636 44884
rect 20692 44828 20702 44884
rect 20860 44828 22204 44884
rect 22260 44828 23548 44884
rect 23884 44884 23940 44940
rect 39788 44884 39844 44940
rect 46732 44884 46788 44940
rect 23884 44828 25060 44884
rect 25218 44828 25228 44884
rect 25284 44828 29596 44884
rect 29652 44828 29662 44884
rect 30034 44828 30044 44884
rect 30100 44828 32004 44884
rect 34738 44828 34748 44884
rect 34804 44828 37324 44884
rect 37380 44828 37390 44884
rect 39106 44828 39116 44884
rect 39172 44828 39228 44884
rect 39284 44828 39294 44884
rect 39788 44828 40012 44884
rect 40068 44828 40796 44884
rect 40852 44828 40862 44884
rect 41010 44828 41020 44884
rect 41076 44828 42028 44884
rect 42084 44828 42094 44884
rect 42364 44828 44884 44884
rect 12348 44772 12404 44828
rect 2034 44716 2044 44772
rect 2100 44716 4172 44772
rect 4228 44716 4238 44772
rect 4946 44716 4956 44772
rect 5012 44716 6300 44772
rect 6356 44716 6366 44772
rect 8082 44716 8092 44772
rect 8148 44716 9436 44772
rect 9492 44716 9502 44772
rect 9660 44716 11004 44772
rect 11060 44716 11070 44772
rect 11330 44716 11340 44772
rect 11396 44716 11564 44772
rect 11620 44716 12348 44772
rect 12404 44716 12414 44772
rect 12786 44716 12796 44772
rect 12852 44716 13356 44772
rect 13412 44716 13422 44772
rect 0 44660 112 44688
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 16828 44660 16884 44828
rect 25004 44772 25060 44828
rect 31948 44772 32004 44828
rect 17042 44716 17052 44772
rect 17108 44716 17276 44772
rect 17332 44716 19796 44772
rect 19954 44716 19964 44772
rect 20020 44716 23660 44772
rect 23716 44716 23726 44772
rect 25004 44716 25900 44772
rect 25956 44716 25966 44772
rect 27570 44716 27580 44772
rect 27636 44716 30716 44772
rect 30772 44716 30782 44772
rect 30930 44716 30940 44772
rect 30996 44716 31164 44772
rect 31220 44716 31230 44772
rect 31378 44716 31388 44772
rect 31444 44716 31724 44772
rect 31780 44716 31790 44772
rect 31948 44716 37660 44772
rect 37716 44716 37726 44772
rect 38658 44716 38668 44772
rect 38724 44716 42140 44772
rect 42196 44716 42206 44772
rect 0 44604 3388 44660
rect 5170 44604 5180 44660
rect 5236 44604 5292 44660
rect 5348 44604 5358 44660
rect 5842 44604 5852 44660
rect 5908 44604 7084 44660
rect 7140 44604 8540 44660
rect 8596 44604 8606 44660
rect 9538 44604 9548 44660
rect 9604 44604 11116 44660
rect 11172 44604 11182 44660
rect 13570 44604 13580 44660
rect 13636 44604 16884 44660
rect 18274 44604 18284 44660
rect 18340 44604 18956 44660
rect 19012 44604 19022 44660
rect 0 44576 112 44604
rect 3332 44548 3388 44604
rect 1922 44492 1932 44548
rect 1988 44492 2156 44548
rect 2212 44492 2222 44548
rect 3332 44492 18172 44548
rect 18228 44492 18238 44548
rect 18386 44492 18396 44548
rect 18452 44492 19292 44548
rect 19348 44492 19358 44548
rect 19740 44436 19796 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 42364 44660 42420 44828
rect 44828 44772 44884 44828
rect 45836 44828 46788 44884
rect 46946 44828 46956 44884
rect 47012 44828 47516 44884
rect 47572 44828 47582 44884
rect 49718 44828 49756 44884
rect 49812 44828 49822 44884
rect 49970 44828 49980 44884
rect 50036 44828 50652 44884
rect 50708 44828 50718 44884
rect 50978 44828 50988 44884
rect 51044 44828 52108 44884
rect 52164 44828 52174 44884
rect 45836 44772 45892 44828
rect 53340 44772 53396 44940
rect 53778 44828 53788 44884
rect 53844 44828 54124 44884
rect 54180 44828 54190 44884
rect 54870 44828 54908 44884
rect 54964 44828 54974 44884
rect 55356 44772 55412 44940
rect 42578 44716 42588 44772
rect 42644 44716 43484 44772
rect 43540 44716 43550 44772
rect 44828 44716 45892 44772
rect 46610 44716 46620 44772
rect 46676 44716 53396 44772
rect 53554 44716 53564 44772
rect 53620 44716 54012 44772
rect 54068 44716 54078 44772
rect 54450 44716 54460 44772
rect 54516 44716 54526 44772
rect 55356 44716 56252 44772
rect 56308 44716 56318 44772
rect 44454 44660 44464 44716
rect 44520 44660 44568 44716
rect 44624 44660 44672 44716
rect 44728 44660 44738 44716
rect 54460 44660 54516 44716
rect 57344 44660 57456 44688
rect 21186 44604 21196 44660
rect 21252 44604 22428 44660
rect 22484 44604 22494 44660
rect 25218 44604 25228 44660
rect 25284 44604 26684 44660
rect 26740 44604 26750 44660
rect 27906 44604 27916 44660
rect 27972 44604 28140 44660
rect 28196 44604 28206 44660
rect 31266 44604 31276 44660
rect 31332 44604 32844 44660
rect 32900 44604 32910 44660
rect 37538 44604 37548 44660
rect 37604 44604 40348 44660
rect 40404 44604 40414 44660
rect 41234 44604 41244 44660
rect 41300 44604 42420 44660
rect 42690 44604 42700 44660
rect 42756 44604 42924 44660
rect 42980 44604 43820 44660
rect 43876 44604 43886 44660
rect 45042 44604 45052 44660
rect 45108 44604 50764 44660
rect 50820 44604 50830 44660
rect 51202 44604 51212 44660
rect 51268 44604 54516 44660
rect 55804 44604 57456 44660
rect 25228 44548 25284 44604
rect 55804 44548 55860 44604
rect 57344 44576 57456 44604
rect 24332 44492 25284 44548
rect 26114 44492 26124 44548
rect 26180 44492 30604 44548
rect 30660 44492 30670 44548
rect 31378 44492 31388 44548
rect 31444 44492 31948 44548
rect 32004 44492 32014 44548
rect 35522 44492 35532 44548
rect 35588 44492 37436 44548
rect 37492 44492 37502 44548
rect 37650 44492 37660 44548
rect 37716 44492 55860 44548
rect 24332 44436 24388 44492
rect 1810 44380 1820 44436
rect 1876 44380 1932 44436
rect 1988 44380 1998 44436
rect 2594 44380 2604 44436
rect 2660 44380 4284 44436
rect 4340 44380 4350 44436
rect 4508 44380 6188 44436
rect 6244 44380 6254 44436
rect 6626 44380 6636 44436
rect 6692 44380 6972 44436
rect 7028 44380 7038 44436
rect 8194 44380 8204 44436
rect 8260 44380 9884 44436
rect 9940 44380 9950 44436
rect 10658 44380 10668 44436
rect 10724 44380 13132 44436
rect 13188 44380 13198 44436
rect 13346 44380 13356 44436
rect 13412 44380 16940 44436
rect 16996 44380 17006 44436
rect 17826 44380 17836 44436
rect 17892 44380 18620 44436
rect 18676 44380 18686 44436
rect 19740 44380 22540 44436
rect 22596 44380 22606 44436
rect 23660 44380 24388 44436
rect 30594 44380 30604 44436
rect 30660 44380 30996 44436
rect 31154 44380 31164 44436
rect 31220 44380 37548 44436
rect 37604 44380 37614 44436
rect 38098 44380 38108 44436
rect 38164 44380 38668 44436
rect 38724 44380 38734 44436
rect 39890 44380 39900 44436
rect 39956 44380 40236 44436
rect 40292 44380 40302 44436
rect 40898 44380 40908 44436
rect 40964 44380 41244 44436
rect 41300 44380 41310 44436
rect 41570 44380 41580 44436
rect 41636 44380 41804 44436
rect 41860 44380 41870 44436
rect 42130 44380 42140 44436
rect 42196 44380 42924 44436
rect 42980 44380 42990 44436
rect 43250 44380 43260 44436
rect 43316 44380 44940 44436
rect 44996 44380 45006 44436
rect 45798 44380 45836 44436
rect 45892 44380 47068 44436
rect 47124 44380 47134 44436
rect 48514 44380 48524 44436
rect 48580 44380 48748 44436
rect 48804 44380 48814 44436
rect 48962 44380 48972 44436
rect 49028 44380 49532 44436
rect 49588 44380 49598 44436
rect 50306 44380 50316 44436
rect 50372 44380 51548 44436
rect 51604 44380 51614 44436
rect 53890 44380 53900 44436
rect 53956 44380 53966 44436
rect 54450 44380 54460 44436
rect 54516 44380 56196 44436
rect 56354 44380 56364 44436
rect 56420 44380 56924 44436
rect 56980 44380 56990 44436
rect 4508 44324 4564 44380
rect 23660 44324 23716 44380
rect 30940 44324 30996 44380
rect 53900 44324 53956 44380
rect 2034 44268 2044 44324
rect 2100 44268 3276 44324
rect 3332 44268 4564 44324
rect 5170 44268 5180 44324
rect 5236 44268 8092 44324
rect 8148 44268 8158 44324
rect 8754 44268 8764 44324
rect 8820 44268 11228 44324
rect 11284 44268 11294 44324
rect 11666 44268 11676 44324
rect 11732 44268 13356 44324
rect 13412 44268 13468 44324
rect 13524 44268 13534 44324
rect 15138 44268 15148 44324
rect 15204 44268 20524 44324
rect 20580 44268 20590 44324
rect 20850 44268 20860 44324
rect 20916 44268 22764 44324
rect 22820 44268 23716 44324
rect 23884 44268 24780 44324
rect 24836 44268 24846 44324
rect 25554 44268 25564 44324
rect 25620 44268 27244 44324
rect 27300 44268 27310 44324
rect 27794 44268 27804 44324
rect 27860 44268 28476 44324
rect 28532 44268 28542 44324
rect 28914 44268 28924 44324
rect 28980 44268 30716 44324
rect 30772 44268 30782 44324
rect 30940 44268 31388 44324
rect 31444 44268 31454 44324
rect 31826 44268 31836 44324
rect 31892 44268 32508 44324
rect 32564 44268 32574 44324
rect 33170 44268 33180 44324
rect 33236 44268 34076 44324
rect 34132 44268 34142 44324
rect 36082 44268 36092 44324
rect 36148 44268 37100 44324
rect 37156 44268 37166 44324
rect 37650 44268 37660 44324
rect 37716 44268 50988 44324
rect 51044 44268 51054 44324
rect 51398 44268 51436 44324
rect 51492 44268 51502 44324
rect 53900 44268 54124 44324
rect 54180 44268 54190 44324
rect 0 44212 112 44240
rect 23884 44212 23940 44268
rect 56140 44212 56196 44380
rect 57344 44212 57456 44240
rect 0 44156 1820 44212
rect 1876 44156 1886 44212
rect 4274 44156 4284 44212
rect 4340 44156 5068 44212
rect 5124 44156 5134 44212
rect 5394 44156 5404 44212
rect 5460 44156 6636 44212
rect 6692 44156 6702 44212
rect 7522 44156 7532 44212
rect 7588 44156 13636 44212
rect 20066 44156 20076 44212
rect 20132 44156 22204 44212
rect 22260 44156 22270 44212
rect 22418 44156 22428 44212
rect 22484 44156 23940 44212
rect 24220 44156 25900 44212
rect 25956 44156 25966 44212
rect 27010 44156 27020 44212
rect 27076 44156 29148 44212
rect 29204 44156 29214 44212
rect 29362 44156 29372 44212
rect 29428 44156 31276 44212
rect 31332 44156 31342 44212
rect 31938 44156 31948 44212
rect 32004 44156 36372 44212
rect 36754 44156 36764 44212
rect 36820 44156 44156 44212
rect 44212 44156 44222 44212
rect 48178 44156 48188 44212
rect 48244 44156 48524 44212
rect 48580 44156 48748 44212
rect 48804 44156 49196 44212
rect 49252 44156 49262 44212
rect 50418 44156 50428 44212
rect 50484 44156 52892 44212
rect 52948 44156 52958 44212
rect 53890 44156 53900 44212
rect 53956 44156 54796 44212
rect 54852 44156 54862 44212
rect 56140 44156 57456 44212
rect 0 44128 112 44156
rect 3668 44044 6860 44100
rect 6916 44044 7364 44100
rect 7522 44044 7532 44100
rect 7588 44044 7980 44100
rect 8036 44044 8046 44100
rect 8194 44044 8204 44100
rect 8260 44044 9772 44100
rect 9828 44044 9838 44100
rect 10322 44044 10332 44100
rect 10388 44044 10780 44100
rect 10836 44044 10846 44100
rect 3668 43988 3724 44044
rect 7308 43988 7364 44044
rect 13580 43988 13636 44156
rect 24220 44100 24276 44156
rect 36316 44100 36372 44156
rect 57344 44128 57456 44156
rect 13794 44044 13804 44100
rect 13860 44044 16156 44100
rect 16212 44044 16222 44100
rect 19058 44044 19068 44100
rect 19124 44044 19628 44100
rect 19684 44044 19694 44100
rect 20962 44044 20972 44100
rect 21028 44044 23996 44100
rect 24052 44044 24062 44100
rect 24210 44044 24220 44100
rect 24276 44044 24286 44100
rect 24770 44044 24780 44100
rect 24836 44044 26684 44100
rect 26740 44044 26750 44100
rect 26898 44044 26908 44100
rect 26964 44044 28980 44100
rect 30594 44044 30604 44100
rect 30660 44044 30940 44100
rect 30996 44044 31006 44100
rect 31490 44044 31500 44100
rect 31556 44044 34076 44100
rect 34132 44044 34142 44100
rect 36316 44044 37436 44100
rect 37492 44044 37502 44100
rect 38658 44044 38668 44100
rect 38724 44044 39228 44100
rect 39284 44044 39294 44100
rect 39778 44044 39788 44100
rect 39844 44044 42812 44100
rect 42868 44044 42878 44100
rect 43036 44044 44660 44100
rect 130 43932 140 43988
rect 196 43932 812 43988
rect 868 43932 878 43988
rect 1586 43932 1596 43988
rect 1652 43932 3724 43988
rect 4162 43932 4172 43988
rect 4228 43932 6804 43988
rect 6934 43932 6972 43988
rect 7028 43932 7038 43988
rect 7308 43932 7868 43988
rect 7924 43932 7934 43988
rect 8418 43932 8428 43988
rect 8484 43932 9828 43988
rect 9986 43932 9996 43988
rect 10052 43932 10668 43988
rect 10724 43932 11116 43988
rect 11172 43932 12236 43988
rect 12292 43932 12302 43988
rect 13580 43932 17276 43988
rect 17332 43932 17342 43988
rect 18498 43932 18508 43988
rect 18564 43932 21308 43988
rect 21364 43932 21374 43988
rect 21532 43932 23548 43988
rect 23604 43932 23614 43988
rect 24882 43932 24892 43988
rect 24948 43932 26124 43988
rect 26180 43932 28700 43988
rect 28756 43932 28766 43988
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 5282 43820 5292 43876
rect 5348 43820 6300 43876
rect 6356 43820 6366 43876
rect 0 43764 112 43792
rect 6748 43764 6804 43932
rect 9772 43876 9828 43932
rect 21532 43876 21588 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 28924 43876 28980 44044
rect 43036 43988 43092 44044
rect 31052 43932 31948 43988
rect 32004 43932 32014 43988
rect 35298 43932 35308 43988
rect 35364 43932 36204 43988
rect 36260 43932 36270 43988
rect 36642 43932 36652 43988
rect 36708 43932 43092 43988
rect 44604 43988 44660 44044
rect 45052 44044 50876 44100
rect 50932 44044 50942 44100
rect 51202 44044 51212 44100
rect 51268 44044 51436 44100
rect 51492 44044 51502 44100
rect 51650 44044 51660 44100
rect 51716 44044 54012 44100
rect 54068 44044 54078 44100
rect 54338 44044 54348 44100
rect 54404 44044 55020 44100
rect 55076 44044 55086 44100
rect 45052 43988 45108 44044
rect 44604 43932 45108 43988
rect 46274 43932 46284 43988
rect 46340 43932 48524 43988
rect 48580 43932 48590 43988
rect 48738 43932 48748 43988
rect 48804 43932 56476 43988
rect 56532 43932 56542 43988
rect 31052 43876 31108 43932
rect 43794 43876 43804 43932
rect 43860 43876 43908 43932
rect 43964 43876 44012 43932
rect 44068 43876 44078 43932
rect 8754 43820 8764 43876
rect 8820 43820 9548 43876
rect 9604 43820 9614 43876
rect 9772 43820 10556 43876
rect 10612 43820 10622 43876
rect 12684 43820 15148 43876
rect 15204 43820 15214 43876
rect 15362 43820 15372 43876
rect 15428 43820 16380 43876
rect 16436 43820 16446 43876
rect 16818 43820 16828 43876
rect 16884 43820 21588 43876
rect 24210 43820 24220 43876
rect 24276 43820 25004 43876
rect 25060 43820 25070 43876
rect 28924 43820 31108 43876
rect 31378 43820 31388 43876
rect 31444 43820 34524 43876
rect 34580 43820 37996 43876
rect 38052 43820 38062 43876
rect 38210 43820 38220 43876
rect 38276 43820 39004 43876
rect 39060 43820 39070 43876
rect 39302 43820 39340 43876
rect 39396 43820 39406 43876
rect 39666 43820 39676 43876
rect 39732 43820 39788 43876
rect 39844 43820 39854 43876
rect 40338 43820 40348 43876
rect 40404 43820 41244 43876
rect 41300 43820 41310 43876
rect 42914 43820 42924 43876
rect 42980 43820 43260 43876
rect 43316 43820 43326 43876
rect 44146 43820 44156 43876
rect 44212 43820 53004 43876
rect 53060 43820 53070 43876
rect 53218 43820 53228 43876
rect 53284 43820 56140 43876
rect 56196 43820 56206 43876
rect 12684 43764 12740 43820
rect 57344 43764 57456 43792
rect 0 43708 140 43764
rect 196 43708 206 43764
rect 3332 43708 5964 43764
rect 6020 43708 6030 43764
rect 6748 43708 11844 43764
rect 12646 43708 12684 43764
rect 12740 43708 12750 43764
rect 12898 43708 12908 43764
rect 12964 43708 20076 43764
rect 20132 43708 20142 43764
rect 20626 43708 20636 43764
rect 20692 43708 22148 43764
rect 22418 43708 22428 43764
rect 22484 43708 26908 43764
rect 26964 43708 26974 43764
rect 29698 43708 29708 43764
rect 29764 43708 32732 43764
rect 32788 43708 32798 43764
rect 33954 43708 33964 43764
rect 34020 43708 36652 43764
rect 36708 43708 36718 43764
rect 37202 43708 37212 43764
rect 37268 43708 38444 43764
rect 38500 43708 41020 43764
rect 41076 43708 41086 43764
rect 41346 43708 41356 43764
rect 41412 43708 43708 43764
rect 43764 43708 43774 43764
rect 43922 43708 43932 43764
rect 43988 43708 50092 43764
rect 50148 43708 50158 43764
rect 51762 43708 51772 43764
rect 51828 43708 52332 43764
rect 52388 43708 52398 43764
rect 53666 43708 53676 43764
rect 53732 43708 54572 43764
rect 54628 43708 54638 43764
rect 54786 43708 54796 43764
rect 54852 43708 54890 43764
rect 57148 43708 57456 43764
rect 0 43680 112 43708
rect 3332 43652 3388 43708
rect 11788 43652 11844 43708
rect 22092 43652 22148 43708
rect 690 43596 700 43652
rect 756 43596 2044 43652
rect 2100 43596 2110 43652
rect 3154 43596 3164 43652
rect 3220 43596 3388 43652
rect 6178 43596 6188 43652
rect 6244 43596 9324 43652
rect 9380 43596 9390 43652
rect 9538 43596 9548 43652
rect 9604 43596 9884 43652
rect 9940 43596 10780 43652
rect 10836 43596 10846 43652
rect 10994 43596 11004 43652
rect 11060 43596 11340 43652
rect 11396 43596 11406 43652
rect 11788 43596 13468 43652
rect 13524 43596 13534 43652
rect 16034 43596 16044 43652
rect 16100 43596 17164 43652
rect 17220 43596 17230 43652
rect 22092 43596 31276 43652
rect 31332 43596 31342 43652
rect 34738 43596 34748 43652
rect 34804 43596 36876 43652
rect 36932 43596 36942 43652
rect 37100 43596 50428 43652
rect 50866 43596 50876 43652
rect 50932 43596 51996 43652
rect 52052 43596 52062 43652
rect 53554 43596 53564 43652
rect 53620 43596 53900 43652
rect 53956 43596 53966 43652
rect 54450 43596 54460 43652
rect 54516 43596 54684 43652
rect 54740 43596 55020 43652
rect 55076 43596 55086 43652
rect 37100 43540 37156 43596
rect 578 43484 588 43540
rect 644 43484 3276 43540
rect 3332 43484 3342 43540
rect 3602 43484 3612 43540
rect 3668 43484 4060 43540
rect 4116 43484 4126 43540
rect 4274 43484 4284 43540
rect 4340 43484 4844 43540
rect 4900 43484 4910 43540
rect 5730 43484 5740 43540
rect 5796 43484 7084 43540
rect 7140 43484 7150 43540
rect 7858 43484 7868 43540
rect 7924 43484 9660 43540
rect 9716 43484 9726 43540
rect 10546 43484 10556 43540
rect 10612 43484 11452 43540
rect 11508 43484 11518 43540
rect 13234 43484 13244 43540
rect 13300 43484 13310 43540
rect 15138 43484 15148 43540
rect 15204 43484 15372 43540
rect 15428 43484 15438 43540
rect 15810 43484 15820 43540
rect 15876 43484 16772 43540
rect 16930 43484 16940 43540
rect 16996 43484 19628 43540
rect 19684 43484 19694 43540
rect 19814 43484 19852 43540
rect 19908 43484 19918 43540
rect 20738 43484 20748 43540
rect 20804 43484 21868 43540
rect 21924 43484 21934 43540
rect 24966 43484 25004 43540
rect 25060 43484 25070 43540
rect 26338 43484 26348 43540
rect 26404 43484 27468 43540
rect 27524 43484 27534 43540
rect 28242 43484 28252 43540
rect 28308 43484 29932 43540
rect 29988 43484 29998 43540
rect 31602 43484 31612 43540
rect 31668 43484 37156 43540
rect 43026 43484 43036 43540
rect 43092 43484 44268 43540
rect 44324 43484 44334 43540
rect 44482 43484 44492 43540
rect 44548 43484 45388 43540
rect 45444 43484 45948 43540
rect 46004 43484 46844 43540
rect 46900 43484 46910 43540
rect 47394 43484 47404 43540
rect 47460 43484 49196 43540
rect 49252 43484 49262 43540
rect 13244 43428 13300 43484
rect 16716 43428 16772 43484
rect 50372 43428 50428 43596
rect 57148 43540 57204 43708
rect 57344 43680 57456 43708
rect 50754 43484 50764 43540
rect 50820 43484 51212 43540
rect 51268 43484 52108 43540
rect 52164 43484 52174 43540
rect 52658 43484 52668 43540
rect 52724 43484 53564 43540
rect 53620 43484 54124 43540
rect 54180 43484 56140 43540
rect 56196 43484 56206 43540
rect 57148 43484 57372 43540
rect 57428 43484 57438 43540
rect 354 43372 364 43428
rect 420 43372 1596 43428
rect 1652 43372 1662 43428
rect 1810 43372 1820 43428
rect 1876 43372 7420 43428
rect 7476 43372 7486 43428
rect 8754 43372 8764 43428
rect 8820 43372 10444 43428
rect 10500 43372 11228 43428
rect 11284 43372 11294 43428
rect 12226 43372 12236 43428
rect 12292 43372 13300 43428
rect 13906 43372 13916 43428
rect 13972 43372 16044 43428
rect 16100 43372 16492 43428
rect 16548 43372 16558 43428
rect 16716 43372 19964 43428
rect 20020 43372 20030 43428
rect 20402 43372 20412 43428
rect 20468 43372 21644 43428
rect 21700 43372 21710 43428
rect 24322 43372 24332 43428
rect 24388 43372 25676 43428
rect 25732 43372 25742 43428
rect 27234 43372 27244 43428
rect 27300 43372 28588 43428
rect 28644 43372 28654 43428
rect 29810 43372 29820 43428
rect 29876 43372 32956 43428
rect 33012 43372 33022 43428
rect 33170 43372 33180 43428
rect 33236 43372 33516 43428
rect 33572 43372 33582 43428
rect 33730 43372 33740 43428
rect 33796 43372 34412 43428
rect 34468 43372 34478 43428
rect 35634 43372 35644 43428
rect 35700 43372 39340 43428
rect 39396 43372 39406 43428
rect 40226 43372 40236 43428
rect 40292 43372 40460 43428
rect 40516 43372 40526 43428
rect 41234 43372 41244 43428
rect 41300 43372 41916 43428
rect 41972 43372 41982 43428
rect 42466 43372 42476 43428
rect 42532 43372 44156 43428
rect 44212 43372 44222 43428
rect 47814 43372 47852 43428
rect 47908 43372 47918 43428
rect 48626 43372 48636 43428
rect 48692 43372 49756 43428
rect 49812 43372 49822 43428
rect 50372 43372 50988 43428
rect 51044 43372 51054 43428
rect 51286 43372 51324 43428
rect 51380 43372 51390 43428
rect 52210 43372 52220 43428
rect 52276 43372 52780 43428
rect 52836 43372 52846 43428
rect 55794 43372 55804 43428
rect 55860 43372 56364 43428
rect 56420 43372 56430 43428
rect 0 43316 112 43344
rect 57344 43316 57456 43344
rect 0 43260 6636 43316
rect 6692 43260 6702 43316
rect 6962 43260 6972 43316
rect 7028 43260 8708 43316
rect 8978 43260 8988 43316
rect 9044 43260 10220 43316
rect 10276 43260 10286 43316
rect 11554 43260 11564 43316
rect 11620 43260 12124 43316
rect 12180 43260 12190 43316
rect 12674 43260 12684 43316
rect 12740 43260 13244 43316
rect 13300 43260 17388 43316
rect 17444 43260 17454 43316
rect 19282 43260 19292 43316
rect 19348 43260 21756 43316
rect 21812 43260 21822 43316
rect 22642 43260 22652 43316
rect 22708 43260 23548 43316
rect 0 43232 112 43260
rect 8652 43204 8708 43260
rect 23492 43204 23548 43260
rect 23660 43260 29372 43316
rect 29428 43260 29438 43316
rect 29586 43260 29596 43316
rect 29652 43260 30268 43316
rect 30324 43260 30334 43316
rect 32274 43260 32284 43316
rect 32340 43260 33180 43316
rect 33236 43260 37100 43316
rect 37156 43260 37324 43316
rect 37380 43260 37390 43316
rect 37734 43260 37772 43316
rect 37828 43260 37838 43316
rect 38882 43260 38892 43316
rect 38948 43260 40908 43316
rect 40964 43260 41804 43316
rect 41860 43260 41870 43316
rect 43586 43260 43596 43316
rect 43652 43260 45724 43316
rect 45780 43260 45790 43316
rect 46610 43260 46620 43316
rect 46676 43260 47180 43316
rect 47236 43260 47246 43316
rect 48402 43260 48412 43316
rect 48468 43260 48860 43316
rect 48916 43260 48926 43316
rect 50530 43260 50540 43316
rect 50596 43260 50764 43316
rect 50820 43260 52556 43316
rect 52612 43260 52622 43316
rect 53526 43260 53564 43316
rect 53620 43260 53630 43316
rect 55458 43260 55468 43316
rect 55524 43260 57456 43316
rect 23660 43204 23716 43260
rect 57344 43232 57456 43260
rect 1138 43148 1148 43204
rect 1204 43148 2940 43204
rect 2996 43148 3006 43204
rect 3378 43148 3388 43204
rect 3444 43148 4284 43204
rect 4340 43148 4350 43204
rect 6738 43148 6748 43204
rect 6804 43148 7196 43204
rect 7252 43148 8428 43204
rect 8484 43148 8494 43204
rect 8652 43148 20972 43204
rect 21028 43148 21038 43204
rect 23492 43148 23716 43204
rect 27234 43148 27244 43204
rect 27300 43148 38556 43204
rect 38612 43148 38622 43204
rect 38770 43148 38780 43204
rect 38836 43148 41020 43204
rect 41076 43148 41086 43204
rect 43138 43148 43148 43204
rect 43204 43148 44268 43204
rect 44324 43148 44334 43204
rect 46162 43148 46172 43204
rect 46228 43148 50372 43204
rect 50428 43148 50438 43204
rect 50652 43148 51660 43204
rect 51716 43148 51996 43204
rect 52052 43148 52062 43204
rect 52220 43148 55020 43204
rect 55076 43148 55086 43204
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 130 43036 140 43092
rect 196 43036 2604 43092
rect 2660 43036 2670 43092
rect 3378 43036 3388 43092
rect 3444 43036 3724 43092
rect 3780 43036 3790 43092
rect 6290 43036 6300 43092
rect 6356 43036 8204 43092
rect 8260 43036 9212 43092
rect 9268 43036 9278 43092
rect 9538 43036 9548 43092
rect 9604 43036 9660 43092
rect 9716 43036 9726 43092
rect 9986 43036 9996 43092
rect 10052 43036 19740 43092
rect 19796 43036 19806 43092
rect 20178 43036 20188 43092
rect 20244 43036 21756 43092
rect 21812 43036 23436 43092
rect 23492 43036 23502 43092
rect 23762 43036 23772 43092
rect 23828 43036 24332 43092
rect 24388 43036 24398 43092
rect 26450 43036 26460 43092
rect 26516 43036 27916 43092
rect 27972 43036 27982 43092
rect 28354 43036 28364 43092
rect 28420 43036 29484 43092
rect 29540 43036 30940 43092
rect 30996 43036 31006 43092
rect 32498 43036 32508 43092
rect 32564 43036 33852 43092
rect 33908 43036 33918 43092
rect 34076 43036 34748 43092
rect 34804 43036 34814 43092
rect 34962 43036 34972 43092
rect 35028 43036 35196 43092
rect 35252 43036 35262 43092
rect 35634 43036 35644 43092
rect 35700 43036 36092 43092
rect 36148 43036 39564 43092
rect 39620 43036 39630 43092
rect 40450 43036 40460 43092
rect 40516 43036 42252 43092
rect 42308 43036 42318 43092
rect 34076 42980 34132 43036
rect 43148 42980 43204 43148
rect 44454 43092 44464 43148
rect 44520 43092 44568 43148
rect 44624 43092 44672 43148
rect 44728 43092 44738 43148
rect 50652 43092 50708 43148
rect 52220 43092 52276 43148
rect 49074 43036 49084 43092
rect 49140 43036 50708 43092
rect 50764 43036 52276 43092
rect 52406 43036 52444 43092
rect 52500 43036 52510 43092
rect 52770 43036 52780 43092
rect 52836 43036 54348 43092
rect 54404 43036 54796 43092
rect 54852 43036 54862 43092
rect 50764 42980 50820 43036
rect 690 42924 700 42980
rect 756 42924 1820 42980
rect 1876 42924 1886 42980
rect 2258 42924 2268 42980
rect 2324 42924 16716 42980
rect 16772 42924 16782 42980
rect 17154 42924 17164 42980
rect 17220 42924 31668 42980
rect 32946 42924 32956 42980
rect 33012 42924 34132 42980
rect 34626 42924 34636 42980
rect 34692 42924 34860 42980
rect 34916 42924 34926 42980
rect 35522 42924 35532 42980
rect 35588 42924 36428 42980
rect 36484 42924 36494 42980
rect 37538 42924 37548 42980
rect 37604 42924 37660 42980
rect 37716 42924 37726 42980
rect 37874 42924 37884 42980
rect 37940 42924 39228 42980
rect 39284 42924 39294 42980
rect 39778 42924 39788 42980
rect 39844 42924 43204 42980
rect 43698 42924 43708 42980
rect 43764 42924 45164 42980
rect 45220 42924 45230 42980
rect 45378 42924 45388 42980
rect 45444 42924 46844 42980
rect 46900 42924 46910 42980
rect 48514 42924 48524 42980
rect 48580 42924 50820 42980
rect 50978 42924 50988 42980
rect 51044 42924 54572 42980
rect 54628 42924 54638 42980
rect 55234 42924 55244 42980
rect 55300 42924 55692 42980
rect 55748 42924 55758 42980
rect 0 42868 112 42896
rect 0 42812 1036 42868
rect 1092 42812 1102 42868
rect 2706 42812 2716 42868
rect 2772 42812 3612 42868
rect 3668 42812 3678 42868
rect 4284 42812 8988 42868
rect 9044 42812 9054 42868
rect 9650 42812 9660 42868
rect 9716 42812 11900 42868
rect 11956 42812 13356 42868
rect 13412 42812 13422 42868
rect 15474 42812 15484 42868
rect 15540 42812 17612 42868
rect 17668 42812 18060 42868
rect 18116 42812 18126 42868
rect 20066 42812 20076 42868
rect 20132 42812 28364 42868
rect 28420 42812 28430 42868
rect 0 42784 112 42812
rect 4284 42756 4340 42812
rect 31612 42756 31668 42924
rect 57344 42868 57456 42896
rect 33618 42812 33628 42868
rect 33684 42812 34412 42868
rect 34468 42812 34478 42868
rect 35746 42812 35756 42868
rect 35812 42812 39676 42868
rect 39732 42812 39742 42868
rect 40338 42812 40348 42868
rect 40404 42812 40908 42868
rect 40964 42812 40974 42868
rect 41206 42812 41244 42868
rect 41300 42812 41310 42868
rect 41458 42812 41468 42868
rect 41524 42812 41580 42868
rect 41636 42812 41646 42868
rect 45266 42812 45276 42868
rect 45332 42812 45724 42868
rect 45780 42812 45790 42868
rect 46610 42812 46620 42868
rect 46676 42812 47292 42868
rect 47348 42812 47358 42868
rect 47842 42812 47852 42868
rect 47908 42812 50204 42868
rect 50260 42812 53676 42868
rect 53732 42812 53742 42868
rect 55020 42812 56028 42868
rect 56084 42812 56094 42868
rect 56476 42812 57456 42868
rect 55020 42756 55076 42812
rect 3266 42700 3276 42756
rect 3332 42700 3500 42756
rect 3556 42700 3566 42756
rect 4274 42700 4284 42756
rect 4340 42700 4350 42756
rect 5954 42700 5964 42756
rect 6020 42700 6412 42756
rect 6468 42700 6478 42756
rect 7298 42700 7308 42756
rect 7364 42700 12124 42756
rect 12180 42700 12190 42756
rect 18508 42700 20860 42756
rect 20916 42700 20926 42756
rect 23090 42700 23100 42756
rect 23156 42700 26348 42756
rect 26404 42700 26414 42756
rect 28690 42700 28700 42756
rect 28756 42700 30044 42756
rect 30100 42700 30110 42756
rect 31612 42700 36316 42756
rect 36372 42700 36382 42756
rect 37090 42700 37100 42756
rect 37156 42700 37884 42756
rect 37940 42700 37950 42756
rect 38210 42700 38220 42756
rect 38276 42700 38668 42756
rect 38724 42700 38734 42756
rect 39330 42700 39340 42756
rect 39396 42700 42252 42756
rect 42308 42700 42318 42756
rect 43922 42700 43932 42756
rect 43988 42700 45052 42756
rect 45108 42700 45118 42756
rect 46274 42700 46284 42756
rect 46340 42700 47068 42756
rect 47124 42700 47134 42756
rect 50530 42700 50540 42756
rect 50596 42700 52108 42756
rect 52164 42700 52174 42756
rect 52434 42700 52444 42756
rect 52500 42700 55076 42756
rect 55234 42700 55244 42756
rect 55300 42700 56252 42756
rect 56308 42700 56318 42756
rect 1922 42588 1932 42644
rect 1988 42588 8092 42644
rect 8148 42588 8158 42644
rect 11778 42588 11788 42644
rect 11844 42588 12236 42644
rect 12292 42588 12302 42644
rect 12450 42588 12460 42644
rect 12516 42588 14588 42644
rect 14644 42588 14924 42644
rect 14980 42588 14990 42644
rect 16034 42588 16044 42644
rect 16100 42588 18284 42644
rect 18340 42588 18350 42644
rect 18508 42532 18564 42700
rect 56476 42644 56532 42812
rect 57344 42784 57456 42812
rect 19618 42588 19628 42644
rect 19684 42588 20524 42644
rect 20580 42588 20590 42644
rect 20962 42588 20972 42644
rect 21028 42588 28476 42644
rect 28532 42588 28542 42644
rect 30716 42588 35420 42644
rect 35476 42588 35486 42644
rect 36642 42588 36652 42644
rect 36708 42588 41132 42644
rect 41188 42588 41198 42644
rect 43362 42588 43372 42644
rect 43428 42588 45164 42644
rect 45220 42588 45724 42644
rect 45780 42588 45836 42644
rect 45892 42588 45902 42644
rect 46050 42588 46060 42644
rect 46116 42588 49196 42644
rect 49252 42588 49262 42644
rect 50204 42588 52892 42644
rect 52948 42588 52958 42644
rect 53442 42588 53452 42644
rect 53508 42588 54460 42644
rect 54516 42588 54526 42644
rect 54786 42588 54796 42644
rect 54852 42588 56532 42644
rect 30716 42532 30772 42588
rect 35420 42532 35476 42588
rect 50204 42532 50260 42588
rect 2258 42476 2268 42532
rect 2324 42476 2660 42532
rect 3350 42476 3388 42532
rect 3444 42476 3454 42532
rect 3938 42476 3948 42532
rect 4004 42476 7364 42532
rect 7522 42476 7532 42532
rect 7588 42476 10108 42532
rect 10164 42476 10556 42532
rect 10612 42476 10622 42532
rect 12114 42476 12124 42532
rect 12180 42476 18564 42532
rect 18946 42476 18956 42532
rect 19012 42476 25228 42532
rect 25284 42476 25294 42532
rect 29110 42476 29148 42532
rect 29204 42476 30772 42532
rect 31378 42476 31388 42532
rect 31444 42476 31948 42532
rect 32004 42476 32014 42532
rect 32946 42476 32956 42532
rect 33012 42476 35084 42532
rect 35140 42476 35150 42532
rect 35420 42476 35980 42532
rect 36036 42476 36046 42532
rect 37202 42476 37212 42532
rect 37268 42476 38668 42532
rect 38724 42476 38734 42532
rect 41346 42476 41356 42532
rect 41412 42476 44212 42532
rect 47730 42476 47740 42532
rect 47796 42476 50260 42532
rect 50418 42476 50428 42532
rect 50484 42476 53228 42532
rect 53284 42476 53294 42532
rect 54562 42476 54572 42532
rect 54628 42476 55244 42532
rect 55300 42476 55310 42532
rect 0 42420 112 42448
rect 2604 42420 2660 42476
rect 7308 42420 7364 42476
rect 44156 42420 44212 42476
rect 57344 42420 57456 42448
rect 0 42364 2380 42420
rect 2436 42364 2446 42420
rect 2604 42364 3500 42420
rect 3556 42364 3566 42420
rect 4834 42364 4844 42420
rect 4900 42364 5740 42420
rect 5796 42364 5806 42420
rect 7308 42364 12572 42420
rect 12628 42364 14700 42420
rect 14756 42364 14766 42420
rect 14914 42364 14924 42420
rect 14980 42364 15820 42420
rect 15876 42364 15886 42420
rect 16034 42364 16044 42420
rect 16100 42364 20300 42420
rect 20356 42364 20366 42420
rect 20626 42364 20636 42420
rect 20692 42364 21308 42420
rect 21364 42364 21374 42420
rect 25218 42364 25228 42420
rect 25284 42364 39676 42420
rect 39732 42364 39742 42420
rect 40898 42364 40908 42420
rect 40964 42364 43372 42420
rect 43428 42364 43438 42420
rect 44156 42364 47908 42420
rect 49746 42364 49756 42420
rect 49812 42364 55580 42420
rect 55636 42364 55646 42420
rect 55794 42364 55804 42420
rect 55860 42364 57456 42420
rect 0 42336 112 42364
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 43794 42308 43804 42364
rect 43860 42308 43908 42364
rect 43964 42308 44012 42364
rect 44068 42308 44078 42364
rect 1250 42252 1260 42308
rect 1316 42252 1484 42308
rect 1540 42252 1550 42308
rect 6290 42252 6300 42308
rect 6356 42252 6860 42308
rect 6916 42252 7084 42308
rect 7140 42252 7150 42308
rect 8418 42252 8428 42308
rect 8484 42252 8876 42308
rect 8932 42252 8942 42308
rect 9090 42252 9100 42308
rect 9156 42252 9324 42308
rect 9380 42252 9390 42308
rect 10108 42252 10892 42308
rect 10948 42252 10958 42308
rect 11106 42252 11116 42308
rect 11172 42252 16268 42308
rect 16324 42252 16334 42308
rect 16818 42252 16828 42308
rect 16884 42252 19740 42308
rect 19796 42252 21980 42308
rect 22036 42252 22046 42308
rect 22306 42252 22316 42308
rect 22372 42252 22764 42308
rect 22820 42252 22830 42308
rect 26450 42252 26460 42308
rect 26516 42252 27468 42308
rect 27524 42252 27692 42308
rect 27748 42252 27758 42308
rect 28354 42252 28364 42308
rect 28420 42252 38220 42308
rect 38276 42252 38286 42308
rect 38658 42252 38668 42308
rect 38724 42252 39564 42308
rect 39620 42252 40572 42308
rect 40628 42252 40638 42308
rect 41010 42252 41020 42308
rect 41076 42252 43484 42308
rect 43540 42252 43550 42308
rect 44146 42252 44156 42308
rect 44212 42252 45388 42308
rect 45444 42252 45454 42308
rect 2930 42140 2940 42196
rect 2996 42140 5348 42196
rect 5506 42140 5516 42196
rect 5572 42140 6188 42196
rect 6244 42140 8988 42196
rect 9044 42140 9054 42196
rect 9314 42140 9324 42196
rect 9380 42140 9548 42196
rect 9604 42140 9614 42196
rect 5292 42084 5348 42140
rect 10108 42084 10164 42252
rect 47852 42196 47908 42364
rect 57344 42336 57456 42364
rect 48066 42252 48076 42308
rect 48132 42252 51772 42308
rect 51828 42252 51838 42308
rect 52546 42252 52556 42308
rect 52612 42252 52668 42308
rect 52724 42252 52734 42308
rect 52882 42252 52892 42308
rect 52948 42252 53788 42308
rect 53844 42252 53854 42308
rect 10546 42140 10556 42196
rect 10612 42140 12796 42196
rect 12852 42140 12862 42196
rect 13010 42140 13020 42196
rect 13076 42140 14812 42196
rect 14868 42140 14878 42196
rect 15810 42140 15820 42196
rect 15876 42140 47628 42196
rect 47684 42140 47694 42196
rect 47852 42140 50204 42196
rect 50260 42140 50270 42196
rect 50418 42140 50428 42196
rect 50484 42140 51436 42196
rect 51492 42140 51502 42196
rect 52098 42140 52108 42196
rect 52164 42140 52444 42196
rect 52500 42140 52510 42196
rect 52658 42140 52668 42196
rect 52724 42140 53452 42196
rect 53508 42140 53518 42196
rect 53778 42140 53788 42196
rect 53844 42140 54572 42196
rect 54628 42140 54638 42196
rect 3154 42028 3164 42084
rect 3220 42028 4284 42084
rect 4340 42028 4350 42084
rect 5292 42028 6636 42084
rect 6692 42028 6702 42084
rect 6962 42028 6972 42084
rect 7028 42028 7420 42084
rect 7476 42028 10164 42084
rect 10434 42028 10444 42084
rect 10500 42028 11788 42084
rect 11844 42028 11854 42084
rect 12002 42028 12012 42084
rect 12068 42028 12106 42084
rect 12338 42028 12348 42084
rect 12404 42028 12908 42084
rect 12964 42028 12974 42084
rect 13458 42028 13468 42084
rect 13524 42028 13580 42084
rect 13636 42028 14924 42084
rect 14980 42028 14990 42084
rect 17612 42028 24220 42084
rect 24276 42028 25452 42084
rect 25508 42028 25518 42084
rect 27234 42028 27244 42084
rect 27300 42028 28700 42084
rect 28756 42028 28766 42084
rect 29362 42028 29372 42084
rect 29428 42028 31388 42084
rect 31444 42028 31454 42084
rect 35074 42028 35084 42084
rect 35140 42028 37100 42084
rect 37156 42028 37166 42084
rect 37426 42028 37436 42084
rect 37492 42028 37772 42084
rect 37828 42028 37838 42084
rect 38098 42028 38108 42084
rect 38164 42028 41580 42084
rect 41636 42028 41646 42084
rect 42242 42028 42252 42084
rect 42308 42028 52332 42084
rect 52388 42028 52398 42084
rect 53778 42028 53788 42084
rect 53844 42028 55020 42084
rect 55076 42028 55086 42084
rect 55346 42028 55356 42084
rect 55412 42028 55580 42084
rect 55636 42028 55646 42084
rect 56102 42028 56140 42084
rect 56196 42028 56206 42084
rect 56774 42028 56812 42084
rect 56868 42028 56878 42084
rect 0 41972 112 42000
rect 17612 41972 17668 42028
rect 57344 41972 57456 42000
rect 0 41916 1708 41972
rect 1764 41916 1774 41972
rect 3490 41916 3500 41972
rect 3556 41916 4060 41972
rect 4116 41916 4126 41972
rect 5618 41916 5628 41972
rect 5684 41916 8764 41972
rect 8820 41916 8830 41972
rect 9314 41916 9324 41972
rect 9380 41916 11004 41972
rect 11060 41916 11070 41972
rect 12114 41916 12124 41972
rect 12180 41916 14812 41972
rect 14868 41916 14878 41972
rect 15474 41916 15484 41972
rect 15540 41916 17612 41972
rect 17668 41916 17678 41972
rect 19058 41916 19068 41972
rect 19124 41916 19516 41972
rect 19572 41916 19582 41972
rect 20178 41916 20188 41972
rect 20244 41916 20860 41972
rect 20916 41916 21980 41972
rect 22036 41916 22316 41972
rect 22372 41916 22382 41972
rect 22530 41916 22540 41972
rect 22596 41916 23324 41972
rect 23380 41916 23390 41972
rect 24210 41916 24220 41972
rect 24276 41916 25004 41972
rect 25060 41916 25070 41972
rect 31154 41916 31164 41972
rect 31220 41916 32060 41972
rect 32116 41916 32126 41972
rect 32386 41916 32396 41972
rect 32452 41916 32620 41972
rect 32676 41916 32686 41972
rect 33618 41916 33628 41972
rect 33684 41916 34076 41972
rect 34132 41916 34142 41972
rect 34514 41916 34524 41972
rect 34580 41916 38220 41972
rect 38276 41916 38286 41972
rect 38546 41916 38556 41972
rect 38612 41916 39788 41972
rect 39844 41916 39854 41972
rect 40338 41916 40348 41972
rect 40404 41916 40572 41972
rect 40628 41916 40638 41972
rect 41010 41916 41020 41972
rect 41076 41916 43652 41972
rect 44930 41916 44940 41972
rect 44996 41916 46508 41972
rect 46564 41916 46574 41972
rect 46722 41916 46732 41972
rect 46788 41916 46956 41972
rect 47012 41916 47022 41972
rect 47394 41916 47404 41972
rect 47460 41916 48524 41972
rect 48580 41916 49420 41972
rect 49476 41916 49486 41972
rect 49858 41916 49868 41972
rect 49924 41916 57456 41972
rect 0 41888 112 41916
rect 43596 41860 43652 41916
rect 57344 41888 57456 41916
rect 1558 41804 1596 41860
rect 1652 41804 1662 41860
rect 2482 41804 2492 41860
rect 2548 41804 3164 41860
rect 3220 41804 3230 41860
rect 3378 41804 3388 41860
rect 3444 41804 4172 41860
rect 4228 41804 4238 41860
rect 5058 41804 5068 41860
rect 5124 41804 5292 41860
rect 5348 41804 5516 41860
rect 5572 41804 5582 41860
rect 7410 41804 7420 41860
rect 7476 41804 8764 41860
rect 8820 41804 8830 41860
rect 10322 41804 10332 41860
rect 10388 41804 13020 41860
rect 13076 41804 13086 41860
rect 13244 41804 13468 41860
rect 13524 41804 14700 41860
rect 14756 41804 14766 41860
rect 15092 41804 18732 41860
rect 18788 41804 18798 41860
rect 21980 41804 25956 41860
rect 26338 41804 26348 41860
rect 26404 41804 29148 41860
rect 29204 41804 29214 41860
rect 30706 41804 30716 41860
rect 30772 41804 31612 41860
rect 31668 41804 31678 41860
rect 35186 41804 35196 41860
rect 35252 41804 35532 41860
rect 35588 41804 37212 41860
rect 37268 41804 37278 41860
rect 37398 41804 37436 41860
rect 37492 41804 37502 41860
rect 38612 41804 40684 41860
rect 40740 41804 40750 41860
rect 41906 41804 41916 41860
rect 41972 41804 42364 41860
rect 42420 41804 42430 41860
rect 42578 41804 42588 41860
rect 42644 41804 43036 41860
rect 43092 41804 43372 41860
rect 43428 41804 43438 41860
rect 43596 41804 55468 41860
rect 55524 41804 55534 41860
rect 13244 41748 13300 41804
rect 15092 41748 15148 41804
rect 21980 41748 22036 41804
rect 25900 41748 25956 41804
rect 38612 41748 38668 41804
rect 2482 41692 2492 41748
rect 2548 41692 2716 41748
rect 2772 41692 2782 41748
rect 3042 41692 3052 41748
rect 3108 41692 9660 41748
rect 9716 41692 9726 41748
rect 11732 41692 13300 41748
rect 13906 41692 13916 41748
rect 13972 41692 15148 41748
rect 16482 41692 16492 41748
rect 16548 41692 18508 41748
rect 18564 41692 18574 41748
rect 21970 41692 21980 41748
rect 22036 41692 22046 41748
rect 22866 41692 22876 41748
rect 22932 41692 24780 41748
rect 24836 41692 24846 41748
rect 25890 41692 25900 41748
rect 25956 41692 29820 41748
rect 29876 41692 29886 41748
rect 30594 41692 30604 41748
rect 30660 41692 33292 41748
rect 33348 41692 33358 41748
rect 34738 41692 34748 41748
rect 34804 41692 38668 41748
rect 38770 41692 38780 41748
rect 38836 41692 39676 41748
rect 39732 41692 41132 41748
rect 41188 41692 41198 41748
rect 43250 41692 43260 41748
rect 43316 41692 44828 41748
rect 44884 41692 44894 41748
rect 45490 41692 45500 41748
rect 45556 41692 47404 41748
rect 47460 41692 47470 41748
rect 47954 41692 47964 41748
rect 48020 41692 48076 41748
rect 48132 41692 48142 41748
rect 49186 41692 49196 41748
rect 49252 41692 50876 41748
rect 50932 41692 50942 41748
rect 51202 41692 51212 41748
rect 51268 41692 52332 41748
rect 52388 41692 52398 41748
rect 52882 41692 52892 41748
rect 52948 41692 53676 41748
rect 53732 41692 53742 41748
rect 55458 41692 55468 41748
rect 55524 41692 55692 41748
rect 55748 41692 55758 41748
rect 802 41580 812 41636
rect 868 41580 4284 41636
rect 4340 41580 4350 41636
rect 6850 41580 6860 41636
rect 6916 41580 8708 41636
rect 8866 41580 8876 41636
rect 8932 41580 10892 41636
rect 10948 41580 11340 41636
rect 11396 41580 11406 41636
rect 0 41524 112 41552
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 8652 41524 8708 41580
rect 11732 41524 11788 41692
rect 40684 41636 40740 41692
rect 55468 41636 55524 41692
rect 12002 41580 12012 41636
rect 12068 41580 16044 41636
rect 16100 41580 16110 41636
rect 16716 41580 20972 41636
rect 21028 41580 21038 41636
rect 23538 41580 23548 41636
rect 23604 41580 24220 41636
rect 24276 41580 24286 41636
rect 26226 41580 26236 41636
rect 26292 41580 28140 41636
rect 28196 41580 28206 41636
rect 28466 41580 28476 41636
rect 28532 41580 40516 41636
rect 40674 41580 40684 41636
rect 40740 41580 40750 41636
rect 41234 41580 41244 41636
rect 41300 41580 44156 41636
rect 44212 41580 44222 41636
rect 45714 41580 45724 41636
rect 45780 41580 49868 41636
rect 49924 41580 49934 41636
rect 50092 41580 52780 41636
rect 52836 41580 52846 41636
rect 53106 41580 53116 41636
rect 53172 41580 55524 41636
rect 56802 41580 56812 41636
rect 56868 41580 57148 41636
rect 57204 41580 57214 41636
rect 16716 41524 16772 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 40460 41524 40516 41580
rect 44454 41524 44464 41580
rect 44520 41524 44568 41580
rect 44624 41524 44672 41580
rect 44728 41524 44738 41580
rect 50092 41524 50148 41580
rect 57344 41524 57456 41552
rect 0 41468 1036 41524
rect 1092 41468 1102 41524
rect 2258 41468 2268 41524
rect 2324 41468 2380 41524
rect 2436 41468 3052 41524
rect 3108 41468 3118 41524
rect 3602 41468 3612 41524
rect 3668 41468 4172 41524
rect 4228 41468 4238 41524
rect 5058 41468 5068 41524
rect 5124 41468 5628 41524
rect 5684 41468 5694 41524
rect 7074 41468 7084 41524
rect 7140 41468 7756 41524
rect 7812 41468 7822 41524
rect 8652 41468 9548 41524
rect 9604 41468 11788 41524
rect 12786 41468 12796 41524
rect 12852 41468 16772 41524
rect 16930 41468 16940 41524
rect 16996 41468 19516 41524
rect 19572 41468 19582 41524
rect 23202 41468 23212 41524
rect 23268 41468 23884 41524
rect 23940 41468 23950 41524
rect 28802 41468 28812 41524
rect 28868 41468 30268 41524
rect 30324 41468 30334 41524
rect 30482 41468 30492 41524
rect 30548 41468 31276 41524
rect 31332 41468 31342 41524
rect 34710 41468 34748 41524
rect 34804 41468 34814 41524
rect 35858 41468 35868 41524
rect 35924 41468 36764 41524
rect 36820 41468 38108 41524
rect 38164 41468 38174 41524
rect 40460 41468 42364 41524
rect 42420 41468 42430 41524
rect 42914 41468 42924 41524
rect 42980 41468 44100 41524
rect 45378 41468 45388 41524
rect 45444 41468 45836 41524
rect 45892 41468 48860 41524
rect 48916 41468 48926 41524
rect 49970 41468 49980 41524
rect 50036 41468 50148 41524
rect 50372 41468 51548 41524
rect 51604 41468 51614 41524
rect 52882 41468 52892 41524
rect 52948 41468 57456 41524
rect 0 41440 112 41468
rect 44044 41412 44100 41468
rect 50372 41412 50428 41468
rect 57344 41440 57456 41468
rect 690 41356 700 41412
rect 756 41356 6972 41412
rect 7028 41356 7038 41412
rect 8082 41356 8092 41412
rect 8148 41356 19292 41412
rect 19348 41356 19358 41412
rect 22316 41356 26908 41412
rect 29810 41356 29820 41412
rect 29876 41356 33404 41412
rect 33460 41356 33470 41412
rect 34626 41356 34636 41412
rect 34692 41356 40236 41412
rect 40292 41356 40302 41412
rect 40898 41356 40908 41412
rect 40964 41356 42588 41412
rect 42644 41356 42654 41412
rect 42802 41356 42812 41412
rect 42868 41356 43820 41412
rect 43876 41356 43886 41412
rect 44044 41356 48972 41412
rect 49028 41356 49038 41412
rect 49410 41356 49420 41412
rect 49476 41356 50428 41412
rect 50754 41356 50764 41412
rect 50820 41356 54908 41412
rect 54964 41356 54974 41412
rect 55346 41356 55356 41412
rect 55412 41356 55916 41412
rect 55972 41356 55982 41412
rect 56326 41356 56364 41412
rect 56420 41356 56430 41412
rect 2380 41244 4508 41300
rect 4564 41244 4574 41300
rect 4834 41244 4844 41300
rect 4900 41244 8372 41300
rect 8530 41244 8540 41300
rect 8596 41244 9660 41300
rect 9716 41244 10332 41300
rect 10388 41244 10398 41300
rect 10658 41244 10668 41300
rect 10724 41244 13580 41300
rect 13636 41244 13646 41300
rect 13794 41244 13804 41300
rect 13860 41244 14364 41300
rect 14420 41244 14812 41300
rect 14868 41244 14878 41300
rect 15250 41244 15260 41300
rect 15316 41244 15596 41300
rect 15652 41244 15662 41300
rect 16034 41244 16044 41300
rect 16100 41244 17388 41300
rect 17444 41244 17454 41300
rect 17714 41244 17724 41300
rect 17780 41244 18508 41300
rect 18564 41244 18574 41300
rect 19282 41244 19292 41300
rect 19348 41244 22092 41300
rect 22148 41244 22158 41300
rect 1698 41132 1708 41188
rect 1764 41132 2044 41188
rect 2100 41132 2110 41188
rect 0 41076 112 41104
rect 0 41020 1708 41076
rect 1764 41020 1774 41076
rect 0 40992 112 41020
rect 2380 40964 2436 41244
rect 8316 41188 8372 41244
rect 22316 41188 22372 41356
rect 26852 41300 26908 41356
rect 22754 41244 22764 41300
rect 22820 41244 26572 41300
rect 26628 41244 26638 41300
rect 26852 41244 31444 41300
rect 32946 41244 32956 41300
rect 33012 41244 34076 41300
rect 34132 41244 34142 41300
rect 34402 41244 34412 41300
rect 34468 41244 35308 41300
rect 35364 41244 35980 41300
rect 36036 41244 36046 41300
rect 38994 41244 39004 41300
rect 39060 41244 41916 41300
rect 41972 41244 41982 41300
rect 43138 41244 43148 41300
rect 43204 41244 48076 41300
rect 48132 41244 48142 41300
rect 48738 41244 48748 41300
rect 48804 41244 49700 41300
rect 49858 41244 49868 41300
rect 49924 41244 51324 41300
rect 51380 41244 51390 41300
rect 52658 41244 52668 41300
rect 52724 41244 53564 41300
rect 53620 41244 53630 41300
rect 54002 41244 54012 41300
rect 54068 41244 54348 41300
rect 54404 41244 54414 41300
rect 31388 41188 31444 41244
rect 49644 41188 49700 41244
rect 2594 41132 2604 41188
rect 2660 41132 5068 41188
rect 5124 41132 5134 41188
rect 5506 41132 5516 41188
rect 5572 41132 5628 41188
rect 5684 41132 5694 41188
rect 6738 41132 6748 41188
rect 6804 41132 7308 41188
rect 7364 41132 7374 41188
rect 8316 41132 8428 41188
rect 8484 41132 8494 41188
rect 8754 41132 8764 41188
rect 8820 41132 9324 41188
rect 9380 41132 9390 41188
rect 9762 41132 9772 41188
rect 9828 41132 9996 41188
rect 10052 41132 10062 41188
rect 12002 41132 12012 41188
rect 12068 41132 12796 41188
rect 12852 41132 12862 41188
rect 13458 41132 13468 41188
rect 13524 41132 22372 41188
rect 22978 41132 22988 41188
rect 23044 41132 23660 41188
rect 23716 41132 23726 41188
rect 25218 41132 25228 41188
rect 25284 41132 26236 41188
rect 26292 41132 26302 41188
rect 26562 41132 26572 41188
rect 26628 41132 28140 41188
rect 28196 41132 28206 41188
rect 28364 41132 29036 41188
rect 29092 41132 29102 41188
rect 29474 41132 29484 41188
rect 29540 41132 30716 41188
rect 30772 41132 30782 41188
rect 30930 41132 30940 41188
rect 30996 41132 31034 41188
rect 31388 41132 36540 41188
rect 36596 41132 36606 41188
rect 38210 41132 38220 41188
rect 38276 41132 40572 41188
rect 40628 41132 40638 41188
rect 43586 41132 43596 41188
rect 43652 41132 44156 41188
rect 44212 41132 44940 41188
rect 44996 41132 45006 41188
rect 45154 41132 45164 41188
rect 45220 41132 46956 41188
rect 47012 41132 47022 41188
rect 48290 41132 48300 41188
rect 48356 41132 49308 41188
rect 49364 41132 49374 41188
rect 49644 41132 50876 41188
rect 50932 41132 50942 41188
rect 51090 41132 51100 41188
rect 51156 41132 51772 41188
rect 51828 41132 51838 41188
rect 52322 41132 52332 41188
rect 52388 41132 52892 41188
rect 52948 41132 55356 41188
rect 55412 41132 55422 41188
rect 55794 41132 55804 41188
rect 55860 41132 55916 41188
rect 55972 41132 55982 41188
rect 56998 41132 57036 41188
rect 57092 41132 57102 41188
rect 5628 41076 5684 41132
rect 28364 41076 28420 41132
rect 57344 41076 57456 41104
rect 2818 41020 2828 41076
rect 2884 41020 3388 41076
rect 3444 41020 3836 41076
rect 3892 41020 3902 41076
rect 4246 41020 4284 41076
rect 4340 41020 4350 41076
rect 5628 41020 10332 41076
rect 10388 41020 10398 41076
rect 13682 41020 13692 41076
rect 13748 41020 18844 41076
rect 18900 41020 18910 41076
rect 19506 41020 19516 41076
rect 19572 41020 23436 41076
rect 23492 41020 23502 41076
rect 24210 41020 24220 41076
rect 24276 41020 28420 41076
rect 28914 41020 28924 41076
rect 28980 41020 31220 41076
rect 31378 41020 31388 41076
rect 31444 41020 33628 41076
rect 33684 41020 33694 41076
rect 33954 41020 33964 41076
rect 34020 41020 35196 41076
rect 35252 41020 35262 41076
rect 35970 41020 35980 41076
rect 36036 41020 37548 41076
rect 37604 41020 37614 41076
rect 38434 41020 38444 41076
rect 38500 41020 42252 41076
rect 42308 41020 42318 41076
rect 43148 41020 49756 41076
rect 49812 41020 49822 41076
rect 49970 41020 49980 41076
rect 50036 41020 50204 41076
rect 50260 41020 50270 41076
rect 50418 41020 50428 41076
rect 50484 41020 52220 41076
rect 52276 41020 52286 41076
rect 52546 41020 52556 41076
rect 52612 41020 53452 41076
rect 53508 41020 53518 41076
rect 56578 41020 56588 41076
rect 56644 41020 57456 41076
rect 28924 40964 28980 41020
rect 31164 40964 31220 41020
rect 2370 40908 2380 40964
rect 2436 40908 2446 40964
rect 3602 40908 3612 40964
rect 3668 40908 7756 40964
rect 7812 40908 7822 40964
rect 8092 40908 8876 40964
rect 8932 40908 8942 40964
rect 9090 40908 9100 40964
rect 9156 40908 9548 40964
rect 9604 40908 9614 40964
rect 11330 40908 11340 40964
rect 11396 40908 14140 40964
rect 14196 40908 14206 40964
rect 16790 40908 16828 40964
rect 16884 40908 16894 40964
rect 17154 40908 17164 40964
rect 17220 40908 17836 40964
rect 17892 40908 17902 40964
rect 18610 40908 18620 40964
rect 18676 40908 22316 40964
rect 22372 40908 22382 40964
rect 23874 40908 23884 40964
rect 23940 40908 25340 40964
rect 25396 40908 25406 40964
rect 26226 40908 26236 40964
rect 26292 40908 28980 40964
rect 29810 40908 29820 40964
rect 29876 40908 29932 40964
rect 29988 40908 30940 40964
rect 30996 40908 31006 40964
rect 31164 40908 33852 40964
rect 33908 40908 33918 40964
rect 35410 40908 35420 40964
rect 35476 40908 36764 40964
rect 36820 40908 36830 40964
rect 39554 40908 39564 40964
rect 39620 40908 40572 40964
rect 40628 40908 40638 40964
rect 8092 40852 8148 40908
rect 3378 40796 3388 40852
rect 3444 40796 3500 40852
rect 3556 40796 3566 40852
rect 4162 40796 4172 40852
rect 4228 40796 4732 40852
rect 4788 40796 4798 40852
rect 4946 40796 4956 40852
rect 5012 40796 6188 40852
rect 6244 40796 6254 40852
rect 6514 40796 6524 40852
rect 6580 40796 6972 40852
rect 7028 40796 8148 40852
rect 8306 40796 8316 40852
rect 8372 40796 18956 40852
rect 19012 40796 19022 40852
rect 24434 40796 24444 40852
rect 24500 40796 34636 40852
rect 34692 40796 34702 40852
rect 35074 40796 35084 40852
rect 35140 40796 37548 40852
rect 37604 40796 37614 40852
rect 37762 40796 37772 40852
rect 37828 40796 38668 40852
rect 39442 40796 39452 40852
rect 39508 40796 40236 40852
rect 40292 40796 42476 40852
rect 42532 40796 42542 40852
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 38612 40740 38668 40796
rect 43148 40740 43204 41020
rect 57344 40992 57456 41020
rect 43362 40908 43372 40964
rect 43428 40908 45500 40964
rect 45556 40908 45566 40964
rect 45938 40908 45948 40964
rect 46004 40908 47964 40964
rect 48020 40908 48030 40964
rect 48402 40908 48412 40964
rect 48468 40908 48972 40964
rect 49028 40908 49038 40964
rect 50306 40908 50316 40964
rect 50372 40908 50428 40964
rect 50484 40908 50494 40964
rect 50652 40908 52444 40964
rect 52500 40908 52510 40964
rect 54338 40908 54348 40964
rect 54404 40908 55804 40964
rect 55860 40908 55870 40964
rect 50652 40852 50708 40908
rect 44146 40796 44156 40852
rect 44212 40796 45276 40852
rect 45332 40796 45342 40852
rect 46834 40796 46844 40852
rect 46900 40796 48748 40852
rect 48804 40796 48814 40852
rect 48972 40796 50708 40852
rect 50764 40796 53340 40852
rect 53396 40796 53406 40852
rect 43794 40740 43804 40796
rect 43860 40740 43908 40796
rect 43964 40740 44012 40796
rect 44068 40740 44078 40796
rect 48972 40740 49028 40796
rect 50764 40740 50820 40796
rect 1922 40684 1932 40740
rect 1988 40684 2156 40740
rect 2212 40684 2222 40740
rect 4162 40684 4172 40740
rect 4228 40684 5180 40740
rect 5236 40684 5246 40740
rect 5394 40684 5404 40740
rect 5460 40684 12236 40740
rect 12292 40684 12302 40740
rect 12450 40684 12460 40740
rect 12516 40684 12554 40740
rect 13346 40684 13356 40740
rect 13412 40684 13916 40740
rect 13972 40684 13982 40740
rect 14130 40684 14140 40740
rect 14196 40684 16268 40740
rect 16324 40684 16334 40740
rect 18834 40684 18844 40740
rect 18900 40684 21980 40740
rect 22036 40684 22316 40740
rect 22372 40684 22382 40740
rect 28690 40684 28700 40740
rect 28756 40684 33964 40740
rect 34020 40684 34030 40740
rect 34262 40684 34300 40740
rect 34356 40684 35196 40740
rect 35252 40684 35262 40740
rect 35634 40684 35644 40740
rect 35700 40684 37940 40740
rect 38612 40684 43204 40740
rect 45154 40684 45164 40740
rect 45220 40684 47740 40740
rect 47796 40684 47806 40740
rect 48962 40684 48972 40740
rect 49028 40684 49038 40740
rect 49196 40684 50820 40740
rect 50978 40684 50988 40740
rect 51044 40684 52220 40740
rect 52276 40684 52444 40740
rect 52500 40684 52510 40740
rect 0 40628 112 40656
rect 37884 40628 37940 40684
rect 49196 40628 49252 40684
rect 57344 40628 57456 40656
rect 0 40572 20972 40628
rect 21028 40572 21038 40628
rect 21634 40572 21644 40628
rect 21700 40572 37660 40628
rect 37716 40572 37726 40628
rect 37884 40572 49252 40628
rect 49858 40572 49868 40628
rect 49924 40572 49934 40628
rect 50530 40572 50540 40628
rect 50596 40572 57456 40628
rect 0 40544 112 40572
rect 49868 40516 49924 40572
rect 57344 40544 57456 40572
rect 1138 40460 1148 40516
rect 1204 40460 3500 40516
rect 3556 40460 3566 40516
rect 4060 40460 5740 40516
rect 5796 40460 5806 40516
rect 6290 40460 6300 40516
rect 6356 40460 9604 40516
rect 10210 40460 10220 40516
rect 10276 40460 12684 40516
rect 12740 40460 12750 40516
rect 13244 40460 13580 40516
rect 13636 40460 13646 40516
rect 14578 40460 14588 40516
rect 14644 40460 22428 40516
rect 22484 40460 22494 40516
rect 22754 40460 22764 40516
rect 22820 40460 23212 40516
rect 23268 40460 23278 40516
rect 23762 40460 23772 40516
rect 23828 40460 28700 40516
rect 28756 40460 28766 40516
rect 29026 40460 29036 40516
rect 29092 40460 31388 40516
rect 31444 40460 31454 40516
rect 32050 40460 32060 40516
rect 32116 40460 32956 40516
rect 33012 40460 33022 40516
rect 33282 40460 33292 40516
rect 33348 40460 35644 40516
rect 35700 40460 36092 40516
rect 36148 40460 36158 40516
rect 37538 40460 37548 40516
rect 37604 40460 42588 40516
rect 42644 40460 42654 40516
rect 42802 40460 42812 40516
rect 42868 40460 44268 40516
rect 44324 40460 44334 40516
rect 44482 40460 44492 40516
rect 44548 40460 46620 40516
rect 46676 40460 46686 40516
rect 48514 40460 48524 40516
rect 48580 40460 49924 40516
rect 50194 40460 50204 40516
rect 50260 40460 51996 40516
rect 52052 40460 52062 40516
rect 53218 40460 53228 40516
rect 53284 40460 53340 40516
rect 53396 40460 55916 40516
rect 55972 40460 55982 40516
rect 4060 40404 4116 40460
rect 9548 40404 9604 40460
rect 1586 40348 1596 40404
rect 1652 40348 2828 40404
rect 2884 40348 2894 40404
rect 3042 40348 3052 40404
rect 3108 40348 4116 40404
rect 4274 40348 4284 40404
rect 4340 40348 5516 40404
rect 5572 40348 5582 40404
rect 8194 40348 8204 40404
rect 8260 40348 9324 40404
rect 9380 40348 9390 40404
rect 9548 40348 10556 40404
rect 10612 40348 10622 40404
rect 11890 40348 11900 40404
rect 11956 40348 12236 40404
rect 12292 40348 12302 40404
rect 13244 40292 13300 40460
rect 1110 40236 1148 40292
rect 1204 40236 1214 40292
rect 1708 40236 12460 40292
rect 12516 40236 12526 40292
rect 13010 40236 13020 40292
rect 13076 40236 13300 40292
rect 13356 40348 13468 40404
rect 13524 40348 13534 40404
rect 14466 40348 14476 40404
rect 14532 40348 15708 40404
rect 15764 40348 16940 40404
rect 16996 40348 17006 40404
rect 19170 40348 19180 40404
rect 19236 40348 19516 40404
rect 19572 40348 19582 40404
rect 19954 40348 19964 40404
rect 20020 40348 21420 40404
rect 21476 40348 22092 40404
rect 22148 40348 23100 40404
rect 23156 40348 23436 40404
rect 23492 40348 23502 40404
rect 25106 40348 25116 40404
rect 25172 40348 26236 40404
rect 26292 40348 26302 40404
rect 27010 40348 27020 40404
rect 27076 40348 33628 40404
rect 33684 40348 33694 40404
rect 33842 40348 33852 40404
rect 33908 40348 33918 40404
rect 35074 40348 35084 40404
rect 35140 40348 36652 40404
rect 36708 40348 36718 40404
rect 38770 40348 38780 40404
rect 38836 40348 39564 40404
rect 39620 40348 39630 40404
rect 41458 40348 41468 40404
rect 41524 40348 42028 40404
rect 42084 40348 42094 40404
rect 43362 40348 43372 40404
rect 43428 40348 48076 40404
rect 48132 40348 48142 40404
rect 49410 40348 49420 40404
rect 49476 40348 49868 40404
rect 49924 40348 49934 40404
rect 50082 40348 50092 40404
rect 50148 40348 50988 40404
rect 51044 40348 51054 40404
rect 0 40180 112 40208
rect 1708 40180 1764 40236
rect 13356 40180 13412 40348
rect 33852 40292 33908 40348
rect 13570 40236 13580 40292
rect 13636 40236 14252 40292
rect 14308 40236 14318 40292
rect 16566 40236 16604 40292
rect 16660 40236 16670 40292
rect 18162 40236 18172 40292
rect 18228 40236 18844 40292
rect 18900 40236 18910 40292
rect 19730 40236 19740 40292
rect 19796 40236 19852 40292
rect 19908 40236 19918 40292
rect 21074 40236 21084 40292
rect 21140 40236 22652 40292
rect 22708 40236 22718 40292
rect 23538 40236 23548 40292
rect 23604 40236 24500 40292
rect 24854 40236 24892 40292
rect 24948 40236 24958 40292
rect 31378 40236 31388 40292
rect 31444 40236 33292 40292
rect 33348 40236 33358 40292
rect 33852 40236 34132 40292
rect 34934 40236 34972 40292
rect 35028 40236 35038 40292
rect 35746 40236 35756 40292
rect 35812 40236 36428 40292
rect 36484 40236 36988 40292
rect 37044 40236 37054 40292
rect 37426 40236 37436 40292
rect 37492 40236 39452 40292
rect 39508 40236 39518 40292
rect 40236 40236 48972 40292
rect 49028 40236 49038 40292
rect 49270 40236 49308 40292
rect 49364 40236 49374 40292
rect 53106 40236 53116 40292
rect 53172 40236 55356 40292
rect 55412 40236 55422 40292
rect 24444 40180 24500 40236
rect 34076 40180 34132 40236
rect 40236 40180 40292 40236
rect 57344 40180 57456 40208
rect 0 40124 1764 40180
rect 2706 40124 2716 40180
rect 2772 40124 5404 40180
rect 5460 40124 5470 40180
rect 5618 40124 5628 40180
rect 5684 40124 7420 40180
rect 7476 40124 7486 40180
rect 8204 40124 10668 40180
rect 10724 40124 10734 40180
rect 10882 40124 10892 40180
rect 10948 40124 11452 40180
rect 11508 40124 11518 40180
rect 13356 40124 13916 40180
rect 13972 40124 13982 40180
rect 15092 40124 15820 40180
rect 15876 40124 15886 40180
rect 16146 40124 16156 40180
rect 16212 40124 24220 40180
rect 24276 40124 24286 40180
rect 24444 40124 24948 40180
rect 26674 40124 26684 40180
rect 26740 40124 26908 40180
rect 26964 40124 26974 40180
rect 27458 40124 27468 40180
rect 27524 40124 28028 40180
rect 28084 40124 28094 40180
rect 28578 40124 28588 40180
rect 28644 40124 30492 40180
rect 30548 40124 30558 40180
rect 32722 40124 32732 40180
rect 32788 40124 33852 40180
rect 33908 40124 33918 40180
rect 34076 40124 35980 40180
rect 36036 40124 36046 40180
rect 37202 40124 37212 40180
rect 37268 40124 37884 40180
rect 37940 40124 37950 40180
rect 38994 40124 39004 40180
rect 39060 40124 40292 40180
rect 41570 40124 41580 40180
rect 41636 40124 44828 40180
rect 44884 40124 44894 40180
rect 45266 40124 45276 40180
rect 45332 40124 47628 40180
rect 47684 40124 47694 40180
rect 50418 40124 50428 40180
rect 50484 40124 51996 40180
rect 52052 40124 52062 40180
rect 53442 40124 53452 40180
rect 53508 40124 57456 40180
rect 0 40096 112 40124
rect 8204 40068 8260 40124
rect 15092 40068 15148 40124
rect 1362 40012 1372 40068
rect 1428 40012 4172 40068
rect 4228 40012 4238 40068
rect 6850 40012 6860 40068
rect 6916 40012 8260 40068
rect 8316 40012 15148 40068
rect 19058 40012 19068 40068
rect 19124 40012 19852 40068
rect 19908 40012 19918 40068
rect 20066 40012 20076 40068
rect 20132 40012 20972 40068
rect 21028 40012 21038 40068
rect 22754 40012 22764 40068
rect 22820 40012 23436 40068
rect 23492 40012 23502 40068
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 2258 39900 2268 39956
rect 2324 39900 2604 39956
rect 2660 39900 2670 39956
rect 3266 39900 3276 39956
rect 3332 39900 4172 39956
rect 4228 39900 4238 39956
rect 7270 39900 7308 39956
rect 7364 39900 7374 39956
rect 8316 39844 8372 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 24892 39956 24948 40124
rect 57344 40096 57456 40124
rect 32274 40012 32284 40068
rect 32340 40012 33068 40068
rect 33124 40012 33964 40068
rect 34020 40012 34030 40068
rect 34738 40012 34748 40068
rect 34804 40012 38444 40068
rect 38500 40012 38510 40068
rect 38612 40012 39228 40068
rect 39284 40012 39294 40068
rect 40002 40012 40012 40068
rect 40068 40012 40124 40068
rect 40180 40012 41020 40068
rect 41076 40012 41086 40068
rect 41234 40012 41244 40068
rect 41300 40012 44156 40068
rect 44212 40012 44222 40068
rect 45154 40012 45164 40068
rect 45220 40012 49756 40068
rect 49812 40012 49822 40068
rect 50418 40012 50428 40068
rect 50484 40012 51660 40068
rect 51716 40012 51726 40068
rect 38612 39956 38668 40012
rect 44454 39956 44464 40012
rect 44520 39956 44568 40012
rect 44624 39956 44672 40012
rect 44728 39956 44738 40012
rect 2034 39788 2044 39844
rect 2100 39788 8372 39844
rect 8428 39900 21028 39956
rect 22306 39900 22316 39956
rect 22372 39900 22540 39956
rect 22596 39900 22606 39956
rect 24892 39900 26796 39956
rect 26852 39900 26862 39956
rect 30818 39900 30828 39956
rect 30884 39900 38668 39956
rect 45378 39900 45388 39956
rect 45444 39900 47068 39956
rect 47124 39900 47134 39956
rect 47506 39900 47516 39956
rect 47572 39900 55692 39956
rect 55748 39900 55758 39956
rect 0 39732 112 39760
rect 8428 39732 8484 39900
rect 20972 39844 21028 39900
rect 8838 39788 8876 39844
rect 8932 39788 9212 39844
rect 9268 39788 9278 39844
rect 9538 39788 9548 39844
rect 9604 39788 10108 39844
rect 10164 39788 10174 39844
rect 10658 39788 10668 39844
rect 10724 39788 13020 39844
rect 13076 39788 13086 39844
rect 13346 39788 13356 39844
rect 13412 39788 16940 39844
rect 16996 39788 17006 39844
rect 20972 39788 35196 39844
rect 35252 39788 35262 39844
rect 35858 39788 35868 39844
rect 35924 39788 41580 39844
rect 41636 39788 41646 39844
rect 42242 39788 42252 39844
rect 42308 39788 45052 39844
rect 45108 39788 45118 39844
rect 45490 39788 45500 39844
rect 45556 39788 47180 39844
rect 47236 39788 47246 39844
rect 47730 39788 47740 39844
rect 47796 39788 52668 39844
rect 52724 39788 52892 39844
rect 52948 39788 52958 39844
rect 10108 39732 10164 39788
rect 57344 39732 57456 39760
rect 0 39676 8484 39732
rect 8540 39676 9492 39732
rect 9762 39676 9772 39732
rect 9828 39676 9884 39732
rect 9940 39676 9950 39732
rect 10108 39676 10668 39732
rect 10724 39676 10734 39732
rect 11778 39676 11788 39732
rect 11844 39676 11900 39732
rect 11956 39676 11966 39732
rect 13580 39676 14140 39732
rect 14196 39676 14206 39732
rect 14578 39676 14588 39732
rect 14644 39676 16268 39732
rect 16324 39676 16334 39732
rect 16706 39676 16716 39732
rect 16772 39676 18844 39732
rect 18900 39676 18910 39732
rect 23202 39676 23212 39732
rect 23268 39676 25228 39732
rect 25284 39676 25294 39732
rect 26226 39676 26236 39732
rect 26292 39676 26796 39732
rect 26852 39676 26862 39732
rect 34178 39676 34188 39732
rect 34244 39676 34524 39732
rect 34580 39676 34590 39732
rect 35410 39676 35420 39732
rect 35476 39676 38668 39732
rect 38724 39676 38734 39732
rect 39218 39676 39228 39732
rect 39284 39676 40236 39732
rect 40292 39676 40302 39732
rect 42578 39676 42588 39732
rect 42644 39676 45164 39732
rect 45220 39676 45230 39732
rect 47394 39676 47404 39732
rect 47460 39676 48188 39732
rect 48244 39676 48254 39732
rect 48524 39676 50316 39732
rect 50372 39676 50382 39732
rect 52546 39676 52556 39732
rect 52612 39676 54796 39732
rect 54852 39676 54862 39732
rect 57250 39676 57260 39732
rect 57316 39676 57456 39732
rect 0 39648 112 39676
rect 8540 39620 8596 39676
rect 1138 39564 1148 39620
rect 1204 39564 3052 39620
rect 3108 39564 3118 39620
rect 3266 39564 3276 39620
rect 3332 39564 5180 39620
rect 5236 39564 5246 39620
rect 5730 39564 5740 39620
rect 5796 39564 6636 39620
rect 6692 39564 8596 39620
rect 9436 39620 9492 39676
rect 13580 39620 13636 39676
rect 48524 39620 48580 39676
rect 57344 39648 57456 39676
rect 9436 39564 13636 39620
rect 14242 39564 14252 39620
rect 14308 39564 22540 39620
rect 22596 39564 24332 39620
rect 24388 39564 24398 39620
rect 26114 39564 26124 39620
rect 26180 39564 26684 39620
rect 26740 39564 27244 39620
rect 27300 39564 27310 39620
rect 30594 39564 30604 39620
rect 30660 39564 33628 39620
rect 33684 39564 33694 39620
rect 34066 39564 34076 39620
rect 34132 39564 35084 39620
rect 35140 39564 39284 39620
rect 42466 39564 42476 39620
rect 42532 39564 45724 39620
rect 45780 39564 45790 39620
rect 47618 39564 47628 39620
rect 47684 39564 48524 39620
rect 48580 39564 48590 39620
rect 48850 39564 48860 39620
rect 48916 39564 50988 39620
rect 51044 39564 53340 39620
rect 53396 39564 53406 39620
rect 53890 39564 53900 39620
rect 53956 39564 54348 39620
rect 54404 39564 54414 39620
rect 56018 39564 56028 39620
rect 56084 39564 56140 39620
rect 56196 39564 56206 39620
rect 39228 39508 39284 39564
rect 2370 39452 2380 39508
rect 2436 39452 3164 39508
rect 3220 39452 3230 39508
rect 3378 39452 3388 39508
rect 3444 39452 7980 39508
rect 8036 39452 8046 39508
rect 8194 39452 8204 39508
rect 8260 39452 9548 39508
rect 9604 39452 9614 39508
rect 12562 39452 12572 39508
rect 12628 39452 13020 39508
rect 13076 39452 13086 39508
rect 13346 39452 13356 39508
rect 13412 39452 13468 39508
rect 13524 39452 13534 39508
rect 14102 39452 14140 39508
rect 14196 39452 14206 39508
rect 15250 39452 15260 39508
rect 15316 39452 16044 39508
rect 16100 39452 16110 39508
rect 16818 39452 16828 39508
rect 16884 39452 23772 39508
rect 23828 39452 23838 39508
rect 24098 39452 24108 39508
rect 24164 39452 26068 39508
rect 26338 39452 26348 39508
rect 26404 39452 26460 39508
rect 26516 39452 26526 39508
rect 26674 39452 26684 39508
rect 26740 39452 35308 39508
rect 35364 39452 35374 39508
rect 35634 39452 35644 39508
rect 35700 39452 36204 39508
rect 36260 39452 36270 39508
rect 39228 39452 40124 39508
rect 40180 39452 40190 39508
rect 41122 39452 41132 39508
rect 41188 39452 42252 39508
rect 42308 39452 42318 39508
rect 43698 39452 43708 39508
rect 43764 39452 44716 39508
rect 44772 39452 44782 39508
rect 45938 39452 45948 39508
rect 46004 39452 54628 39508
rect 55570 39452 55580 39508
rect 55636 39452 56476 39508
rect 56532 39452 56542 39508
rect 26012 39396 26068 39452
rect 3332 39340 24276 39396
rect 25218 39340 25228 39396
rect 25284 39340 25676 39396
rect 25732 39340 25742 39396
rect 26012 39340 28588 39396
rect 28644 39340 28654 39396
rect 31266 39340 31276 39396
rect 31332 39340 44548 39396
rect 45042 39340 45052 39396
rect 45108 39340 46508 39396
rect 46564 39340 46574 39396
rect 47058 39340 47068 39396
rect 47124 39340 48524 39396
rect 48580 39340 48590 39396
rect 51090 39340 51100 39396
rect 51156 39340 52444 39396
rect 52500 39340 52510 39396
rect 52658 39340 52668 39396
rect 52724 39340 53116 39396
rect 53172 39340 53182 39396
rect 53750 39340 53788 39396
rect 53844 39340 53854 39396
rect 0 39284 112 39312
rect 3332 39284 3388 39340
rect 24220 39284 24276 39340
rect 44492 39284 44548 39340
rect 54572 39284 54628 39452
rect 57344 39284 57456 39312
rect 0 39228 3388 39284
rect 4162 39228 4172 39284
rect 4228 39228 10892 39284
rect 10948 39228 10958 39284
rect 11778 39228 11788 39284
rect 11844 39228 12572 39284
rect 12628 39228 12638 39284
rect 13122 39228 13132 39284
rect 13188 39228 15932 39284
rect 15988 39228 15998 39284
rect 24220 39228 30716 39284
rect 30772 39228 30782 39284
rect 34850 39228 34860 39284
rect 34916 39228 37660 39284
rect 37716 39228 37726 39284
rect 38546 39228 38556 39284
rect 38612 39228 38892 39284
rect 38948 39228 39676 39284
rect 39732 39228 39742 39284
rect 40114 39228 40124 39284
rect 40180 39228 41356 39284
rect 41412 39228 41422 39284
rect 44492 39228 50428 39284
rect 50484 39228 50494 39284
rect 50642 39228 50652 39284
rect 50708 39228 50764 39284
rect 50820 39228 50830 39284
rect 50988 39228 52444 39284
rect 52500 39228 52510 39284
rect 53554 39228 53564 39284
rect 53620 39228 54348 39284
rect 54404 39228 54414 39284
rect 54572 39228 57456 39284
rect 0 39200 112 39228
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 43794 39172 43804 39228
rect 43860 39172 43908 39228
rect 43964 39172 44012 39228
rect 44068 39172 44078 39228
rect 50988 39172 51044 39228
rect 57344 39200 57456 39228
rect 242 39116 252 39172
rect 308 39116 1036 39172
rect 1092 39116 1102 39172
rect 4386 39116 4396 39172
rect 4452 39116 4844 39172
rect 4900 39116 4910 39172
rect 5394 39116 5404 39172
rect 5460 39116 6748 39172
rect 6804 39116 6814 39172
rect 8530 39116 8540 39172
rect 8596 39116 11900 39172
rect 11956 39116 11966 39172
rect 12236 39116 12460 39172
rect 12516 39116 13244 39172
rect 13300 39116 13310 39172
rect 14914 39116 14924 39172
rect 14980 39116 15820 39172
rect 15876 39116 15886 39172
rect 16594 39116 16604 39172
rect 16660 39116 23548 39172
rect 23604 39116 23614 39172
rect 26226 39116 26236 39172
rect 26292 39116 26460 39172
rect 26516 39116 26526 39172
rect 26674 39116 26684 39172
rect 26740 39116 27020 39172
rect 27076 39116 27086 39172
rect 28690 39116 28700 39172
rect 28756 39116 29036 39172
rect 29092 39116 29102 39172
rect 33282 39116 33292 39172
rect 33348 39116 35868 39172
rect 35924 39116 35934 39172
rect 37314 39116 37324 39172
rect 37380 39116 39620 39172
rect 39778 39116 39788 39172
rect 39844 39116 41916 39172
rect 41972 39116 41982 39172
rect 42578 39116 42588 39172
rect 42644 39116 43484 39172
rect 43540 39116 43550 39172
rect 44370 39116 44380 39172
rect 44436 39116 45388 39172
rect 45444 39116 45454 39172
rect 45602 39116 45612 39172
rect 45668 39116 49140 39172
rect 49298 39116 49308 39172
rect 49364 39116 49868 39172
rect 49924 39116 49934 39172
rect 50194 39116 50204 39172
rect 50260 39116 51044 39172
rect 51202 39116 51212 39172
rect 51268 39116 52556 39172
rect 52612 39116 52622 39172
rect 52770 39116 52780 39172
rect 52836 39116 53116 39172
rect 53172 39116 55244 39172
rect 55300 39116 55310 39172
rect 1810 39004 1820 39060
rect 1876 39004 2044 39060
rect 2100 39004 2110 39060
rect 3490 39004 3500 39060
rect 3556 39004 6188 39060
rect 6244 39004 6254 39060
rect 7970 39004 7980 39060
rect 8036 39004 11788 39060
rect 11844 39004 11854 39060
rect 12236 38948 12292 39116
rect 12450 39004 12460 39060
rect 12516 39004 25228 39060
rect 25284 39004 25294 39060
rect 25666 39004 25676 39060
rect 25732 39004 39508 39060
rect 466 38892 476 38948
rect 532 38892 1260 38948
rect 1316 38892 2492 38948
rect 2548 38892 2558 38948
rect 3266 38892 3276 38948
rect 3332 38892 9884 38948
rect 9940 38892 9950 38948
rect 10108 38892 12292 38948
rect 12450 38892 12460 38948
rect 12516 38892 16604 38948
rect 16660 38892 16670 38948
rect 21298 38892 21308 38948
rect 21364 38892 23548 38948
rect 23604 38892 25116 38948
rect 25172 38892 25182 38948
rect 25442 38892 25452 38948
rect 25508 38892 28868 38948
rect 29474 38892 29484 38948
rect 29540 38892 30156 38948
rect 30212 38892 30222 38948
rect 31378 38892 31388 38948
rect 31444 38892 34076 38948
rect 34132 38892 34142 38948
rect 35522 38892 35532 38948
rect 35588 38892 35756 38948
rect 35812 38892 35822 38948
rect 36726 38892 36764 38948
rect 36820 38892 36988 38948
rect 37044 38892 37054 38948
rect 37874 38892 37884 38948
rect 37940 38892 38444 38948
rect 38500 38892 38510 38948
rect 0 38836 112 38864
rect 10108 38836 10164 38892
rect 28812 38836 28868 38892
rect 38612 38836 38668 38948
rect 38724 38892 38734 38948
rect 0 38780 700 38836
rect 756 38780 766 38836
rect 2146 38780 2156 38836
rect 2212 38780 3836 38836
rect 3892 38780 3902 38836
rect 4050 38780 4060 38836
rect 4116 38780 4284 38836
rect 4340 38780 4350 38836
rect 4946 38780 4956 38836
rect 5012 38780 5068 38836
rect 5124 38780 5134 38836
rect 5282 38780 5292 38836
rect 5348 38780 7532 38836
rect 7588 38780 7598 38836
rect 7970 38780 7980 38836
rect 8036 38780 8204 38836
rect 8260 38780 8270 38836
rect 8418 38780 8428 38836
rect 8484 38780 10164 38836
rect 10294 38780 10332 38836
rect 10388 38780 10398 38836
rect 10770 38780 10780 38836
rect 10836 38780 12684 38836
rect 12740 38780 12750 38836
rect 12898 38780 12908 38836
rect 12964 38780 13132 38836
rect 13188 38780 13198 38836
rect 14578 38780 14588 38836
rect 14644 38780 14924 38836
rect 14980 38780 14990 38836
rect 15260 38780 23772 38836
rect 23828 38780 23838 38836
rect 23986 38780 23996 38836
rect 24052 38780 25116 38836
rect 25172 38780 25182 38836
rect 26226 38780 26236 38836
rect 26292 38780 28588 38836
rect 28644 38780 28654 38836
rect 28812 38780 36092 38836
rect 36148 38780 36158 38836
rect 36316 38780 38668 38836
rect 39452 38836 39508 39004
rect 39564 38948 39620 39116
rect 49084 39060 49140 39116
rect 40338 39004 40348 39060
rect 40404 39004 47180 39060
rect 47236 39004 47246 39060
rect 49084 39004 50092 39060
rect 50148 39004 50158 39060
rect 50418 39004 50428 39060
rect 50484 39004 50876 39060
rect 50932 39004 50942 39060
rect 51874 39004 51884 39060
rect 51940 39004 53340 39060
rect 53396 39004 53406 39060
rect 54226 39004 54236 39060
rect 54292 39004 55804 39060
rect 55860 39004 55870 39060
rect 39564 38892 39676 38948
rect 39732 38892 40348 38948
rect 40404 38892 40796 38948
rect 40852 38892 40862 38948
rect 41020 38892 50092 38948
rect 50148 38892 50158 38948
rect 50754 38892 50764 38948
rect 50820 38892 52220 38948
rect 52276 38892 53452 38948
rect 53508 38892 53676 38948
rect 53732 38892 53742 38948
rect 54562 38892 54572 38948
rect 54628 38892 55692 38948
rect 55748 38892 55758 38948
rect 41020 38836 41076 38892
rect 57344 38836 57456 38864
rect 39452 38780 41076 38836
rect 42018 38780 42028 38836
rect 42084 38780 45948 38836
rect 46004 38780 46014 38836
rect 46386 38780 46396 38836
rect 46452 38780 46844 38836
rect 46900 38780 46910 38836
rect 47506 38780 47516 38836
rect 47572 38780 50204 38836
rect 50260 38780 50270 38836
rect 50418 38780 50428 38836
rect 50484 38780 52444 38836
rect 52500 38780 52510 38836
rect 54450 38780 54460 38836
rect 54516 38780 55580 38836
rect 55636 38780 55646 38836
rect 55916 38780 57456 38836
rect 0 38752 112 38780
rect 15260 38724 15316 38780
rect 36316 38724 36372 38780
rect 55916 38724 55972 38780
rect 57344 38752 57456 38780
rect 690 38668 700 38724
rect 756 38668 1708 38724
rect 1764 38668 2940 38724
rect 2996 38668 3006 38724
rect 3836 38668 4732 38724
rect 4788 38668 4798 38724
rect 4946 38668 4956 38724
rect 5012 38668 5180 38724
rect 5236 38668 5246 38724
rect 7858 38668 7868 38724
rect 7924 38668 8260 38724
rect 8418 38668 8428 38724
rect 8484 38668 9212 38724
rect 9268 38668 9278 38724
rect 9538 38668 9548 38724
rect 9604 38668 9772 38724
rect 9828 38668 9838 38724
rect 10770 38668 10780 38724
rect 10836 38668 11004 38724
rect 11060 38668 14588 38724
rect 14644 38668 14654 38724
rect 15148 38668 15316 38724
rect 18162 38668 18172 38724
rect 18228 38668 18844 38724
rect 18900 38668 21644 38724
rect 21700 38668 21710 38724
rect 23314 38668 23324 38724
rect 23380 38668 26908 38724
rect 26964 38668 26974 38724
rect 29222 38668 29260 38724
rect 29316 38668 29820 38724
rect 29876 38668 29886 38724
rect 31154 38668 31164 38724
rect 31220 38668 33180 38724
rect 33236 38668 33246 38724
rect 33506 38668 33516 38724
rect 33572 38668 33964 38724
rect 34020 38668 34636 38724
rect 34692 38668 34702 38724
rect 34860 38668 36372 38724
rect 38434 38668 38444 38724
rect 38500 38668 40012 38724
rect 40068 38668 40078 38724
rect 41906 38668 41916 38724
rect 41972 38668 43932 38724
rect 43988 38668 44380 38724
rect 44436 38668 44446 38724
rect 44706 38668 44716 38724
rect 44772 38668 45164 38724
rect 45220 38668 45230 38724
rect 46050 38668 46060 38724
rect 46116 38668 46956 38724
rect 47012 38668 47022 38724
rect 47282 38668 47292 38724
rect 47348 38668 48076 38724
rect 48132 38668 48142 38724
rect 48290 38668 48300 38724
rect 48356 38668 50652 38724
rect 50708 38668 50718 38724
rect 52108 38668 53564 38724
rect 53620 38668 53630 38724
rect 54338 38668 54348 38724
rect 54404 38668 55972 38724
rect 56690 38668 56700 38724
rect 56756 38668 56812 38724
rect 56868 38668 56878 38724
rect 3836 38612 3892 38668
rect 8204 38612 8260 38668
rect 15148 38612 15204 38668
rect 2380 38556 3892 38612
rect 4284 38556 7140 38612
rect 7298 38556 7308 38612
rect 7364 38556 7756 38612
rect 7812 38556 7822 38612
rect 8204 38556 8988 38612
rect 9044 38556 9054 38612
rect 10882 38556 10892 38612
rect 10948 38556 15204 38612
rect 15362 38556 15372 38612
rect 15428 38556 15596 38612
rect 15652 38556 15662 38612
rect 18498 38556 18508 38612
rect 18564 38556 19292 38612
rect 19348 38556 23996 38612
rect 24052 38556 24062 38612
rect 24220 38556 25452 38612
rect 25508 38556 25518 38612
rect 27794 38556 27804 38612
rect 27860 38556 29708 38612
rect 29764 38556 29774 38612
rect 30818 38556 30828 38612
rect 30884 38556 31276 38612
rect 31332 38556 31342 38612
rect 31490 38556 31500 38612
rect 31556 38556 31836 38612
rect 31892 38556 31948 38612
rect 32004 38556 32014 38612
rect 33506 38556 33516 38612
rect 33572 38556 34076 38612
rect 34132 38556 34142 38612
rect 2380 38500 2436 38556
rect 2370 38444 2380 38500
rect 2436 38444 2446 38500
rect 0 38388 112 38416
rect 4284 38388 4340 38556
rect 7084 38500 7140 38556
rect 24220 38500 24276 38556
rect 4834 38444 4844 38500
rect 4900 38444 6860 38500
rect 6916 38444 6926 38500
rect 7084 38444 9548 38500
rect 9604 38444 9614 38500
rect 13570 38444 13580 38500
rect 13636 38444 14252 38500
rect 14308 38444 14318 38500
rect 14578 38444 14588 38500
rect 14644 38444 21252 38500
rect 23762 38444 23772 38500
rect 23828 38444 24276 38500
rect 25442 38444 25452 38500
rect 25508 38444 27972 38500
rect 28130 38444 28140 38500
rect 28196 38444 30156 38500
rect 30212 38444 33516 38500
rect 33572 38444 33582 38500
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 21196 38388 21252 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 27916 38388 27972 38444
rect 34860 38388 34916 38668
rect 52108 38612 52164 38668
rect 39666 38556 39676 38612
rect 39732 38556 42476 38612
rect 42532 38556 42542 38612
rect 43036 38556 52164 38612
rect 52882 38556 52892 38612
rect 52948 38556 53228 38612
rect 53284 38556 53294 38612
rect 54646 38556 54684 38612
rect 54740 38556 55244 38612
rect 55300 38556 55310 38612
rect 55570 38556 55580 38612
rect 55636 38556 56588 38612
rect 56644 38556 56654 38612
rect 43036 38500 43092 38556
rect 35186 38444 35196 38500
rect 35252 38444 41356 38500
rect 41412 38444 41422 38500
rect 41906 38444 41916 38500
rect 41972 38444 43092 38500
rect 44930 38444 44940 38500
rect 44996 38444 47852 38500
rect 47908 38444 47918 38500
rect 51314 38444 51324 38500
rect 51380 38444 54796 38500
rect 54852 38444 54862 38500
rect 56690 38444 56700 38500
rect 56756 38444 57036 38500
rect 57092 38444 57102 38500
rect 44454 38388 44464 38444
rect 44520 38388 44568 38444
rect 44624 38388 44672 38444
rect 44728 38388 44738 38444
rect 57344 38388 57456 38416
rect 0 38332 252 38388
rect 308 38332 318 38388
rect 3602 38332 3612 38388
rect 3668 38332 4340 38388
rect 5058 38332 5068 38388
rect 5124 38332 11340 38388
rect 11396 38332 11406 38388
rect 11900 38332 12684 38388
rect 12740 38332 12750 38388
rect 13794 38332 13804 38388
rect 13860 38332 14476 38388
rect 14532 38332 14542 38388
rect 15250 38332 15260 38388
rect 15316 38332 15372 38388
rect 15428 38332 15438 38388
rect 16258 38332 16268 38388
rect 16324 38332 20972 38388
rect 21028 38332 21038 38388
rect 21196 38332 24220 38388
rect 24276 38332 24286 38388
rect 25106 38332 25116 38388
rect 25172 38332 26236 38388
rect 26292 38332 26302 38388
rect 27916 38332 29372 38388
rect 29428 38332 29438 38388
rect 31042 38332 31052 38388
rect 31108 38332 33740 38388
rect 33796 38332 34916 38388
rect 35858 38332 35868 38388
rect 35924 38332 42140 38388
rect 42196 38332 42206 38388
rect 42924 38332 44268 38388
rect 44324 38332 44334 38388
rect 51538 38332 51548 38388
rect 51604 38332 54572 38388
rect 54628 38332 54638 38388
rect 56354 38332 56364 38388
rect 56420 38332 56588 38388
rect 56644 38332 56654 38388
rect 56802 38332 56812 38388
rect 56868 38332 57456 38388
rect 0 38304 112 38332
rect 11900 38276 11956 38332
rect 42924 38276 42980 38332
rect 57344 38304 57456 38332
rect 2258 38220 2268 38276
rect 2324 38220 3948 38276
rect 4004 38220 4014 38276
rect 6402 38220 6412 38276
rect 6468 38220 7084 38276
rect 7140 38220 7150 38276
rect 7858 38220 7868 38276
rect 7924 38220 11956 38276
rect 12114 38220 12124 38276
rect 12180 38220 14812 38276
rect 14868 38220 14878 38276
rect 27682 38220 27692 38276
rect 27748 38220 28756 38276
rect 29250 38220 29260 38276
rect 29316 38220 30940 38276
rect 30996 38220 31006 38276
rect 39554 38220 39564 38276
rect 39620 38220 41468 38276
rect 41524 38220 41804 38276
rect 41860 38220 41870 38276
rect 42018 38220 42028 38276
rect 42084 38220 42980 38276
rect 43250 38220 43260 38276
rect 43316 38220 44940 38276
rect 44996 38220 45006 38276
rect 45164 38220 47516 38276
rect 47572 38220 47582 38276
rect 48178 38220 48188 38276
rect 48244 38220 48412 38276
rect 48468 38220 49084 38276
rect 49140 38220 49150 38276
rect 49298 38220 49308 38276
rect 49364 38220 53900 38276
rect 53956 38220 53966 38276
rect 55412 38220 56700 38276
rect 56756 38220 56766 38276
rect 28700 38164 28756 38220
rect 45164 38164 45220 38220
rect 55412 38164 55468 38220
rect 1558 38108 1596 38164
rect 1652 38108 1662 38164
rect 3332 38108 6188 38164
rect 6244 38108 6254 38164
rect 7746 38108 7756 38164
rect 7812 38108 8876 38164
rect 8932 38108 8942 38164
rect 9202 38108 9212 38164
rect 9268 38108 9884 38164
rect 9940 38108 9950 38164
rect 10994 38108 11004 38164
rect 11060 38108 11564 38164
rect 11620 38108 13692 38164
rect 13748 38108 13758 38164
rect 14242 38108 14252 38164
rect 14308 38108 18956 38164
rect 19012 38108 19022 38164
rect 19180 38108 23324 38164
rect 23380 38108 23390 38164
rect 23874 38108 23884 38164
rect 23940 38108 25228 38164
rect 25284 38108 25294 38164
rect 28700 38108 30828 38164
rect 30884 38108 31388 38164
rect 31444 38108 31454 38164
rect 34850 38108 34860 38164
rect 34916 38108 37884 38164
rect 37940 38108 39788 38164
rect 39844 38108 39854 38164
rect 41346 38108 41356 38164
rect 41412 38108 45220 38164
rect 46722 38108 46732 38164
rect 46788 38108 47292 38164
rect 47348 38108 48076 38164
rect 48132 38108 48142 38164
rect 48402 38108 48412 38164
rect 48468 38108 49308 38164
rect 49364 38108 49374 38164
rect 49532 38108 55468 38164
rect 56354 38108 56364 38164
rect 56420 38108 56812 38164
rect 56868 38108 56878 38164
rect 3332 38052 3388 38108
rect 2482 37996 2492 38052
rect 2548 37996 3388 38052
rect 3602 37996 3612 38052
rect 3668 37996 5068 38052
rect 5124 37996 5134 38052
rect 5590 37996 5628 38052
rect 5684 37996 5694 38052
rect 8194 37996 8204 38052
rect 8260 37996 9324 38052
rect 9380 37996 9390 38052
rect 10546 37996 10556 38052
rect 10612 37996 13132 38052
rect 13188 37996 13198 38052
rect 14690 37996 14700 38052
rect 14756 37996 15372 38052
rect 15428 37996 15438 38052
rect 0 37940 112 37968
rect 19180 37940 19236 38108
rect 49532 38052 49588 38108
rect 19954 37996 19964 38052
rect 20020 37996 23548 38052
rect 23604 37996 23614 38052
rect 27906 37996 27916 38052
rect 27972 37996 28700 38052
rect 28756 37996 28766 38052
rect 28998 37996 29036 38052
rect 29092 37996 29102 38052
rect 30930 37996 30940 38052
rect 30996 37996 31052 38052
rect 31108 37996 31118 38052
rect 36306 37996 36316 38052
rect 36372 37996 44492 38052
rect 44548 37996 44558 38052
rect 45042 37996 45052 38052
rect 45108 37996 49588 38052
rect 51090 37996 51100 38052
rect 51156 37996 51660 38052
rect 51716 37996 51726 38052
rect 52434 37996 52444 38052
rect 52500 37996 53340 38052
rect 53396 37996 53564 38052
rect 53620 37996 54572 38052
rect 54628 37996 54638 38052
rect 56018 37996 56028 38052
rect 56084 37996 56700 38052
rect 56756 37996 56766 38052
rect 45052 37940 45108 37996
rect 57344 37940 57456 37968
rect 0 37884 2044 37940
rect 2100 37884 2110 37940
rect 2930 37884 2940 37940
rect 2996 37884 5516 37940
rect 5572 37884 5582 37940
rect 5740 37884 19236 37940
rect 19618 37884 19628 37940
rect 19684 37884 21756 37940
rect 21812 37884 22316 37940
rect 22372 37884 22382 37940
rect 22866 37884 22876 37940
rect 22932 37884 24556 37940
rect 24612 37884 24622 37940
rect 38882 37884 38892 37940
rect 38948 37884 42476 37940
rect 42532 37884 45108 37940
rect 45826 37884 45836 37940
rect 45892 37884 45948 37940
rect 46004 37884 46014 37940
rect 46722 37884 46732 37940
rect 46788 37884 49196 37940
rect 49252 37884 49262 37940
rect 50082 37884 50092 37940
rect 50148 37884 57456 37940
rect 0 37856 112 37884
rect 5740 37828 5796 37884
rect 57344 37856 57456 37884
rect 2706 37772 2716 37828
rect 2772 37772 4396 37828
rect 4452 37772 4462 37828
rect 4732 37772 5796 37828
rect 6178 37772 6188 37828
rect 6244 37772 11340 37828
rect 11396 37772 11406 37828
rect 12236 37772 14588 37828
rect 14644 37772 14654 37828
rect 15026 37772 15036 37828
rect 15092 37772 15820 37828
rect 15876 37772 15886 37828
rect 16034 37772 16044 37828
rect 16100 37772 49308 37828
rect 49364 37772 49374 37828
rect 51090 37772 51100 37828
rect 51156 37772 55356 37828
rect 55412 37772 55422 37828
rect 4732 37716 4788 37772
rect 4274 37660 4284 37716
rect 4340 37660 4788 37716
rect 4946 37660 4956 37716
rect 5012 37660 5292 37716
rect 5348 37660 5358 37716
rect 8418 37660 8428 37716
rect 8484 37660 12012 37716
rect 12068 37660 12078 37716
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 12236 37604 12292 37772
rect 12674 37660 12684 37716
rect 12740 37660 16268 37716
rect 16324 37660 16334 37716
rect 17154 37660 17164 37716
rect 17220 37660 18284 37716
rect 18340 37660 18350 37716
rect 24322 37660 24332 37716
rect 24388 37660 26908 37716
rect 26964 37660 26974 37716
rect 28364 37660 38668 37716
rect 40786 37660 40796 37716
rect 40852 37660 41468 37716
rect 41524 37660 41534 37716
rect 41794 37660 41804 37716
rect 41860 37660 42140 37716
rect 42196 37660 42206 37716
rect 44146 37660 44156 37716
rect 44212 37660 44940 37716
rect 44996 37660 45006 37716
rect 47506 37660 47516 37716
rect 47572 37660 48188 37716
rect 48244 37660 48254 37716
rect 48850 37660 48860 37716
rect 48916 37660 49084 37716
rect 49140 37660 51436 37716
rect 51492 37660 52444 37716
rect 52500 37660 52510 37716
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 28364 37604 28420 37660
rect 38612 37604 38668 37660
rect 43794 37604 43804 37660
rect 43860 37604 43908 37660
rect 43964 37604 44012 37660
rect 44068 37604 44078 37660
rect 3378 37548 3388 37604
rect 3444 37548 3500 37604
rect 3556 37548 3566 37604
rect 4162 37548 4172 37604
rect 4228 37548 4956 37604
rect 5012 37548 5022 37604
rect 5170 37548 5180 37604
rect 5236 37548 5964 37604
rect 6020 37548 6030 37604
rect 6514 37548 6524 37604
rect 6580 37548 7868 37604
rect 7924 37548 8316 37604
rect 8372 37548 8382 37604
rect 8530 37548 8540 37604
rect 8596 37548 8876 37604
rect 8932 37548 8942 37604
rect 9650 37548 9660 37604
rect 9716 37548 11228 37604
rect 11284 37548 12292 37604
rect 14466 37548 14476 37604
rect 14532 37548 18060 37604
rect 18116 37548 18126 37604
rect 18386 37548 18396 37604
rect 18452 37548 21084 37604
rect 21140 37548 21150 37604
rect 24210 37548 24220 37604
rect 24276 37548 24892 37604
rect 24948 37548 24958 37604
rect 25106 37548 25116 37604
rect 25172 37548 26012 37604
rect 26068 37548 26078 37604
rect 26898 37548 26908 37604
rect 26964 37548 28420 37604
rect 31826 37548 31836 37604
rect 31892 37548 34468 37604
rect 38612 37548 43260 37604
rect 43316 37548 43326 37604
rect 44482 37548 44492 37604
rect 44548 37548 54348 37604
rect 54404 37548 54414 37604
rect 55122 37548 55132 37604
rect 55188 37548 55356 37604
rect 55412 37548 55422 37604
rect 0 37492 112 37520
rect 34412 37492 34468 37548
rect 57344 37492 57456 37520
rect 0 37436 33628 37492
rect 33684 37436 33694 37492
rect 34412 37436 54124 37492
rect 54180 37436 54190 37492
rect 55234 37436 55244 37492
rect 55300 37436 57456 37492
rect 0 37408 112 37436
rect 57344 37408 57456 37436
rect 2146 37324 2156 37380
rect 2212 37324 5068 37380
rect 5124 37324 5134 37380
rect 5282 37324 5292 37380
rect 5348 37324 19180 37380
rect 19236 37324 19246 37380
rect 22540 37324 25452 37380
rect 25508 37324 25518 37380
rect 27122 37324 27132 37380
rect 27188 37324 28476 37380
rect 28532 37324 28542 37380
rect 30594 37324 30604 37380
rect 30660 37324 34076 37380
rect 34132 37324 34142 37380
rect 36082 37324 36092 37380
rect 36148 37324 37548 37380
rect 37604 37324 37614 37380
rect 40114 37324 40124 37380
rect 40180 37324 41244 37380
rect 41300 37324 41310 37380
rect 41458 37324 41468 37380
rect 41524 37324 41804 37380
rect 41860 37324 41870 37380
rect 42690 37324 42700 37380
rect 42756 37324 42812 37380
rect 42868 37324 42878 37380
rect 43586 37324 43596 37380
rect 43652 37324 45164 37380
rect 45220 37324 45230 37380
rect 46274 37324 46284 37380
rect 46340 37324 47292 37380
rect 47348 37324 47358 37380
rect 49746 37324 49756 37380
rect 49812 37324 50092 37380
rect 50148 37324 51772 37380
rect 51828 37324 51838 37380
rect 53116 37324 53228 37380
rect 53284 37324 53294 37380
rect 55122 37324 55132 37380
rect 55188 37324 56476 37380
rect 56532 37324 56542 37380
rect 1474 37212 1484 37268
rect 1540 37212 5068 37268
rect 5124 37212 5134 37268
rect 8194 37212 8204 37268
rect 8260 37212 9884 37268
rect 9940 37212 10332 37268
rect 10388 37212 13804 37268
rect 13860 37212 13870 37268
rect 14802 37212 14812 37268
rect 14868 37212 15932 37268
rect 15988 37212 15998 37268
rect 17602 37212 17612 37268
rect 17668 37212 17724 37268
rect 17780 37212 17790 37268
rect 22540 37156 22596 37324
rect 53116 37268 53172 37324
rect 22764 37212 24892 37268
rect 24948 37212 24958 37268
rect 25106 37212 25116 37268
rect 25172 37212 25676 37268
rect 25732 37212 25742 37268
rect 27206 37212 27244 37268
rect 27300 37212 27310 37268
rect 28354 37212 28364 37268
rect 28420 37212 31052 37268
rect 31108 37212 31118 37268
rect 31938 37212 31948 37268
rect 32004 37212 33628 37268
rect 33684 37212 33694 37268
rect 34850 37212 34860 37268
rect 34916 37212 36540 37268
rect 36596 37212 36764 37268
rect 36820 37212 36830 37268
rect 37202 37212 37212 37268
rect 37268 37212 37660 37268
rect 37716 37212 39564 37268
rect 39620 37212 39630 37268
rect 39750 37212 39788 37268
rect 39844 37212 39854 37268
rect 41906 37212 41916 37268
rect 41972 37212 43708 37268
rect 43764 37212 43774 37268
rect 44482 37212 44492 37268
rect 44548 37212 50540 37268
rect 50596 37212 50606 37268
rect 51324 37212 53172 37268
rect 53330 37212 53340 37268
rect 53396 37212 53788 37268
rect 53844 37212 53854 37268
rect 54236 37212 57260 37268
rect 57316 37212 57326 37268
rect 2818 37100 2828 37156
rect 2884 37100 3668 37156
rect 4162 37100 4172 37156
rect 4228 37100 4396 37156
rect 4452 37100 4462 37156
rect 4610 37100 4620 37156
rect 4676 37100 4844 37156
rect 4900 37100 4910 37156
rect 5506 37100 5516 37156
rect 5572 37100 6188 37156
rect 6244 37100 6254 37156
rect 6850 37100 6860 37156
rect 6916 37100 10332 37156
rect 10388 37100 10398 37156
rect 13234 37100 13244 37156
rect 13300 37100 14476 37156
rect 14532 37100 14542 37156
rect 15026 37100 15036 37156
rect 15092 37100 17388 37156
rect 17444 37100 18508 37156
rect 18564 37100 18574 37156
rect 19394 37100 19404 37156
rect 19460 37100 22540 37156
rect 22596 37100 22606 37156
rect 0 37044 112 37072
rect 0 36988 3556 37044
rect 3612 36988 3668 37100
rect 22764 37044 22820 37212
rect 51324 37156 51380 37212
rect 54236 37156 54292 37212
rect 23426 37100 23436 37156
rect 23492 37100 24220 37156
rect 24276 37100 24286 37156
rect 24546 37100 24556 37156
rect 24612 37100 26012 37156
rect 26068 37100 26078 37156
rect 26450 37100 26460 37156
rect 26516 37100 27020 37156
rect 27076 37100 27086 37156
rect 28242 37100 28252 37156
rect 28308 37100 29036 37156
rect 29092 37100 29372 37156
rect 29428 37100 29438 37156
rect 29922 37100 29932 37156
rect 29988 37100 33068 37156
rect 33124 37100 33134 37156
rect 33628 37100 34748 37156
rect 34804 37100 34814 37156
rect 35634 37100 35644 37156
rect 35700 37100 35868 37156
rect 35924 37100 35934 37156
rect 36082 37100 36092 37156
rect 36148 37100 44156 37156
rect 44212 37100 44716 37156
rect 44772 37100 44782 37156
rect 50642 37100 50652 37156
rect 50708 37100 51380 37156
rect 51538 37100 51548 37156
rect 51604 37100 54292 37156
rect 55122 37100 55132 37156
rect 55188 37100 55468 37156
rect 55524 37100 55534 37156
rect 33628 37044 33684 37100
rect 57344 37044 57456 37072
rect 3724 36988 3734 37044
rect 5058 36988 5068 37044
rect 5124 36988 7980 37044
rect 8036 36988 8046 37044
rect 8194 36988 8204 37044
rect 8260 36988 9436 37044
rect 9492 36988 9502 37044
rect 9650 36988 9660 37044
rect 9716 36988 10444 37044
rect 10500 36988 10510 37044
rect 12338 36988 12348 37044
rect 12404 36988 12684 37044
rect 12740 36988 12750 37044
rect 15138 36988 15148 37044
rect 15204 36988 15484 37044
rect 15540 36988 15550 37044
rect 15698 36988 15708 37044
rect 15764 36988 16828 37044
rect 16884 36988 16894 37044
rect 17164 36988 18284 37044
rect 18340 36988 21308 37044
rect 21364 36988 21374 37044
rect 22754 36988 22764 37044
rect 22820 36988 22830 37044
rect 23090 36988 23100 37044
rect 23156 36988 25564 37044
rect 25620 36988 25630 37044
rect 25788 36988 32508 37044
rect 32564 36988 32574 37044
rect 33170 36988 33180 37044
rect 33236 36988 33684 37044
rect 33842 36988 33852 37044
rect 33908 36988 36764 37044
rect 36820 36988 36830 37044
rect 38612 36988 42700 37044
rect 42756 36988 42766 37044
rect 43586 36988 43596 37044
rect 43652 36988 49196 37044
rect 49252 36988 49262 37044
rect 49522 36988 49532 37044
rect 49588 36988 50540 37044
rect 50596 36988 50764 37044
rect 50820 36988 50830 37044
rect 52854 36988 52892 37044
rect 52948 36988 52958 37044
rect 53106 36988 53116 37044
rect 53172 36988 53564 37044
rect 53620 36988 53630 37044
rect 53778 36988 53788 37044
rect 53844 36988 54124 37044
rect 54180 36988 54190 37044
rect 54450 36988 54460 37044
rect 54516 36988 55132 37044
rect 55188 36988 55198 37044
rect 57250 36988 57260 37044
rect 57316 36988 57456 37044
rect 0 36960 112 36988
rect 3500 36932 3556 36988
rect 5068 36932 5124 36988
rect 3500 36876 4284 36932
rect 4340 36876 4350 36932
rect 4834 36876 4844 36932
rect 4900 36876 5124 36932
rect 7858 36876 7868 36932
rect 7924 36876 9324 36932
rect 9380 36876 9390 36932
rect 9762 36876 9772 36932
rect 9828 36876 9996 36932
rect 10052 36876 10062 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 17164 36820 17220 36988
rect 25788 36932 25844 36988
rect 38612 36932 38668 36988
rect 57344 36960 57456 36988
rect 17378 36876 17388 36932
rect 17444 36876 18844 36932
rect 18900 36876 18910 36932
rect 25442 36876 25452 36932
rect 25508 36876 25844 36932
rect 26786 36876 26796 36932
rect 26852 36876 29148 36932
rect 29204 36876 29214 36932
rect 29922 36876 29932 36932
rect 29988 36876 35196 36932
rect 35252 36876 35262 36932
rect 37660 36876 38668 36932
rect 40562 36876 40572 36932
rect 40628 36876 41356 36932
rect 41412 36876 41422 36932
rect 41682 36876 41692 36932
rect 41748 36876 41804 36932
rect 41860 36876 41870 36932
rect 42466 36876 42476 36932
rect 42532 36876 44156 36932
rect 44212 36876 44222 36932
rect 49970 36876 49980 36932
rect 50036 36876 51660 36932
rect 51716 36876 51726 36932
rect 52546 36876 52556 36932
rect 52612 36876 55692 36932
rect 55748 36876 55758 36932
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 37660 36820 37716 36876
rect 44454 36820 44464 36876
rect 44520 36820 44568 36876
rect 44624 36820 44672 36876
rect 44728 36820 44738 36876
rect 578 36764 588 36820
rect 644 36764 1596 36820
rect 1652 36764 1662 36820
rect 2146 36764 2156 36820
rect 2212 36764 2716 36820
rect 2772 36764 2782 36820
rect 5058 36764 5068 36820
rect 5124 36764 6300 36820
rect 6356 36764 6366 36820
rect 6636 36764 7756 36820
rect 7812 36764 7822 36820
rect 8082 36764 8092 36820
rect 8148 36764 9660 36820
rect 9716 36764 9726 36820
rect 10098 36764 10108 36820
rect 10164 36764 11340 36820
rect 11396 36764 11406 36820
rect 12562 36764 12572 36820
rect 12628 36764 13132 36820
rect 13188 36764 14476 36820
rect 14532 36764 17220 36820
rect 17490 36764 17500 36820
rect 17556 36764 17836 36820
rect 17892 36764 20972 36820
rect 21028 36764 21038 36820
rect 21858 36764 21868 36820
rect 21924 36764 22204 36820
rect 22260 36764 22270 36820
rect 23762 36764 23772 36820
rect 23828 36764 24220 36820
rect 24276 36764 24286 36820
rect 24882 36764 24892 36820
rect 24948 36764 30940 36820
rect 30996 36764 31006 36820
rect 32834 36764 32844 36820
rect 32900 36764 34860 36820
rect 34916 36764 34926 36820
rect 35298 36764 35308 36820
rect 35364 36764 37716 36820
rect 38612 36764 41244 36820
rect 41300 36764 44156 36820
rect 44212 36764 44222 36820
rect 46498 36764 46508 36820
rect 46564 36764 46732 36820
rect 46788 36764 46798 36820
rect 47394 36764 47404 36820
rect 47460 36764 50372 36820
rect 52434 36764 52444 36820
rect 52500 36764 56252 36820
rect 56308 36764 56318 36820
rect 57026 36764 57036 36820
rect 57092 36764 57260 36820
rect 57316 36764 57326 36820
rect 6636 36708 6692 36764
rect 38612 36708 38668 36764
rect 50316 36708 50372 36764
rect 2034 36652 2044 36708
rect 2100 36652 6692 36708
rect 6822 36652 6860 36708
rect 6916 36652 6926 36708
rect 7186 36652 7196 36708
rect 7252 36652 8596 36708
rect 9202 36652 9212 36708
rect 9268 36652 13356 36708
rect 13412 36652 13422 36708
rect 13570 36652 13580 36708
rect 13636 36652 37436 36708
rect 37492 36652 38668 36708
rect 40562 36652 40572 36708
rect 40628 36652 41244 36708
rect 41300 36652 41310 36708
rect 42242 36652 42252 36708
rect 42308 36652 42476 36708
rect 42532 36652 42542 36708
rect 43362 36652 43372 36708
rect 43428 36652 50092 36708
rect 50148 36652 50158 36708
rect 50316 36652 52388 36708
rect 52658 36652 52668 36708
rect 52724 36652 53116 36708
rect 53172 36652 53182 36708
rect 53666 36652 53676 36708
rect 53732 36652 53900 36708
rect 53956 36652 53966 36708
rect 0 36596 112 36624
rect 8540 36596 8596 36652
rect 0 36540 7140 36596
rect 7298 36540 7308 36596
rect 7364 36540 8316 36596
rect 8372 36540 8382 36596
rect 8540 36540 9660 36596
rect 9716 36540 9726 36596
rect 10108 36540 13580 36596
rect 13636 36540 13646 36596
rect 14886 36540 14924 36596
rect 14980 36540 14990 36596
rect 15092 36540 33964 36596
rect 34020 36540 34030 36596
rect 35186 36540 35196 36596
rect 35252 36540 38052 36596
rect 38182 36540 38220 36596
rect 38276 36540 42700 36596
rect 42756 36540 42766 36596
rect 43372 36540 51772 36596
rect 51828 36540 51838 36596
rect 0 36512 112 36540
rect 7084 36484 7140 36540
rect 2818 36428 2828 36484
rect 2884 36428 4732 36484
rect 4788 36428 5852 36484
rect 5908 36428 5918 36484
rect 7084 36428 9436 36484
rect 9492 36428 9502 36484
rect 10108 36372 10164 36540
rect 15092 36484 15148 36540
rect 37996 36484 38052 36540
rect 43372 36484 43428 36540
rect 52332 36484 52388 36652
rect 57344 36596 57456 36624
rect 52770 36540 52780 36596
rect 52836 36540 55916 36596
rect 55972 36540 55982 36596
rect 56914 36540 56924 36596
rect 56980 36540 57456 36596
rect 57344 36512 57456 36540
rect 10994 36428 11004 36484
rect 11060 36428 14700 36484
rect 14756 36428 14766 36484
rect 14924 36428 15148 36484
rect 19730 36428 19740 36484
rect 19796 36428 20860 36484
rect 20916 36428 20926 36484
rect 22082 36428 22092 36484
rect 22148 36428 23548 36484
rect 23604 36428 24892 36484
rect 24948 36428 24958 36484
rect 26786 36428 26796 36484
rect 26852 36428 27468 36484
rect 27524 36428 27534 36484
rect 29474 36428 29484 36484
rect 29540 36428 30044 36484
rect 30100 36428 30110 36484
rect 32946 36428 32956 36484
rect 33012 36428 33180 36484
rect 33236 36428 33246 36484
rect 34738 36428 34748 36484
rect 34804 36428 35532 36484
rect 35588 36428 35598 36484
rect 37426 36428 37436 36484
rect 37492 36428 37548 36484
rect 37604 36428 37614 36484
rect 37996 36428 43204 36484
rect 43362 36428 43372 36484
rect 43428 36428 43438 36484
rect 46050 36428 46060 36484
rect 46116 36428 46956 36484
rect 47012 36428 47964 36484
rect 48020 36428 48030 36484
rect 48738 36428 48748 36484
rect 48804 36428 51044 36484
rect 51314 36428 51324 36484
rect 51380 36428 52108 36484
rect 52164 36428 52174 36484
rect 52332 36428 53340 36484
rect 53396 36428 53406 36484
rect 54338 36428 54348 36484
rect 54404 36428 54684 36484
rect 54740 36428 54750 36484
rect 54898 36428 54908 36484
rect 54964 36428 56252 36484
rect 56308 36428 56318 36484
rect 14924 36372 14980 36428
rect 43148 36372 43204 36428
rect 50988 36372 51044 36428
rect 2930 36316 2940 36372
rect 2996 36316 3052 36372
rect 3108 36316 3276 36372
rect 3332 36316 3342 36372
rect 4050 36316 4060 36372
rect 4116 36316 4508 36372
rect 4564 36316 4574 36372
rect 5954 36316 5964 36372
rect 6020 36316 8204 36372
rect 8260 36316 8270 36372
rect 8642 36316 8652 36372
rect 8708 36316 8876 36372
rect 8932 36316 8942 36372
rect 9538 36316 9548 36372
rect 9604 36316 10108 36372
rect 10164 36316 10174 36372
rect 13458 36316 13468 36372
rect 13524 36316 14980 36372
rect 15586 36316 15596 36372
rect 15652 36316 21756 36372
rect 21812 36316 22204 36372
rect 22260 36316 22988 36372
rect 23044 36316 24724 36372
rect 27122 36316 27132 36372
rect 27188 36316 29932 36372
rect 29988 36316 29998 36372
rect 30370 36316 30380 36372
rect 30436 36316 35980 36372
rect 36036 36316 36046 36372
rect 36530 36316 36540 36372
rect 36596 36316 37884 36372
rect 37940 36316 37950 36372
rect 41094 36316 41132 36372
rect 41188 36316 41692 36372
rect 41748 36316 41758 36372
rect 43148 36316 43484 36372
rect 43540 36316 43550 36372
rect 43698 36316 43708 36372
rect 43764 36316 45388 36372
rect 45444 36316 49084 36372
rect 49140 36316 50764 36372
rect 50820 36316 50830 36372
rect 50988 36316 54796 36372
rect 54852 36316 54862 36372
rect 55346 36316 55356 36372
rect 55412 36316 55804 36372
rect 55860 36316 56140 36372
rect 56196 36316 56206 36372
rect 1474 36204 1484 36260
rect 1540 36204 2492 36260
rect 2548 36204 2558 36260
rect 3332 36204 14924 36260
rect 14980 36204 14990 36260
rect 15810 36204 15820 36260
rect 15876 36204 23660 36260
rect 23716 36204 23726 36260
rect 0 36148 112 36176
rect 3332 36148 3388 36204
rect 24668 36148 24724 36316
rect 43484 36260 43540 36316
rect 24882 36204 24892 36260
rect 24948 36204 41356 36260
rect 41412 36204 41422 36260
rect 43484 36204 46508 36260
rect 46564 36204 46574 36260
rect 46946 36204 46956 36260
rect 47012 36204 48860 36260
rect 48916 36204 48926 36260
rect 49074 36204 49084 36260
rect 49140 36204 52108 36260
rect 52164 36204 52174 36260
rect 52770 36204 52780 36260
rect 52836 36204 56252 36260
rect 56308 36204 56318 36260
rect 57344 36148 57456 36176
rect 0 36092 3388 36148
rect 4386 36092 4396 36148
rect 4452 36092 5068 36148
rect 5124 36092 5134 36148
rect 5730 36092 5740 36148
rect 5796 36092 6188 36148
rect 6244 36092 6972 36148
rect 7028 36092 7038 36148
rect 7410 36092 7420 36148
rect 7476 36092 10444 36148
rect 10500 36092 10510 36148
rect 12338 36092 12348 36148
rect 12404 36092 13580 36148
rect 13636 36092 13646 36148
rect 15250 36092 15260 36148
rect 15316 36092 15372 36148
rect 15428 36092 15438 36148
rect 16818 36092 16828 36148
rect 16884 36092 17948 36148
rect 18004 36092 18014 36148
rect 18498 36092 18508 36148
rect 18564 36092 19404 36148
rect 19460 36092 21084 36148
rect 21140 36092 21150 36148
rect 24668 36092 25228 36148
rect 25284 36092 25294 36148
rect 26674 36092 26684 36148
rect 26740 36092 31612 36148
rect 31668 36092 31678 36148
rect 33282 36092 33292 36148
rect 33348 36092 35196 36148
rect 35252 36092 35262 36148
rect 35858 36092 35868 36148
rect 35924 36092 37996 36148
rect 38052 36092 38062 36148
rect 47506 36092 47516 36148
rect 47572 36092 49196 36148
rect 49252 36092 49262 36148
rect 51426 36092 51436 36148
rect 51492 36092 51772 36148
rect 51828 36092 51838 36148
rect 56466 36092 56476 36148
rect 56532 36092 57456 36148
rect 0 36064 112 36092
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 26684 36036 26740 36092
rect 43794 36036 43804 36092
rect 43860 36036 43908 36092
rect 43964 36036 44012 36092
rect 44068 36036 44078 36092
rect 57344 36064 57456 36092
rect 4498 35980 4508 36036
rect 4564 35980 8988 36036
rect 9044 35980 9054 36036
rect 9212 35980 22428 36036
rect 22484 35980 22494 36036
rect 23314 35980 23324 36036
rect 23380 35980 23660 36036
rect 23716 35980 23726 36036
rect 24210 35980 24220 36036
rect 24276 35980 24892 36036
rect 24948 35980 24958 36036
rect 25218 35980 25228 36036
rect 25284 35980 26740 36036
rect 27346 35980 27356 36036
rect 27412 35980 30044 36036
rect 30100 35980 30110 36036
rect 31378 35980 31388 36036
rect 31444 35980 33740 36036
rect 33796 35980 33806 36036
rect 33954 35980 33964 36036
rect 34020 35980 40124 36036
rect 40180 35980 40190 36036
rect 41356 35980 43596 36036
rect 43652 35980 43662 36036
rect 44370 35980 44380 36036
rect 44436 35980 46732 36036
rect 46788 35980 47628 36036
rect 47684 35980 47694 36036
rect 48178 35980 48188 36036
rect 48244 35980 49420 36036
rect 49476 35980 49486 36036
rect 50372 35980 52668 36036
rect 52724 35980 52734 36036
rect 54786 35980 54796 36036
rect 54852 35980 55468 36036
rect 55524 35980 55534 36036
rect 3490 35868 3500 35924
rect 3556 35868 3948 35924
rect 4004 35868 4284 35924
rect 4340 35868 5292 35924
rect 5348 35868 5358 35924
rect 6066 35868 6076 35924
rect 6132 35868 7868 35924
rect 7924 35868 7934 35924
rect 8642 35868 8652 35924
rect 8708 35868 8876 35924
rect 8932 35868 8942 35924
rect 3378 35756 3388 35812
rect 3444 35756 4956 35812
rect 5012 35756 5022 35812
rect 5702 35756 5740 35812
rect 5796 35756 8428 35812
rect 8484 35756 8494 35812
rect 0 35700 112 35728
rect 9212 35700 9268 35980
rect 41356 35924 41412 35980
rect 50372 35924 50428 35980
rect 9426 35868 9436 35924
rect 9492 35868 41412 35924
rect 41570 35868 41580 35924
rect 41636 35868 44268 35924
rect 44324 35868 44334 35924
rect 44492 35868 50428 35924
rect 51538 35868 51548 35924
rect 51604 35868 51996 35924
rect 52052 35868 52062 35924
rect 52434 35868 52444 35924
rect 52500 35868 55804 35924
rect 55860 35868 55870 35924
rect 44492 35812 44548 35868
rect 9426 35756 9436 35812
rect 9492 35756 10556 35812
rect 10612 35756 10622 35812
rect 11778 35756 11788 35812
rect 11844 35756 11900 35812
rect 11956 35756 11966 35812
rect 12114 35756 12124 35812
rect 12180 35756 41916 35812
rect 41972 35756 41982 35812
rect 43474 35756 43484 35812
rect 43540 35756 44548 35812
rect 45490 35756 45500 35812
rect 45556 35756 46732 35812
rect 46788 35756 46956 35812
rect 47012 35756 47022 35812
rect 47506 35756 47516 35812
rect 47572 35756 49868 35812
rect 49924 35756 52556 35812
rect 52612 35756 52622 35812
rect 54786 35756 54796 35812
rect 54852 35756 56476 35812
rect 56532 35756 56542 35812
rect 57344 35700 57456 35728
rect 0 35644 9268 35700
rect 12786 35644 12796 35700
rect 12852 35644 13916 35700
rect 13972 35644 14756 35700
rect 14914 35644 14924 35700
rect 14980 35644 15820 35700
rect 15876 35644 15886 35700
rect 17266 35644 17276 35700
rect 17332 35644 17388 35700
rect 17444 35644 17454 35700
rect 22418 35644 22428 35700
rect 22484 35644 26124 35700
rect 26180 35644 26908 35700
rect 30034 35644 30044 35700
rect 30100 35644 31052 35700
rect 31108 35644 31118 35700
rect 33254 35644 33292 35700
rect 33348 35644 33358 35700
rect 33618 35644 33628 35700
rect 33684 35644 39116 35700
rect 39172 35644 39182 35700
rect 39778 35644 39788 35700
rect 39844 35644 40236 35700
rect 40292 35644 40302 35700
rect 40870 35644 40908 35700
rect 40964 35644 40974 35700
rect 43586 35644 43596 35700
rect 43652 35644 45276 35700
rect 45332 35644 45948 35700
rect 46004 35644 46014 35700
rect 46610 35644 46620 35700
rect 46676 35644 48412 35700
rect 48468 35644 48478 35700
rect 50418 35644 50428 35700
rect 50484 35644 52108 35700
rect 52164 35644 52174 35700
rect 52322 35644 52332 35700
rect 52388 35644 54124 35700
rect 54180 35644 54190 35700
rect 55234 35644 55244 35700
rect 55300 35644 55356 35700
rect 55412 35644 55422 35700
rect 55570 35644 55580 35700
rect 55636 35644 57456 35700
rect 0 35616 112 35644
rect 14700 35588 14756 35644
rect 26852 35588 26908 35644
rect 57344 35616 57456 35644
rect 3826 35532 3836 35588
rect 3892 35532 4508 35588
rect 4564 35532 4574 35588
rect 5842 35532 5852 35588
rect 5908 35532 6412 35588
rect 6468 35532 6478 35588
rect 6636 35532 8428 35588
rect 8484 35532 8494 35588
rect 8978 35532 8988 35588
rect 9044 35532 9436 35588
rect 9492 35532 9502 35588
rect 14326 35532 14364 35588
rect 14420 35532 14430 35588
rect 14700 35532 15596 35588
rect 15652 35532 15662 35588
rect 17378 35532 17388 35588
rect 17444 35532 17612 35588
rect 17668 35532 17678 35588
rect 18050 35532 18060 35588
rect 18116 35532 19740 35588
rect 19796 35532 19806 35588
rect 21858 35532 21868 35588
rect 21924 35532 22092 35588
rect 22148 35532 22158 35588
rect 22978 35532 22988 35588
rect 23044 35532 23324 35588
rect 23380 35532 23390 35588
rect 23762 35532 23772 35588
rect 23828 35532 26012 35588
rect 26068 35532 26078 35588
rect 26852 35532 31164 35588
rect 31220 35532 31230 35588
rect 31826 35532 31836 35588
rect 31892 35532 33180 35588
rect 33236 35532 38780 35588
rect 38836 35532 38846 35588
rect 39666 35532 39676 35588
rect 39732 35532 42364 35588
rect 42420 35532 42430 35588
rect 42914 35532 42924 35588
rect 42980 35532 43036 35588
rect 43092 35532 43148 35588
rect 43204 35532 43214 35588
rect 43698 35532 43708 35588
rect 43764 35532 53116 35588
rect 53172 35532 55132 35588
rect 55188 35532 55198 35588
rect 6636 35476 6692 35532
rect 2370 35420 2380 35476
rect 2436 35420 5964 35476
rect 6020 35420 6030 35476
rect 6290 35420 6300 35476
rect 6356 35420 6636 35476
rect 6692 35420 6702 35476
rect 7858 35420 7868 35476
rect 7924 35420 7980 35476
rect 8036 35420 13244 35476
rect 13300 35420 13310 35476
rect 14578 35420 14588 35476
rect 14644 35420 22708 35476
rect 22866 35420 22876 35476
rect 22932 35420 23100 35476
rect 23156 35420 23166 35476
rect 23650 35420 23660 35476
rect 23716 35420 24220 35476
rect 24276 35420 24444 35476
rect 24500 35420 24510 35476
rect 24658 35420 24668 35476
rect 24724 35420 25116 35476
rect 25172 35420 25182 35476
rect 25554 35420 25564 35476
rect 25620 35420 28700 35476
rect 28756 35420 28766 35476
rect 29110 35420 29148 35476
rect 29204 35420 29820 35476
rect 29876 35420 29886 35476
rect 30258 35420 30268 35476
rect 30324 35420 31276 35476
rect 31332 35420 31342 35476
rect 34150 35420 34188 35476
rect 34244 35420 34254 35476
rect 35970 35420 35980 35476
rect 36036 35420 36540 35476
rect 36596 35420 36606 35476
rect 37202 35420 37212 35476
rect 37268 35420 37548 35476
rect 37604 35420 37614 35476
rect 39890 35420 39900 35476
rect 39956 35420 41468 35476
rect 41524 35420 41534 35476
rect 42242 35420 42252 35476
rect 42308 35420 45500 35476
rect 45556 35420 45566 35476
rect 46386 35420 46396 35476
rect 46452 35420 47292 35476
rect 47348 35420 47358 35476
rect 47506 35420 47516 35476
rect 47572 35420 49084 35476
rect 49140 35420 49150 35476
rect 50082 35420 50092 35476
rect 50148 35420 50988 35476
rect 51044 35420 51054 35476
rect 51986 35420 51996 35476
rect 52052 35420 52892 35476
rect 52948 35420 52958 35476
rect 54114 35420 54124 35476
rect 54180 35420 56140 35476
rect 56196 35420 56206 35476
rect 22652 35364 22708 35420
rect 1698 35308 1708 35364
rect 1764 35308 3836 35364
rect 3892 35308 3902 35364
rect 4844 35308 5292 35364
rect 5348 35308 5358 35364
rect 5506 35308 5516 35364
rect 5572 35308 6020 35364
rect 6962 35308 6972 35364
rect 7028 35308 7196 35364
rect 7252 35308 7262 35364
rect 7410 35308 7420 35364
rect 7476 35308 11116 35364
rect 11172 35308 11182 35364
rect 11330 35308 11340 35364
rect 11396 35308 18620 35364
rect 18676 35308 18686 35364
rect 19730 35308 19740 35364
rect 19796 35308 19806 35364
rect 22652 35308 24388 35364
rect 25106 35308 25116 35364
rect 25172 35308 31836 35364
rect 31892 35308 31902 35364
rect 35410 35308 35420 35364
rect 35476 35308 37100 35364
rect 37156 35308 37166 35364
rect 39218 35308 39228 35364
rect 39284 35308 43372 35364
rect 43428 35308 43438 35364
rect 44818 35308 44828 35364
rect 44884 35308 44894 35364
rect 46386 35308 46396 35364
rect 46452 35308 48524 35364
rect 48580 35308 48590 35364
rect 48748 35308 49532 35364
rect 49588 35308 49598 35364
rect 50372 35308 51548 35364
rect 51604 35308 51614 35364
rect 51874 35308 51884 35364
rect 51940 35308 53676 35364
rect 53732 35308 53742 35364
rect 0 35252 112 35280
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 4844 35252 4900 35308
rect 5964 35252 6020 35308
rect 19740 35252 19796 35308
rect 0 35196 2604 35252
rect 2660 35196 2670 35252
rect 3042 35196 3052 35252
rect 3108 35196 3724 35252
rect 3780 35196 3790 35252
rect 4844 35196 5068 35252
rect 5124 35196 5740 35252
rect 5796 35196 5806 35252
rect 5954 35196 5964 35252
rect 6020 35196 6030 35252
rect 6188 35196 13020 35252
rect 13076 35196 13086 35252
rect 14690 35196 14700 35252
rect 14756 35196 17164 35252
rect 17220 35196 17230 35252
rect 18498 35196 18508 35252
rect 18564 35196 19796 35252
rect 20188 35196 22764 35252
rect 22820 35196 23772 35252
rect 23828 35196 23838 35252
rect 0 35168 112 35196
rect 6188 35140 6244 35196
rect 3490 35084 3500 35140
rect 3556 35084 4844 35140
rect 4900 35084 4910 35140
rect 5068 35084 5516 35140
rect 5572 35084 5582 35140
rect 6066 35084 6076 35140
rect 6132 35084 6244 35140
rect 7186 35084 7196 35140
rect 7252 35084 16156 35140
rect 16212 35084 16222 35140
rect 16818 35084 16828 35140
rect 16884 35084 18620 35140
rect 18676 35084 18686 35140
rect 19170 35084 19180 35140
rect 19236 35084 19404 35140
rect 19460 35084 19470 35140
rect 5068 35028 5124 35084
rect 20188 35028 20244 35196
rect 24332 35140 24388 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 44454 35252 44464 35308
rect 44520 35252 44568 35308
rect 44624 35252 44672 35308
rect 44728 35252 44738 35308
rect 44828 35252 44884 35308
rect 48748 35252 48804 35308
rect 27570 35196 27580 35252
rect 27636 35196 28700 35252
rect 28756 35196 28766 35252
rect 29586 35196 29596 35252
rect 29652 35196 38444 35252
rect 38500 35196 38510 35252
rect 38658 35196 38668 35252
rect 38724 35196 39004 35252
rect 39060 35196 42812 35252
rect 42868 35196 43596 35252
rect 43652 35196 43662 35252
rect 44828 35196 45948 35252
rect 46004 35196 46014 35252
rect 46162 35196 46172 35252
rect 46228 35196 47740 35252
rect 47796 35196 48804 35252
rect 20598 35084 20636 35140
rect 20692 35084 20702 35140
rect 21410 35084 21420 35140
rect 21476 35084 21644 35140
rect 21700 35084 21710 35140
rect 24332 35084 25564 35140
rect 25620 35084 25630 35140
rect 28802 35084 28812 35140
rect 28868 35084 29820 35140
rect 29876 35084 33460 35140
rect 33618 35084 33628 35140
rect 33684 35084 38444 35140
rect 38500 35084 38510 35140
rect 38658 35084 38668 35140
rect 38724 35084 38836 35140
rect 40786 35084 40796 35140
rect 40852 35084 41468 35140
rect 41524 35084 42028 35140
rect 42084 35084 42094 35140
rect 42690 35084 42700 35140
rect 42756 35084 44828 35140
rect 44884 35084 44894 35140
rect 45042 35084 45052 35140
rect 45108 35084 45836 35140
rect 45892 35084 46284 35140
rect 46340 35084 46350 35140
rect 46498 35084 46508 35140
rect 46564 35084 47180 35140
rect 47236 35084 47246 35140
rect 33404 35028 33460 35084
rect 38780 35028 38836 35084
rect 50372 35028 50428 35308
rect 57344 35252 57456 35280
rect 50866 35196 50876 35252
rect 50932 35196 51100 35252
rect 51156 35196 51166 35252
rect 51762 35196 51772 35252
rect 51828 35196 53452 35252
rect 53508 35196 53518 35252
rect 53778 35196 53788 35252
rect 53844 35196 54684 35252
rect 54740 35196 54750 35252
rect 57250 35196 57260 35252
rect 57316 35196 57456 35252
rect 57344 35168 57456 35196
rect 50978 35084 50988 35140
rect 51044 35084 51212 35140
rect 51268 35084 51278 35140
rect 52770 35084 52780 35140
rect 52836 35084 53340 35140
rect 53396 35084 53406 35140
rect 2818 34972 2828 35028
rect 2884 34972 5124 35028
rect 5282 34972 5292 35028
rect 5348 34972 8092 35028
rect 8148 34972 8158 35028
rect 10444 34972 12348 35028
rect 12404 34972 12414 35028
rect 13570 34972 13580 35028
rect 13636 34972 14812 35028
rect 14868 34972 14878 35028
rect 15092 34972 17724 35028
rect 17780 34972 17790 35028
rect 18050 34972 18060 35028
rect 18116 34972 20244 35028
rect 20402 34972 20412 35028
rect 20468 34972 20972 35028
rect 21028 34972 22204 35028
rect 22260 34972 22270 35028
rect 22418 34972 22428 35028
rect 22484 34972 31836 35028
rect 31892 34972 31902 35028
rect 33404 34972 33964 35028
rect 34020 34972 34030 35028
rect 35970 34972 35980 35028
rect 36036 34972 36988 35028
rect 37044 34972 37054 35028
rect 37650 34972 37660 35028
rect 37716 34972 38220 35028
rect 38276 34972 38286 35028
rect 38780 34972 50428 35028
rect 50652 34972 53564 35028
rect 53620 34972 53630 35028
rect 54674 34972 54684 35028
rect 54740 34972 56140 35028
rect 56196 34972 56206 35028
rect 10444 34916 10500 34972
rect 15092 34916 15148 34972
rect 2706 34860 2716 34916
rect 2772 34860 3500 34916
rect 3556 34860 3566 34916
rect 3714 34860 3724 34916
rect 3780 34860 7756 34916
rect 7812 34860 7822 34916
rect 8418 34860 8428 34916
rect 8484 34860 10500 34916
rect 11442 34860 11452 34916
rect 11508 34860 13020 34916
rect 13076 34860 15148 34916
rect 15362 34860 15372 34916
rect 15428 34860 20524 34916
rect 20580 34860 20590 34916
rect 23762 34860 23772 34916
rect 23828 34860 25676 34916
rect 25732 34860 27692 34916
rect 27748 34860 27758 34916
rect 28018 34860 28028 34916
rect 28084 34860 28924 34916
rect 28980 34860 28990 34916
rect 29474 34860 29484 34916
rect 29540 34860 30156 34916
rect 30212 34860 30222 34916
rect 30370 34860 30380 34916
rect 30436 34860 30940 34916
rect 30996 34860 31500 34916
rect 31556 34860 31566 34916
rect 32274 34860 32284 34916
rect 32340 34860 39900 34916
rect 39956 34860 39966 34916
rect 41132 34860 48300 34916
rect 48356 34860 48366 34916
rect 0 34804 112 34832
rect 0 34748 6468 34804
rect 6626 34748 6636 34804
rect 6692 34748 7980 34804
rect 8036 34748 8046 34804
rect 8754 34748 8764 34804
rect 8820 34748 9324 34804
rect 9380 34748 9390 34804
rect 9958 34748 9996 34804
rect 10052 34748 10062 34804
rect 14802 34748 14812 34804
rect 14868 34748 19852 34804
rect 19908 34748 19918 34804
rect 20738 34748 20748 34804
rect 20804 34748 21532 34804
rect 21588 34748 25116 34804
rect 25172 34748 25182 34804
rect 25330 34748 25340 34804
rect 25396 34748 25452 34804
rect 25508 34748 25518 34804
rect 26852 34748 29260 34804
rect 29316 34748 31164 34804
rect 31220 34748 31230 34804
rect 32834 34748 32844 34804
rect 32900 34748 33180 34804
rect 33236 34748 33246 34804
rect 33618 34748 33628 34804
rect 33684 34748 34860 34804
rect 34916 34748 34926 34804
rect 35522 34748 35532 34804
rect 35588 34748 37156 34804
rect 38770 34748 38780 34804
rect 38836 34748 39676 34804
rect 39732 34748 39742 34804
rect 0 34720 112 34748
rect 6412 34692 6468 34748
rect 26852 34692 26908 34748
rect 37100 34692 37156 34748
rect 3612 34636 3724 34692
rect 3780 34636 3790 34692
rect 3938 34636 3948 34692
rect 4004 34636 5068 34692
rect 5124 34636 5134 34692
rect 6412 34636 13468 34692
rect 13524 34636 13534 34692
rect 13682 34636 13692 34692
rect 13748 34636 13916 34692
rect 13972 34636 13982 34692
rect 14130 34636 14140 34692
rect 14196 34636 15372 34692
rect 15428 34636 15438 34692
rect 15586 34636 15596 34692
rect 15652 34636 16716 34692
rect 16772 34636 16782 34692
rect 19058 34636 19068 34692
rect 19124 34636 19628 34692
rect 19684 34636 19694 34692
rect 23874 34636 23884 34692
rect 23940 34636 26908 34692
rect 27122 34636 27132 34692
rect 27188 34636 27244 34692
rect 27300 34636 27310 34692
rect 31938 34636 31948 34692
rect 32004 34636 36876 34692
rect 36932 34636 36942 34692
rect 37100 34636 40348 34692
rect 40404 34636 40414 34692
rect 40674 34636 40684 34692
rect 40740 34636 40750 34692
rect 3612 34468 3668 34636
rect 40684 34580 40740 34636
rect 4274 34524 4284 34580
rect 4340 34524 5292 34580
rect 5348 34524 5358 34580
rect 5842 34524 5852 34580
rect 5908 34524 6076 34580
rect 6132 34524 6142 34580
rect 6402 34524 6412 34580
rect 6468 34524 7756 34580
rect 7812 34524 7822 34580
rect 8418 34524 8428 34580
rect 8484 34524 12012 34580
rect 12068 34524 15708 34580
rect 15764 34524 16492 34580
rect 16548 34524 16558 34580
rect 16716 34524 21420 34580
rect 21476 34524 21486 34580
rect 24546 34524 24556 34580
rect 24612 34524 29820 34580
rect 29876 34524 38892 34580
rect 38948 34524 38958 34580
rect 39554 34524 39564 34580
rect 39620 34524 40740 34580
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 16716 34468 16772 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 3602 34412 3612 34468
rect 3668 34412 3678 34468
rect 4386 34412 4396 34468
rect 4452 34412 4956 34468
rect 5012 34412 8764 34468
rect 8820 34412 8830 34468
rect 8978 34412 8988 34468
rect 9044 34412 14252 34468
rect 14308 34412 14318 34468
rect 16146 34412 16156 34468
rect 16212 34412 16772 34468
rect 19058 34412 19068 34468
rect 19124 34412 19516 34468
rect 19572 34412 19582 34468
rect 19730 34412 19740 34468
rect 19796 34412 23436 34468
rect 23492 34412 23660 34468
rect 23716 34412 23726 34468
rect 24882 34412 24892 34468
rect 24948 34412 29372 34468
rect 29428 34412 29438 34468
rect 30594 34412 30604 34468
rect 30660 34412 31052 34468
rect 31108 34412 31118 34468
rect 31826 34412 31836 34468
rect 31892 34412 33740 34468
rect 33796 34412 33806 34468
rect 34290 34412 34300 34468
rect 34356 34412 34636 34468
rect 34692 34412 34702 34468
rect 35410 34412 35420 34468
rect 35476 34412 36540 34468
rect 36596 34412 36606 34468
rect 37314 34412 37324 34468
rect 37380 34412 38220 34468
rect 38276 34412 38286 34468
rect 40338 34412 40348 34468
rect 40404 34412 40684 34468
rect 40740 34412 40750 34468
rect 0 34356 112 34384
rect 41132 34356 41188 34860
rect 41682 34748 41692 34804
rect 41748 34748 44716 34804
rect 44772 34748 44782 34804
rect 46498 34748 46508 34804
rect 46564 34748 46732 34804
rect 46788 34748 46798 34804
rect 47282 34748 47292 34804
rect 47348 34748 50204 34804
rect 50260 34748 50270 34804
rect 50652 34692 50708 34972
rect 50866 34860 50876 34916
rect 50932 34860 55916 34916
rect 55972 34860 55982 34916
rect 57344 34804 57456 34832
rect 43250 34636 43260 34692
rect 43316 34636 46620 34692
rect 46676 34636 46686 34692
rect 46946 34636 46956 34692
rect 47012 34636 47404 34692
rect 47460 34636 47470 34692
rect 47618 34636 47628 34692
rect 47684 34636 50708 34692
rect 50764 34748 52780 34804
rect 52836 34748 53900 34804
rect 53956 34748 54348 34804
rect 54404 34748 54414 34804
rect 55010 34748 55020 34804
rect 55076 34748 56140 34804
rect 56196 34748 56206 34804
rect 57138 34748 57148 34804
rect 57204 34748 57456 34804
rect 50764 34580 50820 34748
rect 57344 34720 57456 34748
rect 51650 34636 51660 34692
rect 51716 34636 55916 34692
rect 55972 34636 55982 34692
rect 42018 34524 42028 34580
rect 42084 34524 43372 34580
rect 43428 34524 43438 34580
rect 45490 34524 45500 34580
rect 45556 34524 50316 34580
rect 50372 34524 50382 34580
rect 50754 34524 50764 34580
rect 50820 34524 50830 34580
rect 50988 34524 52108 34580
rect 52164 34524 52892 34580
rect 52948 34524 52958 34580
rect 43794 34468 43804 34524
rect 43860 34468 43908 34524
rect 43964 34468 44012 34524
rect 44068 34468 44078 34524
rect 41570 34412 41580 34468
rect 41636 34412 43260 34468
rect 43316 34412 43326 34468
rect 44492 34412 50652 34468
rect 50708 34412 50718 34468
rect 44492 34356 44548 34412
rect 0 34300 1036 34356
rect 1092 34300 1102 34356
rect 1484 34300 41188 34356
rect 41346 34300 41356 34356
rect 41412 34300 44548 34356
rect 45602 34300 45612 34356
rect 45668 34300 46956 34356
rect 47012 34300 47022 34356
rect 47170 34300 47180 34356
rect 47236 34300 47516 34356
rect 47572 34300 47582 34356
rect 0 34272 112 34300
rect 690 34076 700 34132
rect 756 34076 1260 34132
rect 1316 34076 1326 34132
rect 0 33908 112 33936
rect 1484 33908 1540 34300
rect 50988 34244 51044 34524
rect 57344 34356 57456 34384
rect 51762 34300 51772 34356
rect 51828 34300 57456 34356
rect 57344 34272 57456 34300
rect 2594 34188 2604 34244
rect 2660 34188 5516 34244
rect 5572 34188 5582 34244
rect 5852 34188 9772 34244
rect 9828 34188 9996 34244
rect 10052 34188 10062 34244
rect 10546 34188 10556 34244
rect 10612 34188 12460 34244
rect 12516 34188 14140 34244
rect 14196 34188 14206 34244
rect 15362 34188 15372 34244
rect 15428 34188 18060 34244
rect 18116 34188 18126 34244
rect 18274 34188 18284 34244
rect 18340 34188 24892 34244
rect 24948 34188 24958 34244
rect 26572 34188 26684 34244
rect 26740 34188 32284 34244
rect 32340 34188 32350 34244
rect 32498 34188 32508 34244
rect 32564 34188 33628 34244
rect 33684 34188 33694 34244
rect 34290 34188 34300 34244
rect 34356 34188 35308 34244
rect 35364 34188 35374 34244
rect 35634 34188 35644 34244
rect 35700 34188 35868 34244
rect 35924 34188 35934 34244
rect 36082 34188 36092 34244
rect 36148 34188 36764 34244
rect 36820 34188 36830 34244
rect 37762 34188 37772 34244
rect 37828 34188 38108 34244
rect 38164 34188 38174 34244
rect 38322 34188 38332 34244
rect 38388 34188 40796 34244
rect 40852 34188 40862 34244
rect 41794 34188 41804 34244
rect 41860 34188 46340 34244
rect 46498 34188 46508 34244
rect 46564 34188 46956 34244
rect 47012 34188 47022 34244
rect 47282 34188 47292 34244
rect 47348 34188 47964 34244
rect 48020 34188 48030 34244
rect 48290 34188 48300 34244
rect 48356 34188 48860 34244
rect 48916 34188 49532 34244
rect 49588 34188 49598 34244
rect 50642 34188 50652 34244
rect 50708 34188 51044 34244
rect 52546 34188 52556 34244
rect 52612 34188 52892 34244
rect 52948 34188 55692 34244
rect 55748 34188 55758 34244
rect 5852 34132 5908 34188
rect 26572 34132 26628 34188
rect 46284 34132 46340 34188
rect 3042 34076 3052 34132
rect 3108 34076 3948 34132
rect 4004 34076 4014 34132
rect 4274 34076 4284 34132
rect 4340 34076 5908 34132
rect 6066 34076 6076 34132
rect 6132 34076 6142 34132
rect 6290 34076 6300 34132
rect 6356 34076 6692 34132
rect 8082 34076 8092 34132
rect 8148 34076 11004 34132
rect 11060 34076 11070 34132
rect 13682 34076 13692 34132
rect 13748 34076 14252 34132
rect 14308 34076 14318 34132
rect 14578 34076 14588 34132
rect 14644 34076 14812 34132
rect 14868 34076 14878 34132
rect 15092 34076 17052 34132
rect 17108 34076 17118 34132
rect 18610 34076 18620 34132
rect 18676 34076 18844 34132
rect 18900 34076 19628 34132
rect 19684 34076 19694 34132
rect 19954 34076 19964 34132
rect 20020 34076 20524 34132
rect 20580 34076 20590 34132
rect 20850 34076 20860 34132
rect 20916 34076 21756 34132
rect 21812 34076 21822 34132
rect 22866 34076 22876 34132
rect 22932 34076 26628 34132
rect 26786 34076 26796 34132
rect 26852 34076 30268 34132
rect 30324 34076 30334 34132
rect 30930 34076 30940 34132
rect 30996 34076 32060 34132
rect 32116 34076 33292 34132
rect 33348 34076 33358 34132
rect 33730 34076 33740 34132
rect 33796 34076 34524 34132
rect 34580 34076 39004 34132
rect 39060 34076 39070 34132
rect 40310 34076 40348 34132
rect 40404 34076 40414 34132
rect 40898 34076 40908 34132
rect 40964 34076 44380 34132
rect 44436 34076 44446 34132
rect 44818 34076 44828 34132
rect 44884 34076 46060 34132
rect 46116 34076 46126 34132
rect 46284 34076 46396 34132
rect 46452 34076 46462 34132
rect 47842 34076 47852 34132
rect 47908 34076 48076 34132
rect 48132 34076 48142 34132
rect 51874 34076 51884 34132
rect 51940 34076 53228 34132
rect 53284 34076 53294 34132
rect 53554 34076 53564 34132
rect 53620 34076 54124 34132
rect 54180 34076 54190 34132
rect 54338 34076 54348 34132
rect 54404 34076 55244 34132
rect 55300 34076 55310 34132
rect 6076 34020 6132 34076
rect 6636 34020 6692 34076
rect 15092 34020 15148 34076
rect 2482 33964 2492 34020
rect 2548 33964 4116 34020
rect 4386 33964 4396 34020
rect 4452 33964 5292 34020
rect 5348 33964 5358 34020
rect 6076 33964 6412 34020
rect 6468 33964 6478 34020
rect 6636 33964 8428 34020
rect 8484 33964 8494 34020
rect 9090 33964 9100 34020
rect 9156 33964 15148 34020
rect 15260 33964 17388 34020
rect 17444 33964 17454 34020
rect 18498 33964 18508 34020
rect 18564 33964 20748 34020
rect 20804 33964 20814 34020
rect 21634 33964 21644 34020
rect 21700 33964 23268 34020
rect 23426 33964 23436 34020
rect 23492 33964 24892 34020
rect 24948 33964 24958 34020
rect 28802 33964 28812 34020
rect 28868 33964 32508 34020
rect 32564 33964 32574 34020
rect 33842 33964 33852 34020
rect 33908 33964 36316 34020
rect 36372 33964 36382 34020
rect 37426 33964 37436 34020
rect 37492 33964 39676 34020
rect 39732 33964 39742 34020
rect 43026 33964 43036 34020
rect 43092 33964 46284 34020
rect 46340 33964 46350 34020
rect 47282 33964 47292 34020
rect 47348 33964 47684 34020
rect 48598 33964 48636 34020
rect 48692 33964 48702 34020
rect 50754 33964 50764 34020
rect 50820 33964 50830 34020
rect 50978 33964 50988 34020
rect 51044 33964 52836 34020
rect 52994 33964 53004 34020
rect 53060 33964 54012 34020
rect 54068 33964 54078 34020
rect 54450 33964 54460 34020
rect 54516 33964 55020 34020
rect 55076 33964 55086 34020
rect 4060 33908 4116 33964
rect 15260 33908 15316 33964
rect 23212 33908 23268 33964
rect 47628 33908 47684 33964
rect 50764 33908 50820 33964
rect 0 33852 1540 33908
rect 1698 33852 1708 33908
rect 1764 33852 1932 33908
rect 1988 33852 3836 33908
rect 3892 33852 3902 33908
rect 4060 33852 7196 33908
rect 7252 33852 7262 33908
rect 7420 33852 9996 33908
rect 10052 33852 10062 33908
rect 10966 33852 11004 33908
rect 11060 33852 11070 33908
rect 11778 33852 11788 33908
rect 11844 33852 13356 33908
rect 13412 33852 15316 33908
rect 15586 33852 15596 33908
rect 15652 33852 22876 33908
rect 22932 33852 22942 33908
rect 23212 33852 23884 33908
rect 23940 33852 23950 33908
rect 24098 33852 24108 33908
rect 24164 33852 26908 33908
rect 27010 33852 27020 33908
rect 27076 33852 27356 33908
rect 27412 33852 27422 33908
rect 27570 33852 27580 33908
rect 27636 33852 31836 33908
rect 31892 33852 32844 33908
rect 32900 33852 32910 33908
rect 33058 33852 33068 33908
rect 33124 33852 33628 33908
rect 33684 33852 33694 33908
rect 35298 33852 35308 33908
rect 35364 33852 36092 33908
rect 36148 33852 36158 33908
rect 36866 33852 36876 33908
rect 36932 33852 37212 33908
rect 37268 33852 37884 33908
rect 37940 33852 37950 33908
rect 38098 33852 38108 33908
rect 38164 33852 38500 33908
rect 38994 33852 39004 33908
rect 39060 33852 40460 33908
rect 40516 33852 40526 33908
rect 42364 33852 47180 33908
rect 47236 33852 47246 33908
rect 47618 33852 47628 33908
rect 47684 33852 47694 33908
rect 49858 33852 49868 33908
rect 49924 33852 50820 33908
rect 52780 33908 52836 33964
rect 57344 33908 57456 33936
rect 52780 33852 53788 33908
rect 53844 33852 53854 33908
rect 56354 33852 56364 33908
rect 56420 33852 57456 33908
rect 0 33824 112 33852
rect 7420 33796 7476 33852
rect 26852 33796 26908 33852
rect 38444 33796 38500 33852
rect 2258 33740 2268 33796
rect 2324 33740 3500 33796
rect 3556 33740 4284 33796
rect 4340 33740 4350 33796
rect 4834 33740 4844 33796
rect 4900 33740 5740 33796
rect 5796 33740 7476 33796
rect 7746 33740 7756 33796
rect 7812 33740 8652 33796
rect 8708 33740 8718 33796
rect 9874 33740 9884 33796
rect 9940 33740 14028 33796
rect 14084 33740 14094 33796
rect 14242 33740 14252 33796
rect 14308 33740 15372 33796
rect 15428 33740 15438 33796
rect 15586 33740 15596 33796
rect 15652 33740 16828 33796
rect 16884 33740 16894 33796
rect 17154 33740 17164 33796
rect 17220 33740 17612 33796
rect 17668 33740 18956 33796
rect 19012 33740 19022 33796
rect 19842 33740 19852 33796
rect 19908 33740 20188 33796
rect 20244 33740 20254 33796
rect 20626 33740 20636 33796
rect 20692 33740 24332 33796
rect 24388 33740 24398 33796
rect 24882 33740 24892 33796
rect 24948 33740 25116 33796
rect 25172 33740 25182 33796
rect 26852 33740 27132 33796
rect 27188 33740 27198 33796
rect 30156 33740 38108 33796
rect 38164 33740 38174 33796
rect 38434 33740 38444 33796
rect 38500 33740 38510 33796
rect 38882 33740 38892 33796
rect 38948 33740 40236 33796
rect 40292 33740 41244 33796
rect 41300 33740 41310 33796
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 1810 33628 1820 33684
rect 1876 33628 4340 33684
rect 5282 33628 5292 33684
rect 5348 33628 6524 33684
rect 6580 33628 6590 33684
rect 11788 33628 21868 33684
rect 21924 33628 21934 33684
rect 24892 33628 27580 33684
rect 27636 33628 27646 33684
rect 28242 33628 28252 33684
rect 28308 33628 28476 33684
rect 28532 33628 28542 33684
rect 28914 33628 28924 33684
rect 28980 33628 29484 33684
rect 29540 33628 29550 33684
rect 4284 33572 4340 33628
rect 1362 33516 1372 33572
rect 1428 33516 2716 33572
rect 2772 33516 2782 33572
rect 3154 33516 3164 33572
rect 3220 33516 3948 33572
rect 4004 33516 4014 33572
rect 4284 33516 5404 33572
rect 5460 33516 5470 33572
rect 5618 33516 5628 33572
rect 5684 33516 10780 33572
rect 10836 33516 10846 33572
rect 0 33460 112 33488
rect 0 33404 1652 33460
rect 2006 33404 2044 33460
rect 2100 33404 2110 33460
rect 2482 33404 2492 33460
rect 2548 33404 2828 33460
rect 2884 33404 6636 33460
rect 6692 33404 6702 33460
rect 7522 33404 7532 33460
rect 7588 33404 9884 33460
rect 9940 33404 9950 33460
rect 0 33376 112 33404
rect 1596 33236 1652 33404
rect 4722 33292 4732 33348
rect 4788 33292 7084 33348
rect 7140 33292 7150 33348
rect 7970 33292 7980 33348
rect 8036 33292 11452 33348
rect 11508 33292 11518 33348
rect 4060 33236 4564 33238
rect 11788 33236 11844 33628
rect 24892 33572 24948 33628
rect 30156 33572 30212 33740
rect 42364 33684 42420 33852
rect 57344 33824 57456 33852
rect 43362 33740 43372 33796
rect 43428 33740 44268 33796
rect 44324 33740 44334 33796
rect 45042 33740 45052 33796
rect 45108 33740 45836 33796
rect 45892 33740 46956 33796
rect 47012 33740 47022 33796
rect 47954 33740 47964 33796
rect 48020 33740 50932 33796
rect 51090 33740 51100 33796
rect 51156 33740 51194 33796
rect 44454 33684 44464 33740
rect 44520 33684 44568 33740
rect 44624 33684 44672 33740
rect 44728 33684 44738 33740
rect 30482 33628 30492 33684
rect 30548 33628 37324 33684
rect 37380 33628 37390 33684
rect 37762 33628 37772 33684
rect 37828 33628 39340 33684
rect 39396 33628 39406 33684
rect 39666 33628 39676 33684
rect 39732 33628 42420 33684
rect 43250 33628 43260 33684
rect 43316 33628 44324 33684
rect 44818 33628 44828 33684
rect 44884 33628 47292 33684
rect 47348 33628 47358 33684
rect 47842 33628 47852 33684
rect 47908 33628 47964 33684
rect 48020 33628 48030 33684
rect 49970 33628 49980 33684
rect 50036 33628 50540 33684
rect 50596 33628 50606 33684
rect 50876 33628 50932 33740
rect 52770 33628 52780 33684
rect 52836 33628 53116 33684
rect 53172 33628 53182 33684
rect 53330 33628 53340 33684
rect 53396 33628 53844 33684
rect 56578 33628 56588 33684
rect 56644 33628 57372 33684
rect 57428 33628 57438 33684
rect 44268 33572 44324 33628
rect 47506 33572 47516 33628
rect 47572 33572 47628 33628
rect 47684 33572 47694 33628
rect 50866 33572 50876 33628
rect 50932 33572 50942 33628
rect 12114 33516 12124 33572
rect 12180 33516 13244 33572
rect 13300 33516 13310 33572
rect 13878 33516 13916 33572
rect 13972 33516 13982 33572
rect 16034 33516 16044 33572
rect 16100 33516 22652 33572
rect 22708 33516 24948 33572
rect 25106 33516 25116 33572
rect 25172 33516 30212 33572
rect 30370 33516 30380 33572
rect 30436 33516 30604 33572
rect 30660 33516 30670 33572
rect 31154 33516 31164 33572
rect 31220 33516 31500 33572
rect 31556 33516 31566 33572
rect 33058 33516 33068 33572
rect 33124 33516 33516 33572
rect 33572 33516 33582 33572
rect 34402 33516 34412 33572
rect 34468 33516 43932 33572
rect 43988 33516 43998 33572
rect 44268 33516 45052 33572
rect 45108 33516 45118 33572
rect 45602 33516 45612 33572
rect 45668 33516 45948 33572
rect 46004 33516 46014 33572
rect 46386 33516 46396 33572
rect 46452 33516 46732 33572
rect 46788 33516 46798 33572
rect 48402 33516 48412 33572
rect 48468 33516 48636 33572
rect 48692 33516 48702 33572
rect 49298 33516 49308 33572
rect 49364 33516 49420 33572
rect 49476 33516 49486 33572
rect 49858 33516 49868 33572
rect 49924 33516 50540 33572
rect 50596 33516 50606 33572
rect 51090 33516 51100 33572
rect 51156 33516 51436 33572
rect 51492 33516 51502 33572
rect 51650 33516 51660 33572
rect 51716 33516 51884 33572
rect 51940 33516 51950 33572
rect 52210 33516 52220 33572
rect 52276 33516 52286 33572
rect 30380 33460 30436 33516
rect 52220 33460 52276 33516
rect 53788 33460 53844 33628
rect 57344 33460 57456 33488
rect 13794 33404 13804 33460
rect 13860 33404 15372 33460
rect 15428 33404 15438 33460
rect 16482 33404 16492 33460
rect 16548 33404 19516 33460
rect 19572 33404 19582 33460
rect 19740 33404 21420 33460
rect 21476 33404 23212 33460
rect 23268 33404 23278 33460
rect 23874 33404 23884 33460
rect 23940 33404 30436 33460
rect 30706 33404 30716 33460
rect 30772 33404 35532 33460
rect 35588 33404 35598 33460
rect 36876 33404 37660 33460
rect 37716 33404 37726 33460
rect 38434 33404 38444 33460
rect 38500 33404 39956 33460
rect 40114 33404 40124 33460
rect 40180 33404 46900 33460
rect 47506 33404 47516 33460
rect 47572 33404 50204 33460
rect 50260 33404 50270 33460
rect 50642 33404 50652 33460
rect 50708 33404 51212 33460
rect 51268 33404 52276 33460
rect 52658 33404 52668 33460
rect 52724 33404 52892 33460
rect 52948 33404 52958 33460
rect 53778 33404 53788 33460
rect 53844 33404 53854 33460
rect 54226 33404 54236 33460
rect 54292 33404 57456 33460
rect 19740 33348 19796 33404
rect 36876 33348 36932 33404
rect 39900 33348 39956 33404
rect 13458 33292 13468 33348
rect 13524 33292 14924 33348
rect 14980 33292 14990 33348
rect 15138 33292 15148 33348
rect 15204 33292 16324 33348
rect 17378 33292 17388 33348
rect 17444 33292 19796 33348
rect 19954 33292 19964 33348
rect 20020 33292 21084 33348
rect 21140 33292 21150 33348
rect 21746 33292 21756 33348
rect 21812 33292 22540 33348
rect 22596 33292 25116 33348
rect 25172 33292 25182 33348
rect 26114 33292 26124 33348
rect 26180 33292 33516 33348
rect 33572 33292 33582 33348
rect 33842 33292 33852 33348
rect 33908 33292 36932 33348
rect 37090 33292 37100 33348
rect 37156 33292 38108 33348
rect 38164 33292 38174 33348
rect 38332 33292 39676 33348
rect 39732 33292 39742 33348
rect 39900 33292 40740 33348
rect 40898 33292 40908 33348
rect 40964 33292 41468 33348
rect 41524 33292 41534 33348
rect 42690 33292 42700 33348
rect 42756 33292 43596 33348
rect 43652 33292 43662 33348
rect 43922 33292 43932 33348
rect 43988 33292 44380 33348
rect 44436 33292 45836 33348
rect 45892 33292 45902 33348
rect 16268 33236 16324 33292
rect 21756 33236 21812 33292
rect 38332 33236 38388 33292
rect 1596 33182 11844 33236
rect 1596 33180 4116 33182
rect 4508 33180 11844 33182
rect 13244 33180 16044 33236
rect 16100 33180 16110 33236
rect 16268 33180 21812 33236
rect 21970 33180 21980 33236
rect 22036 33180 31052 33236
rect 31108 33180 31118 33236
rect 31826 33180 31836 33236
rect 31892 33180 38388 33236
rect 13244 33124 13300 33180
rect 40684 33124 40740 33292
rect 46844 33236 46900 33404
rect 57344 33376 57456 33404
rect 47058 33292 47068 33348
rect 47124 33292 48748 33348
rect 48804 33292 49084 33348
rect 49140 33292 49150 33348
rect 50082 33292 50092 33348
rect 50148 33292 52780 33348
rect 52836 33292 52846 33348
rect 53106 33292 53116 33348
rect 53172 33292 53900 33348
rect 53956 33292 53966 33348
rect 42690 33180 42700 33236
rect 42756 33180 46620 33236
rect 46676 33180 46686 33236
rect 46844 33180 49980 33236
rect 50036 33180 50046 33236
rect 50194 33180 50204 33236
rect 50260 33180 50652 33236
rect 50708 33180 50718 33236
rect 50866 33180 50876 33236
rect 50932 33180 55916 33236
rect 55972 33180 55982 33236
rect 1810 33068 1820 33124
rect 1876 33068 4060 33124
rect 4116 33068 4126 33124
rect 5058 33068 5068 33124
rect 5124 33068 5964 33124
rect 6020 33068 6030 33124
rect 8418 33068 8428 33124
rect 8484 33068 11004 33124
rect 11060 33068 12908 33124
rect 12964 33068 12974 33124
rect 13234 33068 13244 33124
rect 13300 33068 13310 33124
rect 14476 33068 18508 33124
rect 18564 33068 18574 33124
rect 20738 33068 20748 33124
rect 20804 33068 22988 33124
rect 23044 33068 23054 33124
rect 23650 33068 23660 33124
rect 23716 33068 25452 33124
rect 25508 33068 25518 33124
rect 25890 33068 25900 33124
rect 25956 33068 26572 33124
rect 26628 33068 26638 33124
rect 27906 33068 27916 33124
rect 27972 33068 31948 33124
rect 32004 33068 32014 33124
rect 33058 33068 33068 33124
rect 33124 33068 33516 33124
rect 33572 33068 33582 33124
rect 34178 33068 34188 33124
rect 34244 33068 34860 33124
rect 34916 33068 34926 33124
rect 36642 33068 36652 33124
rect 36708 33068 38892 33124
rect 38948 33068 38958 33124
rect 40684 33068 45332 33124
rect 45602 33068 45612 33124
rect 45668 33068 53004 33124
rect 53060 33068 53070 33124
rect 53330 33068 53340 33124
rect 53396 33068 54012 33124
rect 54068 33068 54078 33124
rect 0 33012 112 33040
rect 14476 33012 14532 33068
rect 45276 33012 45332 33068
rect 57344 33012 57456 33040
rect 0 32956 588 33012
rect 644 32956 654 33012
rect 1474 32956 1484 33012
rect 1540 32956 2044 33012
rect 2100 32956 2110 33012
rect 4274 32956 4284 33012
rect 4340 32956 4620 33012
rect 4676 32956 4686 33012
rect 4834 32956 4844 33012
rect 4900 32956 6636 33012
rect 6692 32956 6702 33012
rect 7074 32956 7084 33012
rect 7140 32956 8428 33012
rect 8484 32956 8494 33012
rect 8652 32956 10276 33012
rect 10546 32956 10556 33012
rect 10612 32956 11340 33012
rect 11396 32956 14532 33012
rect 15250 32956 15260 33012
rect 15316 32956 23548 33012
rect 24210 32956 24220 33012
rect 24276 32956 25004 33012
rect 25060 32956 25070 33012
rect 25330 32956 25340 33012
rect 25396 32956 40348 33012
rect 40404 32956 41244 33012
rect 41300 32956 41310 33012
rect 41570 32956 41580 33012
rect 41636 32956 41916 33012
rect 41972 32956 41982 33012
rect 42466 32956 42476 33012
rect 42532 32956 42700 33012
rect 42756 32956 43148 33012
rect 43204 32956 43214 33012
rect 44258 32956 44268 33012
rect 44324 32956 45052 33012
rect 45108 32956 45118 33012
rect 45276 32956 46228 33012
rect 46722 32956 46732 33012
rect 46788 32956 50652 33012
rect 50708 32956 50718 33012
rect 50978 32956 50988 33012
rect 51044 32956 51100 33012
rect 51156 32956 51166 33012
rect 52210 32956 52220 33012
rect 52276 32956 57456 33012
rect 0 32928 112 32956
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 8652 32900 8708 32956
rect 10220 32900 10276 32956
rect 4274 32844 4284 32900
rect 4340 32844 4396 32900
rect 4452 32844 4462 32900
rect 4732 32844 6860 32900
rect 6916 32844 8708 32900
rect 8866 32844 8876 32900
rect 8932 32844 10164 32900
rect 10220 32844 11340 32900
rect 11396 32844 11406 32900
rect 12002 32844 12012 32900
rect 12068 32844 20636 32900
rect 20692 32844 22876 32900
rect 22932 32844 22942 32900
rect 914 32732 924 32788
rect 980 32732 1484 32788
rect 1540 32732 1550 32788
rect 2594 32732 2604 32788
rect 2660 32732 3612 32788
rect 3668 32732 3678 32788
rect 4732 32676 4788 32844
rect 10108 32788 10164 32844
rect 23492 32788 23548 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 43794 32900 43804 32956
rect 43860 32900 43908 32956
rect 43964 32900 44012 32956
rect 44068 32900 44078 32956
rect 24882 32844 24892 32900
rect 24948 32844 26516 32900
rect 27570 32844 27580 32900
rect 27636 32844 39228 32900
rect 39284 32844 39294 32900
rect 41122 32844 41132 32900
rect 41188 32844 43372 32900
rect 43428 32844 43438 32900
rect 26460 32788 26516 32844
rect 46172 32788 46228 32956
rect 57344 32928 57456 32956
rect 46498 32844 46508 32900
rect 46564 32844 52276 32900
rect 52434 32844 52444 32900
rect 52500 32844 53900 32900
rect 53956 32844 53966 32900
rect 52220 32788 52276 32844
rect 7970 32732 7980 32788
rect 8036 32732 9212 32788
rect 9268 32732 9884 32788
rect 9940 32732 9950 32788
rect 10108 32732 15260 32788
rect 15316 32732 15326 32788
rect 15474 32732 15484 32788
rect 15540 32732 15708 32788
rect 15764 32732 15774 32788
rect 16930 32732 16940 32788
rect 16996 32732 18620 32788
rect 18676 32732 18686 32788
rect 18946 32732 18956 32788
rect 19012 32732 21868 32788
rect 21924 32732 22316 32788
rect 22372 32732 22382 32788
rect 23492 32732 25900 32788
rect 25956 32732 25966 32788
rect 26460 32732 30380 32788
rect 30436 32732 30604 32788
rect 30660 32732 30670 32788
rect 32386 32732 32396 32788
rect 32452 32732 34076 32788
rect 34132 32732 34142 32788
rect 35298 32732 35308 32788
rect 35364 32732 36204 32788
rect 36260 32732 36270 32788
rect 39106 32732 39116 32788
rect 39172 32732 44940 32788
rect 44996 32732 45006 32788
rect 45266 32732 45276 32788
rect 45332 32732 45948 32788
rect 46004 32732 46014 32788
rect 46172 32732 48188 32788
rect 48244 32732 48636 32788
rect 48692 32732 48702 32788
rect 49410 32732 49420 32788
rect 49476 32732 50260 32788
rect 50204 32676 50260 32732
rect 50652 32732 51436 32788
rect 51492 32732 51502 32788
rect 52220 32732 54684 32788
rect 54740 32732 54750 32788
rect 50652 32676 50708 32732
rect 1026 32620 1036 32676
rect 1092 32620 3948 32676
rect 4004 32620 4014 32676
rect 4162 32620 4172 32676
rect 4228 32620 4788 32676
rect 4956 32620 18284 32676
rect 18340 32620 18350 32676
rect 18834 32620 18844 32676
rect 18900 32620 21420 32676
rect 21476 32620 21644 32676
rect 21700 32620 21710 32676
rect 21858 32620 21868 32676
rect 21924 32620 27300 32676
rect 29362 32620 29372 32676
rect 29428 32620 33348 32676
rect 33506 32620 33516 32676
rect 33572 32620 34748 32676
rect 34804 32620 35196 32676
rect 35252 32620 35262 32676
rect 35830 32620 35868 32676
rect 35924 32620 35934 32676
rect 36642 32620 36652 32676
rect 36708 32620 36876 32676
rect 36932 32620 37996 32676
rect 38052 32620 38062 32676
rect 38210 32620 38220 32676
rect 38276 32620 47180 32676
rect 47236 32620 47246 32676
rect 49858 32620 49868 32676
rect 49924 32620 49980 32676
rect 50036 32620 50046 32676
rect 50204 32620 50708 32676
rect 51538 32620 51548 32676
rect 51604 32620 52388 32676
rect 52854 32620 52892 32676
rect 52948 32620 52958 32676
rect 0 32564 112 32592
rect 0 32508 924 32564
rect 980 32508 990 32564
rect 1138 32508 1148 32564
rect 1204 32508 4620 32564
rect 4676 32508 4686 32564
rect 0 32480 112 32508
rect 4956 32452 5012 32620
rect 27244 32564 27300 32620
rect 33292 32564 33348 32620
rect 52332 32564 52388 32620
rect 57344 32564 57456 32592
rect 5506 32508 5516 32564
rect 5572 32508 6524 32564
rect 6580 32508 6590 32564
rect 7186 32508 7196 32564
rect 7252 32508 8988 32564
rect 9044 32508 9212 32564
rect 9268 32508 9278 32564
rect 11414 32508 11452 32564
rect 11508 32508 11900 32564
rect 11956 32508 11966 32564
rect 12226 32508 12236 32564
rect 12292 32508 13916 32564
rect 13972 32508 14700 32564
rect 14756 32508 14766 32564
rect 15026 32508 15036 32564
rect 15092 32508 15820 32564
rect 15876 32508 15886 32564
rect 16230 32508 16268 32564
rect 16324 32508 16334 32564
rect 16594 32508 16604 32564
rect 16660 32508 16828 32564
rect 16884 32508 18508 32564
rect 18564 32508 18574 32564
rect 19506 32508 19516 32564
rect 19572 32508 24892 32564
rect 24948 32508 24958 32564
rect 27244 32508 31724 32564
rect 31780 32508 31790 32564
rect 32498 32508 32508 32564
rect 32564 32508 33068 32564
rect 33124 32508 33134 32564
rect 33292 32508 37436 32564
rect 37492 32508 37502 32564
rect 38210 32508 38220 32564
rect 38276 32508 41468 32564
rect 41524 32508 41534 32564
rect 43474 32508 43484 32564
rect 43540 32508 44268 32564
rect 44324 32508 44334 32564
rect 44482 32508 44492 32564
rect 44548 32508 44940 32564
rect 44996 32508 45612 32564
rect 45668 32508 45678 32564
rect 47282 32508 47292 32564
rect 47348 32508 50428 32564
rect 50484 32508 50494 32564
rect 51762 32508 51772 32564
rect 51828 32508 51884 32564
rect 51940 32508 51950 32564
rect 52332 32508 53564 32564
rect 53620 32508 53630 32564
rect 57026 32508 57036 32564
rect 57092 32508 57456 32564
rect 44492 32452 44548 32508
rect 57344 32480 57456 32508
rect 1250 32396 1260 32452
rect 1316 32396 1708 32452
rect 1764 32396 1774 32452
rect 3378 32396 3388 32452
rect 3444 32396 3612 32452
rect 3668 32396 3678 32452
rect 4050 32396 4060 32452
rect 4116 32396 5012 32452
rect 5954 32396 5964 32452
rect 6020 32396 7532 32452
rect 7588 32396 7980 32452
rect 8036 32396 8046 32452
rect 8418 32396 8428 32452
rect 8484 32396 9436 32452
rect 9492 32396 9502 32452
rect 9762 32396 9772 32452
rect 9828 32396 12236 32452
rect 12292 32396 12302 32452
rect 13458 32396 13468 32452
rect 13524 32396 14476 32452
rect 14532 32396 14542 32452
rect 16034 32396 16044 32452
rect 16100 32396 16940 32452
rect 16996 32396 17006 32452
rect 17350 32396 17388 32452
rect 17444 32396 17454 32452
rect 21270 32396 21308 32452
rect 21364 32396 25676 32452
rect 25732 32396 25742 32452
rect 27458 32396 27468 32452
rect 27524 32396 28140 32452
rect 28196 32396 28206 32452
rect 29362 32396 29372 32452
rect 29428 32396 32956 32452
rect 33012 32396 33022 32452
rect 33394 32396 33404 32452
rect 33460 32396 34300 32452
rect 34356 32396 34366 32452
rect 35270 32396 35308 32452
rect 35364 32396 35374 32452
rect 35858 32396 35868 32452
rect 35924 32396 36764 32452
rect 36820 32396 38780 32452
rect 38836 32396 38846 32452
rect 39218 32396 39228 32452
rect 39284 32396 43260 32452
rect 43316 32396 43326 32452
rect 43586 32396 43596 32452
rect 43652 32396 44548 32452
rect 44930 32396 44940 32452
rect 44996 32396 46508 32452
rect 46564 32396 46574 32452
rect 46722 32396 46732 32452
rect 46788 32396 46956 32452
rect 47012 32396 47022 32452
rect 50764 32396 55692 32452
rect 55748 32396 55758 32452
rect 50764 32340 50820 32396
rect 802 32284 812 32340
rect 868 32284 1372 32340
rect 1428 32284 1596 32340
rect 1652 32284 1662 32340
rect 3602 32284 3612 32340
rect 3668 32284 4172 32340
rect 4228 32284 4238 32340
rect 5506 32284 5516 32340
rect 5572 32284 5582 32340
rect 7074 32284 7084 32340
rect 7140 32284 7756 32340
rect 7812 32284 8204 32340
rect 8260 32284 8270 32340
rect 8418 32284 8428 32340
rect 8484 32284 13692 32340
rect 13748 32284 13758 32340
rect 13906 32284 13916 32340
rect 13972 32284 14140 32340
rect 14196 32284 14700 32340
rect 14756 32284 14766 32340
rect 14924 32284 15484 32340
rect 15540 32284 15550 32340
rect 16482 32284 16492 32340
rect 16548 32284 27356 32340
rect 27412 32284 27422 32340
rect 28914 32284 28924 32340
rect 28980 32284 29148 32340
rect 29204 32284 29214 32340
rect 29362 32284 29372 32340
rect 29428 32284 29708 32340
rect 29764 32284 29774 32340
rect 30034 32284 30044 32340
rect 30100 32284 37100 32340
rect 37156 32284 37166 32340
rect 37426 32284 37436 32340
rect 37492 32284 37548 32340
rect 37604 32284 37614 32340
rect 37986 32284 37996 32340
rect 38052 32284 40404 32340
rect 41346 32284 41356 32340
rect 41412 32284 44884 32340
rect 49186 32284 49196 32340
rect 49252 32284 50820 32340
rect 51538 32284 51548 32340
rect 51604 32284 54236 32340
rect 54292 32284 54302 32340
rect 55122 32284 55132 32340
rect 55188 32284 56476 32340
rect 56532 32284 56542 32340
rect 5516 32228 5572 32284
rect 14924 32228 14980 32284
rect 40348 32228 40404 32284
rect 2706 32172 2716 32228
rect 2772 32172 3836 32228
rect 3892 32172 3902 32228
rect 4844 32172 5572 32228
rect 7634 32172 7644 32228
rect 7700 32172 8764 32228
rect 8820 32172 9212 32228
rect 9268 32172 9278 32228
rect 9538 32172 9548 32228
rect 9604 32172 14980 32228
rect 15092 32172 23660 32228
rect 23716 32172 23726 32228
rect 24994 32172 25004 32228
rect 25060 32172 34860 32228
rect 34916 32172 34926 32228
rect 35298 32172 35308 32228
rect 35364 32172 38220 32228
rect 38276 32172 38286 32228
rect 38994 32172 39004 32228
rect 39060 32172 39116 32228
rect 39172 32172 39182 32228
rect 40348 32172 41580 32228
rect 41636 32172 41646 32228
rect 42242 32172 42252 32228
rect 42308 32172 44156 32228
rect 44212 32172 44222 32228
rect 0 32116 112 32144
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 0 32060 812 32116
rect 868 32060 878 32116
rect 2818 32060 2828 32116
rect 2884 32060 3500 32116
rect 3556 32060 3566 32116
rect 3938 32060 3948 32116
rect 4004 32060 4340 32116
rect 0 32032 112 32060
rect 4284 32004 4340 32060
rect 4844 32004 4900 32172
rect 9212 32116 9268 32172
rect 15092 32116 15148 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 44454 32116 44464 32172
rect 44520 32116 44568 32172
rect 44624 32116 44672 32172
rect 44728 32116 44738 32172
rect 44828 32116 44884 32284
rect 45042 32172 45052 32228
rect 45108 32172 46620 32228
rect 46676 32172 47964 32228
rect 48020 32172 48030 32228
rect 50082 32172 50092 32228
rect 50148 32172 50988 32228
rect 51044 32172 51436 32228
rect 51492 32172 53340 32228
rect 53396 32172 54012 32228
rect 54068 32172 55244 32228
rect 55300 32172 55310 32228
rect 57344 32116 57456 32144
rect 5282 32060 5292 32116
rect 5348 32060 6412 32116
rect 6468 32060 6478 32116
rect 7858 32060 7868 32116
rect 7924 32060 7980 32116
rect 8036 32060 8046 32116
rect 9212 32060 10332 32116
rect 10388 32060 10398 32116
rect 10882 32060 10892 32116
rect 10948 32060 15148 32116
rect 17462 32060 17500 32116
rect 17556 32060 17566 32116
rect 22866 32060 22876 32116
rect 22932 32060 23884 32116
rect 23940 32060 23950 32116
rect 26226 32060 26236 32116
rect 26292 32060 26572 32116
rect 26628 32060 30380 32116
rect 30436 32060 30446 32116
rect 30930 32060 30940 32116
rect 30996 32060 32676 32116
rect 33170 32060 33180 32116
rect 33236 32060 35644 32116
rect 35700 32060 35710 32116
rect 37314 32060 37324 32116
rect 37380 32060 39228 32116
rect 39284 32060 39294 32116
rect 39452 32060 43596 32116
rect 43652 32060 43662 32116
rect 44828 32060 50652 32116
rect 50708 32060 51884 32116
rect 51940 32060 51950 32116
rect 52546 32060 52556 32116
rect 52612 32060 54180 32116
rect 55346 32060 55356 32116
rect 55412 32060 55422 32116
rect 57250 32060 57260 32116
rect 57316 32060 57456 32116
rect 32620 32004 32676 32060
rect 39452 32004 39508 32060
rect 4284 31948 4900 32004
rect 5292 31948 5740 32004
rect 5796 31948 5806 32004
rect 6178 31948 6188 32004
rect 6244 31948 10780 32004
rect 10836 31948 11788 32004
rect 11890 31948 11900 32004
rect 11956 31948 12236 32004
rect 12292 31948 12302 32004
rect 12562 31948 12572 32004
rect 12628 31948 18452 32004
rect 21158 31948 21196 32004
rect 21252 31948 21262 32004
rect 24546 31948 24556 32004
rect 24612 31948 25676 32004
rect 25732 31948 25742 32004
rect 25890 31948 25900 32004
rect 25956 31948 28812 32004
rect 28868 31948 28878 32004
rect 29586 31948 29596 32004
rect 29652 31948 30492 32004
rect 30548 31948 30558 32004
rect 31602 31948 31612 32004
rect 31668 31948 32396 32004
rect 32452 31948 32462 32004
rect 32620 31948 39508 32004
rect 39666 31948 39676 32004
rect 39732 31948 41020 32004
rect 41076 31948 41086 32004
rect 45612 31948 47628 32004
rect 47684 31948 47694 32004
rect 50418 31948 50428 32004
rect 50484 31948 51548 32004
rect 51604 31948 51614 32004
rect 51762 31948 51772 32004
rect 51828 31948 52556 32004
rect 52612 31948 52622 32004
rect 53106 31948 53116 32004
rect 53172 31948 53788 32004
rect 53844 31948 53854 32004
rect 5292 31892 5348 31948
rect 11732 31892 11788 31948
rect 18396 31892 18452 31948
rect 45612 31892 45668 31948
rect 54124 31892 54180 32060
rect 354 31836 364 31892
rect 420 31836 2156 31892
rect 2212 31836 2222 31892
rect 3350 31836 3388 31892
rect 3444 31836 3454 31892
rect 3602 31836 3612 31892
rect 3668 31836 5348 31892
rect 5618 31836 5628 31892
rect 5684 31836 7308 31892
rect 7364 31836 7374 31892
rect 7970 31836 7980 31892
rect 8036 31836 9324 31892
rect 9380 31836 9390 31892
rect 9650 31836 9660 31892
rect 9716 31836 9726 31892
rect 11732 31836 13188 31892
rect 14914 31836 14924 31892
rect 14980 31836 15484 31892
rect 15540 31836 15550 31892
rect 16678 31836 16716 31892
rect 16772 31836 16782 31892
rect 18396 31836 21980 31892
rect 22036 31836 22046 31892
rect 22418 31836 22428 31892
rect 22484 31836 25228 31892
rect 25284 31836 25294 31892
rect 26226 31836 26236 31892
rect 26292 31836 26572 31892
rect 26628 31836 32060 31892
rect 32116 31836 32126 31892
rect 32946 31836 32956 31892
rect 33012 31836 33068 31892
rect 33124 31836 33134 31892
rect 34962 31836 34972 31892
rect 35028 31836 35532 31892
rect 35588 31836 35598 31892
rect 36530 31836 36540 31892
rect 36596 31836 36876 31892
rect 36932 31836 36942 31892
rect 37324 31836 38892 31892
rect 38948 31836 38958 31892
rect 39330 31836 39340 31892
rect 39396 31836 40908 31892
rect 40964 31836 40974 31892
rect 43586 31836 43596 31892
rect 43652 31836 44436 31892
rect 45378 31836 45388 31892
rect 45444 31836 45668 31892
rect 47058 31836 47068 31892
rect 47124 31836 51772 31892
rect 51828 31836 51838 31892
rect 52322 31836 52332 31892
rect 52388 31836 53732 31892
rect 54086 31836 54124 31892
rect 54180 31836 54190 31892
rect 9660 31780 9716 31836
rect 13132 31780 13188 31836
rect 37324 31780 37380 31836
rect 44380 31780 44436 31836
rect 53676 31780 53732 31836
rect 55356 31780 55412 32060
rect 57344 32032 57456 32060
rect 3266 31724 3276 31780
rect 3332 31724 3612 31780
rect 3668 31724 3678 31780
rect 4274 31724 4284 31780
rect 4340 31724 4378 31780
rect 4834 31724 4844 31780
rect 4900 31724 5180 31780
rect 5236 31724 9716 31780
rect 9874 31724 9884 31780
rect 9940 31724 12012 31780
rect 12068 31724 12078 31780
rect 12338 31724 12348 31780
rect 12404 31724 12908 31780
rect 12964 31724 12974 31780
rect 13122 31724 13132 31780
rect 13188 31724 13916 31780
rect 13972 31724 17836 31780
rect 17892 31724 17902 31780
rect 18246 31724 18284 31780
rect 18340 31724 18350 31780
rect 18956 31724 23100 31780
rect 23156 31724 23166 31780
rect 23874 31724 23884 31780
rect 23940 31724 26908 31780
rect 26964 31724 26974 31780
rect 28914 31724 28924 31780
rect 28980 31724 34636 31780
rect 34692 31724 34702 31780
rect 35298 31724 35308 31780
rect 35364 31724 37380 31780
rect 37650 31724 37660 31780
rect 37716 31724 37996 31780
rect 38052 31724 38062 31780
rect 38658 31724 38668 31780
rect 38724 31724 39340 31780
rect 39396 31724 39406 31780
rect 41122 31724 41132 31780
rect 41188 31724 41692 31780
rect 41748 31724 42028 31780
rect 42084 31724 42094 31780
rect 42466 31724 42476 31780
rect 42532 31724 43260 31780
rect 43316 31724 43326 31780
rect 44380 31724 45836 31780
rect 45892 31724 45948 31780
rect 46004 31724 46014 31780
rect 47506 31724 47516 31780
rect 47572 31724 48412 31780
rect 48468 31724 48478 31780
rect 50418 31724 50428 31780
rect 50484 31724 53452 31780
rect 53508 31724 53518 31780
rect 53676 31724 55412 31780
rect 0 31668 112 31696
rect 18956 31668 19012 31724
rect 57344 31668 57456 31696
rect 0 31612 9604 31668
rect 10294 31612 10332 31668
rect 10388 31612 10398 31668
rect 12226 31612 12236 31668
rect 12292 31612 18732 31668
rect 18788 31612 19012 31668
rect 23538 31612 23548 31668
rect 23604 31612 24668 31668
rect 24724 31612 24734 31668
rect 26002 31612 26012 31668
rect 26068 31612 27916 31668
rect 27972 31612 27982 31668
rect 28690 31612 28700 31668
rect 28756 31612 29484 31668
rect 29540 31612 29550 31668
rect 32050 31612 32060 31668
rect 32116 31612 32956 31668
rect 33012 31612 33022 31668
rect 36306 31612 36316 31668
rect 36372 31612 36428 31668
rect 36484 31612 36494 31668
rect 36866 31612 36876 31668
rect 36932 31612 49084 31668
rect 49140 31612 49150 31668
rect 49634 31612 49644 31668
rect 49700 31612 50316 31668
rect 50372 31612 50382 31668
rect 50540 31612 51100 31668
rect 51156 31612 51166 31668
rect 51314 31612 51324 31668
rect 51380 31612 52220 31668
rect 52276 31612 52286 31668
rect 52770 31612 52780 31668
rect 52836 31612 54348 31668
rect 54404 31612 54414 31668
rect 57138 31612 57148 31668
rect 57204 31612 57456 31668
rect 0 31584 112 31612
rect 9548 31556 9604 31612
rect 50540 31556 50596 31612
rect 57344 31584 57456 31612
rect 3154 31500 3164 31556
rect 3220 31500 5180 31556
rect 5236 31500 5246 31556
rect 5506 31500 5516 31556
rect 5572 31500 7644 31556
rect 7700 31500 7710 31556
rect 7970 31500 7980 31556
rect 8036 31500 8316 31556
rect 8372 31500 8382 31556
rect 9548 31500 12572 31556
rect 12628 31500 12638 31556
rect 19170 31500 19180 31556
rect 19236 31500 20748 31556
rect 20804 31500 20814 31556
rect 21308 31500 44324 31556
rect 44482 31500 44492 31556
rect 44548 31500 46620 31556
rect 46676 31500 47404 31556
rect 47460 31500 47470 31556
rect 47842 31500 47852 31556
rect 47908 31500 48300 31556
rect 48356 31500 48524 31556
rect 48580 31500 48590 31556
rect 50194 31500 50204 31556
rect 50260 31500 50596 31556
rect 50754 31500 50764 31556
rect 50820 31500 51548 31556
rect 51604 31500 51614 31556
rect 51762 31500 51772 31556
rect 51828 31500 56028 31556
rect 56084 31500 56094 31556
rect 21308 31444 21364 31500
rect 44268 31444 44324 31500
rect 700 31388 3612 31444
rect 3668 31388 3678 31444
rect 4274 31388 4284 31444
rect 4340 31388 5068 31444
rect 5124 31388 5134 31444
rect 6178 31388 6188 31444
rect 6244 31388 6300 31444
rect 6356 31388 6366 31444
rect 8194 31388 8204 31444
rect 8260 31388 9548 31444
rect 9604 31388 9614 31444
rect 9986 31388 9996 31444
rect 10052 31388 12124 31444
rect 12180 31388 12190 31444
rect 12674 31388 12684 31444
rect 12740 31388 14252 31444
rect 14308 31388 14318 31444
rect 15092 31388 21364 31444
rect 24882 31388 24892 31444
rect 24948 31388 26124 31444
rect 26180 31388 26190 31444
rect 29026 31388 29036 31444
rect 29092 31388 29484 31444
rect 29540 31388 32172 31444
rect 32228 31388 32238 31444
rect 32834 31388 32844 31444
rect 32900 31388 34076 31444
rect 34132 31388 34142 31444
rect 34738 31388 34748 31444
rect 34804 31388 35420 31444
rect 35476 31388 35644 31444
rect 35700 31388 37884 31444
rect 37940 31388 37950 31444
rect 38098 31388 38108 31444
rect 38164 31388 38780 31444
rect 38836 31388 38846 31444
rect 40226 31388 40236 31444
rect 40292 31388 43260 31444
rect 43316 31388 43326 31444
rect 44268 31388 49196 31444
rect 49252 31388 49262 31444
rect 49410 31388 49420 31444
rect 49476 31388 51156 31444
rect 51874 31388 51884 31444
rect 51940 31388 53060 31444
rect 54338 31388 54348 31444
rect 54404 31388 54460 31444
rect 54516 31388 54526 31444
rect 0 31220 112 31248
rect 700 31220 756 31388
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 12684 31332 12740 31388
rect 3042 31276 3052 31332
rect 3108 31276 3612 31332
rect 3668 31276 3678 31332
rect 4498 31276 4508 31332
rect 4564 31276 6076 31332
rect 6132 31276 6142 31332
rect 6962 31276 6972 31332
rect 7028 31276 8540 31332
rect 8596 31276 8606 31332
rect 8866 31276 8876 31332
rect 8932 31276 9100 31332
rect 9156 31276 9166 31332
rect 10770 31276 10780 31332
rect 10836 31276 12740 31332
rect 13010 31276 13020 31332
rect 13076 31276 14588 31332
rect 14644 31276 14654 31332
rect 15092 31220 15148 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 43794 31332 43804 31388
rect 43860 31332 43908 31388
rect 43964 31332 44012 31388
rect 44068 31332 44078 31388
rect 51100 31332 51156 31388
rect 53004 31332 53060 31388
rect 16930 31276 16940 31332
rect 16996 31276 17836 31332
rect 17892 31276 17902 31332
rect 20626 31276 20636 31332
rect 20692 31276 23660 31332
rect 23716 31276 23726 31332
rect 27020 31276 29596 31332
rect 29652 31276 29662 31332
rect 29810 31276 29820 31332
rect 29876 31276 33740 31332
rect 33796 31276 35308 31332
rect 35364 31276 35374 31332
rect 35746 31276 35756 31332
rect 35812 31276 38444 31332
rect 38500 31276 38510 31332
rect 44146 31276 44156 31332
rect 44212 31276 45500 31332
rect 45556 31276 45566 31332
rect 45826 31276 45836 31332
rect 45892 31276 49588 31332
rect 49746 31276 49756 31332
rect 49812 31276 50764 31332
rect 50820 31276 50830 31332
rect 51100 31276 52780 31332
rect 52836 31276 52846 31332
rect 52994 31276 53004 31332
rect 53060 31276 53070 31332
rect 53218 31276 53228 31332
rect 53284 31276 54236 31332
rect 54292 31276 54302 31332
rect 27020 31220 27076 31276
rect 0 31164 756 31220
rect 914 31164 924 31220
rect 980 31164 15148 31220
rect 17938 31164 17948 31220
rect 18004 31164 18844 31220
rect 18900 31164 18910 31220
rect 20514 31164 20524 31220
rect 20580 31164 21420 31220
rect 21476 31164 21486 31220
rect 22418 31164 22428 31220
rect 22484 31164 24556 31220
rect 24612 31164 24622 31220
rect 25554 31164 25564 31220
rect 25620 31164 26124 31220
rect 26180 31164 26190 31220
rect 26898 31164 26908 31220
rect 26964 31164 27076 31220
rect 27244 31164 27916 31220
rect 27972 31164 29260 31220
rect 29316 31164 30156 31220
rect 30212 31164 30222 31220
rect 30706 31164 30716 31220
rect 30772 31164 33068 31220
rect 33124 31164 33134 31220
rect 33618 31164 33628 31220
rect 33684 31164 34244 31220
rect 35074 31164 35084 31220
rect 35140 31164 37100 31220
rect 37156 31164 37166 31220
rect 37426 31164 37436 31220
rect 37492 31164 37884 31220
rect 37940 31164 37950 31220
rect 38612 31164 42084 31220
rect 42242 31164 42252 31220
rect 42308 31164 43484 31220
rect 43540 31164 47292 31220
rect 47348 31164 47358 31220
rect 47506 31164 47516 31220
rect 47572 31164 48300 31220
rect 48356 31164 48366 31220
rect 48514 31164 48524 31220
rect 48580 31164 49308 31220
rect 49364 31164 49374 31220
rect 0 31136 112 31164
rect 27244 31108 27300 31164
rect 34188 31108 34244 31164
rect 38612 31108 38668 31164
rect 3388 31052 4508 31108
rect 4564 31052 4574 31108
rect 4722 31052 4732 31108
rect 4788 31052 5068 31108
rect 5124 31052 5134 31108
rect 6178 31052 6188 31108
rect 6244 31052 6412 31108
rect 6468 31052 6478 31108
rect 7298 31052 7308 31108
rect 7364 31052 20188 31108
rect 20244 31052 20254 31108
rect 20850 31052 20860 31108
rect 20916 31052 21756 31108
rect 21812 31052 21822 31108
rect 22642 31052 22652 31108
rect 22708 31052 26460 31108
rect 26516 31052 26526 31108
rect 26786 31052 26796 31108
rect 26852 31052 27300 31108
rect 28354 31052 28364 31108
rect 28420 31052 30380 31108
rect 30436 31052 30446 31108
rect 32386 31052 32396 31108
rect 32452 31052 33964 31108
rect 34020 31052 34030 31108
rect 34188 31052 38668 31108
rect 3388 30996 3444 31052
rect 42028 30996 42084 31164
rect 49532 31108 49588 31276
rect 57344 31220 57456 31248
rect 49858 31164 49868 31220
rect 49924 31164 51156 31220
rect 51314 31164 51324 31220
rect 51380 31164 51884 31220
rect 51940 31164 54796 31220
rect 54852 31164 54862 31220
rect 56914 31164 56924 31220
rect 56980 31164 57456 31220
rect 51100 31108 51156 31164
rect 57344 31136 57456 31164
rect 44146 31052 44156 31108
rect 44212 31052 48804 31108
rect 49046 31052 49084 31108
rect 49140 31052 49150 31108
rect 49532 31052 50764 31108
rect 50820 31052 50830 31108
rect 51100 31052 53676 31108
rect 53732 31052 53742 31108
rect 3266 30940 3276 30996
rect 3332 30940 3444 30996
rect 3938 30940 3948 30996
rect 4004 30940 5292 30996
rect 5348 30940 5358 30996
rect 5954 30940 5964 30996
rect 6020 30940 7196 30996
rect 7252 30940 7262 30996
rect 8530 30940 8540 30996
rect 8596 30940 9212 30996
rect 9268 30940 9278 30996
rect 9874 30940 9884 30996
rect 9940 30940 10220 30996
rect 10276 30940 10286 30996
rect 10434 30940 10444 30996
rect 10500 30940 14140 30996
rect 14196 30940 14206 30996
rect 14354 30940 14364 30996
rect 14420 30940 16940 30996
rect 16996 30940 17500 30996
rect 17556 30940 17566 30996
rect 17714 30940 17724 30996
rect 17780 30940 18396 30996
rect 18452 30940 18844 30996
rect 18900 30940 18910 30996
rect 19842 30940 19852 30996
rect 19908 30940 22092 30996
rect 22148 30940 22158 30996
rect 23062 30940 23100 30996
rect 23156 30940 23166 30996
rect 23650 30940 23660 30996
rect 23716 30940 23884 30996
rect 23940 30940 23950 30996
rect 25218 30940 25228 30996
rect 25284 30940 25452 30996
rect 25508 30940 25518 30996
rect 27132 30940 27468 30996
rect 27524 30940 28028 30996
rect 28084 30940 28094 30996
rect 29138 30940 29148 30996
rect 29204 30940 29820 30996
rect 29876 30940 29886 30996
rect 30034 30940 30044 30996
rect 30100 30940 30138 30996
rect 31154 30940 31164 30996
rect 31220 30940 32284 30996
rect 32340 30940 32350 30996
rect 32694 30940 32732 30996
rect 32788 30940 32798 30996
rect 35252 30940 37100 30996
rect 37156 30940 37166 30996
rect 37314 30940 37324 30996
rect 37380 30940 38220 30996
rect 38276 30940 38286 30996
rect 40450 30940 40460 30996
rect 40516 30940 41132 30996
rect 41188 30940 41198 30996
rect 42028 30940 45612 30996
rect 45668 30940 45678 30996
rect 47030 30940 47068 30996
rect 47124 30940 47134 30996
rect 47618 30940 47628 30996
rect 47684 30940 48524 30996
rect 48580 30940 48590 30996
rect 3602 30828 3612 30884
rect 3668 30828 10668 30884
rect 10724 30828 11788 30884
rect 13094 30828 13132 30884
rect 13188 30828 13198 30884
rect 13346 30828 13356 30884
rect 13412 30828 16828 30884
rect 16884 30828 16894 30884
rect 19618 30828 19628 30884
rect 19684 30828 20076 30884
rect 20132 30828 20142 30884
rect 20290 30828 20300 30884
rect 20356 30828 21532 30884
rect 21588 30828 24892 30884
rect 24948 30828 24958 30884
rect 25106 30828 25116 30884
rect 25172 30828 25564 30884
rect 25620 30828 25630 30884
rect 0 30772 112 30800
rect 11732 30772 11788 30828
rect 27132 30772 27188 30940
rect 35252 30884 35308 30940
rect 48748 30884 48804 31052
rect 50372 30940 51212 30996
rect 51268 30940 51278 30996
rect 52210 30940 52220 30996
rect 52276 30940 53676 30996
rect 53732 30940 54348 30996
rect 54404 30940 54414 30996
rect 50372 30884 50428 30940
rect 0 30716 3612 30772
rect 3668 30716 7308 30772
rect 7364 30716 7374 30772
rect 8194 30716 8204 30772
rect 8260 30716 8876 30772
rect 8932 30716 8942 30772
rect 9650 30716 9660 30772
rect 9716 30716 9884 30772
rect 9940 30716 9950 30772
rect 11732 30716 14364 30772
rect 14420 30716 14430 30772
rect 15092 30716 27188 30772
rect 27468 30828 34412 30884
rect 34468 30828 35308 30884
rect 36194 30828 36204 30884
rect 36260 30828 36652 30884
rect 36708 30828 36718 30884
rect 36978 30828 36988 30884
rect 37044 30828 41580 30884
rect 41636 30828 41646 30884
rect 42578 30828 42588 30884
rect 42644 30828 44156 30884
rect 44212 30828 44222 30884
rect 44706 30828 44716 30884
rect 44772 30828 47516 30884
rect 47572 30828 47582 30884
rect 48748 30828 50428 30884
rect 51324 30828 51660 30884
rect 51716 30828 51726 30884
rect 52658 30828 52668 30884
rect 52724 30828 52780 30884
rect 52836 30828 53116 30884
rect 53172 30828 53182 30884
rect 0 30688 112 30716
rect 15092 30660 15148 30716
rect 27468 30660 27524 30828
rect 51324 30772 51380 30828
rect 57344 30772 57456 30800
rect 27794 30716 27804 30772
rect 27860 30716 28812 30772
rect 28868 30716 28878 30772
rect 29250 30716 29260 30772
rect 29316 30716 30044 30772
rect 30100 30716 30110 30772
rect 31490 30716 31500 30772
rect 31556 30716 32732 30772
rect 32788 30716 33404 30772
rect 33460 30716 34076 30772
rect 34132 30716 34142 30772
rect 34626 30716 34636 30772
rect 34692 30716 35084 30772
rect 35140 30716 35150 30772
rect 36194 30716 36204 30772
rect 36260 30716 36876 30772
rect 36932 30716 36988 30772
rect 37044 30716 37054 30772
rect 38098 30716 38108 30772
rect 38164 30716 38444 30772
rect 38500 30716 39228 30772
rect 39284 30716 39294 30772
rect 43586 30716 43596 30772
rect 43652 30716 51324 30772
rect 51380 30716 51390 30772
rect 51510 30716 51548 30772
rect 51604 30716 53676 30772
rect 53732 30716 53742 30772
rect 57250 30716 57260 30772
rect 57316 30716 57456 30772
rect 57344 30688 57456 30716
rect 3378 30604 3388 30660
rect 3444 30604 4060 30660
rect 4116 30604 4126 30660
rect 4946 30604 4956 30660
rect 5012 30604 5964 30660
rect 6020 30604 6030 30660
rect 6626 30604 6636 30660
rect 6692 30604 7980 30660
rect 8036 30604 8428 30660
rect 8484 30604 8494 30660
rect 8754 30604 8764 30660
rect 8820 30604 15148 30660
rect 15922 30604 15932 30660
rect 15988 30604 19852 30660
rect 19908 30604 19918 30660
rect 21634 30604 21644 30660
rect 21700 30604 23548 30660
rect 23604 30604 23614 30660
rect 25442 30604 25452 30660
rect 25508 30604 27524 30660
rect 27682 30604 27692 30660
rect 27748 30604 44156 30660
rect 44212 30604 44222 30660
rect 46162 30604 46172 30660
rect 46228 30604 46732 30660
rect 46788 30604 46798 30660
rect 48850 30604 48860 30660
rect 48916 30604 49644 30660
rect 49700 30604 49868 30660
rect 49924 30604 49934 30660
rect 50754 30604 50764 30660
rect 50820 30604 55580 30660
rect 55636 30604 55646 30660
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 44454 30548 44464 30604
rect 44520 30548 44568 30604
rect 44624 30548 44672 30604
rect 44728 30548 44738 30604
rect 2706 30492 2716 30548
rect 2772 30492 4172 30548
rect 4228 30492 4238 30548
rect 4834 30492 4844 30548
rect 4900 30492 8988 30548
rect 9044 30492 9054 30548
rect 9398 30492 9436 30548
rect 9492 30492 13076 30548
rect 14914 30492 14924 30548
rect 14980 30492 18844 30548
rect 18900 30492 18910 30548
rect 21298 30492 21308 30548
rect 21364 30492 22652 30548
rect 22708 30492 22718 30548
rect 29036 30492 34188 30548
rect 34244 30492 34254 30548
rect 34626 30492 34636 30548
rect 34692 30492 44212 30548
rect 45602 30492 45612 30548
rect 45668 30492 47404 30548
rect 47460 30492 47470 30548
rect 48290 30492 48300 30548
rect 48356 30492 54908 30548
rect 54964 30492 54974 30548
rect 578 30380 588 30436
rect 644 30380 6860 30436
rect 6916 30380 6926 30436
rect 7858 30380 7868 30436
rect 7924 30380 9324 30436
rect 9380 30380 9390 30436
rect 10322 30380 10332 30436
rect 10388 30380 10892 30436
rect 10948 30380 10958 30436
rect 0 30324 112 30352
rect 10332 30324 10388 30380
rect 13020 30324 13076 30492
rect 13794 30380 13804 30436
rect 13860 30380 14588 30436
rect 14644 30380 14654 30436
rect 16706 30380 16716 30436
rect 16772 30380 17276 30436
rect 17332 30380 17342 30436
rect 18498 30380 18508 30436
rect 18564 30380 19068 30436
rect 19124 30380 19964 30436
rect 20020 30380 20030 30436
rect 21522 30380 21532 30436
rect 21588 30380 21644 30436
rect 21700 30380 21710 30436
rect 22978 30380 22988 30436
rect 23044 30380 26684 30436
rect 26740 30380 26750 30436
rect 26852 30380 28364 30436
rect 28420 30380 28430 30436
rect 26852 30324 26908 30380
rect 29036 30324 29092 30492
rect 44156 30436 44212 30492
rect 29474 30380 29484 30436
rect 29540 30380 32844 30436
rect 32900 30380 32910 30436
rect 33058 30380 33068 30436
rect 33124 30380 36988 30436
rect 37044 30380 37548 30436
rect 37604 30380 37614 30436
rect 37874 30380 37884 30436
rect 37940 30380 42588 30436
rect 42644 30380 42654 30436
rect 44156 30380 46284 30436
rect 46340 30380 46956 30436
rect 47012 30380 47022 30436
rect 48514 30380 48524 30436
rect 48580 30380 50092 30436
rect 50148 30380 50158 30436
rect 50306 30380 50316 30436
rect 50372 30380 53844 30436
rect 56130 30380 56140 30436
rect 56196 30380 56476 30436
rect 56532 30380 56542 30436
rect 0 30268 2492 30324
rect 2548 30268 2558 30324
rect 2706 30268 2716 30324
rect 2772 30268 7084 30324
rect 7140 30268 7150 30324
rect 8754 30268 8764 30324
rect 8820 30268 10388 30324
rect 12226 30268 12236 30324
rect 12292 30268 12460 30324
rect 12516 30268 12526 30324
rect 12646 30268 12684 30324
rect 12740 30268 12750 30324
rect 13020 30268 18956 30324
rect 19012 30268 19022 30324
rect 19730 30268 19740 30324
rect 19796 30268 24892 30324
rect 24948 30268 24958 30324
rect 25116 30268 25676 30324
rect 25732 30268 25742 30324
rect 26114 30268 26124 30324
rect 26180 30268 26908 30324
rect 27010 30268 27020 30324
rect 27076 30268 29092 30324
rect 29250 30268 29260 30324
rect 29316 30268 31948 30324
rect 32004 30268 32014 30324
rect 32946 30268 32956 30324
rect 33012 30268 34580 30324
rect 34850 30268 34860 30324
rect 34916 30268 36428 30324
rect 36484 30268 39676 30324
rect 39732 30268 39742 30324
rect 40012 30268 40852 30324
rect 41122 30268 41132 30324
rect 41188 30268 44492 30324
rect 44548 30268 45164 30324
rect 45220 30268 45230 30324
rect 47030 30268 47068 30324
rect 47124 30268 47134 30324
rect 47282 30268 47292 30324
rect 47348 30268 48300 30324
rect 48356 30268 48366 30324
rect 48962 30268 48972 30324
rect 49028 30268 50204 30324
rect 50260 30268 50270 30324
rect 51202 30268 51212 30324
rect 51268 30268 52108 30324
rect 52164 30268 52174 30324
rect 0 30240 112 30268
rect 25116 30212 25172 30268
rect 34524 30212 34580 30268
rect 40012 30212 40068 30268
rect 2930 30156 2940 30212
rect 2996 30156 4060 30212
rect 4116 30156 4284 30212
rect 4340 30156 4350 30212
rect 4498 30156 4508 30212
rect 4564 30156 4844 30212
rect 4900 30156 4910 30212
rect 5590 30156 5628 30212
rect 5684 30156 6076 30212
rect 6132 30156 6142 30212
rect 6626 30156 6636 30212
rect 6692 30156 7084 30212
rect 7140 30156 7420 30212
rect 7476 30156 7486 30212
rect 7746 30156 7756 30212
rect 7812 30156 9268 30212
rect 9762 30156 9772 30212
rect 9828 30156 10220 30212
rect 10276 30156 10286 30212
rect 10434 30156 10444 30212
rect 10500 30156 12796 30212
rect 12852 30156 12862 30212
rect 13234 30156 13244 30212
rect 13300 30156 13804 30212
rect 13860 30156 13870 30212
rect 14242 30156 14252 30212
rect 14308 30156 14476 30212
rect 14532 30156 14542 30212
rect 15250 30156 15260 30212
rect 15316 30156 15596 30212
rect 15652 30156 15662 30212
rect 16034 30156 16044 30212
rect 16100 30156 17164 30212
rect 17220 30156 19628 30212
rect 19684 30156 20972 30212
rect 21028 30156 21038 30212
rect 21186 30156 21196 30212
rect 21252 30156 21644 30212
rect 21700 30156 21812 30212
rect 23314 30156 23324 30212
rect 23380 30156 24332 30212
rect 24388 30156 25172 30212
rect 25442 30156 25452 30212
rect 25508 30156 27468 30212
rect 27524 30156 27534 30212
rect 27794 30156 27804 30212
rect 27860 30156 27916 30212
rect 27972 30156 27982 30212
rect 29026 30156 29036 30212
rect 29092 30156 29484 30212
rect 29540 30156 30380 30212
rect 30436 30156 30446 30212
rect 31490 30156 31500 30212
rect 31556 30156 33404 30212
rect 33460 30156 33470 30212
rect 33618 30156 33628 30212
rect 33684 30156 33964 30212
rect 34020 30156 34030 30212
rect 34524 30156 35644 30212
rect 35700 30156 35710 30212
rect 36054 30156 36092 30212
rect 36148 30156 36158 30212
rect 36306 30156 36316 30212
rect 36372 30156 37660 30212
rect 37716 30156 37726 30212
rect 39554 30156 39564 30212
rect 39620 30156 40068 30212
rect 40198 30156 40236 30212
rect 40292 30156 40302 30212
rect 9212 30100 9268 30156
rect 3490 30044 3500 30100
rect 3556 30044 4396 30100
rect 4452 30044 4462 30100
rect 5282 30044 5292 30100
rect 5348 30044 6300 30100
rect 6356 30044 6366 30100
rect 8194 30044 8204 30100
rect 8260 30044 8988 30100
rect 9044 30044 9054 30100
rect 9212 30044 10332 30100
rect 10388 30044 10398 30100
rect 10658 30044 10668 30100
rect 10724 30044 10892 30100
rect 10948 30044 14588 30100
rect 14644 30044 14654 30100
rect 18050 30044 18060 30100
rect 18116 30044 19852 30100
rect 19908 30044 19918 30100
rect 20178 30044 20188 30100
rect 20244 30044 21700 30100
rect 3052 29932 6972 29988
rect 7028 29932 7038 29988
rect 8306 29932 8316 29988
rect 8372 29932 10556 29988
rect 10612 29932 10622 29988
rect 13570 29932 13580 29988
rect 13636 29932 14364 29988
rect 14420 29932 14430 29988
rect 15810 29932 15820 29988
rect 15876 29932 19180 29988
rect 19236 29932 19246 29988
rect 19506 29932 19516 29988
rect 19572 29932 20076 29988
rect 20132 29932 20142 29988
rect 20402 29932 20412 29988
rect 20468 29932 21196 29988
rect 21252 29932 21262 29988
rect 0 29876 112 29904
rect 3052 29876 3108 29932
rect 0 29820 3052 29876
rect 3108 29820 3118 29876
rect 4386 29820 4396 29876
rect 4452 29820 5292 29876
rect 5348 29820 5358 29876
rect 6066 29820 6076 29876
rect 6132 29820 6412 29876
rect 6468 29820 7420 29876
rect 7476 29820 7486 29876
rect 7858 29820 7868 29876
rect 7924 29820 8092 29876
rect 8148 29820 9660 29876
rect 9716 29820 9726 29876
rect 10882 29820 10892 29876
rect 10948 29820 13692 29876
rect 13748 29820 13758 29876
rect 14466 29820 14476 29876
rect 14532 29820 16940 29876
rect 16996 29820 17388 29876
rect 17444 29820 17454 29876
rect 19292 29820 21420 29876
rect 21476 29820 21486 29876
rect 0 29792 112 29820
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 19292 29764 19348 29820
rect 690 29708 700 29764
rect 756 29708 2604 29764
rect 2660 29708 2670 29764
rect 4274 29708 4284 29764
rect 4340 29708 5068 29764
rect 5124 29708 5134 29764
rect 5506 29708 5516 29764
rect 5572 29708 8204 29764
rect 8260 29708 8270 29764
rect 8754 29708 8764 29764
rect 8820 29708 19348 29764
rect 20066 29708 20076 29764
rect 20132 29708 21140 29764
rect 4050 29596 4060 29652
rect 4116 29596 5180 29652
rect 5236 29596 5246 29652
rect 9314 29596 9324 29652
rect 9380 29596 11788 29652
rect 11844 29596 11854 29652
rect 12226 29596 12236 29652
rect 12292 29596 12460 29652
rect 12516 29596 12526 29652
rect 12898 29596 12908 29652
rect 12964 29596 13468 29652
rect 13524 29596 13534 29652
rect 13682 29596 13692 29652
rect 13748 29596 21028 29652
rect 1922 29484 1932 29540
rect 1988 29484 2492 29540
rect 2548 29484 2558 29540
rect 3266 29484 3276 29540
rect 3332 29484 5404 29540
rect 5460 29484 5470 29540
rect 5954 29484 5964 29540
rect 6020 29484 15820 29540
rect 15876 29484 15886 29540
rect 16044 29484 19068 29540
rect 19124 29484 19134 29540
rect 0 29428 112 29456
rect 0 29372 140 29428
rect 196 29372 206 29428
rect 2818 29372 2828 29428
rect 2884 29372 3836 29428
rect 3892 29372 5964 29428
rect 6020 29372 6030 29428
rect 8978 29372 8988 29428
rect 9044 29372 9884 29428
rect 9940 29372 9950 29428
rect 11218 29372 11228 29428
rect 11284 29372 11676 29428
rect 11732 29372 11742 29428
rect 12012 29372 15148 29428
rect 0 29344 112 29372
rect 12012 29316 12068 29372
rect 1362 29260 1372 29316
rect 1428 29260 1596 29316
rect 1652 29260 1662 29316
rect 2566 29260 2604 29316
rect 2660 29260 2670 29316
rect 3154 29260 3164 29316
rect 3220 29260 4956 29316
rect 5012 29260 5022 29316
rect 5170 29260 5180 29316
rect 5236 29260 6524 29316
rect 6580 29260 12068 29316
rect 12226 29260 12236 29316
rect 12292 29260 14700 29316
rect 14756 29260 14766 29316
rect 15092 29204 15148 29372
rect 16044 29204 16100 29484
rect 17798 29372 17836 29428
rect 17892 29372 17902 29428
rect 18498 29372 18508 29428
rect 18564 29372 18844 29428
rect 18900 29372 19180 29428
rect 19236 29372 19246 29428
rect 19058 29260 19068 29316
rect 19124 29260 20636 29316
rect 20692 29260 20702 29316
rect 20972 29204 21028 29596
rect 21084 29428 21140 29708
rect 21644 29652 21700 30044
rect 21756 29988 21812 30156
rect 40236 30100 40292 30156
rect 22306 30044 22316 30100
rect 22372 30044 22876 30100
rect 22932 30044 25676 30100
rect 25732 30044 26124 30100
rect 26180 30044 26190 30100
rect 27234 30044 27244 30100
rect 27300 30044 27356 30100
rect 27412 30044 27422 30100
rect 27906 30044 27916 30100
rect 27972 30044 29820 30100
rect 29876 30044 29886 30100
rect 30034 30044 30044 30100
rect 30100 30044 32396 30100
rect 32452 30044 40292 30100
rect 40796 30100 40852 30268
rect 53788 30212 53844 30380
rect 57344 30324 57456 30352
rect 56802 30268 56812 30324
rect 56868 30268 57456 30324
rect 57344 30240 57456 30268
rect 40982 30156 41020 30212
rect 41076 30156 41086 30212
rect 41234 30156 41244 30212
rect 41300 30156 44268 30212
rect 44324 30156 44334 30212
rect 44940 30156 45612 30212
rect 45668 30156 45678 30212
rect 46162 30156 46172 30212
rect 46228 30156 46620 30212
rect 46676 30156 47180 30212
rect 47236 30156 47246 30212
rect 47394 30156 47404 30212
rect 47460 30156 48076 30212
rect 48132 30156 48142 30212
rect 48402 30156 48412 30212
rect 48468 30156 49532 30212
rect 49588 30156 49598 30212
rect 50754 30156 50764 30212
rect 50820 30156 51660 30212
rect 51716 30156 51726 30212
rect 53788 30156 55804 30212
rect 55860 30156 55870 30212
rect 44940 30100 44996 30156
rect 40796 30044 44996 30100
rect 45154 30044 45164 30100
rect 45220 30044 46172 30100
rect 46228 30044 46238 30100
rect 47404 29988 47460 30156
rect 47954 30044 47964 30100
rect 48020 30044 52668 30100
rect 52724 30044 52734 30100
rect 53218 30044 53228 30100
rect 53284 30044 53900 30100
rect 53956 30044 53966 30100
rect 21756 29932 27748 29988
rect 27906 29932 27916 29988
rect 27972 29932 28364 29988
rect 28420 29932 28430 29988
rect 30828 29932 33180 29988
rect 33236 29932 33628 29988
rect 33684 29932 33694 29988
rect 34290 29932 34300 29988
rect 34356 29932 34972 29988
rect 35028 29932 35532 29988
rect 35588 29932 35598 29988
rect 37202 29932 37212 29988
rect 37268 29932 37772 29988
rect 37828 29932 37838 29988
rect 38322 29932 38332 29988
rect 38388 29932 44212 29988
rect 44902 29932 44940 29988
rect 44996 29932 45006 29988
rect 45266 29932 45276 29988
rect 45332 29932 47460 29988
rect 48626 29932 48636 29988
rect 48692 29932 49532 29988
rect 49588 29932 49598 29988
rect 49746 29932 49756 29988
rect 49812 29932 50764 29988
rect 50820 29932 54236 29988
rect 54292 29932 54302 29988
rect 27692 29876 27748 29932
rect 30828 29876 30884 29932
rect 44156 29876 44212 29932
rect 57344 29876 57456 29904
rect 27692 29820 30884 29876
rect 31042 29820 31052 29876
rect 31108 29820 33964 29876
rect 34020 29820 34030 29876
rect 34178 29820 34188 29876
rect 34244 29820 34692 29876
rect 34850 29820 34860 29876
rect 34916 29820 35420 29876
rect 35476 29820 35486 29876
rect 38612 29820 42476 29876
rect 42532 29820 42542 29876
rect 44156 29820 52948 29876
rect 53330 29820 53340 29876
rect 53396 29820 53900 29876
rect 53956 29820 53966 29876
rect 56578 29820 56588 29876
rect 56644 29820 57456 29876
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 34636 29764 34692 29820
rect 38612 29764 38668 29820
rect 43794 29764 43804 29820
rect 43860 29764 43908 29820
rect 43964 29764 44012 29820
rect 44068 29764 44078 29820
rect 52892 29764 52948 29820
rect 57344 29792 57456 29820
rect 31042 29708 31052 29764
rect 31108 29708 32956 29764
rect 33012 29708 33022 29764
rect 33730 29708 33740 29764
rect 33796 29708 34412 29764
rect 34468 29708 34478 29764
rect 34626 29708 34636 29764
rect 34692 29708 38668 29764
rect 38770 29708 38780 29764
rect 38836 29708 40460 29764
rect 40516 29708 40526 29764
rect 44146 29708 44156 29764
rect 44212 29708 48524 29764
rect 48580 29708 48860 29764
rect 48916 29708 48926 29764
rect 49074 29708 49084 29764
rect 49140 29708 52332 29764
rect 52388 29708 52398 29764
rect 52892 29708 55020 29764
rect 55076 29708 55086 29764
rect 21644 29596 29260 29652
rect 29316 29596 29326 29652
rect 31826 29596 31836 29652
rect 31892 29596 34748 29652
rect 34804 29596 34814 29652
rect 36530 29596 36540 29652
rect 36596 29596 37324 29652
rect 37380 29596 37390 29652
rect 38882 29596 38892 29652
rect 38948 29596 48748 29652
rect 48804 29596 48814 29652
rect 50082 29596 50092 29652
rect 50148 29596 54908 29652
rect 54964 29596 54974 29652
rect 21858 29484 21868 29540
rect 21924 29484 23436 29540
rect 23492 29484 23996 29540
rect 24052 29484 26236 29540
rect 26292 29484 27916 29540
rect 27972 29484 27982 29540
rect 28578 29484 28588 29540
rect 28644 29484 31108 29540
rect 31266 29484 31276 29540
rect 31332 29484 32620 29540
rect 32676 29484 35532 29540
rect 35588 29484 35598 29540
rect 36166 29484 36204 29540
rect 36260 29484 36270 29540
rect 36978 29484 36988 29540
rect 37044 29484 45948 29540
rect 46004 29484 46014 29540
rect 46834 29484 46844 29540
rect 46900 29484 48188 29540
rect 48244 29484 48254 29540
rect 50194 29484 50204 29540
rect 50260 29484 51660 29540
rect 51716 29484 51726 29540
rect 53330 29484 53340 29540
rect 53396 29484 53452 29540
rect 53508 29484 53518 29540
rect 31052 29428 31108 29484
rect 57344 29428 57456 29456
rect 21084 29372 26908 29428
rect 28242 29372 28252 29428
rect 28308 29372 30828 29428
rect 30884 29372 30894 29428
rect 31052 29372 38780 29428
rect 38836 29372 40236 29428
rect 40292 29372 40302 29428
rect 44258 29372 44268 29428
rect 44324 29372 44334 29428
rect 47506 29372 47516 29428
rect 47572 29372 48412 29428
rect 48468 29372 48478 29428
rect 49522 29372 49532 29428
rect 49588 29372 50316 29428
rect 50372 29372 50382 29428
rect 52770 29372 52780 29428
rect 52836 29372 56028 29428
rect 56084 29372 56094 29428
rect 56354 29372 56364 29428
rect 56420 29372 57456 29428
rect 26852 29316 26908 29372
rect 44268 29316 44324 29372
rect 57344 29344 57456 29372
rect 22054 29260 22092 29316
rect 22148 29260 23100 29316
rect 23156 29260 23166 29316
rect 24434 29260 24444 29316
rect 24500 29260 25228 29316
rect 25284 29260 26684 29316
rect 26740 29260 26750 29316
rect 26852 29260 31892 29316
rect 32162 29260 32172 29316
rect 32228 29260 32396 29316
rect 32452 29260 32462 29316
rect 32946 29260 32956 29316
rect 33012 29260 34300 29316
rect 34356 29260 34366 29316
rect 35186 29260 35196 29316
rect 35252 29260 36820 29316
rect 40338 29260 40348 29316
rect 40404 29260 40908 29316
rect 40964 29260 40974 29316
rect 44268 29260 46956 29316
rect 47012 29260 47022 29316
rect 49858 29260 49868 29316
rect 49924 29260 50764 29316
rect 50820 29260 50830 29316
rect 53890 29260 53900 29316
rect 53956 29260 54348 29316
rect 54404 29260 54414 29316
rect 31836 29204 31892 29260
rect 36764 29204 36820 29260
rect 2146 29148 2156 29204
rect 2212 29148 5964 29204
rect 6020 29148 6030 29204
rect 8978 29148 8988 29204
rect 9044 29148 12348 29204
rect 12404 29148 12414 29204
rect 12562 29148 12572 29204
rect 12628 29148 14476 29204
rect 14532 29148 14542 29204
rect 15092 29148 16100 29204
rect 16818 29148 16828 29204
rect 16884 29148 19180 29204
rect 19236 29148 19246 29204
rect 19842 29148 19852 29204
rect 19908 29148 20916 29204
rect 20972 29148 31052 29204
rect 31108 29148 31118 29204
rect 31836 29148 34972 29204
rect 35028 29148 35420 29204
rect 35476 29148 35486 29204
rect 36754 29148 36764 29204
rect 36820 29148 42700 29204
rect 42756 29148 42766 29204
rect 44930 29148 44940 29204
rect 44996 29148 46060 29204
rect 46116 29148 46126 29204
rect 48514 29148 48524 29204
rect 48580 29148 49084 29204
rect 49140 29148 49150 29204
rect 49746 29148 49756 29204
rect 49812 29148 52556 29204
rect 52612 29148 52622 29204
rect 53666 29148 53676 29204
rect 53732 29148 55916 29204
rect 55972 29148 55982 29204
rect 20860 29092 20916 29148
rect 2706 29036 2716 29092
rect 2772 29036 4172 29092
rect 4228 29036 4238 29092
rect 4946 29036 4956 29092
rect 5012 29036 12908 29092
rect 12964 29036 12974 29092
rect 13682 29036 13692 29092
rect 13748 29036 13916 29092
rect 13972 29036 13982 29092
rect 16482 29036 16492 29092
rect 16548 29036 16716 29092
rect 16772 29036 20076 29092
rect 20132 29036 20142 29092
rect 20860 29036 23660 29092
rect 23716 29036 23726 29092
rect 25106 29036 25116 29092
rect 25172 29036 28252 29092
rect 28308 29036 28318 29092
rect 28476 29036 29204 29092
rect 32722 29036 32732 29092
rect 32788 29036 33516 29092
rect 33572 29036 33582 29092
rect 33954 29036 33964 29092
rect 34020 29036 35196 29092
rect 35252 29036 35262 29092
rect 37650 29036 37660 29092
rect 37716 29036 39340 29092
rect 39396 29036 43484 29092
rect 43540 29036 43550 29092
rect 48402 29036 48412 29092
rect 48468 29036 49700 29092
rect 49970 29036 49980 29092
rect 50036 29036 50316 29092
rect 50372 29036 50382 29092
rect 52322 29036 52332 29092
rect 52388 29036 53340 29092
rect 53396 29036 55132 29092
rect 55188 29036 55198 29092
rect 0 28980 112 29008
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 28476 28980 28532 29036
rect 29148 28980 29204 29036
rect 44454 28980 44464 29036
rect 44520 28980 44568 29036
rect 44624 28980 44672 29036
rect 44728 28980 44738 29036
rect 49644 28980 49700 29036
rect 57344 28980 57456 29008
rect 0 28924 2604 28980
rect 2660 28924 2670 28980
rect 3378 28924 3388 28980
rect 3444 28924 3500 28980
rect 3556 28924 3566 28980
rect 5842 28924 5852 28980
rect 5908 28924 7196 28980
rect 7252 28924 7262 28980
rect 7410 28924 7420 28980
rect 7476 28924 10780 28980
rect 10836 28924 10846 28980
rect 11442 28924 11452 28980
rect 11508 28924 15932 28980
rect 15988 28924 15998 28980
rect 16156 28924 18172 28980
rect 18228 28924 18238 28980
rect 18610 28924 18620 28980
rect 18676 28924 23660 28980
rect 23716 28924 23726 28980
rect 26450 28924 26460 28980
rect 26516 28924 28532 28980
rect 29138 28924 29148 28980
rect 29204 28924 32284 28980
rect 32340 28924 32350 28980
rect 34738 28924 34748 28980
rect 34804 28924 36204 28980
rect 36260 28924 36652 28980
rect 36708 28924 36718 28980
rect 36866 28924 36876 28980
rect 36932 28924 40236 28980
rect 40292 28924 40302 28980
rect 41010 28924 41020 28980
rect 41076 28924 42140 28980
rect 42196 28924 43148 28980
rect 43204 28924 43214 28980
rect 43362 28924 43372 28980
rect 43428 28924 44156 28980
rect 44212 28924 44222 28980
rect 45490 28924 45500 28980
rect 45556 28924 49308 28980
rect 49364 28924 49420 28980
rect 49476 28924 49486 28980
rect 49634 28924 49644 28980
rect 49700 28924 49710 28980
rect 51090 28924 51100 28980
rect 51156 28924 53788 28980
rect 53844 28924 53854 28980
rect 56354 28924 56364 28980
rect 56420 28924 57456 28980
rect 0 28896 112 28924
rect 16156 28868 16212 28924
rect 57344 28896 57456 28924
rect 2818 28812 2828 28868
rect 2884 28812 3276 28868
rect 3332 28812 3342 28868
rect 3602 28812 3612 28868
rect 3668 28812 4956 28868
rect 5012 28812 5022 28868
rect 6626 28812 6636 28868
rect 6692 28812 9044 28868
rect 10882 28812 10892 28868
rect 10948 28812 16212 28868
rect 16370 28812 16380 28868
rect 16436 28812 18508 28868
rect 18564 28812 18574 28868
rect 19058 28812 19068 28868
rect 19124 28812 20748 28868
rect 20804 28812 20814 28868
rect 23538 28812 23548 28868
rect 23604 28812 25508 28868
rect 25666 28812 25676 28868
rect 25732 28812 26012 28868
rect 26068 28812 26460 28868
rect 26516 28812 26526 28868
rect 27356 28812 27916 28868
rect 27972 28812 27982 28868
rect 28998 28812 29036 28868
rect 29092 28812 29820 28868
rect 29876 28812 29886 28868
rect 31714 28812 31724 28868
rect 31780 28812 33068 28868
rect 33124 28812 34860 28868
rect 34916 28812 34926 28868
rect 35830 28812 35868 28868
rect 35924 28812 40908 28868
rect 40964 28812 42252 28868
rect 42308 28812 44268 28868
rect 44324 28812 44334 28868
rect 45714 28812 45724 28868
rect 45780 28812 46172 28868
rect 46228 28812 46238 28868
rect 47068 28812 52108 28868
rect 52164 28812 52174 28868
rect 52546 28812 52556 28868
rect 52612 28812 53004 28868
rect 53060 28812 55020 28868
rect 55076 28812 55086 28868
rect 55878 28812 55916 28868
rect 55972 28812 55982 28868
rect 8988 28756 9044 28812
rect 25452 28756 25508 28812
rect 27356 28756 27412 28812
rect 45948 28756 46004 28812
rect 3612 28700 4956 28756
rect 5012 28700 5022 28756
rect 5954 28700 5964 28756
rect 6020 28700 6076 28756
rect 6132 28700 6142 28756
rect 7196 28700 8764 28756
rect 8820 28700 8830 28756
rect 8988 28700 12460 28756
rect 12516 28700 12526 28756
rect 13468 28700 20636 28756
rect 20692 28700 20702 28756
rect 20962 28700 20972 28756
rect 21028 28700 22204 28756
rect 22260 28700 22270 28756
rect 23650 28700 23660 28756
rect 23716 28700 25116 28756
rect 25172 28700 25182 28756
rect 25452 28700 27412 28756
rect 27570 28700 27580 28756
rect 27636 28700 28364 28756
rect 28420 28700 28430 28756
rect 28914 28700 28924 28756
rect 28980 28700 29708 28756
rect 29764 28700 29774 28756
rect 31602 28700 31612 28756
rect 31668 28700 35308 28756
rect 35364 28700 35374 28756
rect 37174 28700 37212 28756
rect 37268 28700 37278 28756
rect 37874 28700 37884 28756
rect 37940 28700 38668 28756
rect 38724 28700 38734 28756
rect 38994 28700 39004 28756
rect 39060 28700 39844 28756
rect 41906 28700 41916 28756
rect 41972 28700 43708 28756
rect 43764 28700 45276 28756
rect 45332 28700 45342 28756
rect 45938 28700 45948 28756
rect 46004 28700 46014 28756
rect 3612 28644 3668 28700
rect 3602 28588 3612 28644
rect 3668 28588 3678 28644
rect 3938 28588 3948 28644
rect 4004 28588 6748 28644
rect 6804 28588 6814 28644
rect 0 28532 112 28560
rect 7196 28532 7252 28700
rect 7970 28588 7980 28644
rect 8036 28588 8204 28644
rect 8260 28588 8270 28644
rect 9660 28588 12348 28644
rect 12404 28588 12414 28644
rect 12534 28588 12572 28644
rect 12628 28588 12638 28644
rect 9660 28532 9716 28588
rect 13468 28532 13524 28700
rect 39788 28644 39844 28700
rect 13692 28588 15260 28644
rect 15316 28588 15326 28644
rect 15586 28588 15596 28644
rect 15652 28588 15932 28644
rect 15988 28588 15998 28644
rect 18498 28588 18508 28644
rect 18564 28588 19516 28644
rect 19572 28588 20860 28644
rect 20916 28588 20926 28644
rect 21186 28588 21196 28644
rect 21252 28588 22092 28644
rect 22148 28588 22158 28644
rect 22306 28588 22316 28644
rect 22372 28588 22540 28644
rect 22596 28588 28980 28644
rect 29698 28588 29708 28644
rect 29764 28588 30268 28644
rect 30324 28588 30334 28644
rect 31938 28588 31948 28644
rect 32004 28588 33180 28644
rect 33236 28588 33246 28644
rect 33394 28588 33404 28644
rect 33460 28588 35252 28644
rect 35522 28588 35532 28644
rect 35588 28588 35644 28644
rect 35700 28588 35710 28644
rect 36754 28588 36764 28644
rect 36820 28588 39564 28644
rect 39620 28588 39630 28644
rect 39778 28588 39788 28644
rect 39844 28588 45724 28644
rect 45780 28588 45790 28644
rect 13692 28532 13748 28588
rect 28924 28532 28980 28588
rect 35196 28532 35252 28588
rect 47068 28532 47124 28812
rect 47618 28700 47628 28756
rect 47684 28700 51996 28756
rect 52052 28700 52062 28756
rect 52854 28700 52892 28756
rect 52948 28700 54348 28756
rect 54404 28700 54414 28756
rect 47506 28588 47516 28644
rect 47572 28588 48188 28644
rect 48244 28588 48254 28644
rect 49718 28588 49756 28644
rect 49812 28588 49822 28644
rect 50978 28588 50988 28644
rect 51044 28588 54796 28644
rect 54852 28588 54862 28644
rect 55570 28588 55580 28644
rect 55636 28588 55916 28644
rect 55972 28588 55982 28644
rect 57344 28532 57456 28560
rect 0 28476 7252 28532
rect 7522 28476 7532 28532
rect 7588 28476 8092 28532
rect 8148 28476 8158 28532
rect 8876 28476 9716 28532
rect 9874 28476 9884 28532
rect 9940 28476 10332 28532
rect 10388 28476 10556 28532
rect 10612 28476 10622 28532
rect 10770 28476 10780 28532
rect 10836 28476 13244 28532
rect 13300 28476 13524 28532
rect 13682 28476 13692 28532
rect 13748 28476 13758 28532
rect 15362 28476 15372 28532
rect 15428 28476 17164 28532
rect 17220 28476 17230 28532
rect 18946 28476 18956 28532
rect 19012 28476 19292 28532
rect 19348 28476 19358 28532
rect 20066 28476 20076 28532
rect 20132 28476 20524 28532
rect 20580 28476 20590 28532
rect 21186 28476 21196 28532
rect 21252 28476 21308 28532
rect 21364 28476 21374 28532
rect 21522 28476 21532 28532
rect 21588 28476 24332 28532
rect 24388 28476 24398 28532
rect 24882 28476 24892 28532
rect 24948 28476 26012 28532
rect 26068 28476 26236 28532
rect 26292 28476 26302 28532
rect 26908 28476 28476 28532
rect 28532 28476 28542 28532
rect 28924 28476 30604 28532
rect 30660 28476 33516 28532
rect 33572 28476 33582 28532
rect 33964 28476 34412 28532
rect 34468 28476 34478 28532
rect 35196 28476 35756 28532
rect 35812 28476 35822 28532
rect 38770 28476 38780 28532
rect 38836 28476 39676 28532
rect 39732 28476 39742 28532
rect 43362 28476 43372 28532
rect 43428 28476 44268 28532
rect 44324 28476 44334 28532
rect 44594 28476 44604 28532
rect 44660 28476 47124 28532
rect 47954 28476 47964 28532
rect 48020 28476 48636 28532
rect 48692 28476 51996 28532
rect 52052 28476 52062 28532
rect 54002 28476 54012 28532
rect 54068 28476 56140 28532
rect 56196 28476 56206 28532
rect 56466 28476 56476 28532
rect 56532 28476 57456 28532
rect 0 28448 112 28476
rect 466 28364 476 28420
rect 532 28364 1036 28420
rect 1092 28364 1102 28420
rect 3266 28364 3276 28420
rect 3332 28364 4228 28420
rect 4386 28364 4396 28420
rect 4452 28364 4844 28420
rect 4900 28364 4910 28420
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 4172 28196 4228 28364
rect 8876 28308 8932 28476
rect 26908 28420 26964 28476
rect 33964 28420 34020 28476
rect 57344 28448 57456 28476
rect 10098 28364 10108 28420
rect 10164 28364 14364 28420
rect 14420 28364 14430 28420
rect 16482 28364 16492 28420
rect 16548 28364 26964 28420
rect 27122 28364 27132 28420
rect 27188 28364 28364 28420
rect 28420 28364 28430 28420
rect 31602 28364 31612 28420
rect 31668 28378 33684 28420
rect 31668 28364 33796 28378
rect 33954 28364 33964 28420
rect 34020 28364 34030 28420
rect 34402 28364 34412 28420
rect 34468 28364 35308 28420
rect 35410 28364 35420 28420
rect 35476 28364 38444 28420
rect 38500 28364 38510 28420
rect 38854 28364 38892 28420
rect 38948 28364 38958 28420
rect 39778 28364 39788 28420
rect 39844 28364 43596 28420
rect 43652 28364 43662 28420
rect 44258 28364 44268 28420
rect 44324 28364 45052 28420
rect 45108 28364 45118 28420
rect 47394 28364 47404 28420
rect 47460 28364 48524 28420
rect 48580 28364 48590 28420
rect 52210 28364 52220 28420
rect 52276 28364 52556 28420
rect 52612 28364 52622 28420
rect 33628 28322 33796 28364
rect 33740 28308 33796 28322
rect 5842 28252 5852 28308
rect 5908 28252 8932 28308
rect 9090 28252 9100 28308
rect 9156 28252 9996 28308
rect 10052 28252 10062 28308
rect 10658 28252 10668 28308
rect 10724 28252 10892 28308
rect 10948 28252 10958 28308
rect 11330 28252 11340 28308
rect 11396 28252 12796 28308
rect 12852 28252 12862 28308
rect 13010 28252 13020 28308
rect 13076 28252 15036 28308
rect 15092 28252 16268 28308
rect 16324 28252 23548 28308
rect 24210 28252 24220 28308
rect 24276 28252 31276 28308
rect 31332 28252 31342 28308
rect 33740 28252 34076 28308
rect 34132 28252 34188 28308
rect 34244 28252 34254 28308
rect 35252 28252 35308 28364
rect 35364 28252 35374 28308
rect 36306 28252 36316 28308
rect 36372 28252 36764 28308
rect 36820 28252 36830 28308
rect 36978 28252 36988 28308
rect 37044 28252 38108 28308
rect 38164 28252 38174 28308
rect 42354 28252 42364 28308
rect 42420 28252 42476 28308
rect 42532 28252 42542 28308
rect 45154 28252 45164 28308
rect 45220 28252 47852 28308
rect 47908 28252 53340 28308
rect 53396 28252 53406 28308
rect 53554 28252 53564 28308
rect 53620 28252 54908 28308
rect 54964 28252 54974 28308
rect 4162 28140 4172 28196
rect 4228 28140 4238 28196
rect 4722 28140 4732 28196
rect 4788 28140 4956 28196
rect 5012 28140 5022 28196
rect 6066 28140 6076 28196
rect 6132 28140 6300 28196
rect 6356 28140 6366 28196
rect 7522 28140 7532 28196
rect 7588 28140 7980 28196
rect 8036 28140 8046 28196
rect 8530 28140 8540 28196
rect 8596 28140 11340 28196
rect 11396 28140 11406 28196
rect 12338 28140 12348 28196
rect 12404 28140 17052 28196
rect 17108 28140 17118 28196
rect 17378 28140 17388 28196
rect 17444 28140 22316 28196
rect 22372 28140 22382 28196
rect 0 28084 112 28112
rect 0 28028 1204 28084
rect 2370 28028 2380 28084
rect 2436 28028 3388 28084
rect 4386 28028 4396 28084
rect 4452 28028 5068 28084
rect 5124 28028 5134 28084
rect 6300 28028 13020 28084
rect 13076 28028 13086 28084
rect 13318 28028 13356 28084
rect 13412 28028 13422 28084
rect 20514 28028 20524 28084
rect 20580 28028 21756 28084
rect 21812 28028 21822 28084
rect 0 28000 112 28028
rect 1148 27972 1204 28028
rect 3332 27972 3388 28028
rect 6300 27972 6356 28028
rect 23492 27972 23548 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 43794 28196 43804 28252
rect 43860 28196 43908 28252
rect 43964 28196 44012 28252
rect 44068 28196 44078 28252
rect 26226 28140 26236 28196
rect 26292 28140 28700 28196
rect 28756 28140 32956 28196
rect 33012 28140 33022 28196
rect 33618 28140 33628 28196
rect 33684 28140 34300 28196
rect 34356 28140 34366 28196
rect 34524 28140 38668 28196
rect 39554 28140 39564 28196
rect 39620 28140 40796 28196
rect 40852 28140 40862 28196
rect 44706 28140 44716 28196
rect 44772 28140 45388 28196
rect 45444 28140 45454 28196
rect 47282 28140 47292 28196
rect 47348 28140 52108 28196
rect 52164 28140 52174 28196
rect 53900 28140 54124 28196
rect 54180 28140 54190 28196
rect 34524 28084 34580 28140
rect 38612 28084 38668 28140
rect 53900 28084 53956 28140
rect 57344 28084 57456 28112
rect 24770 28028 24780 28084
rect 24836 28028 26852 28084
rect 27010 28028 27020 28084
rect 27076 28028 27580 28084
rect 27636 28028 27646 28084
rect 28130 28028 28140 28084
rect 28196 28028 31052 28084
rect 31108 28028 31118 28084
rect 31714 28028 31724 28084
rect 31780 28028 34580 28084
rect 35186 28028 35196 28084
rect 35252 28028 36876 28084
rect 36932 28028 36942 28084
rect 38612 28028 39228 28084
rect 39284 28028 39294 28084
rect 39442 28028 39452 28084
rect 39508 28028 39788 28084
rect 39844 28028 39854 28084
rect 40002 28028 40012 28084
rect 40068 28028 40124 28084
rect 40180 28028 40190 28084
rect 40674 28028 40684 28084
rect 40740 28028 42140 28084
rect 42196 28028 42206 28084
rect 42578 28028 42588 28084
rect 42644 28028 44492 28084
rect 44548 28028 50204 28084
rect 50260 28028 50270 28084
rect 51314 28028 51324 28084
rect 51380 28028 53340 28084
rect 53396 28028 53406 28084
rect 53890 28028 53900 28084
rect 53956 28028 53966 28084
rect 55458 28028 55468 28084
rect 55524 28028 57456 28084
rect 26796 27972 26852 28028
rect 57344 28000 57456 28028
rect 1148 27916 2492 27972
rect 2548 27916 2558 27972
rect 3332 27916 6300 27972
rect 6356 27916 6366 27972
rect 7858 27916 7868 27972
rect 7924 27916 8876 27972
rect 8932 27916 8942 27972
rect 16930 27916 16940 27972
rect 16996 27916 17500 27972
rect 17556 27916 17566 27972
rect 17938 27916 17948 27972
rect 18004 27916 19180 27972
rect 19236 27916 19246 27972
rect 19394 27916 19404 27972
rect 19460 27916 20412 27972
rect 20468 27916 21532 27972
rect 21588 27916 21598 27972
rect 21858 27916 21868 27972
rect 21924 27916 22092 27972
rect 22148 27916 22158 27972
rect 23492 27916 26460 27972
rect 26516 27916 26526 27972
rect 26796 27916 42476 27972
rect 42532 27916 42542 27972
rect 43138 27916 43148 27972
rect 43204 27916 45164 27972
rect 45220 27916 45230 27972
rect 1250 27804 1260 27860
rect 1316 27804 1372 27860
rect 1428 27804 1438 27860
rect 2146 27804 2156 27860
rect 2212 27804 2716 27860
rect 2772 27804 2782 27860
rect 3490 27804 3500 27860
rect 3556 27804 3724 27860
rect 3780 27804 3790 27860
rect 3938 27804 3948 27860
rect 4004 27804 5292 27860
rect 5348 27804 5358 27860
rect 6850 27804 6860 27860
rect 6916 27804 7756 27860
rect 7812 27804 7822 27860
rect 9986 27804 9996 27860
rect 10052 27804 12796 27860
rect 12852 27804 12862 27860
rect 13122 27804 13132 27860
rect 13188 27804 14028 27860
rect 14084 27804 14094 27860
rect 14550 27804 14588 27860
rect 14644 27804 18508 27860
rect 18564 27804 18574 27860
rect 19058 27804 19068 27860
rect 19124 27804 19628 27860
rect 19684 27804 20636 27860
rect 20692 27804 20702 27860
rect 20860 27804 23100 27860
rect 23156 27804 23166 27860
rect 23426 27804 23436 27860
rect 23492 27804 24220 27860
rect 24276 27804 24286 27860
rect 28914 27804 28924 27860
rect 28980 27804 29484 27860
rect 29540 27804 29550 27860
rect 29922 27804 29932 27860
rect 29988 27804 30828 27860
rect 30884 27804 30894 27860
rect 31714 27804 31724 27860
rect 31780 27804 35196 27860
rect 35252 27804 35262 27860
rect 38322 27804 38332 27860
rect 38388 27804 39564 27860
rect 39620 27804 39630 27860
rect 40002 27804 40012 27860
rect 40068 27804 40236 27860
rect 40292 27804 44716 27860
rect 44772 27804 44782 27860
rect 45042 27804 45052 27860
rect 45108 27804 52556 27860
rect 52612 27804 52622 27860
rect 53330 27804 53340 27860
rect 53396 27804 55076 27860
rect 20860 27748 20916 27804
rect 55020 27748 55076 27804
rect 2930 27692 2940 27748
rect 2996 27692 4396 27748
rect 4452 27692 4462 27748
rect 4620 27692 6972 27748
rect 7028 27692 7038 27748
rect 7196 27692 8540 27748
rect 8596 27692 8606 27748
rect 8866 27692 8876 27748
rect 8932 27692 10332 27748
rect 10388 27692 10398 27748
rect 12114 27692 12124 27748
rect 12180 27692 13020 27748
rect 13076 27692 13086 27748
rect 14242 27692 14252 27748
rect 14308 27692 15148 27748
rect 15204 27692 15214 27748
rect 16034 27692 16044 27748
rect 16100 27692 20916 27748
rect 22194 27692 22204 27748
rect 22260 27692 24780 27748
rect 24836 27692 24846 27748
rect 27906 27692 27916 27748
rect 27972 27692 40964 27748
rect 41570 27692 41580 27748
rect 41636 27692 43372 27748
rect 43428 27692 43438 27748
rect 43586 27692 43596 27748
rect 43652 27692 48860 27748
rect 48916 27692 48926 27748
rect 51874 27692 51884 27748
rect 51940 27692 53340 27748
rect 53396 27692 53406 27748
rect 55010 27692 55020 27748
rect 55076 27692 55132 27748
rect 55188 27692 55198 27748
rect 0 27636 112 27664
rect 4620 27636 4676 27692
rect 7196 27636 7252 27692
rect 40908 27636 40964 27692
rect 57344 27636 57456 27664
rect 0 27580 4676 27636
rect 5506 27580 5516 27636
rect 5572 27580 5964 27636
rect 6020 27580 6030 27636
rect 6178 27580 6188 27636
rect 6244 27580 7252 27636
rect 8418 27580 8428 27636
rect 8484 27580 10892 27636
rect 10948 27580 10958 27636
rect 11218 27580 11228 27636
rect 11284 27580 14140 27636
rect 14196 27580 14206 27636
rect 14354 27580 14364 27636
rect 14420 27580 16604 27636
rect 16660 27580 16670 27636
rect 17378 27580 17388 27636
rect 17444 27580 17948 27636
rect 18004 27580 19404 27636
rect 19460 27580 19470 27636
rect 19628 27580 29596 27636
rect 29652 27580 29662 27636
rect 31826 27580 31836 27636
rect 31892 27580 34524 27636
rect 34580 27580 35420 27636
rect 35476 27580 35486 27636
rect 40562 27580 40572 27636
rect 40628 27580 40684 27636
rect 40740 27580 40750 27636
rect 40908 27580 56028 27636
rect 56084 27580 56094 27636
rect 57138 27580 57148 27636
rect 57204 27580 57456 27636
rect 0 27552 112 27580
rect 19628 27524 19684 27580
rect 57344 27552 57456 27580
rect 1558 27468 1596 27524
rect 1652 27468 1662 27524
rect 4946 27468 4956 27524
rect 5012 27468 5740 27524
rect 5796 27468 7084 27524
rect 7140 27468 7150 27524
rect 7970 27468 7980 27524
rect 8036 27468 9660 27524
rect 9716 27468 9726 27524
rect 11666 27468 11676 27524
rect 11732 27468 19684 27524
rect 20038 27468 20076 27524
rect 20132 27468 20142 27524
rect 21298 27468 21308 27524
rect 21364 27468 21756 27524
rect 21812 27468 21822 27524
rect 23090 27468 23100 27524
rect 23156 27468 24220 27524
rect 24276 27468 24286 27524
rect 24882 27468 24892 27524
rect 24948 27468 25508 27524
rect 26898 27468 26908 27524
rect 26964 27468 27132 27524
rect 27188 27468 27198 27524
rect 30258 27468 30268 27524
rect 30324 27468 31388 27524
rect 31444 27468 31454 27524
rect 33730 27468 33740 27524
rect 33796 27468 35868 27524
rect 35924 27468 35934 27524
rect 36316 27468 41132 27524
rect 41188 27468 41198 27524
rect 43474 27468 43484 27524
rect 43540 27468 44156 27524
rect 44212 27468 44222 27524
rect 45602 27468 45612 27524
rect 45668 27468 46284 27524
rect 46340 27468 46350 27524
rect 47282 27468 47292 27524
rect 47348 27468 52780 27524
rect 52836 27468 52846 27524
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 25452 27412 25508 27468
rect 588 27356 3724 27412
rect 3780 27356 4340 27412
rect 4946 27356 4956 27412
rect 5012 27356 5292 27412
rect 5348 27356 5358 27412
rect 7158 27356 7196 27412
rect 7252 27356 10892 27412
rect 10948 27356 10958 27412
rect 11890 27356 11900 27412
rect 11956 27356 13020 27412
rect 13076 27356 13086 27412
rect 18386 27356 18396 27412
rect 18452 27356 20524 27412
rect 20580 27356 20590 27412
rect 20962 27356 20972 27412
rect 21028 27356 21532 27412
rect 21588 27356 21598 27412
rect 22082 27356 22092 27412
rect 22148 27356 22316 27412
rect 22372 27356 22988 27412
rect 23044 27356 23054 27412
rect 23202 27356 23212 27412
rect 23268 27356 23884 27412
rect 23940 27356 24332 27412
rect 24388 27356 24398 27412
rect 24882 27356 24892 27412
rect 24948 27356 25228 27412
rect 25284 27356 25294 27412
rect 25452 27356 28924 27412
rect 28980 27356 28990 27412
rect 30258 27356 30268 27412
rect 30324 27356 35532 27412
rect 35588 27356 35598 27412
rect 0 27188 112 27216
rect 588 27188 644 27356
rect 4284 27300 4340 27356
rect 36316 27300 36372 27468
rect 44454 27412 44464 27468
rect 44520 27412 44568 27468
rect 44624 27412 44672 27468
rect 44728 27412 44738 27468
rect 36530 27356 36540 27412
rect 36596 27356 37100 27412
rect 37156 27356 41804 27412
rect 41860 27356 41870 27412
rect 42130 27356 42140 27412
rect 42196 27356 44324 27412
rect 44268 27300 44324 27356
rect 44828 27356 49084 27412
rect 49140 27356 49150 27412
rect 49410 27356 49420 27412
rect 49476 27356 50876 27412
rect 50932 27356 50988 27412
rect 51044 27356 51054 27412
rect 51212 27356 53228 27412
rect 53284 27356 53294 27412
rect 53778 27356 53788 27412
rect 53844 27356 54348 27412
rect 54404 27356 54414 27412
rect 44828 27300 44884 27356
rect 51212 27300 51268 27356
rect 3042 27244 3052 27300
rect 3108 27244 3948 27300
rect 4004 27244 4014 27300
rect 4284 27244 6860 27300
rect 6916 27244 6926 27300
rect 7084 27244 10108 27300
rect 10164 27244 10780 27300
rect 10836 27244 10846 27300
rect 12226 27244 12236 27300
rect 12292 27244 13916 27300
rect 13972 27244 13982 27300
rect 17042 27244 17052 27300
rect 17108 27244 25116 27300
rect 25172 27244 25182 27300
rect 26338 27244 26348 27300
rect 26404 27244 28980 27300
rect 30370 27244 30380 27300
rect 30436 27244 36372 27300
rect 38658 27244 38668 27300
rect 38724 27244 38892 27300
rect 38948 27244 40236 27300
rect 40292 27244 40302 27300
rect 41122 27244 41132 27300
rect 41188 27244 43876 27300
rect 44268 27244 44884 27300
rect 45154 27244 45164 27300
rect 45220 27244 45500 27300
rect 45556 27244 45566 27300
rect 45714 27244 45724 27300
rect 45780 27244 46172 27300
rect 46228 27244 46238 27300
rect 49858 27244 49868 27300
rect 49924 27244 51268 27300
rect 53218 27244 53228 27300
rect 53284 27244 55020 27300
rect 55076 27244 55086 27300
rect 7084 27188 7140 27244
rect 28924 27188 28980 27244
rect 43820 27188 43876 27244
rect 57344 27188 57456 27216
rect 0 27132 644 27188
rect 1698 27132 1708 27188
rect 1764 27132 3164 27188
rect 3220 27132 3230 27188
rect 3602 27132 3612 27188
rect 3668 27132 4956 27188
rect 5012 27132 5022 27188
rect 6290 27132 6300 27188
rect 6356 27132 7140 27188
rect 7970 27132 7980 27188
rect 8036 27132 8988 27188
rect 9044 27132 9054 27188
rect 11890 27132 11900 27188
rect 11956 27132 12460 27188
rect 12516 27132 12526 27188
rect 12786 27132 12796 27188
rect 12852 27132 16380 27188
rect 16436 27132 16446 27188
rect 16594 27132 16604 27188
rect 16660 27132 17164 27188
rect 17220 27132 17230 27188
rect 18946 27132 18956 27188
rect 19012 27132 19852 27188
rect 19908 27132 19918 27188
rect 20514 27132 20524 27188
rect 20580 27132 21308 27188
rect 21364 27132 21532 27188
rect 21588 27132 21598 27188
rect 21858 27132 21868 27188
rect 21924 27132 22316 27188
rect 22372 27132 22382 27188
rect 22978 27132 22988 27188
rect 23044 27132 25004 27188
rect 25060 27132 25070 27188
rect 25340 27132 26124 27188
rect 26180 27132 26190 27188
rect 26562 27132 26572 27188
rect 26628 27132 27580 27188
rect 27636 27132 28700 27188
rect 28756 27132 28766 27188
rect 28924 27132 30940 27188
rect 30996 27132 31006 27188
rect 31714 27132 31724 27188
rect 31780 27132 32508 27188
rect 32564 27132 32574 27188
rect 32946 27132 32956 27188
rect 33012 27132 34188 27188
rect 34244 27132 34254 27188
rect 34738 27132 34748 27188
rect 34804 27132 35196 27188
rect 35252 27132 35262 27188
rect 36316 27132 38220 27188
rect 38276 27132 38286 27188
rect 38434 27132 38444 27188
rect 38500 27132 39564 27188
rect 39620 27132 39630 27188
rect 40562 27132 40572 27188
rect 40628 27132 41468 27188
rect 41524 27132 42252 27188
rect 42308 27132 42318 27188
rect 43250 27132 43260 27188
rect 43316 27132 43596 27188
rect 43652 27132 43662 27188
rect 43820 27132 51772 27188
rect 51828 27132 51838 27188
rect 52658 27132 52668 27188
rect 52724 27132 53116 27188
rect 53172 27132 53182 27188
rect 53554 27132 53564 27188
rect 53620 27132 54236 27188
rect 54292 27132 54302 27188
rect 57026 27132 57036 27188
rect 57092 27132 57456 27188
rect 0 27104 112 27132
rect 25340 27076 25396 27132
rect 36316 27076 36372 27132
rect 57344 27104 57456 27132
rect 1026 27020 1036 27076
rect 1092 27020 4340 27076
rect 4610 27020 4620 27076
rect 4676 27020 4844 27076
rect 4900 27020 6412 27076
rect 6468 27020 6478 27076
rect 6962 27020 6972 27076
rect 7028 27020 7868 27076
rect 7924 27020 7934 27076
rect 9538 27020 9548 27076
rect 9604 27020 10668 27076
rect 10724 27020 10734 27076
rect 11442 27020 11452 27076
rect 11508 27020 12908 27076
rect 12964 27020 12974 27076
rect 13570 27020 13580 27076
rect 13636 27020 17612 27076
rect 17668 27020 17678 27076
rect 18050 27020 18060 27076
rect 18116 27020 18284 27076
rect 18340 27020 18732 27076
rect 18788 27020 18798 27076
rect 19170 27020 19180 27076
rect 19236 27020 25396 27076
rect 25554 27020 25564 27076
rect 25620 27020 26908 27076
rect 26964 27020 26974 27076
rect 29586 27020 29596 27076
rect 29652 27020 31836 27076
rect 31892 27020 31902 27076
rect 33506 27020 33516 27076
rect 33572 27020 36372 27076
rect 39554 27020 39564 27076
rect 39620 27020 40236 27076
rect 40292 27020 40302 27076
rect 40674 27020 40684 27076
rect 40740 27020 41132 27076
rect 41188 27020 41198 27076
rect 41682 27020 41692 27076
rect 41748 27020 42028 27076
rect 42084 27020 42094 27076
rect 42802 27020 42812 27076
rect 42868 27020 45500 27076
rect 45556 27020 45612 27076
rect 45668 27020 45678 27076
rect 49410 27020 49420 27076
rect 49476 27020 51100 27076
rect 51156 27020 51166 27076
rect 55234 27020 55244 27076
rect 55300 27020 56140 27076
rect 56196 27020 56206 27076
rect 3938 26908 3948 26964
rect 4004 26908 4228 26964
rect 2818 26796 2828 26852
rect 2884 26796 3836 26852
rect 3892 26796 3902 26852
rect 0 26740 112 26768
rect 4172 26740 4228 26908
rect 4284 26852 4340 27020
rect 4946 26908 4956 26964
rect 5012 26908 5180 26964
rect 5236 26908 5246 26964
rect 5394 26908 5404 26964
rect 5460 26908 10444 26964
rect 10500 26908 10510 26964
rect 10770 26908 10780 26964
rect 10836 26908 13972 26964
rect 14354 26908 14364 26964
rect 14420 26908 16156 26964
rect 16212 26908 16222 26964
rect 16828 26908 18396 26964
rect 18452 26908 18462 26964
rect 20514 26908 20524 26964
rect 20580 26908 21700 26964
rect 22306 26908 22316 26964
rect 22372 26908 23660 26964
rect 23716 26908 23726 26964
rect 24892 26908 26348 26964
rect 26404 26908 26414 26964
rect 27346 26908 27356 26964
rect 27412 26908 29708 26964
rect 29764 26908 29774 26964
rect 31378 26908 31388 26964
rect 31444 26908 31948 26964
rect 32722 26908 32732 26964
rect 32788 26908 34076 26964
rect 34132 26908 34142 26964
rect 34402 26908 34412 26964
rect 34468 26908 34748 26964
rect 34804 26908 34814 26964
rect 35746 26908 35756 26964
rect 35812 26908 38556 26964
rect 38612 26908 38622 26964
rect 38882 26908 38892 26964
rect 38948 26908 39228 26964
rect 39284 26908 39294 26964
rect 39890 26908 39900 26964
rect 39956 26908 40124 26964
rect 40180 26908 40190 26964
rect 41346 26908 41356 26964
rect 41412 26908 43260 26964
rect 43316 26908 43326 26964
rect 43586 26908 43596 26964
rect 43652 26908 44100 26964
rect 45378 26908 45388 26964
rect 45444 26908 48188 26964
rect 48244 26908 48254 26964
rect 50428 26908 53452 26964
rect 53508 26908 53518 26964
rect 55346 26908 55356 26964
rect 55412 26908 55916 26964
rect 55972 26908 55982 26964
rect 13916 26852 13972 26908
rect 4284 26796 6636 26852
rect 6692 26796 6702 26852
rect 7746 26796 7756 26852
rect 7812 26796 11676 26852
rect 11732 26796 11742 26852
rect 12114 26796 12124 26852
rect 12180 26796 12460 26852
rect 12516 26796 12526 26852
rect 12898 26796 12908 26852
rect 12964 26796 13244 26852
rect 13300 26796 13310 26852
rect 13916 26796 14924 26852
rect 14980 26796 15036 26852
rect 15092 26796 15102 26852
rect 16828 26740 16884 26908
rect 21644 26852 21812 26908
rect 24892 26852 24948 26908
rect 31892 26852 31948 26908
rect 44044 26852 44100 26908
rect 50428 26852 50484 26908
rect 17378 26796 17388 26852
rect 17444 26796 21308 26852
rect 21364 26796 21374 26852
rect 21756 26796 24948 26852
rect 25106 26796 25116 26852
rect 25172 26796 30268 26852
rect 30324 26796 30334 26852
rect 31892 26796 33852 26852
rect 33908 26796 33918 26852
rect 34850 26796 34860 26852
rect 34916 26796 34972 26852
rect 35028 26796 35038 26852
rect 35634 26796 35644 26852
rect 35700 26796 39004 26852
rect 39060 26796 39070 26852
rect 39330 26796 39340 26852
rect 39396 26796 39676 26852
rect 39732 26796 39742 26852
rect 40450 26796 40460 26852
rect 40516 26796 43148 26852
rect 43204 26796 43214 26852
rect 44044 26796 50484 26852
rect 50642 26796 50652 26852
rect 50708 26796 54012 26852
rect 54068 26796 54078 26852
rect 57344 26740 57456 26768
rect 0 26684 3388 26740
rect 4172 26684 5180 26740
rect 5236 26684 5246 26740
rect 6850 26684 6860 26740
rect 6916 26684 7140 26740
rect 7298 26684 7308 26740
rect 7364 26684 7644 26740
rect 7700 26684 9548 26740
rect 9604 26684 9614 26740
rect 10546 26684 10556 26740
rect 10612 26684 13132 26740
rect 13188 26684 16884 26740
rect 17602 26684 17612 26740
rect 17668 26684 20524 26740
rect 20580 26684 20590 26740
rect 20962 26684 20972 26740
rect 21028 26684 21756 26740
rect 21812 26684 21822 26740
rect 24882 26684 24892 26740
rect 24948 26684 28476 26740
rect 28532 26684 28542 26740
rect 28690 26684 28700 26740
rect 28756 26684 31276 26740
rect 31332 26684 31342 26740
rect 31490 26684 31500 26740
rect 31556 26684 32844 26740
rect 32900 26684 38108 26740
rect 38164 26684 38174 26740
rect 38882 26684 38892 26740
rect 38948 26684 39228 26740
rect 39284 26684 39294 26740
rect 39442 26684 39452 26740
rect 39508 26684 40572 26740
rect 40628 26684 40638 26740
rect 45378 26684 45388 26740
rect 45444 26684 53676 26740
rect 53732 26684 53742 26740
rect 54450 26684 54460 26740
rect 54516 26684 55244 26740
rect 55300 26684 55310 26740
rect 56578 26684 56588 26740
rect 56644 26684 57456 26740
rect 0 26656 112 26684
rect 3332 26516 3388 26684
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 7084 26628 7140 26684
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 43794 26628 43804 26684
rect 43860 26628 43908 26684
rect 43964 26628 44012 26684
rect 44068 26628 44078 26684
rect 57344 26656 57456 26684
rect 3490 26572 3500 26628
rect 3556 26572 3594 26628
rect 4386 26572 4396 26628
rect 4452 26572 5348 26628
rect 7084 26572 8540 26628
rect 8596 26572 13580 26628
rect 13636 26572 13646 26628
rect 14130 26572 14140 26628
rect 14196 26572 15820 26628
rect 15876 26572 15886 26628
rect 17602 26572 17612 26628
rect 17668 26572 22260 26628
rect 24210 26572 24220 26628
rect 24276 26572 25900 26628
rect 25956 26572 25966 26628
rect 29026 26572 29036 26628
rect 29092 26572 29540 26628
rect 29698 26572 29708 26628
rect 29764 26572 31612 26628
rect 31668 26572 36092 26628
rect 36148 26572 38556 26628
rect 38612 26572 38622 26628
rect 38994 26572 39004 26628
rect 39060 26572 41468 26628
rect 41524 26572 41534 26628
rect 44258 26572 44268 26628
rect 44324 26572 44660 26628
rect 44930 26572 44940 26628
rect 44996 26572 45276 26628
rect 45332 26572 45342 26628
rect 46610 26572 46620 26628
rect 46676 26572 52220 26628
rect 52276 26572 52286 26628
rect 52434 26572 52444 26628
rect 52500 26572 52556 26628
rect 52612 26572 52622 26628
rect 52882 26572 52892 26628
rect 52948 26572 55580 26628
rect 55636 26572 55646 26628
rect 3332 26460 4956 26516
rect 5012 26460 5022 26516
rect 5292 26404 5348 26572
rect 7186 26460 7196 26516
rect 7252 26460 7868 26516
rect 7924 26460 7934 26516
rect 8418 26460 8428 26516
rect 8484 26460 9772 26516
rect 9828 26460 9838 26516
rect 10658 26460 10668 26516
rect 10724 26460 16044 26516
rect 16100 26460 16110 26516
rect 16258 26460 16268 26516
rect 16324 26460 18956 26516
rect 19012 26460 19022 26516
rect 20850 26460 20860 26516
rect 20916 26460 21196 26516
rect 21252 26460 21262 26516
rect 22204 26404 22260 26572
rect 29484 26516 29540 26572
rect 44604 26516 44660 26572
rect 29484 26460 29820 26516
rect 29876 26460 29886 26516
rect 33842 26460 33852 26516
rect 33908 26460 35420 26516
rect 35476 26460 35486 26516
rect 38098 26460 38108 26516
rect 38164 26460 40404 26516
rect 40786 26460 40796 26516
rect 40852 26460 41524 26516
rect 43586 26460 43596 26516
rect 43652 26460 44380 26516
rect 44436 26460 44446 26516
rect 44604 26460 46508 26516
rect 46564 26460 46574 26516
rect 47618 26460 47628 26516
rect 47684 26460 48188 26516
rect 48244 26460 48254 26516
rect 48412 26460 49308 26516
rect 49364 26460 53788 26516
rect 53844 26460 53854 26516
rect 33852 26404 33908 26460
rect 3042 26348 3052 26404
rect 3108 26348 4956 26404
rect 5012 26348 5022 26404
rect 5292 26348 5628 26404
rect 5684 26348 6188 26404
rect 6244 26348 6254 26404
rect 6850 26348 6860 26404
rect 6916 26348 19740 26404
rect 19796 26348 19806 26404
rect 20066 26348 20076 26404
rect 20132 26348 21868 26404
rect 21924 26348 21934 26404
rect 22204 26348 25564 26404
rect 25620 26348 25630 26404
rect 31892 26348 33908 26404
rect 34178 26348 34188 26404
rect 34244 26348 36932 26404
rect 37874 26348 37884 26404
rect 37940 26348 39676 26404
rect 39732 26348 39742 26404
rect 0 26292 112 26320
rect 31892 26292 31948 26348
rect 0 26236 2716 26292
rect 2772 26236 2782 26292
rect 4386 26236 4396 26292
rect 4452 26236 5068 26292
rect 5124 26236 5134 26292
rect 5842 26236 5852 26292
rect 5908 26236 8092 26292
rect 8148 26236 8158 26292
rect 8306 26236 8316 26292
rect 8372 26236 9660 26292
rect 9716 26236 9726 26292
rect 12674 26236 12684 26292
rect 12740 26236 13244 26292
rect 13300 26236 13310 26292
rect 15362 26236 15372 26292
rect 15428 26236 16828 26292
rect 16884 26236 16894 26292
rect 21186 26236 21196 26292
rect 21252 26236 21644 26292
rect 21700 26236 21710 26292
rect 21858 26236 21868 26292
rect 21924 26236 26908 26292
rect 27794 26236 27804 26292
rect 27860 26236 29036 26292
rect 29092 26236 29102 26292
rect 29698 26236 29708 26292
rect 29764 26236 31948 26292
rect 32386 26236 32396 26292
rect 32452 26236 32732 26292
rect 32788 26236 32798 26292
rect 32946 26236 32956 26292
rect 33012 26236 34412 26292
rect 34468 26236 34478 26292
rect 35298 26236 35308 26292
rect 35364 26236 36540 26292
rect 36596 26236 36606 26292
rect 0 26208 112 26236
rect 26852 26180 26908 26236
rect 36876 26180 36932 26348
rect 40348 26292 40404 26460
rect 41468 26404 41524 26460
rect 48412 26404 48468 26460
rect 41458 26348 41468 26404
rect 41524 26348 41534 26404
rect 44146 26348 44156 26404
rect 44212 26348 44940 26404
rect 44996 26348 45006 26404
rect 45332 26348 48468 26404
rect 52546 26348 52556 26404
rect 52612 26348 54796 26404
rect 54852 26348 54862 26404
rect 45332 26292 45388 26348
rect 57344 26292 57456 26320
rect 37202 26236 37212 26292
rect 37268 26236 40124 26292
rect 40180 26236 40190 26292
rect 40348 26236 42700 26292
rect 42756 26236 44604 26292
rect 44660 26236 44670 26292
rect 44818 26236 44828 26292
rect 44884 26236 45388 26292
rect 45602 26236 45612 26292
rect 45668 26236 47180 26292
rect 47236 26236 47246 26292
rect 52658 26236 52668 26292
rect 52724 26236 53900 26292
rect 53956 26236 53966 26292
rect 55570 26236 55580 26292
rect 55636 26236 56140 26292
rect 56196 26236 56206 26292
rect 56914 26236 56924 26292
rect 56980 26236 57456 26292
rect 57344 26208 57456 26236
rect 2482 26124 2492 26180
rect 2548 26124 7196 26180
rect 7252 26124 7262 26180
rect 7410 26124 7420 26180
rect 7476 26124 8764 26180
rect 8820 26124 8830 26180
rect 8978 26124 8988 26180
rect 9044 26124 9772 26180
rect 9828 26124 10332 26180
rect 10388 26124 10398 26180
rect 12226 26124 12236 26180
rect 12292 26124 12572 26180
rect 12628 26124 12638 26180
rect 13570 26124 13580 26180
rect 13636 26124 17612 26180
rect 17668 26124 17678 26180
rect 17938 26124 17948 26180
rect 18004 26124 22988 26180
rect 23044 26124 23054 26180
rect 23426 26124 23436 26180
rect 23492 26124 24220 26180
rect 24276 26124 24286 26180
rect 24434 26124 24444 26180
rect 24500 26124 25004 26180
rect 25060 26124 25070 26180
rect 26226 26124 26236 26180
rect 26292 26124 26572 26180
rect 26628 26124 26638 26180
rect 26852 26124 30044 26180
rect 30100 26124 30110 26180
rect 31154 26124 31164 26180
rect 31220 26124 35644 26180
rect 35700 26124 35710 26180
rect 35970 26124 35980 26180
rect 36036 26124 36652 26180
rect 36708 26124 36718 26180
rect 36876 26124 36988 26180
rect 37044 26124 38108 26180
rect 38164 26124 38174 26180
rect 38322 26124 38332 26180
rect 38388 26124 39004 26180
rect 39060 26124 39070 26180
rect 41234 26124 41244 26180
rect 41300 26124 41692 26180
rect 41748 26124 43372 26180
rect 43428 26124 43438 26180
rect 43698 26124 43708 26180
rect 43764 26124 50092 26180
rect 50148 26124 50158 26180
rect 50372 26124 52556 26180
rect 52612 26124 52622 26180
rect 53554 26124 53564 26180
rect 53620 26124 54236 26180
rect 54292 26124 54302 26180
rect 1362 26012 1372 26068
rect 1428 26012 1708 26068
rect 1764 26012 1774 26068
rect 2706 26012 2716 26068
rect 2772 26012 8036 26068
rect 9538 26012 9548 26068
rect 9604 26012 13132 26068
rect 13188 26012 13198 26068
rect 15250 26012 15260 26068
rect 15316 26012 16604 26068
rect 16660 26012 16670 26068
rect 17490 26012 17500 26068
rect 17556 26012 19516 26068
rect 19572 26012 19582 26068
rect 19730 26012 19740 26068
rect 19796 26012 30156 26068
rect 30212 26012 30222 26068
rect 30930 26012 30940 26068
rect 30996 26012 33068 26068
rect 33124 26012 33134 26068
rect 33282 26012 33292 26068
rect 33348 26012 35196 26068
rect 35252 26012 35262 26068
rect 38882 26012 38892 26068
rect 38948 26012 39284 26068
rect 40450 26012 40460 26068
rect 40516 26012 43260 26068
rect 43316 26012 43326 26068
rect 43474 26012 43484 26068
rect 43540 26012 48188 26068
rect 48244 26012 48254 26068
rect 3042 25900 3052 25956
rect 3108 25900 3276 25956
rect 3332 25900 3342 25956
rect 4946 25900 4956 25956
rect 5012 25900 5516 25956
rect 5572 25900 5582 25956
rect 6066 25900 6076 25956
rect 6132 25900 7084 25956
rect 7140 25900 7150 25956
rect 0 25844 112 25872
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 7980 25844 8036 26012
rect 30940 25956 30996 26012
rect 8194 25900 8204 25956
rect 8260 25900 10108 25956
rect 10164 25900 10174 25956
rect 10770 25900 10780 25956
rect 10836 25900 11676 25956
rect 11732 25900 14364 25956
rect 14420 25900 14430 25956
rect 14588 25900 15596 25956
rect 15652 25900 15662 25956
rect 16818 25900 16828 25956
rect 16884 25900 20748 25956
rect 20804 25900 21308 25956
rect 21364 25900 21374 25956
rect 22194 25900 22204 25956
rect 22260 25900 23436 25956
rect 23492 25900 23502 25956
rect 28578 25900 28588 25956
rect 28644 25900 30996 25956
rect 39228 25956 39284 26012
rect 50372 25956 50428 26124
rect 52210 26012 52220 26068
rect 52276 26012 54348 26068
rect 54404 26012 54414 26068
rect 39228 25900 43708 25956
rect 43764 25900 43774 25956
rect 44828 25900 50428 25956
rect 14588 25844 14644 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 44454 25844 44464 25900
rect 44520 25844 44568 25900
rect 44624 25844 44672 25900
rect 44728 25844 44738 25900
rect 0 25788 3388 25844
rect 3826 25788 3836 25844
rect 3892 25788 4284 25844
rect 4340 25788 4350 25844
rect 4834 25788 4844 25844
rect 4900 25788 5404 25844
rect 5460 25788 5470 25844
rect 5618 25788 5628 25844
rect 5684 25788 7308 25844
rect 7364 25788 7374 25844
rect 7522 25788 7532 25844
rect 7588 25788 7756 25844
rect 7812 25788 7822 25844
rect 7980 25788 11900 25844
rect 11956 25788 11966 25844
rect 12786 25788 12796 25844
rect 12852 25788 13244 25844
rect 13300 25788 13310 25844
rect 13458 25788 13468 25844
rect 13524 25788 14644 25844
rect 15092 25788 21868 25844
rect 21924 25788 21934 25844
rect 22306 25788 22316 25844
rect 22372 25788 22428 25844
rect 22484 25788 22494 25844
rect 23090 25788 23100 25844
rect 23156 25788 24332 25844
rect 24388 25788 24398 25844
rect 28018 25788 28028 25844
rect 28084 25788 31500 25844
rect 31556 25788 31566 25844
rect 32274 25788 32284 25844
rect 32340 25788 33740 25844
rect 33796 25788 34748 25844
rect 34804 25788 34814 25844
rect 35186 25788 35196 25844
rect 35252 25788 36092 25844
rect 36148 25788 36316 25844
rect 36372 25788 36382 25844
rect 39666 25788 39676 25844
rect 39732 25788 40124 25844
rect 40180 25788 40190 25844
rect 40450 25788 40460 25844
rect 40516 25788 41468 25844
rect 41524 25788 41534 25844
rect 0 25760 112 25788
rect 3332 25732 3388 25788
rect 15092 25732 15148 25788
rect 44828 25732 44884 25900
rect 57344 25844 57456 25872
rect 45350 25788 45388 25844
rect 45444 25788 45454 25844
rect 50306 25788 50316 25844
rect 50372 25788 54796 25844
rect 54852 25788 54862 25844
rect 55682 25788 55692 25844
rect 55748 25788 57456 25844
rect 57344 25760 57456 25788
rect 802 25676 812 25732
rect 868 25676 878 25732
rect 1698 25676 1708 25732
rect 1764 25676 1820 25732
rect 1876 25676 1886 25732
rect 3332 25676 15148 25732
rect 16034 25676 16044 25732
rect 16100 25676 17052 25732
rect 17108 25676 17118 25732
rect 18498 25676 18508 25732
rect 18564 25676 20412 25732
rect 20468 25676 20478 25732
rect 20626 25676 20636 25732
rect 20692 25676 24780 25732
rect 24836 25676 24846 25732
rect 25890 25676 25900 25732
rect 25956 25676 26796 25732
rect 26852 25676 26862 25732
rect 29250 25676 29260 25732
rect 29316 25676 29372 25732
rect 29428 25676 33628 25732
rect 33684 25676 33694 25732
rect 33842 25676 33852 25732
rect 33908 25676 35308 25732
rect 35364 25676 35374 25732
rect 36530 25676 36540 25732
rect 36596 25676 38780 25732
rect 38836 25676 38846 25732
rect 40674 25676 40684 25732
rect 40740 25676 41804 25732
rect 41860 25676 41870 25732
rect 42018 25676 42028 25732
rect 42084 25676 42476 25732
rect 42532 25676 42542 25732
rect 43362 25676 43372 25732
rect 43428 25676 44884 25732
rect 45490 25676 45500 25732
rect 45556 25676 49308 25732
rect 49364 25676 49644 25732
rect 49700 25676 49868 25732
rect 49924 25676 49934 25732
rect 50306 25676 50316 25732
rect 50372 25676 50540 25732
rect 50596 25676 53564 25732
rect 53620 25676 53630 25732
rect 812 25620 868 25676
rect 812 25564 4452 25620
rect 4610 25564 4620 25620
rect 4676 25564 5292 25620
rect 5348 25564 5358 25620
rect 6290 25564 6300 25620
rect 6356 25564 6972 25620
rect 7028 25564 7868 25620
rect 7924 25564 7934 25620
rect 8866 25564 8876 25620
rect 8932 25564 9884 25620
rect 9940 25564 9950 25620
rect 11554 25564 11564 25620
rect 11620 25564 13356 25620
rect 13412 25564 13422 25620
rect 13906 25564 13916 25620
rect 13972 25564 14364 25620
rect 14420 25564 14700 25620
rect 14756 25564 14766 25620
rect 16146 25564 16156 25620
rect 16212 25564 17724 25620
rect 17780 25564 17790 25620
rect 19954 25564 19964 25620
rect 20020 25564 20972 25620
rect 21028 25564 21038 25620
rect 21186 25564 21196 25620
rect 21252 25564 22876 25620
rect 22932 25564 22942 25620
rect 23650 25564 23660 25620
rect 23716 25564 28252 25620
rect 28308 25564 28318 25620
rect 28690 25564 28700 25620
rect 28756 25564 29036 25620
rect 29092 25564 29102 25620
rect 31500 25564 32396 25620
rect 32452 25564 32462 25620
rect 32946 25564 32956 25620
rect 33012 25564 33180 25620
rect 33236 25564 33516 25620
rect 33572 25564 33582 25620
rect 34822 25564 34860 25620
rect 34916 25564 34926 25620
rect 35410 25564 35420 25620
rect 35476 25564 36764 25620
rect 36820 25564 36830 25620
rect 37202 25564 37212 25620
rect 37268 25564 37548 25620
rect 37604 25564 37614 25620
rect 38444 25564 39620 25620
rect 40114 25564 40124 25620
rect 40180 25564 40796 25620
rect 40852 25564 40862 25620
rect 41010 25564 41020 25620
rect 41076 25564 42700 25620
rect 42756 25564 42766 25620
rect 44034 25564 44044 25620
rect 44100 25564 53004 25620
rect 53060 25564 53070 25620
rect 53862 25564 53900 25620
rect 53956 25564 53966 25620
rect 4396 25508 4452 25564
rect 802 25452 812 25508
rect 868 25452 1260 25508
rect 1316 25452 1326 25508
rect 3378 25452 3388 25508
rect 3444 25452 4172 25508
rect 4228 25452 4238 25508
rect 4396 25452 4956 25508
rect 5012 25452 5022 25508
rect 5170 25452 5180 25508
rect 5236 25452 7420 25508
rect 7476 25452 7486 25508
rect 8754 25452 8764 25508
rect 8820 25452 9996 25508
rect 10052 25452 10062 25508
rect 11750 25452 11788 25508
rect 11844 25452 11854 25508
rect 12002 25452 12012 25508
rect 12068 25452 12106 25508
rect 12236 25452 16492 25508
rect 16548 25452 16558 25508
rect 17154 25452 17164 25508
rect 17220 25452 17500 25508
rect 17556 25452 17566 25508
rect 19394 25452 19404 25508
rect 19460 25452 19740 25508
rect 19796 25452 19806 25508
rect 19964 25452 20636 25508
rect 20692 25452 20702 25508
rect 21074 25452 21084 25508
rect 21140 25452 25228 25508
rect 25284 25452 25294 25508
rect 26674 25452 26684 25508
rect 26740 25452 28588 25508
rect 28644 25452 28654 25508
rect 0 25396 112 25424
rect 0 25340 2716 25396
rect 2772 25340 2782 25396
rect 3602 25340 3612 25396
rect 3668 25340 5628 25396
rect 5684 25340 5694 25396
rect 6066 25340 6076 25396
rect 6132 25340 7532 25396
rect 7588 25340 7598 25396
rect 7970 25340 7980 25396
rect 8036 25340 9548 25396
rect 9604 25340 9614 25396
rect 9762 25340 9772 25396
rect 9828 25340 11004 25396
rect 11060 25340 11070 25396
rect 0 25312 112 25340
rect 1586 25228 1596 25284
rect 1652 25228 4452 25284
rect 5506 25228 5516 25284
rect 5572 25228 7756 25284
rect 7812 25228 7822 25284
rect 8418 25228 8428 25284
rect 8484 25228 8540 25284
rect 8596 25228 8606 25284
rect 9202 25228 9212 25284
rect 9268 25228 9884 25284
rect 9940 25228 11340 25284
rect 11396 25228 11406 25284
rect 4396 25172 4452 25228
rect 12236 25172 12292 25452
rect 19964 25396 20020 25452
rect 31500 25396 31556 25564
rect 38444 25508 38500 25564
rect 39564 25508 39620 25564
rect 31714 25452 31724 25508
rect 31780 25452 32620 25508
rect 32676 25452 33740 25508
rect 33796 25452 35084 25508
rect 35140 25452 35150 25508
rect 36530 25452 36540 25508
rect 36596 25452 36988 25508
rect 37044 25452 37324 25508
rect 37380 25452 38500 25508
rect 39106 25452 39116 25508
rect 39172 25452 39340 25508
rect 39396 25452 39406 25508
rect 39564 25452 40292 25508
rect 40450 25452 40460 25508
rect 40516 25452 41244 25508
rect 41300 25452 41310 25508
rect 42578 25452 42588 25508
rect 42644 25452 43036 25508
rect 43092 25452 43102 25508
rect 43250 25452 43260 25508
rect 43316 25452 44156 25508
rect 44212 25452 45612 25508
rect 45668 25452 45678 25508
rect 49746 25452 49756 25508
rect 49812 25452 50540 25508
rect 50596 25452 50606 25508
rect 50978 25452 50988 25508
rect 51044 25452 51100 25508
rect 51156 25452 51166 25508
rect 40236 25396 40292 25452
rect 57344 25396 57456 25424
rect 12450 25340 12460 25396
rect 12516 25340 13244 25396
rect 13300 25340 13692 25396
rect 13748 25340 13758 25396
rect 18946 25340 18956 25396
rect 19012 25340 19404 25396
rect 19460 25340 20020 25396
rect 20514 25340 20524 25396
rect 20580 25340 25004 25396
rect 25060 25340 25070 25396
rect 26226 25340 26236 25396
rect 26292 25340 31556 25396
rect 31826 25340 31836 25396
rect 31892 25340 33628 25396
rect 33684 25340 34860 25396
rect 34916 25340 34926 25396
rect 35186 25340 35196 25396
rect 35252 25340 36428 25396
rect 36484 25340 36494 25396
rect 38098 25340 38108 25396
rect 38164 25340 39788 25396
rect 39844 25340 39854 25396
rect 40236 25340 41020 25396
rect 41076 25340 41086 25396
rect 41570 25340 41580 25396
rect 41636 25340 42700 25396
rect 42756 25340 42766 25396
rect 42914 25340 42924 25396
rect 42980 25340 45276 25396
rect 45332 25340 45342 25396
rect 47292 25340 50540 25396
rect 50596 25340 51772 25396
rect 51828 25340 51838 25396
rect 52098 25340 52108 25396
rect 52164 25340 55916 25396
rect 55972 25340 55982 25396
rect 57250 25340 57260 25396
rect 57316 25340 57456 25396
rect 13122 25228 13132 25284
rect 13188 25228 28644 25284
rect 28802 25228 28812 25284
rect 28868 25228 30828 25284
rect 30884 25228 30894 25284
rect 31714 25228 31724 25284
rect 31780 25228 34524 25284
rect 34580 25228 34590 25284
rect 34738 25228 34748 25284
rect 34804 25228 38332 25284
rect 38388 25228 38398 25284
rect 39302 25228 39340 25284
rect 39396 25228 39406 25284
rect 41794 25228 41804 25284
rect 41860 25228 47068 25284
rect 47124 25228 47134 25284
rect 28588 25172 28644 25228
rect 47292 25172 47348 25340
rect 57344 25312 57456 25340
rect 48178 25228 48188 25284
rect 48244 25228 50204 25284
rect 50260 25228 50270 25284
rect 51314 25228 51324 25284
rect 51380 25228 53732 25284
rect 55458 25228 55468 25284
rect 55524 25228 55804 25284
rect 55860 25228 55870 25284
rect 53676 25172 53732 25228
rect 2258 25116 2268 25172
rect 2324 25116 3388 25172
rect 3444 25116 3454 25172
rect 4396 25116 5852 25172
rect 5908 25116 5918 25172
rect 6076 25116 12292 25172
rect 15586 25116 15596 25172
rect 15652 25116 16492 25172
rect 16548 25116 16558 25172
rect 22642 25116 22652 25172
rect 22708 25116 23324 25172
rect 23380 25116 23390 25172
rect 24434 25116 24444 25172
rect 24500 25116 25228 25172
rect 25284 25116 26124 25172
rect 26180 25116 26190 25172
rect 28588 25116 29540 25172
rect 30146 25116 30156 25172
rect 30212 25116 38220 25172
rect 38276 25116 38286 25172
rect 44146 25116 44156 25172
rect 44212 25116 44940 25172
rect 44996 25116 45006 25172
rect 45378 25116 45388 25172
rect 45444 25116 45948 25172
rect 46004 25116 46014 25172
rect 46172 25116 47348 25172
rect 49410 25116 49420 25172
rect 49476 25116 51548 25172
rect 51604 25116 51614 25172
rect 53676 25116 54012 25172
rect 54068 25116 54078 25172
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 6076 25060 6132 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 4946 25004 4956 25060
rect 5012 25004 5292 25060
rect 5348 25004 5358 25060
rect 5506 25004 5516 25060
rect 5572 25004 6132 25060
rect 6402 25004 6412 25060
rect 6468 25004 10220 25060
rect 10276 25004 10286 25060
rect 11666 25004 11676 25060
rect 11732 25004 15148 25060
rect 15204 25004 15214 25060
rect 16370 25004 16380 25060
rect 16436 25004 23548 25060
rect 23604 25004 23614 25060
rect 28690 25004 28700 25060
rect 28756 25004 29260 25060
rect 29316 25004 29326 25060
rect 0 24948 112 24976
rect 28700 24948 28756 25004
rect 0 24892 15148 24948
rect 18834 24892 18844 24948
rect 18900 24892 19852 24948
rect 19908 24892 19918 24948
rect 20514 24892 20524 24948
rect 20580 24892 22092 24948
rect 22148 24892 22158 24948
rect 22306 24892 22316 24948
rect 22372 24892 22540 24948
rect 22596 24892 22606 24948
rect 22754 24892 22764 24948
rect 22820 24892 28756 24948
rect 0 24864 112 24892
rect 15092 24836 15148 24892
rect 29484 24836 29540 25116
rect 43794 25060 43804 25116
rect 43860 25060 43908 25116
rect 43964 25060 44012 25116
rect 44068 25060 44078 25116
rect 46172 25060 46228 25116
rect 30034 25004 30044 25060
rect 30100 25004 30716 25060
rect 30772 25004 30782 25060
rect 32246 25004 32284 25060
rect 32340 25004 32350 25060
rect 32946 25004 32956 25060
rect 33012 25004 34076 25060
rect 34132 25004 34972 25060
rect 35028 25004 35038 25060
rect 39638 25004 39676 25060
rect 39732 25004 39742 25060
rect 41570 25004 41580 25060
rect 41636 25004 41692 25060
rect 41748 25004 41758 25060
rect 42130 25004 42140 25060
rect 42196 25004 43260 25060
rect 43316 25004 43326 25060
rect 44146 25004 44156 25060
rect 44212 25004 46228 25060
rect 46386 25004 46396 25060
rect 46452 25004 52108 25060
rect 52164 25004 52174 25060
rect 57344 24948 57456 24976
rect 30482 24892 30492 24948
rect 30548 24892 44268 24948
rect 44324 24892 44334 24948
rect 50278 24892 50316 24948
rect 50372 24892 50382 24948
rect 50642 24892 50652 24948
rect 50708 24892 50988 24948
rect 51044 24892 52444 24948
rect 52500 24892 52510 24948
rect 56802 24892 56812 24948
rect 56868 24892 57456 24948
rect 57344 24864 57456 24892
rect 1698 24780 1708 24836
rect 1764 24780 5628 24836
rect 5684 24780 6188 24836
rect 6244 24780 6254 24836
rect 6850 24780 6860 24836
rect 6916 24780 9604 24836
rect 9762 24780 9772 24836
rect 9828 24780 11788 24836
rect 11844 24780 12236 24836
rect 12292 24780 12302 24836
rect 15092 24780 24892 24836
rect 24948 24780 24958 24836
rect 26114 24780 26124 24836
rect 26180 24780 29260 24836
rect 29316 24780 29326 24836
rect 29484 24780 33740 24836
rect 33796 24780 33806 24836
rect 34066 24780 34076 24836
rect 34132 24780 36540 24836
rect 36596 24780 36606 24836
rect 36754 24780 36764 24836
rect 36820 24780 37884 24836
rect 37940 24780 37950 24836
rect 38210 24780 38220 24836
rect 38276 24780 41580 24836
rect 41636 24780 41646 24836
rect 41906 24780 41916 24836
rect 41972 24780 42476 24836
rect 42532 24780 42542 24836
rect 43260 24780 44156 24836
rect 44212 24780 44222 24836
rect 47394 24780 47404 24836
rect 47460 24780 49756 24836
rect 49812 24780 49822 24836
rect 51090 24780 51100 24836
rect 51156 24780 53228 24836
rect 53284 24780 53294 24836
rect 54562 24780 54572 24836
rect 54628 24780 55244 24836
rect 55300 24780 55310 24836
rect 2118 24668 2156 24724
rect 2212 24668 2222 24724
rect 3266 24668 3276 24724
rect 3332 24668 3388 24724
rect 3444 24668 3454 24724
rect 3612 24668 4956 24724
rect 5012 24668 5022 24724
rect 5506 24668 5516 24724
rect 5572 24668 5964 24724
rect 6020 24668 7644 24724
rect 7700 24668 7710 24724
rect 3612 24612 3668 24668
rect 9548 24612 9604 24780
rect 43260 24724 43316 24780
rect 12898 24668 12908 24724
rect 12964 24668 16828 24724
rect 16884 24668 16894 24724
rect 19506 24668 19516 24724
rect 19572 24668 19628 24724
rect 19684 24668 19694 24724
rect 19954 24668 19964 24724
rect 20020 24668 22764 24724
rect 22820 24668 22830 24724
rect 24434 24668 24444 24724
rect 24500 24668 25340 24724
rect 25396 24668 26124 24724
rect 26180 24668 26190 24724
rect 27906 24668 27916 24724
rect 27972 24668 29036 24724
rect 29092 24668 31276 24724
rect 31332 24668 31342 24724
rect 31462 24668 31500 24724
rect 31556 24668 31566 24724
rect 32162 24668 32172 24724
rect 32228 24668 33740 24724
rect 33796 24668 33806 24724
rect 34710 24668 34748 24724
rect 34804 24668 34814 24724
rect 35186 24668 35196 24724
rect 35252 24668 36316 24724
rect 36372 24668 36382 24724
rect 37314 24668 37324 24724
rect 37380 24668 37660 24724
rect 37716 24668 43316 24724
rect 43586 24668 43596 24724
rect 43652 24668 50204 24724
rect 50260 24668 50652 24724
rect 50708 24668 51660 24724
rect 51716 24668 51726 24724
rect 1138 24556 1148 24612
rect 1204 24556 2492 24612
rect 2548 24556 2558 24612
rect 3154 24556 3164 24612
rect 3220 24556 3668 24612
rect 3938 24556 3948 24612
rect 4004 24556 5292 24612
rect 5348 24556 5358 24612
rect 5506 24556 5516 24612
rect 5572 24556 7756 24612
rect 7812 24556 7822 24612
rect 9548 24556 21028 24612
rect 21522 24556 21532 24612
rect 21588 24556 21644 24612
rect 21700 24556 21710 24612
rect 21858 24556 21868 24612
rect 21924 24556 24556 24612
rect 24612 24556 24622 24612
rect 24882 24556 24892 24612
rect 24948 24556 27356 24612
rect 27412 24556 27422 24612
rect 27794 24556 27804 24612
rect 27860 24556 29932 24612
rect 29988 24556 29998 24612
rect 32050 24556 32060 24612
rect 32116 24556 32284 24612
rect 32340 24556 32350 24612
rect 33058 24556 33068 24612
rect 33124 24556 33516 24612
rect 33572 24556 34412 24612
rect 34468 24556 34478 24612
rect 34626 24556 34636 24612
rect 34692 24556 34972 24612
rect 35028 24556 41356 24612
rect 41412 24556 41422 24612
rect 41570 24556 41580 24612
rect 41636 24556 41972 24612
rect 42242 24556 42252 24612
rect 42308 24556 45276 24612
rect 45332 24556 47684 24612
rect 47842 24556 47852 24612
rect 47908 24556 51212 24612
rect 51268 24556 51278 24612
rect 51650 24556 51660 24612
rect 51716 24556 54236 24612
rect 54292 24556 54302 24612
rect 0 24500 112 24528
rect 20972 24500 21028 24556
rect 41916 24500 41972 24556
rect 47628 24500 47684 24556
rect 57344 24500 57456 24528
rect 0 24444 15148 24500
rect 15698 24444 15708 24500
rect 15764 24444 16268 24500
rect 16324 24444 17052 24500
rect 17108 24444 17118 24500
rect 17826 24444 17836 24500
rect 17892 24444 19740 24500
rect 19796 24444 19806 24500
rect 20972 24444 24948 24500
rect 26646 24444 26684 24500
rect 26740 24444 26750 24500
rect 26852 24444 27916 24500
rect 27972 24444 27982 24500
rect 28130 24444 28140 24500
rect 28196 24444 38220 24500
rect 38276 24444 38286 24500
rect 41122 24444 41132 24500
rect 41188 24444 41692 24500
rect 41748 24444 41758 24500
rect 41916 24444 44884 24500
rect 45378 24444 45388 24500
rect 45444 24444 45836 24500
rect 45892 24444 45902 24500
rect 46834 24444 46844 24500
rect 46900 24444 46956 24500
rect 47012 24444 47022 24500
rect 47628 24444 49644 24500
rect 49700 24444 49710 24500
rect 55010 24444 55020 24500
rect 55076 24444 55468 24500
rect 55524 24444 55534 24500
rect 56466 24444 56476 24500
rect 56532 24444 57456 24500
rect 0 24416 112 24444
rect 15092 24388 15148 24444
rect 24892 24388 24948 24444
rect 26852 24388 26908 24444
rect 1810 24332 1820 24388
rect 1876 24332 1932 24388
rect 1988 24332 1998 24388
rect 4834 24332 4844 24388
rect 4900 24332 5068 24388
rect 5124 24332 5134 24388
rect 5282 24332 5292 24388
rect 5348 24332 7980 24388
rect 8036 24332 8046 24388
rect 8194 24332 8204 24388
rect 8260 24332 13132 24388
rect 13188 24332 13198 24388
rect 14242 24332 14252 24388
rect 14308 24332 14588 24388
rect 14644 24332 14654 24388
rect 15092 24332 17612 24388
rect 17668 24332 17678 24388
rect 19282 24332 19292 24388
rect 19348 24332 21196 24388
rect 21252 24332 21262 24388
rect 21634 24332 21644 24388
rect 21700 24332 21868 24388
rect 21924 24332 21934 24388
rect 22082 24332 22092 24388
rect 22148 24332 23100 24388
rect 23156 24332 23166 24388
rect 24892 24332 26908 24388
rect 27458 24332 27468 24388
rect 27524 24332 27692 24388
rect 27748 24332 27758 24388
rect 27906 24332 27916 24388
rect 27972 24332 28476 24388
rect 28532 24332 28542 24388
rect 29026 24332 29036 24388
rect 29092 24332 29484 24388
rect 29540 24332 32116 24388
rect 32498 24332 32508 24388
rect 32564 24332 33292 24388
rect 33348 24332 33358 24388
rect 34402 24332 34412 24388
rect 34468 24332 34636 24388
rect 34692 24332 34702 24388
rect 35252 24332 37660 24388
rect 37716 24332 37726 24388
rect 37986 24332 37996 24388
rect 38052 24332 43596 24388
rect 43652 24332 43662 24388
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 32060 24276 32116 24332
rect 35252 24276 35308 24332
rect 44454 24276 44464 24332
rect 44520 24276 44568 24332
rect 44624 24276 44672 24332
rect 44728 24276 44738 24332
rect 44828 24276 44884 24444
rect 57344 24416 57456 24444
rect 45714 24332 45724 24388
rect 45780 24332 46396 24388
rect 46452 24332 46462 24388
rect 49298 24332 49308 24388
rect 49364 24332 51324 24388
rect 51380 24332 52556 24388
rect 52612 24332 52622 24388
rect 53330 24332 53340 24388
rect 53396 24332 53452 24388
rect 53508 24332 53518 24388
rect 56364 24332 57148 24388
rect 57204 24332 57214 24388
rect 3378 24220 3388 24276
rect 3444 24220 3948 24276
rect 4004 24220 4014 24276
rect 4946 24220 4956 24276
rect 5012 24220 9772 24276
rect 9828 24220 9838 24276
rect 12674 24220 12684 24276
rect 12740 24220 20076 24276
rect 20132 24220 20142 24276
rect 21298 24220 21308 24276
rect 21364 24220 22428 24276
rect 22484 24220 22494 24276
rect 23538 24220 23548 24276
rect 23604 24220 24220 24276
rect 24276 24220 24286 24276
rect 26450 24220 26460 24276
rect 26516 24220 28700 24276
rect 28756 24220 28766 24276
rect 29810 24220 29820 24276
rect 29876 24220 31724 24276
rect 31780 24220 31790 24276
rect 32060 24220 35308 24276
rect 36194 24220 36204 24276
rect 36260 24220 39228 24276
rect 39284 24220 39294 24276
rect 39638 24220 39676 24276
rect 39732 24220 39742 24276
rect 40226 24220 40236 24276
rect 40292 24220 41468 24276
rect 41524 24220 41534 24276
rect 41682 24220 41692 24276
rect 41748 24220 44156 24276
rect 44212 24220 44222 24276
rect 44828 24220 56140 24276
rect 56196 24220 56206 24276
rect 56364 24164 56420 24332
rect 2594 24108 2604 24164
rect 2660 24108 3724 24164
rect 3780 24108 3790 24164
rect 5058 24108 5068 24164
rect 5124 24108 5180 24164
rect 5236 24108 5246 24164
rect 5394 24108 5404 24164
rect 5460 24108 6076 24164
rect 6132 24108 6142 24164
rect 6514 24108 6524 24164
rect 6580 24108 8988 24164
rect 9044 24108 9054 24164
rect 9212 24108 21700 24164
rect 0 24052 112 24080
rect 9212 24052 9268 24108
rect 21644 24052 21700 24108
rect 22092 24108 28476 24164
rect 28532 24108 28542 24164
rect 32386 24108 32396 24164
rect 32452 24108 32844 24164
rect 32900 24108 32910 24164
rect 33590 24108 33628 24164
rect 33684 24108 36988 24164
rect 37044 24108 37996 24164
rect 38052 24108 38062 24164
rect 38210 24108 38220 24164
rect 38276 24108 39004 24164
rect 39060 24108 39070 24164
rect 41010 24108 41020 24164
rect 41076 24108 41916 24164
rect 41972 24108 41982 24164
rect 44258 24108 44268 24164
rect 44324 24108 56420 24164
rect 22092 24052 22148 24108
rect 57344 24052 57456 24080
rect 0 23996 9268 24052
rect 9986 23996 9996 24052
rect 10052 23996 11676 24052
rect 11732 23996 11742 24052
rect 15092 23996 18508 24052
rect 18564 23996 18574 24052
rect 20850 23996 20860 24052
rect 20916 23996 21420 24052
rect 21476 23996 21486 24052
rect 21644 23996 22148 24052
rect 24546 23996 24556 24052
rect 24612 23996 30044 24052
rect 30100 23996 30110 24052
rect 31154 23996 31164 24052
rect 31220 23996 31500 24052
rect 31556 23996 31566 24052
rect 33058 23996 33068 24052
rect 33124 23996 35644 24052
rect 35700 23996 41804 24052
rect 41860 23996 41870 24052
rect 43138 23996 43148 24052
rect 43204 23996 44380 24052
rect 44436 23996 47852 24052
rect 47908 23996 47918 24052
rect 48850 23996 48860 24052
rect 48916 23996 52108 24052
rect 52164 23996 52174 24052
rect 52994 23996 53004 24052
rect 53060 23996 53228 24052
rect 53284 23996 53294 24052
rect 56802 23996 56812 24052
rect 56868 23996 57456 24052
rect 0 23968 112 23996
rect 15092 23940 15148 23996
rect 57344 23968 57456 23996
rect 3378 23884 3388 23940
rect 3444 23884 3836 23940
rect 3892 23884 3902 23940
rect 5590 23884 5628 23940
rect 5684 23884 5694 23940
rect 6962 23884 6972 23940
rect 7028 23884 7420 23940
rect 7476 23884 7486 23940
rect 7858 23884 7868 23940
rect 7924 23884 9324 23940
rect 9380 23884 9390 23940
rect 11106 23884 11116 23940
rect 11172 23884 12684 23940
rect 12740 23884 14700 23940
rect 14756 23884 15148 23940
rect 17266 23884 17276 23940
rect 17332 23884 17500 23940
rect 17556 23884 17612 23940
rect 17668 23884 17678 23940
rect 18172 23884 19180 23940
rect 19236 23884 19246 23940
rect 19730 23884 19740 23940
rect 19796 23884 22316 23940
rect 22372 23884 22382 23940
rect 23874 23884 23884 23940
rect 23940 23884 25900 23940
rect 25956 23884 25966 23940
rect 26310 23884 26348 23940
rect 26404 23884 26414 23940
rect 27682 23884 27692 23940
rect 27748 23884 27916 23940
rect 27972 23884 27982 23940
rect 28690 23884 28700 23940
rect 28756 23884 29036 23940
rect 29092 23884 29102 23940
rect 30258 23884 30268 23940
rect 30324 23884 33852 23940
rect 33908 23884 33918 23940
rect 34290 23884 34300 23940
rect 34356 23884 37268 23940
rect 37426 23884 37436 23940
rect 37492 23884 38724 23940
rect 39330 23884 39340 23940
rect 39396 23884 40012 23940
rect 40068 23884 40078 23940
rect 41458 23884 41468 23940
rect 41524 23884 41692 23940
rect 41748 23884 41758 23940
rect 42018 23884 42028 23940
rect 42084 23884 46508 23940
rect 46564 23884 46574 23940
rect 53218 23884 53228 23940
rect 53284 23884 54012 23940
rect 54068 23884 54078 23940
rect 56578 23884 56588 23940
rect 56644 23884 56812 23940
rect 56868 23884 56878 23940
rect 18172 23828 18228 23884
rect 1698 23772 1708 23828
rect 1764 23772 5068 23828
rect 5124 23772 5292 23828
rect 5348 23772 5358 23828
rect 5954 23772 5964 23828
rect 6020 23772 10444 23828
rect 10500 23772 10510 23828
rect 12226 23772 12236 23828
rect 12292 23772 13468 23828
rect 13524 23772 13534 23828
rect 13682 23772 13692 23828
rect 13748 23772 18228 23828
rect 18722 23772 18732 23828
rect 18788 23772 20636 23828
rect 20692 23772 20702 23828
rect 20962 23772 20972 23828
rect 21028 23772 21084 23828
rect 21140 23772 21150 23828
rect 21298 23772 21308 23828
rect 21364 23772 21868 23828
rect 21924 23772 21934 23828
rect 22204 23772 24556 23828
rect 24612 23772 24622 23828
rect 25218 23772 25228 23828
rect 25284 23772 36428 23828
rect 36484 23772 36494 23828
rect 36642 23772 36652 23828
rect 36708 23772 36988 23828
rect 37044 23772 37054 23828
rect 22204 23716 22260 23772
rect 1586 23660 1596 23716
rect 1652 23660 2380 23716
rect 2436 23660 2446 23716
rect 3332 23660 4228 23716
rect 6738 23660 6748 23716
rect 6804 23660 7308 23716
rect 7364 23660 7868 23716
rect 7924 23660 7934 23716
rect 9090 23660 9100 23716
rect 9156 23660 9324 23716
rect 9380 23660 9390 23716
rect 9986 23660 9996 23716
rect 10052 23660 12572 23716
rect 12628 23660 12638 23716
rect 15922 23660 15932 23716
rect 15988 23660 17276 23716
rect 17332 23660 18172 23716
rect 18228 23660 18238 23716
rect 20402 23660 20412 23716
rect 20468 23660 21196 23716
rect 21252 23660 21262 23716
rect 21494 23660 21532 23716
rect 21588 23660 21598 23716
rect 21858 23660 21868 23716
rect 21924 23660 22260 23716
rect 22978 23660 22988 23716
rect 23044 23660 25676 23716
rect 25732 23660 25844 23716
rect 27682 23660 27692 23716
rect 27748 23660 31612 23716
rect 31668 23660 34860 23716
rect 34916 23660 34926 23716
rect 0 23604 112 23632
rect 3332 23604 3388 23660
rect 4172 23604 4228 23660
rect 25788 23604 25844 23660
rect 36428 23604 36484 23772
rect 37212 23716 37268 23884
rect 38668 23828 38724 23884
rect 37650 23772 37660 23828
rect 37716 23772 38444 23828
rect 38500 23772 38510 23828
rect 38668 23772 49868 23828
rect 49924 23772 49934 23828
rect 51538 23772 51548 23828
rect 51604 23772 54236 23828
rect 54292 23772 54302 23828
rect 56690 23772 56700 23828
rect 56756 23772 57260 23828
rect 57316 23772 57326 23828
rect 36754 23660 36764 23716
rect 36820 23660 37268 23716
rect 39554 23660 39564 23716
rect 39620 23660 44212 23716
rect 46498 23660 46508 23716
rect 46564 23660 48300 23716
rect 48356 23660 48366 23716
rect 56242 23660 56252 23716
rect 56308 23660 56812 23716
rect 56868 23660 56878 23716
rect 44156 23604 44212 23660
rect 57344 23604 57456 23632
rect 0 23548 3388 23604
rect 3602 23548 3612 23604
rect 3668 23548 3678 23604
rect 4172 23548 6692 23604
rect 6850 23548 6860 23604
rect 6916 23548 7756 23604
rect 7812 23548 9548 23604
rect 9604 23548 9614 23604
rect 11788 23548 17948 23604
rect 18004 23548 18014 23604
rect 22754 23548 22764 23604
rect 22820 23548 23100 23604
rect 23156 23548 23166 23604
rect 25526 23548 25564 23604
rect 25620 23548 25630 23604
rect 25788 23548 29036 23604
rect 29092 23548 29102 23604
rect 29250 23548 29260 23604
rect 29316 23548 30156 23604
rect 30212 23548 30222 23604
rect 31042 23548 31052 23604
rect 31108 23548 32564 23604
rect 0 23520 112 23548
rect 3612 23492 3668 23548
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 6636 23492 6692 23548
rect 11788 23492 11844 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 32508 23492 32564 23548
rect 32732 23548 33404 23604
rect 33460 23548 33470 23604
rect 33842 23548 33852 23604
rect 33908 23548 34636 23604
rect 34692 23548 34702 23604
rect 36428 23548 40796 23604
rect 40852 23548 41020 23604
rect 41076 23548 41086 23604
rect 41346 23548 41356 23604
rect 41412 23548 43484 23604
rect 43540 23548 43550 23604
rect 44156 23548 46844 23604
rect 46900 23548 46910 23604
rect 47058 23548 47068 23604
rect 47124 23548 55468 23604
rect 56354 23548 56364 23604
rect 56420 23548 57456 23604
rect 32732 23492 32788 23548
rect 43794 23492 43804 23548
rect 43860 23492 43908 23548
rect 43964 23492 44012 23548
rect 44068 23492 44078 23548
rect 55412 23492 55468 23548
rect 57344 23520 57456 23548
rect 3266 23436 3276 23492
rect 3332 23436 3668 23492
rect 4274 23436 4284 23492
rect 4340 23436 4732 23492
rect 4788 23436 4798 23492
rect 6636 23436 9212 23492
rect 9268 23436 9278 23492
rect 9762 23436 9772 23492
rect 9828 23436 11844 23492
rect 12562 23436 12572 23492
rect 12628 23436 13804 23492
rect 13860 23436 13870 23492
rect 14130 23436 14140 23492
rect 14196 23436 14476 23492
rect 14532 23436 15372 23492
rect 15428 23436 16884 23492
rect 17042 23436 17052 23492
rect 17108 23436 17276 23492
rect 17332 23436 17342 23492
rect 18050 23436 18060 23492
rect 18116 23436 18732 23492
rect 18788 23436 18798 23492
rect 21298 23436 21308 23492
rect 21364 23436 21588 23492
rect 22082 23436 22092 23492
rect 22148 23436 23436 23492
rect 23492 23436 23502 23492
rect 24210 23436 24220 23492
rect 24276 23436 25452 23492
rect 25508 23436 25518 23492
rect 26674 23436 26684 23492
rect 26740 23436 26908 23492
rect 26964 23436 32060 23492
rect 32116 23436 32172 23492
rect 32228 23436 32238 23492
rect 32498 23436 32508 23492
rect 32564 23436 32574 23492
rect 32722 23436 32732 23492
rect 32788 23436 32798 23492
rect 32946 23436 32956 23492
rect 33012 23436 34076 23492
rect 34132 23436 34142 23492
rect 35410 23436 35420 23492
rect 35476 23436 36988 23492
rect 37044 23436 37054 23492
rect 37202 23436 37212 23492
rect 37268 23436 37306 23492
rect 38546 23436 38556 23492
rect 38612 23436 39116 23492
rect 39172 23436 39182 23492
rect 39890 23436 39900 23492
rect 39956 23436 40236 23492
rect 40292 23436 40302 23492
rect 40684 23436 41580 23492
rect 41636 23436 41646 23492
rect 41906 23436 41916 23492
rect 41972 23436 42700 23492
rect 42756 23436 42766 23492
rect 44146 23436 44156 23492
rect 44212 23436 49812 23492
rect 55412 23436 55916 23492
rect 55972 23436 55982 23492
rect 3602 23324 3612 23380
rect 3668 23324 13692 23380
rect 13748 23324 13758 23380
rect 16828 23268 16884 23436
rect 21532 23380 21588 23436
rect 40684 23380 40740 23436
rect 17826 23324 17836 23380
rect 17892 23324 19404 23380
rect 19460 23324 19470 23380
rect 19730 23324 19740 23380
rect 19796 23324 21252 23380
rect 21532 23324 21868 23380
rect 21924 23324 21934 23380
rect 22306 23324 22316 23380
rect 22372 23324 22428 23380
rect 22484 23324 22494 23380
rect 23090 23324 23100 23380
rect 23156 23324 25116 23380
rect 25172 23324 25182 23380
rect 25340 23324 39676 23380
rect 39732 23324 39742 23380
rect 40012 23324 40740 23380
rect 49756 23380 49812 23436
rect 49756 23324 54796 23380
rect 54852 23324 54862 23380
rect 21196 23268 21252 23324
rect 914 23212 924 23268
rect 980 23212 3108 23268
rect 4050 23212 4060 23268
rect 4116 23212 6412 23268
rect 6468 23212 6478 23268
rect 6962 23212 6972 23268
rect 7028 23212 9996 23268
rect 10052 23212 10062 23268
rect 10994 23212 11004 23268
rect 11060 23212 12012 23268
rect 12068 23212 12078 23268
rect 13794 23212 13804 23268
rect 13860 23212 14476 23268
rect 14532 23212 14542 23268
rect 15026 23212 15036 23268
rect 15092 23212 16772 23268
rect 16828 23212 20972 23268
rect 21028 23212 21038 23268
rect 21196 23212 21868 23268
rect 21924 23212 21934 23268
rect 23314 23212 23324 23268
rect 23380 23212 25004 23268
rect 25060 23212 25070 23268
rect 0 23156 112 23184
rect 0 23100 2828 23156
rect 2884 23100 2894 23156
rect 0 23072 112 23100
rect 3052 23044 3108 23212
rect 4834 23100 4844 23156
rect 4900 23100 4956 23156
rect 5012 23100 5022 23156
rect 5170 23100 5180 23156
rect 5236 23100 6524 23156
rect 6580 23100 6590 23156
rect 7186 23100 7196 23156
rect 7252 23100 7420 23156
rect 7476 23100 7486 23156
rect 7970 23100 7980 23156
rect 8036 23100 8876 23156
rect 8932 23100 8942 23156
rect 9762 23100 9772 23156
rect 9828 23100 10780 23156
rect 10836 23100 10846 23156
rect 15148 23100 16492 23156
rect 16548 23100 16558 23156
rect 15148 23044 15204 23100
rect 16716 23044 16772 23212
rect 25340 23156 25396 23324
rect 40012 23268 40068 23324
rect 26114 23212 26124 23268
rect 26180 23212 28700 23268
rect 28756 23212 30268 23268
rect 30324 23212 30334 23268
rect 31378 23212 31388 23268
rect 31444 23212 33852 23268
rect 33908 23212 33918 23268
rect 34178 23212 34188 23268
rect 34244 23212 34524 23268
rect 34580 23212 34590 23268
rect 36306 23212 36316 23268
rect 36372 23212 36876 23268
rect 36932 23212 36942 23268
rect 37090 23212 37100 23268
rect 37156 23212 38444 23268
rect 38500 23212 40068 23268
rect 42466 23212 42476 23268
rect 42532 23212 44156 23268
rect 44212 23212 44222 23268
rect 45154 23212 45164 23268
rect 45220 23212 48748 23268
rect 48804 23212 48814 23268
rect 49634 23212 49644 23268
rect 49700 23212 50428 23268
rect 50484 23212 50764 23268
rect 50820 23212 52220 23268
rect 52276 23212 52892 23268
rect 52948 23212 53564 23268
rect 53620 23212 53630 23268
rect 53778 23212 53788 23268
rect 53844 23212 54460 23268
rect 54516 23212 54526 23268
rect 56242 23212 56252 23268
rect 56308 23212 56812 23268
rect 56868 23212 56878 23268
rect 57344 23156 57456 23184
rect 16930 23100 16940 23156
rect 16996 23100 18060 23156
rect 18116 23100 18126 23156
rect 18834 23100 18844 23156
rect 18900 23100 18956 23156
rect 19012 23100 19022 23156
rect 19394 23100 19404 23156
rect 19460 23100 19740 23156
rect 19796 23100 19806 23156
rect 20290 23100 20300 23156
rect 20356 23100 20524 23156
rect 20580 23100 20590 23156
rect 20738 23100 20748 23156
rect 20804 23100 20842 23156
rect 22530 23100 22540 23156
rect 22596 23100 22876 23156
rect 22932 23100 22942 23156
rect 23090 23100 23100 23156
rect 23156 23100 23884 23156
rect 23940 23100 23950 23156
rect 24210 23100 24220 23156
rect 24276 23100 25396 23156
rect 28578 23100 28588 23156
rect 28644 23100 29484 23156
rect 29540 23100 29550 23156
rect 30594 23100 30604 23156
rect 30660 23100 32620 23156
rect 32676 23100 32686 23156
rect 33282 23100 33292 23156
rect 33348 23100 34468 23156
rect 35298 23100 35308 23156
rect 35364 23100 36652 23156
rect 36708 23100 37212 23156
rect 37268 23100 37278 23156
rect 39666 23100 39676 23156
rect 39732 23100 40236 23156
rect 40292 23100 40572 23156
rect 40628 23100 40638 23156
rect 41570 23100 41580 23156
rect 41636 23100 41916 23156
rect 41972 23100 41982 23156
rect 43586 23100 43596 23156
rect 43652 23100 45052 23156
rect 45108 23100 45118 23156
rect 45724 23100 46060 23156
rect 46116 23100 46126 23156
rect 46470 23100 46508 23156
rect 46564 23100 46574 23156
rect 47814 23100 47852 23156
rect 47908 23100 47918 23156
rect 48962 23100 48972 23156
rect 49028 23100 57456 23156
rect 34412 23044 34468 23100
rect 45724 23044 45780 23100
rect 57344 23072 57456 23100
rect 3052 22988 6524 23044
rect 6580 22988 6590 23044
rect 8530 22988 8540 23044
rect 8596 22988 9884 23044
rect 9940 22988 9950 23044
rect 11218 22988 11228 23044
rect 11284 22988 11564 23044
rect 11620 22988 15148 23044
rect 15204 22988 15214 23044
rect 15474 22988 15484 23044
rect 15540 22988 16492 23044
rect 16548 22988 16558 23044
rect 16716 22988 18732 23044
rect 18788 22988 21812 23044
rect 23538 22988 23548 23044
rect 23604 22988 24892 23044
rect 24948 22988 25508 23044
rect 26674 22988 26684 23044
rect 26740 22988 30268 23044
rect 30324 22988 30334 23044
rect 31126 22988 31164 23044
rect 31220 22988 31230 23044
rect 32274 22988 32284 23044
rect 32340 22988 33068 23044
rect 33124 22988 33134 23044
rect 33282 22988 33292 23044
rect 33348 22988 34356 23044
rect 34412 22988 41580 23044
rect 41636 22988 42924 23044
rect 42980 22988 42990 23044
rect 44146 22988 44156 23044
rect 44212 22988 45780 23044
rect 45938 22988 45948 23044
rect 46004 22988 48748 23044
rect 48804 22988 48814 23044
rect 49074 22988 49084 23044
rect 49140 22988 50428 23044
rect 50866 22988 50876 23044
rect 50932 22988 52332 23044
rect 52388 22988 52398 23044
rect 52630 22988 52668 23044
rect 52724 22988 52734 23044
rect 21756 22932 21812 22988
rect 25452 22932 25508 22988
rect 34300 22932 34356 22988
rect 50372 22932 50428 22988
rect 578 22876 588 22932
rect 644 22876 3388 22932
rect 3444 22876 3454 22932
rect 4162 22876 4172 22932
rect 4228 22876 8092 22932
rect 8148 22876 8158 22932
rect 8530 22876 8540 22932
rect 8596 22876 15148 22932
rect 15250 22876 15260 22932
rect 15316 22876 17052 22932
rect 17108 22876 19292 22932
rect 19348 22876 19358 22932
rect 19730 22876 19740 22932
rect 19796 22876 19964 22932
rect 20020 22876 20030 22932
rect 20738 22876 20748 22932
rect 20804 22876 21532 22932
rect 21588 22876 21598 22932
rect 21756 22876 21924 22932
rect 22530 22876 22540 22932
rect 22596 22876 24220 22932
rect 24276 22876 24286 22932
rect 24770 22876 24780 22932
rect 24836 22876 25228 22932
rect 25284 22876 25294 22932
rect 25452 22876 33404 22932
rect 33460 22876 33470 22932
rect 34290 22876 34300 22932
rect 34356 22876 35308 22932
rect 35364 22876 35374 22932
rect 36418 22876 36428 22932
rect 36484 22876 36540 22932
rect 36596 22876 36606 22932
rect 36978 22876 36988 22932
rect 37044 22876 38892 22932
rect 38948 22876 38958 22932
rect 39218 22876 39228 22932
rect 39284 22876 47180 22932
rect 47236 22876 47246 22932
rect 49970 22876 49980 22932
rect 50036 22876 50092 22932
rect 50148 22876 50158 22932
rect 50372 22876 51100 22932
rect 51156 22876 51166 22932
rect 53106 22876 53116 22932
rect 53172 22876 54908 22932
rect 54964 22876 54974 22932
rect 15092 22820 15148 22876
rect 21868 22820 21924 22876
rect 7186 22764 7196 22820
rect 7252 22764 14980 22820
rect 15092 22764 19740 22820
rect 19796 22764 19806 22820
rect 21868 22764 22316 22820
rect 22372 22764 22382 22820
rect 26348 22764 29036 22820
rect 29092 22764 29708 22820
rect 29764 22764 30828 22820
rect 30884 22764 30894 22820
rect 31042 22764 31052 22820
rect 31108 22764 34188 22820
rect 34244 22764 34254 22820
rect 34626 22764 34636 22820
rect 34692 22764 34860 22820
rect 34916 22764 34926 22820
rect 35074 22764 35084 22820
rect 35140 22764 35196 22820
rect 35252 22764 43148 22820
rect 43204 22764 43214 22820
rect 44828 22764 47628 22820
rect 47684 22764 49700 22820
rect 50194 22764 50204 22820
rect 50260 22764 54684 22820
rect 54740 22764 54750 22820
rect 0 22708 112 22736
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 14924 22708 14980 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 26348 22708 26404 22764
rect 44454 22708 44464 22764
rect 44520 22708 44568 22764
rect 44624 22708 44672 22764
rect 44728 22708 44738 22764
rect 0 22652 2716 22708
rect 2772 22652 2782 22708
rect 4834 22652 4844 22708
rect 4900 22652 5068 22708
rect 5124 22652 8092 22708
rect 8148 22652 8158 22708
rect 9650 22652 9660 22708
rect 9716 22652 9772 22708
rect 9828 22652 9838 22708
rect 10210 22652 10220 22708
rect 10276 22652 10892 22708
rect 10948 22652 14140 22708
rect 14196 22652 14206 22708
rect 14924 22652 16156 22708
rect 16212 22652 16222 22708
rect 16482 22652 16492 22708
rect 16548 22652 16828 22708
rect 16884 22652 16894 22708
rect 17378 22652 17388 22708
rect 17444 22652 17612 22708
rect 17668 22652 17678 22708
rect 18050 22652 18060 22708
rect 18116 22652 18396 22708
rect 18452 22652 21308 22708
rect 21364 22652 21374 22708
rect 21522 22652 21532 22708
rect 21588 22652 22764 22708
rect 22820 22652 22830 22708
rect 25778 22652 25788 22708
rect 25844 22652 26404 22708
rect 27468 22652 36932 22708
rect 37090 22652 37100 22708
rect 37156 22652 39228 22708
rect 39284 22652 39294 22708
rect 40562 22652 40572 22708
rect 40628 22652 41580 22708
rect 41636 22652 41646 22708
rect 41906 22652 41916 22708
rect 41972 22652 44156 22708
rect 44212 22652 44222 22708
rect 0 22624 112 22652
rect 27468 22596 27524 22652
rect 36876 22596 36932 22652
rect 44828 22596 44884 22764
rect 49644 22708 49700 22764
rect 57344 22708 57456 22736
rect 46834 22652 46844 22708
rect 46900 22652 49588 22708
rect 49644 22652 51100 22708
rect 51156 22652 51166 22708
rect 57250 22652 57260 22708
rect 57316 22652 57456 22708
rect 49532 22596 49588 22652
rect 57344 22624 57456 22652
rect 2370 22540 2380 22596
rect 2436 22540 2492 22596
rect 2548 22540 2558 22596
rect 3378 22540 3388 22596
rect 3444 22540 4956 22596
rect 5012 22540 7532 22596
rect 7588 22540 7598 22596
rect 7746 22540 7756 22596
rect 7812 22540 11788 22596
rect 11844 22540 11854 22596
rect 12338 22540 12348 22596
rect 12404 22540 20972 22596
rect 21028 22540 24332 22596
rect 24388 22540 27524 22596
rect 27682 22540 27692 22596
rect 27748 22540 28812 22596
rect 28868 22540 28878 22596
rect 30258 22540 30268 22596
rect 30324 22540 32060 22596
rect 32116 22540 32284 22596
rect 32340 22540 32350 22596
rect 33282 22540 33292 22596
rect 33348 22540 36540 22596
rect 36596 22540 36606 22596
rect 36876 22540 37212 22596
rect 37268 22540 37278 22596
rect 40338 22540 40348 22596
rect 40404 22540 44156 22596
rect 44212 22540 44222 22596
rect 44370 22540 44380 22596
rect 44436 22540 44884 22596
rect 47394 22540 47404 22596
rect 47460 22540 47740 22596
rect 47796 22540 47806 22596
rect 48514 22540 48524 22596
rect 48580 22540 49308 22596
rect 49364 22540 49374 22596
rect 49532 22540 50876 22596
rect 50932 22540 50942 22596
rect 51762 22540 51772 22596
rect 51828 22540 54124 22596
rect 54180 22540 54190 22596
rect 2482 22428 2492 22484
rect 2548 22428 13804 22484
rect 13860 22428 13870 22484
rect 15250 22428 15260 22484
rect 15316 22428 17892 22484
rect 19282 22428 19292 22484
rect 19348 22428 19628 22484
rect 19684 22428 19694 22484
rect 20514 22428 20524 22484
rect 20580 22428 21980 22484
rect 22036 22428 26908 22484
rect 28102 22428 28140 22484
rect 28196 22428 28206 22484
rect 29138 22428 29148 22484
rect 29204 22428 30604 22484
rect 30660 22428 30670 22484
rect 30818 22428 30828 22484
rect 30884 22428 32172 22484
rect 32228 22428 32238 22484
rect 33394 22428 33404 22484
rect 33460 22428 40460 22484
rect 40516 22428 42028 22484
rect 42084 22428 42094 22484
rect 43474 22428 43484 22484
rect 43540 22428 45164 22484
rect 45220 22428 45230 22484
rect 46050 22428 46060 22484
rect 46116 22428 48188 22484
rect 48244 22428 48254 22484
rect 17836 22372 17892 22428
rect 26852 22372 26908 22428
rect 1922 22316 1932 22372
rect 1988 22316 3724 22372
rect 3780 22316 3790 22372
rect 3938 22316 3948 22372
rect 4004 22316 4014 22372
rect 4946 22316 4956 22372
rect 5012 22316 9660 22372
rect 9716 22316 9726 22372
rect 10434 22316 10444 22372
rect 10500 22316 11004 22372
rect 11060 22316 11070 22372
rect 11330 22316 11340 22372
rect 11396 22316 12124 22372
rect 12180 22316 12190 22372
rect 13682 22316 13692 22372
rect 13748 22316 14812 22372
rect 14868 22316 15372 22372
rect 15428 22316 15708 22372
rect 15764 22316 15774 22372
rect 16930 22316 16940 22372
rect 16996 22316 17276 22372
rect 17332 22316 17342 22372
rect 17836 22316 19348 22372
rect 19506 22316 19516 22372
rect 19572 22316 21420 22372
rect 21476 22316 21486 22372
rect 22950 22316 22988 22372
rect 23044 22316 23054 22372
rect 26002 22316 26012 22372
rect 26068 22316 26124 22372
rect 26180 22316 26190 22372
rect 26852 22316 30268 22372
rect 30324 22316 30334 22372
rect 30930 22316 30940 22372
rect 30996 22316 31164 22372
rect 31220 22316 31230 22372
rect 33842 22316 33852 22372
rect 33908 22316 34188 22372
rect 34244 22316 34254 22372
rect 34514 22316 34524 22372
rect 34580 22316 34860 22372
rect 34916 22316 34926 22372
rect 37538 22316 37548 22372
rect 37604 22316 42588 22372
rect 42644 22316 42654 22372
rect 42812 22316 45500 22372
rect 45556 22316 45566 22372
rect 47842 22316 47852 22372
rect 47908 22316 48412 22372
rect 48468 22316 48478 22372
rect 49074 22316 49084 22372
rect 49140 22316 49644 22372
rect 49700 22316 50988 22372
rect 51044 22316 51054 22372
rect 0 22260 112 22288
rect 3948 22260 4004 22316
rect 19292 22260 19348 22316
rect 42812 22260 42868 22316
rect 57344 22260 57456 22288
rect 0 22204 700 22260
rect 756 22204 766 22260
rect 2370 22204 2380 22260
rect 2436 22204 2716 22260
rect 2772 22204 2782 22260
rect 3948 22204 16268 22260
rect 16324 22204 16334 22260
rect 17938 22204 17948 22260
rect 18004 22204 18396 22260
rect 18452 22204 18462 22260
rect 19292 22204 20748 22260
rect 20804 22204 20814 22260
rect 21084 22204 42868 22260
rect 43026 22204 43036 22260
rect 43092 22204 50428 22260
rect 50530 22204 50540 22260
rect 50596 22204 57456 22260
rect 0 22176 112 22204
rect 21084 22148 21140 22204
rect 2818 22092 2828 22148
rect 2884 22092 5404 22148
rect 5460 22092 5470 22148
rect 7634 22092 7644 22148
rect 7700 22092 9548 22148
rect 9604 22092 9614 22148
rect 9874 22092 9884 22148
rect 9940 22092 12348 22148
rect 12404 22092 12414 22148
rect 12786 22092 12796 22148
rect 12852 22092 21140 22148
rect 21522 22092 21532 22148
rect 21588 22092 22540 22148
rect 22596 22092 22606 22148
rect 23660 22092 33292 22148
rect 33348 22092 33358 22148
rect 33618 22092 33628 22148
rect 33684 22092 33964 22148
rect 34020 22092 37436 22148
rect 37492 22092 37502 22148
rect 38612 22092 45892 22148
rect 46050 22092 46060 22148
rect 46116 22092 49644 22148
rect 49700 22092 49710 22148
rect 7074 21980 7084 22036
rect 7140 21980 9436 22036
rect 9492 21980 9502 22036
rect 9986 21980 9996 22036
rect 10052 21980 10556 22036
rect 10612 21980 10622 22036
rect 13794 21980 13804 22036
rect 13860 21980 23436 22036
rect 23492 21980 23502 22036
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 23660 21924 23716 22092
rect 38612 22036 38668 22092
rect 24546 21980 24556 22036
rect 24612 21980 26796 22036
rect 26852 21980 26862 22036
rect 30146 21980 30156 22036
rect 30212 21980 30940 22036
rect 30996 21980 31006 22036
rect 32498 21980 32508 22036
rect 32564 21980 38668 22036
rect 45836 22036 45892 22092
rect 50372 22036 50428 22204
rect 57344 22176 57456 22204
rect 52994 22092 53004 22148
rect 53060 22092 54012 22148
rect 54068 22092 54078 22148
rect 55234 22092 55244 22148
rect 55300 22092 56028 22148
rect 56084 22092 56094 22148
rect 45836 21980 46396 22036
rect 46452 21980 46462 22036
rect 46722 21980 46732 22036
rect 46788 21980 47404 22036
rect 47460 21980 47470 22036
rect 50372 21980 55356 22036
rect 55412 21980 55422 22036
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 43794 21924 43804 21980
rect 43860 21924 43908 21980
rect 43964 21924 44012 21980
rect 44068 21924 44078 21980
rect 1596 21868 3388 21924
rect 3444 21868 3454 21924
rect 5058 21868 5068 21924
rect 5124 21868 7812 21924
rect 8306 21868 8316 21924
rect 8372 21868 12236 21924
rect 12292 21868 12302 21924
rect 12450 21868 12460 21924
rect 12516 21868 23716 21924
rect 26236 21868 27020 21924
rect 27076 21868 27086 21924
rect 27794 21868 27804 21924
rect 27860 21868 30212 21924
rect 34290 21868 34300 21924
rect 34356 21868 34748 21924
rect 34804 21868 35420 21924
rect 35476 21868 35486 21924
rect 38210 21868 38220 21924
rect 38276 21868 38444 21924
rect 38500 21868 38510 21924
rect 38658 21868 38668 21924
rect 38724 21868 39340 21924
rect 39396 21868 39406 21924
rect 39554 21868 39564 21924
rect 39620 21868 40012 21924
rect 40068 21868 40078 21924
rect 40422 21868 40460 21924
rect 40516 21868 40526 21924
rect 40786 21868 40796 21924
rect 40852 21868 42140 21924
rect 42196 21868 42206 21924
rect 43026 21868 43036 21924
rect 43092 21868 43484 21924
rect 43540 21868 43550 21924
rect 45938 21868 45948 21924
rect 46004 21868 51212 21924
rect 51268 21868 51278 21924
rect 55654 21868 55692 21924
rect 55748 21868 55758 21924
rect 0 21812 112 21840
rect 1596 21812 1652 21868
rect 7756 21812 7812 21868
rect 0 21756 1652 21812
rect 1708 21756 4172 21812
rect 4228 21756 4238 21812
rect 5394 21756 5404 21812
rect 5460 21756 5470 21812
rect 7746 21756 7756 21812
rect 7812 21756 7822 21812
rect 8642 21756 8652 21812
rect 8708 21756 11116 21812
rect 11172 21756 11182 21812
rect 12114 21756 12124 21812
rect 12180 21756 13132 21812
rect 13188 21756 13198 21812
rect 13878 21756 13916 21812
rect 13972 21756 13982 21812
rect 14214 21756 14252 21812
rect 14308 21756 14318 21812
rect 15810 21756 15820 21812
rect 15876 21756 16156 21812
rect 16212 21756 17164 21812
rect 17220 21756 17230 21812
rect 17490 21756 17500 21812
rect 17556 21756 18508 21812
rect 18564 21756 18574 21812
rect 18722 21756 18732 21812
rect 18788 21756 21532 21812
rect 21588 21756 22204 21812
rect 22260 21756 22270 21812
rect 22418 21756 22428 21812
rect 22484 21756 25452 21812
rect 25508 21756 25518 21812
rect 0 21728 112 21756
rect 1708 21700 1764 21756
rect 5404 21700 5460 21756
rect 26236 21700 26292 21868
rect 30156 21812 30212 21868
rect 57344 21812 57456 21840
rect 26450 21756 26460 21812
rect 26516 21756 29148 21812
rect 29204 21756 29214 21812
rect 30156 21756 33964 21812
rect 34020 21756 34030 21812
rect 34188 21756 35532 21812
rect 35588 21756 35598 21812
rect 36754 21756 36764 21812
rect 36820 21756 37772 21812
rect 37828 21756 37838 21812
rect 38668 21756 40572 21812
rect 40628 21756 40638 21812
rect 41346 21756 41356 21812
rect 41412 21756 41916 21812
rect 41972 21756 42140 21812
rect 42196 21756 42206 21812
rect 42354 21756 42364 21812
rect 42420 21756 42700 21812
rect 42756 21756 42766 21812
rect 43362 21756 43372 21812
rect 43428 21756 44380 21812
rect 44436 21756 44446 21812
rect 44818 21756 44828 21812
rect 44884 21756 45948 21812
rect 46004 21756 46014 21812
rect 46620 21756 46956 21812
rect 47012 21756 47068 21812
rect 47124 21756 48860 21812
rect 48916 21756 48926 21812
rect 51874 21756 51884 21812
rect 51940 21756 52668 21812
rect 52724 21756 52734 21812
rect 52882 21756 52892 21812
rect 52948 21756 53564 21812
rect 53620 21756 53630 21812
rect 54114 21756 54124 21812
rect 54180 21756 54236 21812
rect 54292 21756 54684 21812
rect 54740 21756 54750 21812
rect 55412 21756 57456 21812
rect 34188 21700 34244 21756
rect 38668 21700 38724 21756
rect 46620 21700 46676 21756
rect 55412 21700 55468 21756
rect 57344 21728 57456 21756
rect 1362 21644 1372 21700
rect 1428 21644 1764 21700
rect 2706 21644 2716 21700
rect 2772 21644 4116 21700
rect 4274 21644 4284 21700
rect 4340 21644 8204 21700
rect 8260 21644 8270 21700
rect 10546 21644 10556 21700
rect 10612 21644 12012 21700
rect 12068 21644 12078 21700
rect 13766 21644 13804 21700
rect 13860 21644 13870 21700
rect 16258 21644 16268 21700
rect 16324 21644 26292 21700
rect 26450 21644 26460 21700
rect 26516 21644 27804 21700
rect 27860 21644 27870 21700
rect 28242 21644 28252 21700
rect 28308 21644 28476 21700
rect 28532 21644 28542 21700
rect 31714 21644 31724 21700
rect 31780 21644 34244 21700
rect 35522 21644 35532 21700
rect 35588 21644 38724 21700
rect 38882 21644 38892 21700
rect 38948 21644 39620 21700
rect 40002 21644 40012 21700
rect 40068 21644 40348 21700
rect 40404 21644 40414 21700
rect 40898 21644 40908 21700
rect 40964 21644 41580 21700
rect 41636 21644 46676 21700
rect 46834 21644 46844 21700
rect 46900 21644 55468 21700
rect 55682 21644 55692 21700
rect 55748 21644 55758 21700
rect 4060 21588 4116 21644
rect 39564 21588 39620 21644
rect 55692 21588 55748 21644
rect 466 21532 476 21588
rect 532 21532 3500 21588
rect 3556 21532 3566 21588
rect 4060 21532 5180 21588
rect 5236 21532 5246 21588
rect 6178 21532 6188 21588
rect 6244 21532 7532 21588
rect 7588 21532 7598 21588
rect 8754 21532 8764 21588
rect 8820 21532 8876 21588
rect 8932 21532 8942 21588
rect 9538 21532 9548 21588
rect 9604 21532 9772 21588
rect 9828 21532 9838 21588
rect 10882 21532 10892 21588
rect 10948 21532 15148 21588
rect 15810 21532 15820 21588
rect 15876 21532 20804 21588
rect 20962 21532 20972 21588
rect 21028 21532 23100 21588
rect 23156 21532 23166 21588
rect 23324 21532 24556 21588
rect 24612 21532 24622 21588
rect 24770 21532 24780 21588
rect 24836 21532 28588 21588
rect 28644 21532 28812 21588
rect 28868 21532 28878 21588
rect 29036 21532 36204 21588
rect 36260 21532 36270 21588
rect 37762 21532 37772 21588
rect 37828 21532 39228 21588
rect 39284 21532 39294 21588
rect 39554 21532 39564 21588
rect 39620 21532 39630 21588
rect 40684 21532 46508 21588
rect 46564 21532 46574 21588
rect 46722 21532 46732 21588
rect 46788 21532 49308 21588
rect 49364 21532 49374 21588
rect 49858 21532 49868 21588
rect 49924 21532 53788 21588
rect 53844 21532 53854 21588
rect 54002 21532 54012 21588
rect 54068 21532 55748 21588
rect 15092 21476 15148 21532
rect 20748 21476 20804 21532
rect 23324 21476 23380 21532
rect 29036 21476 29092 21532
rect 40684 21476 40740 21532
rect 1362 21420 1372 21476
rect 1428 21420 1708 21476
rect 1764 21420 1774 21476
rect 5842 21420 5852 21476
rect 5908 21420 6748 21476
rect 6804 21420 7644 21476
rect 7700 21420 7710 21476
rect 7858 21420 7868 21476
rect 7924 21420 10332 21476
rect 10388 21420 10398 21476
rect 11890 21420 11900 21476
rect 11956 21420 14924 21476
rect 14980 21420 14990 21476
rect 15092 21420 18060 21476
rect 18116 21420 18126 21476
rect 19618 21420 19628 21476
rect 19684 21420 20412 21476
rect 20468 21420 20478 21476
rect 20748 21420 23380 21476
rect 23510 21420 23548 21476
rect 23604 21420 23614 21476
rect 23884 21420 24500 21476
rect 24882 21420 24892 21476
rect 24948 21420 25340 21476
rect 25396 21420 25406 21476
rect 26114 21420 26124 21476
rect 26180 21420 26908 21476
rect 26964 21420 26974 21476
rect 27682 21420 27692 21476
rect 27748 21420 29092 21476
rect 30258 21420 30268 21476
rect 30324 21420 40740 21476
rect 40898 21420 40908 21476
rect 40964 21420 41132 21476
rect 41188 21420 41198 21476
rect 41346 21420 41356 21476
rect 41412 21420 41580 21476
rect 41636 21420 41646 21476
rect 43138 21420 43148 21476
rect 43204 21420 47516 21476
rect 47572 21420 47582 21476
rect 47730 21420 47740 21476
rect 47796 21420 47964 21476
rect 48020 21420 48030 21476
rect 48626 21420 48636 21476
rect 48692 21420 48748 21476
rect 48804 21420 50428 21476
rect 50754 21420 50764 21476
rect 50820 21420 56420 21476
rect 0 21364 112 21392
rect 23884 21364 23940 21420
rect 0 21308 1036 21364
rect 1092 21308 1102 21364
rect 1810 21308 1820 21364
rect 1876 21308 2268 21364
rect 2324 21308 6972 21364
rect 7028 21308 7038 21364
rect 7186 21308 7196 21364
rect 7252 21308 8092 21364
rect 8148 21308 8158 21364
rect 9202 21308 9212 21364
rect 9268 21308 17220 21364
rect 17378 21308 17388 21364
rect 17444 21308 17612 21364
rect 17668 21308 17678 21364
rect 17938 21308 17948 21364
rect 18004 21308 18620 21364
rect 18676 21308 18686 21364
rect 18834 21308 18844 21364
rect 18900 21308 21700 21364
rect 23090 21308 23100 21364
rect 23156 21308 23940 21364
rect 24444 21364 24500 21420
rect 50372 21364 50428 21420
rect 56364 21364 56420 21420
rect 57344 21364 57456 21392
rect 24444 21308 25060 21364
rect 25666 21308 25676 21364
rect 25732 21308 26348 21364
rect 26404 21308 26414 21364
rect 26572 21308 28252 21364
rect 28308 21308 28318 21364
rect 28578 21308 28588 21364
rect 28644 21308 29036 21364
rect 29092 21308 29102 21364
rect 30706 21308 30716 21364
rect 30772 21308 32396 21364
rect 32452 21308 32462 21364
rect 32610 21308 32620 21364
rect 32676 21308 44828 21364
rect 44884 21308 44894 21364
rect 46722 21308 46732 21364
rect 46788 21308 47628 21364
rect 47684 21308 47694 21364
rect 47842 21308 47852 21364
rect 47908 21308 48188 21364
rect 48244 21308 48254 21364
rect 50372 21308 52332 21364
rect 52388 21308 52398 21364
rect 52546 21308 52556 21364
rect 52612 21308 56028 21364
rect 56084 21308 56094 21364
rect 56364 21308 57456 21364
rect 0 21280 112 21308
rect 17164 21252 17220 21308
rect 21644 21252 21700 21308
rect 4844 21196 9828 21252
rect 10322 21196 10332 21252
rect 10388 21196 11452 21252
rect 11508 21196 11518 21252
rect 12758 21196 12796 21252
rect 12852 21196 12862 21252
rect 13010 21196 13020 21252
rect 13076 21196 15708 21252
rect 15764 21196 16940 21252
rect 16996 21196 17006 21252
rect 17164 21196 20076 21252
rect 20132 21196 20142 21252
rect 20290 21196 20300 21252
rect 20356 21196 20524 21252
rect 20580 21196 20590 21252
rect 20738 21196 20748 21252
rect 20804 21196 21420 21252
rect 21476 21196 21486 21252
rect 21644 21196 24332 21252
rect 24388 21196 24398 21252
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 1362 21084 1372 21140
rect 1428 21084 3052 21140
rect 3108 21084 3118 21140
rect 3490 21084 3500 21140
rect 3556 21084 4060 21140
rect 4116 21084 4126 21140
rect 4844 21028 4900 21196
rect 9772 21140 9828 21196
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 25004 21140 25060 21308
rect 26572 21252 26628 21308
rect 57344 21280 57456 21308
rect 25554 21196 25564 21252
rect 25620 21196 26628 21252
rect 27458 21196 27468 21252
rect 27524 21196 33180 21252
rect 33236 21196 33246 21252
rect 33394 21196 33404 21252
rect 33460 21196 42924 21252
rect 42980 21196 42990 21252
rect 45938 21196 45948 21252
rect 46004 21196 48916 21252
rect 49186 21196 49196 21252
rect 49252 21196 52780 21252
rect 52836 21196 52846 21252
rect 55654 21196 55692 21252
rect 55748 21196 55758 21252
rect 44454 21140 44464 21196
rect 44520 21140 44568 21196
rect 44624 21140 44672 21196
rect 44728 21140 44738 21196
rect 48860 21140 48916 21196
rect 5170 21084 5180 21140
rect 5236 21084 9548 21140
rect 9604 21084 9614 21140
rect 9772 21084 16380 21140
rect 16436 21084 16446 21140
rect 18162 21084 18172 21140
rect 18228 21084 22988 21140
rect 23044 21084 23054 21140
rect 25004 21084 26460 21140
rect 26516 21084 26526 21140
rect 26674 21084 26684 21140
rect 26740 21084 29036 21140
rect 29092 21084 29102 21140
rect 31266 21084 31276 21140
rect 31332 21084 36428 21140
rect 36484 21084 36494 21140
rect 39190 21084 39228 21140
rect 39284 21084 39294 21140
rect 40460 21084 41132 21140
rect 41188 21084 41198 21140
rect 41570 21084 41580 21140
rect 41636 21084 41804 21140
rect 41860 21084 41870 21140
rect 44828 21084 48636 21140
rect 48692 21084 48702 21140
rect 48860 21084 51884 21140
rect 51940 21084 51950 21140
rect 52322 21084 52332 21140
rect 52388 21084 52892 21140
rect 52948 21084 52958 21140
rect 1586 20972 1596 21028
rect 1652 20972 1708 21028
rect 1764 20972 1774 21028
rect 3490 20972 3500 21028
rect 3556 20972 4900 21028
rect 5282 20972 5292 21028
rect 5348 20972 32620 21028
rect 32676 20972 32686 21028
rect 36642 20972 36652 21028
rect 36708 20972 36764 21028
rect 36820 20972 36830 21028
rect 37650 20972 37660 21028
rect 37716 20972 38668 21028
rect 38724 20972 39116 21028
rect 39172 20972 39182 21028
rect 0 20916 112 20944
rect 40460 20916 40516 21084
rect 41804 21028 41860 21084
rect 44828 21028 44884 21084
rect 40786 20972 40796 21028
rect 40852 20972 41468 21028
rect 41524 20972 41534 21028
rect 41804 20972 44884 21028
rect 46610 20972 46620 21028
rect 46676 20972 47180 21028
rect 47236 20972 47246 21028
rect 48738 20972 48748 21028
rect 48804 20972 49756 21028
rect 49812 20972 49822 21028
rect 50166 20972 50204 21028
rect 50260 20972 50270 21028
rect 55570 20972 55580 21028
rect 55636 20972 56364 21028
rect 56420 20972 56430 21028
rect 57344 20916 57456 20944
rect 0 20860 812 20916
rect 868 20860 878 20916
rect 2828 20860 3052 20916
rect 3108 20860 4732 20916
rect 4788 20860 4798 20916
rect 5292 20860 9660 20916
rect 9716 20860 9726 20916
rect 10658 20860 10668 20916
rect 10724 20860 11340 20916
rect 11396 20860 11406 20916
rect 13794 20860 13804 20916
rect 13860 20860 14812 20916
rect 14868 20860 14878 20916
rect 17938 20860 17948 20916
rect 18004 20860 18172 20916
rect 18228 20860 18238 20916
rect 18610 20860 18620 20916
rect 18676 20860 23100 20916
rect 23156 20860 23166 20916
rect 23538 20860 23548 20916
rect 23604 20860 24220 20916
rect 24276 20860 24286 20916
rect 25302 20860 25340 20916
rect 25396 20860 25406 20916
rect 32620 20860 40516 20916
rect 40674 20860 40684 20916
rect 40740 20860 43036 20916
rect 43092 20860 43102 20916
rect 43586 20860 43596 20916
rect 43652 20860 45948 20916
rect 46004 20860 46014 20916
rect 46834 20860 46844 20916
rect 46900 20860 57456 20916
rect 0 20832 112 20860
rect 2828 20804 2884 20860
rect 5292 20804 5348 20860
rect 2818 20748 2828 20804
rect 2884 20748 2894 20804
rect 3042 20748 3052 20804
rect 3108 20748 5348 20804
rect 5478 20748 5516 20804
rect 5572 20748 5582 20804
rect 6066 20748 6076 20804
rect 6132 20748 6300 20804
rect 6356 20748 6366 20804
rect 6514 20748 6524 20804
rect 6580 20748 8764 20804
rect 8820 20748 8830 20804
rect 9314 20748 9324 20804
rect 9380 20748 11116 20804
rect 11172 20748 11182 20804
rect 14578 20748 14588 20804
rect 14644 20748 16828 20804
rect 16884 20748 16894 20804
rect 17826 20748 17836 20804
rect 17892 20748 19124 20804
rect 19842 20748 19852 20804
rect 19908 20748 23660 20804
rect 23716 20748 23726 20804
rect 23874 20748 23884 20804
rect 23940 20748 26124 20804
rect 26180 20748 26190 20804
rect 29474 20748 29484 20804
rect 29540 20748 31276 20804
rect 31332 20748 31342 20804
rect 19068 20692 19124 20748
rect 32620 20692 32676 20860
rect 57344 20832 57456 20860
rect 34290 20748 34300 20804
rect 34356 20748 34412 20804
rect 34468 20748 34860 20804
rect 34916 20748 34926 20804
rect 35970 20748 35980 20804
rect 36036 20748 38892 20804
rect 38948 20748 38958 20804
rect 39666 20748 39676 20804
rect 39732 20748 40348 20804
rect 40404 20748 40414 20804
rect 40758 20748 40796 20804
rect 40852 20748 40862 20804
rect 41458 20748 41468 20804
rect 41524 20748 42364 20804
rect 42420 20748 42430 20804
rect 42578 20748 42588 20804
rect 42644 20748 43316 20804
rect 43474 20748 43484 20804
rect 43540 20748 46620 20804
rect 46676 20748 46686 20804
rect 48636 20748 49532 20804
rect 49588 20748 49598 20804
rect 51622 20748 51660 20804
rect 51716 20748 51726 20804
rect 52546 20748 52556 20804
rect 52612 20748 54460 20804
rect 54516 20748 54526 20804
rect 43260 20692 43316 20748
rect 48636 20692 48692 20748
rect 2370 20636 2380 20692
rect 2436 20636 3164 20692
rect 3220 20636 3230 20692
rect 5394 20636 5404 20692
rect 5460 20636 8092 20692
rect 8148 20636 8158 20692
rect 9202 20636 9212 20692
rect 9268 20636 9772 20692
rect 9828 20636 9838 20692
rect 11218 20636 11228 20692
rect 11284 20636 11788 20692
rect 11844 20636 11854 20692
rect 12674 20636 12684 20692
rect 12740 20636 18844 20692
rect 18900 20636 18910 20692
rect 19068 20636 20860 20692
rect 20916 20636 21084 20692
rect 21140 20636 22316 20692
rect 22372 20636 23212 20692
rect 23268 20636 23278 20692
rect 23426 20636 23436 20692
rect 23492 20636 24556 20692
rect 24612 20636 24622 20692
rect 24770 20636 24780 20692
rect 24836 20636 26684 20692
rect 26740 20636 26750 20692
rect 27794 20636 27804 20692
rect 27860 20636 28364 20692
rect 28420 20636 28700 20692
rect 28756 20636 28766 20692
rect 29138 20636 29148 20692
rect 29204 20636 32676 20692
rect 35970 20636 35980 20692
rect 36036 20636 36204 20692
rect 36260 20636 36540 20692
rect 36596 20636 36606 20692
rect 39106 20636 39116 20692
rect 39172 20636 39564 20692
rect 39620 20636 40236 20692
rect 40292 20636 40572 20692
rect 40628 20636 41020 20692
rect 41076 20636 42812 20692
rect 42868 20636 42878 20692
rect 43260 20636 45388 20692
rect 45444 20636 47068 20692
rect 48626 20636 48636 20692
rect 48692 20636 48702 20692
rect 52994 20636 53004 20692
rect 53060 20636 54124 20692
rect 54180 20636 54190 20692
rect 47012 20580 47068 20636
rect 2034 20524 2044 20580
rect 2100 20524 13580 20580
rect 13636 20524 13646 20580
rect 14242 20524 14252 20580
rect 14308 20524 17948 20580
rect 18004 20524 18014 20580
rect 18274 20524 18284 20580
rect 18340 20524 21868 20580
rect 21924 20524 22204 20580
rect 22260 20524 22270 20580
rect 22642 20524 22652 20580
rect 22708 20524 24892 20580
rect 24948 20524 24958 20580
rect 25106 20524 25116 20580
rect 25172 20524 25210 20580
rect 26226 20524 26236 20580
rect 26292 20524 28700 20580
rect 28756 20524 29372 20580
rect 29428 20524 29438 20580
rect 31602 20524 31612 20580
rect 31668 20524 31724 20580
rect 31780 20524 31790 20580
rect 33170 20524 33180 20580
rect 33236 20524 33852 20580
rect 33908 20524 33918 20580
rect 39218 20524 39228 20580
rect 39284 20524 40908 20580
rect 40964 20524 40974 20580
rect 41234 20524 41244 20580
rect 41300 20524 46508 20580
rect 46564 20524 46574 20580
rect 47012 20524 49868 20580
rect 49924 20524 49934 20580
rect 51538 20524 51548 20580
rect 51604 20524 51996 20580
rect 52052 20524 52062 20580
rect 0 20468 112 20496
rect 57344 20468 57456 20496
rect 0 20412 3276 20468
rect 3332 20412 3342 20468
rect 4946 20412 4956 20468
rect 5012 20412 5964 20468
rect 6020 20412 6030 20468
rect 6290 20412 6300 20468
rect 6356 20412 6412 20468
rect 6468 20412 10556 20468
rect 10612 20412 10622 20468
rect 10770 20412 10780 20468
rect 10836 20412 11452 20468
rect 11508 20412 11518 20468
rect 11890 20412 11900 20468
rect 11956 20412 15820 20468
rect 15876 20412 15886 20468
rect 16146 20412 16156 20468
rect 16212 20412 16492 20468
rect 16548 20412 16558 20468
rect 17266 20412 17276 20468
rect 17332 20412 18620 20468
rect 18676 20412 19964 20468
rect 20020 20412 20748 20468
rect 20804 20412 20814 20468
rect 20962 20412 20972 20468
rect 21028 20412 22876 20468
rect 22932 20412 22942 20468
rect 24546 20412 24556 20468
rect 24612 20412 27132 20468
rect 27188 20412 28028 20468
rect 28084 20412 28094 20468
rect 30034 20412 30044 20468
rect 30100 20412 32284 20468
rect 32340 20412 32350 20468
rect 32498 20412 32508 20468
rect 32564 20412 35308 20468
rect 35364 20412 35374 20468
rect 41010 20412 41020 20468
rect 41076 20412 41580 20468
rect 41636 20412 41646 20468
rect 42018 20412 42028 20468
rect 42084 20412 43596 20468
rect 43652 20412 43662 20468
rect 47170 20412 47180 20468
rect 47236 20412 57456 20468
rect 0 20384 112 20412
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 43794 20356 43804 20412
rect 43860 20356 43908 20412
rect 43964 20356 44012 20412
rect 44068 20356 44078 20412
rect 57344 20384 57456 20412
rect 1810 20300 1820 20356
rect 1876 20300 2716 20356
rect 2772 20300 3052 20356
rect 3108 20300 3118 20356
rect 5180 20300 21028 20356
rect 23426 20300 23436 20356
rect 23492 20300 23660 20356
rect 23716 20300 23726 20356
rect 24210 20300 24220 20356
rect 24276 20300 25228 20356
rect 25284 20300 25294 20356
rect 25778 20300 25788 20356
rect 25844 20300 27468 20356
rect 27524 20300 27534 20356
rect 28466 20300 28476 20356
rect 28532 20300 33068 20356
rect 33124 20300 33134 20356
rect 34290 20300 34300 20356
rect 34356 20300 37436 20356
rect 37492 20300 37548 20356
rect 37604 20300 37614 20356
rect 38546 20300 38556 20356
rect 38612 20300 38892 20356
rect 38948 20300 38958 20356
rect 41122 20300 41132 20356
rect 41188 20300 41916 20356
rect 41972 20300 41982 20356
rect 45826 20300 45836 20356
rect 45892 20300 46844 20356
rect 46900 20300 46910 20356
rect 47618 20300 47628 20356
rect 47684 20300 52444 20356
rect 52500 20300 52510 20356
rect 1250 20188 1260 20244
rect 1316 20188 2772 20244
rect 2716 20132 2772 20188
rect 5180 20132 5236 20300
rect 20972 20244 21028 20300
rect 6178 20188 6188 20244
rect 6244 20188 8540 20244
rect 8596 20188 8606 20244
rect 8764 20188 12684 20244
rect 12740 20188 12750 20244
rect 14102 20188 14140 20244
rect 14196 20188 18284 20244
rect 18340 20188 18350 20244
rect 18498 20188 18508 20244
rect 18564 20188 20468 20244
rect 20972 20188 50428 20244
rect 50484 20188 50494 20244
rect 51314 20188 51324 20244
rect 51380 20188 51884 20244
rect 51940 20188 51950 20244
rect 54450 20188 54460 20244
rect 54516 20188 55020 20244
rect 55076 20188 55086 20244
rect 55346 20188 55356 20244
rect 55412 20188 56140 20244
rect 56196 20188 56206 20244
rect 8764 20132 8820 20188
rect 20412 20132 20468 20188
rect 1586 20076 1596 20132
rect 1652 20076 1932 20132
rect 1988 20076 1998 20132
rect 2706 20076 2716 20132
rect 2772 20076 2782 20132
rect 3602 20076 3612 20132
rect 3668 20076 5236 20132
rect 7634 20076 7644 20132
rect 7700 20076 8820 20132
rect 9202 20076 9212 20132
rect 9268 20076 9884 20132
rect 9940 20076 11004 20132
rect 11060 20076 11070 20132
rect 14466 20076 14476 20132
rect 14532 20076 17164 20132
rect 17220 20076 17230 20132
rect 17602 20076 17612 20132
rect 17668 20076 19628 20132
rect 19684 20076 19694 20132
rect 20412 20076 25396 20132
rect 25554 20076 25564 20132
rect 25620 20076 26684 20132
rect 26740 20076 26908 20132
rect 29810 20076 29820 20132
rect 29876 20076 30380 20132
rect 30436 20076 30446 20132
rect 31266 20076 31276 20132
rect 31332 20076 33292 20132
rect 33348 20076 33358 20132
rect 35298 20076 35308 20132
rect 35364 20076 44268 20132
rect 44324 20076 44334 20132
rect 45602 20076 45612 20132
rect 45668 20076 48636 20132
rect 48692 20076 48702 20132
rect 48850 20076 48860 20132
rect 48916 20076 50092 20132
rect 50148 20076 54460 20132
rect 54516 20076 54526 20132
rect 0 20020 112 20048
rect 25340 20020 25396 20076
rect 26852 20020 26908 20076
rect 57344 20020 57456 20048
rect 0 19964 3948 20020
rect 4004 19964 4014 20020
rect 4386 19964 4396 20020
rect 4452 19964 4844 20020
rect 4900 19964 4910 20020
rect 5702 19964 5740 20020
rect 5796 19964 6300 20020
rect 6356 19964 6366 20020
rect 6626 19964 6636 20020
rect 6692 19964 9436 20020
rect 9492 19964 10108 20020
rect 10164 19964 13580 20020
rect 13636 19964 13646 20020
rect 14802 19964 14812 20020
rect 14868 19964 15484 20020
rect 15540 19964 18060 20020
rect 18116 19964 18126 20020
rect 18284 19964 21532 20020
rect 21588 19964 21598 20020
rect 22418 19964 22428 20020
rect 22484 19964 23436 20020
rect 23492 19964 23502 20020
rect 23650 19964 23660 20020
rect 23716 19964 25004 20020
rect 25060 19964 25070 20020
rect 25340 19964 25452 20020
rect 25508 19964 25518 20020
rect 26226 19964 26236 20020
rect 26292 19964 26460 20020
rect 26516 19964 26526 20020
rect 26852 19964 29876 20020
rect 30034 19964 30044 20020
rect 30100 19964 30940 20020
rect 30996 19964 31052 20020
rect 31108 19964 31118 20020
rect 31490 19964 31500 20020
rect 31556 19964 32284 20020
rect 32340 19964 32350 20020
rect 37090 19964 37100 20020
rect 37156 19964 39340 20020
rect 39396 19964 40572 20020
rect 40628 19964 40638 20020
rect 41346 19964 41356 20020
rect 41412 19964 42700 20020
rect 42756 19964 42766 20020
rect 43362 19964 43372 20020
rect 43428 19964 45332 20020
rect 46386 19964 46396 20020
rect 46452 19964 47068 20020
rect 47124 19964 47134 20020
rect 47394 19964 47404 20020
rect 47460 19964 47964 20020
rect 48020 19964 48030 20020
rect 48402 19964 48412 20020
rect 48468 19964 57456 20020
rect 0 19936 112 19964
rect 18284 19908 18340 19964
rect 29820 19908 29876 19964
rect 45276 19908 45332 19964
rect 57344 19936 57456 19964
rect 3378 19852 3388 19908
rect 3444 19852 4844 19908
rect 4900 19852 9884 19908
rect 9940 19852 9950 19908
rect 10658 19852 10668 19908
rect 10724 19852 10780 19908
rect 10836 19852 10846 19908
rect 11106 19852 11116 19908
rect 11172 19852 11788 19908
rect 11844 19852 11854 19908
rect 12226 19852 12236 19908
rect 12292 19852 13580 19908
rect 13636 19852 13646 19908
rect 15362 19852 15372 19908
rect 15428 19852 15596 19908
rect 15652 19852 15662 19908
rect 16482 19852 16492 19908
rect 16548 19852 16716 19908
rect 16772 19852 18340 19908
rect 18946 19852 18956 19908
rect 19012 19852 22316 19908
rect 22372 19852 22382 19908
rect 23090 19852 23100 19908
rect 23156 19852 23436 19908
rect 23492 19852 23502 19908
rect 24210 19852 24220 19908
rect 24276 19852 25116 19908
rect 25172 19852 25182 19908
rect 25330 19852 25340 19908
rect 25396 19852 26572 19908
rect 26628 19852 26638 19908
rect 29138 19852 29148 19908
rect 29204 19852 29596 19908
rect 29652 19852 29662 19908
rect 29820 19852 31556 19908
rect 33842 19852 33852 19908
rect 33908 19852 34972 19908
rect 35028 19852 35038 19908
rect 36866 19852 36876 19908
rect 36932 19852 39788 19908
rect 39844 19852 39854 19908
rect 41122 19852 41132 19908
rect 41188 19852 43148 19908
rect 43204 19852 43214 19908
rect 44258 19852 44268 19908
rect 44324 19852 45052 19908
rect 45108 19852 45118 19908
rect 45276 19852 46508 19908
rect 46564 19852 46574 19908
rect 47394 19852 47404 19908
rect 47460 19852 50428 19908
rect 50866 19852 50876 19908
rect 50932 19852 52108 19908
rect 52164 19852 52174 19908
rect 52630 19852 52668 19908
rect 52724 19852 52734 19908
rect 53218 19852 53228 19908
rect 53284 19852 53452 19908
rect 53508 19852 53676 19908
rect 53732 19852 53900 19908
rect 53956 19852 53966 19908
rect 31500 19796 31556 19852
rect 50372 19796 50428 19852
rect 1138 19740 1148 19796
rect 1204 19740 1484 19796
rect 1540 19740 1550 19796
rect 3332 19740 4396 19796
rect 4452 19740 4462 19796
rect 5730 19740 5740 19796
rect 5796 19740 6300 19796
rect 6356 19740 6366 19796
rect 7186 19740 7196 19796
rect 7252 19740 7756 19796
rect 7812 19740 9772 19796
rect 9828 19740 9838 19796
rect 10322 19740 10332 19796
rect 10388 19740 11004 19796
rect 11060 19740 12012 19796
rect 12068 19740 12078 19796
rect 13570 19740 13580 19796
rect 13636 19740 25396 19796
rect 26226 19740 26236 19796
rect 26292 19740 29708 19796
rect 29764 19740 29774 19796
rect 31490 19740 31500 19796
rect 31556 19740 32844 19796
rect 32900 19740 33292 19796
rect 33348 19740 33358 19796
rect 33506 19740 33516 19796
rect 33572 19740 34300 19796
rect 34356 19740 34366 19796
rect 35522 19740 35532 19796
rect 35588 19740 38556 19796
rect 38612 19740 38622 19796
rect 42914 19740 42924 19796
rect 42980 19740 45164 19796
rect 45220 19740 45836 19796
rect 45892 19740 45902 19796
rect 46050 19740 46060 19796
rect 46116 19740 47068 19796
rect 47124 19740 47134 19796
rect 50372 19740 54348 19796
rect 54404 19740 54414 19796
rect 54562 19740 54572 19796
rect 54628 19740 55468 19796
rect 55524 19740 55534 19796
rect 0 19572 112 19600
rect 3332 19572 3388 19740
rect 25340 19684 25396 19740
rect 5842 19628 5852 19684
rect 5908 19628 18284 19684
rect 18340 19628 18350 19684
rect 18498 19628 18508 19684
rect 18564 19628 24220 19684
rect 24276 19628 24286 19684
rect 25330 19628 25340 19684
rect 25396 19628 25406 19684
rect 27878 19628 27916 19684
rect 27972 19628 28420 19684
rect 33394 19628 33404 19684
rect 33460 19628 41132 19684
rect 41188 19628 41198 19684
rect 42130 19628 42140 19684
rect 42196 19628 44156 19684
rect 44212 19628 44222 19684
rect 44828 19628 55916 19684
rect 55972 19628 55982 19684
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 28364 19572 28420 19628
rect 44454 19572 44464 19628
rect 44520 19572 44568 19628
rect 44624 19572 44672 19628
rect 44728 19572 44738 19628
rect 0 19516 3388 19572
rect 5058 19516 5068 19572
rect 5124 19516 6132 19572
rect 6290 19516 6300 19572
rect 6356 19516 15876 19572
rect 16258 19516 16268 19572
rect 16324 19516 16604 19572
rect 16660 19516 16670 19572
rect 18050 19516 18060 19572
rect 18116 19516 19740 19572
rect 19796 19516 19806 19572
rect 20066 19516 20076 19572
rect 20132 19516 21308 19572
rect 21364 19516 21374 19572
rect 21522 19516 21532 19572
rect 21588 19516 24108 19572
rect 24164 19516 24174 19572
rect 24994 19516 25004 19572
rect 25060 19516 27692 19572
rect 27748 19516 27758 19572
rect 28364 19516 44268 19572
rect 44324 19516 44334 19572
rect 0 19488 112 19516
rect 6076 19460 6132 19516
rect 2370 19404 2380 19460
rect 2436 19404 5852 19460
rect 5908 19404 5918 19460
rect 6076 19404 9044 19460
rect 9202 19404 9212 19460
rect 9268 19404 11004 19460
rect 11060 19404 11070 19460
rect 12002 19404 12012 19460
rect 12068 19404 13356 19460
rect 13412 19404 13422 19460
rect 8988 19348 9044 19404
rect 15820 19348 15876 19516
rect 16034 19404 16044 19460
rect 16100 19404 16828 19460
rect 16884 19404 16894 19460
rect 17154 19404 17164 19460
rect 17220 19404 18396 19460
rect 18452 19404 19292 19460
rect 19348 19404 19358 19460
rect 20290 19404 20300 19460
rect 20356 19404 35084 19460
rect 35140 19404 35150 19460
rect 37538 19404 37548 19460
rect 37604 19404 41020 19460
rect 41076 19404 41086 19460
rect 41570 19404 41580 19460
rect 41636 19404 42140 19460
rect 42196 19404 42206 19460
rect 42354 19404 42364 19460
rect 42420 19404 42812 19460
rect 42868 19404 42878 19460
rect 43026 19404 43036 19460
rect 43092 19404 43596 19460
rect 43652 19404 43662 19460
rect 44828 19348 44884 19628
rect 57344 19572 57456 19600
rect 45490 19516 45500 19572
rect 45556 19516 48860 19572
rect 48916 19516 48926 19572
rect 50418 19516 50428 19572
rect 50484 19516 51884 19572
rect 51940 19516 51950 19572
rect 52770 19516 52780 19572
rect 52836 19516 57456 19572
rect 57344 19488 57456 19516
rect 45126 19404 45164 19460
rect 45220 19404 45230 19460
rect 49186 19404 49196 19460
rect 49252 19404 50540 19460
rect 50596 19404 50606 19460
rect 50988 19404 54516 19460
rect 54674 19404 54684 19460
rect 54740 19404 56028 19460
rect 56084 19404 56094 19460
rect 56354 19404 56364 19460
rect 56420 19404 57148 19460
rect 57204 19404 57214 19460
rect 50988 19348 51044 19404
rect 54460 19348 54516 19404
rect 1474 19292 1484 19348
rect 1540 19292 5964 19348
rect 6020 19292 6030 19348
rect 8988 19292 9884 19348
rect 9940 19292 9950 19348
rect 10770 19292 10780 19348
rect 10836 19292 13468 19348
rect 13524 19292 13534 19348
rect 15820 19292 18956 19348
rect 19012 19292 19022 19348
rect 19394 19292 19404 19348
rect 19460 19292 20748 19348
rect 20804 19292 20814 19348
rect 23650 19292 23660 19348
rect 23716 19292 26348 19348
rect 26404 19292 26414 19348
rect 29474 19292 29484 19348
rect 29540 19292 31836 19348
rect 31892 19292 35308 19348
rect 35364 19292 35374 19348
rect 40236 19292 44884 19348
rect 45266 19292 45276 19348
rect 45332 19292 46620 19348
rect 46676 19292 46686 19348
rect 49634 19292 49644 19348
rect 49700 19292 51044 19348
rect 51874 19292 51884 19348
rect 51940 19292 53228 19348
rect 53284 19292 53294 19348
rect 53554 19292 53564 19348
rect 53620 19292 54236 19348
rect 54292 19292 54302 19348
rect 54460 19292 54572 19348
rect 54628 19292 54638 19348
rect 56700 19292 56924 19348
rect 56980 19292 56990 19348
rect 2370 19180 2380 19236
rect 2436 19180 6076 19236
rect 6132 19180 6142 19236
rect 7158 19180 7196 19236
rect 7252 19180 7262 19236
rect 8194 19180 8204 19236
rect 8260 19180 9324 19236
rect 9380 19180 9390 19236
rect 11554 19180 11564 19236
rect 11620 19180 12796 19236
rect 12852 19180 12862 19236
rect 13010 19180 13020 19236
rect 13076 19180 14252 19236
rect 14308 19180 14476 19236
rect 14532 19180 14542 19236
rect 14812 19180 15092 19236
rect 19058 19180 19068 19236
rect 19124 19180 20076 19236
rect 20132 19180 20142 19236
rect 21382 19180 21420 19236
rect 21476 19180 21486 19236
rect 21746 19180 21756 19236
rect 21812 19180 24332 19236
rect 24388 19180 26236 19236
rect 26292 19180 26302 19236
rect 26450 19180 26460 19236
rect 26516 19180 27244 19236
rect 27300 19180 27310 19236
rect 27794 19180 27804 19236
rect 27860 19180 28364 19236
rect 28420 19180 28430 19236
rect 28886 19180 28924 19236
rect 28980 19180 29596 19236
rect 29652 19180 29662 19236
rect 29894 19180 29932 19236
rect 29988 19180 29998 19236
rect 33058 19180 33068 19236
rect 33124 19180 34188 19236
rect 34244 19180 34636 19236
rect 34692 19180 34702 19236
rect 34962 19180 34972 19236
rect 35028 19180 36988 19236
rect 37044 19180 37054 19236
rect 38434 19180 38444 19236
rect 38500 19180 38892 19236
rect 38948 19180 38958 19236
rect 0 19124 112 19152
rect 14812 19124 14868 19180
rect 0 19068 812 19124
rect 868 19068 878 19124
rect 2146 19068 2156 19124
rect 2212 19068 7644 19124
rect 7700 19068 7710 19124
rect 10210 19068 10220 19124
rect 10276 19068 10668 19124
rect 10724 19068 10734 19124
rect 10994 19068 11004 19124
rect 11060 19068 14868 19124
rect 15036 19124 15092 19180
rect 40236 19124 40292 19292
rect 56700 19236 56756 19292
rect 40450 19180 40460 19236
rect 40516 19180 42588 19236
rect 42644 19180 42654 19236
rect 43698 19180 43708 19236
rect 43764 19180 45052 19236
rect 45108 19180 45612 19236
rect 45668 19180 45678 19236
rect 45826 19180 45836 19236
rect 45892 19180 46620 19236
rect 46676 19180 46686 19236
rect 47842 19180 47852 19236
rect 47908 19180 47964 19236
rect 48020 19180 48030 19236
rect 48962 19180 48972 19236
rect 49028 19180 53452 19236
rect 53508 19180 53518 19236
rect 54450 19180 54460 19236
rect 54516 19180 56252 19236
rect 56308 19180 56318 19236
rect 56690 19180 56700 19236
rect 56756 19180 56766 19236
rect 57344 19124 57456 19152
rect 15036 19068 25564 19124
rect 25620 19068 25630 19124
rect 28690 19068 28700 19124
rect 28756 19068 30716 19124
rect 30772 19068 30782 19124
rect 31798 19068 31836 19124
rect 31892 19068 31902 19124
rect 33730 19068 33740 19124
rect 33796 19068 40292 19124
rect 40534 19068 40572 19124
rect 40628 19068 40638 19124
rect 41122 19068 41132 19124
rect 41188 19068 42028 19124
rect 42084 19068 42094 19124
rect 42354 19068 42364 19124
rect 42420 19068 42700 19124
rect 42756 19068 42766 19124
rect 44258 19068 44268 19124
rect 44324 19068 50316 19124
rect 50372 19068 50382 19124
rect 53106 19068 53116 19124
rect 53172 19068 55356 19124
rect 55412 19068 55422 19124
rect 56914 19068 56924 19124
rect 56980 19068 57456 19124
rect 0 19040 112 19068
rect 57344 19040 57456 19068
rect 242 18956 252 19012
rect 308 18956 6300 19012
rect 6356 18956 6366 19012
rect 6514 18956 6524 19012
rect 6580 18956 13580 19012
rect 13636 18956 14252 19012
rect 14308 18956 14318 19012
rect 20860 18956 32228 19012
rect 34850 18956 34860 19012
rect 34916 18956 34972 19012
rect 35028 18956 35038 19012
rect 37986 18956 37996 19012
rect 38052 18956 38668 19012
rect 38724 18956 38734 19012
rect 41122 18956 41132 19012
rect 41188 18956 41804 19012
rect 41860 18956 41870 19012
rect 42588 18956 48076 19012
rect 48132 18956 48142 19012
rect 50194 18956 50204 19012
rect 50260 18956 51996 19012
rect 52052 18956 52062 19012
rect 20860 18900 20916 18956
rect 32172 18900 32228 18956
rect 690 18844 700 18900
rect 756 18844 1484 18900
rect 1540 18844 1550 18900
rect 2034 18844 2044 18900
rect 2100 18844 2492 18900
rect 2548 18844 2558 18900
rect 4274 18844 4284 18900
rect 4340 18844 20916 18900
rect 24210 18844 24220 18900
rect 24276 18844 30940 18900
rect 30996 18844 31006 18900
rect 32172 18844 41244 18900
rect 41300 18844 41310 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 2492 18732 2716 18788
rect 2772 18732 2782 18788
rect 4610 18732 4620 18788
rect 4676 18732 6076 18788
rect 6132 18732 6142 18788
rect 6300 18732 7644 18788
rect 7700 18732 7710 18788
rect 9650 18732 9660 18788
rect 9716 18732 9996 18788
rect 10052 18732 10062 18788
rect 14242 18732 14252 18788
rect 14308 18732 16268 18788
rect 16324 18732 16334 18788
rect 18274 18732 18284 18788
rect 18340 18732 20412 18788
rect 20468 18732 23716 18788
rect 0 18676 112 18704
rect 2492 18676 2548 18732
rect 6300 18676 6356 18732
rect 23660 18676 23716 18732
rect 24220 18732 25004 18788
rect 25060 18732 25070 18788
rect 26338 18732 26348 18788
rect 26404 18732 26796 18788
rect 26852 18732 26862 18788
rect 30818 18732 30828 18788
rect 30884 18732 31612 18788
rect 31668 18732 32508 18788
rect 32564 18732 34188 18788
rect 34244 18732 34860 18788
rect 34916 18732 34926 18788
rect 35074 18732 35084 18788
rect 35140 18732 39340 18788
rect 39396 18732 39406 18788
rect 40982 18732 41020 18788
rect 41076 18732 41086 18788
rect 24220 18676 24276 18732
rect 0 18620 252 18676
rect 308 18620 318 18676
rect 2482 18620 2492 18676
rect 2548 18620 2558 18676
rect 3154 18620 3164 18676
rect 3220 18620 6356 18676
rect 6514 18620 6524 18676
rect 6580 18620 23548 18676
rect 23660 18620 24276 18676
rect 24332 18620 38668 18676
rect 39666 18620 39676 18676
rect 39732 18620 40572 18676
rect 40628 18620 40638 18676
rect 0 18592 112 18620
rect 23492 18564 23548 18620
rect 24332 18564 24388 18620
rect 38612 18564 38668 18620
rect 42588 18564 42644 18956
rect 44146 18844 44156 18900
rect 44212 18844 46396 18900
rect 46452 18844 46462 18900
rect 46620 18844 48244 18900
rect 49746 18844 49756 18900
rect 49812 18844 50428 18900
rect 50484 18844 50494 18900
rect 51202 18844 51212 18900
rect 51268 18844 53452 18900
rect 53508 18844 53518 18900
rect 43794 18788 43804 18844
rect 43860 18788 43908 18844
rect 43964 18788 44012 18844
rect 44068 18788 44078 18844
rect 46620 18788 46676 18844
rect 48188 18788 48244 18844
rect 45332 18732 46676 18788
rect 47282 18732 47292 18788
rect 47348 18732 47964 18788
rect 48020 18732 48030 18788
rect 48188 18732 50316 18788
rect 50372 18732 50382 18788
rect 51650 18732 51660 18788
rect 51716 18732 55468 18788
rect 45332 18676 45388 18732
rect 55412 18676 55468 18732
rect 57344 18676 57456 18704
rect 42802 18620 42812 18676
rect 42868 18620 43932 18676
rect 43988 18620 43998 18676
rect 44604 18620 45388 18676
rect 45602 18620 45612 18676
rect 45668 18620 45836 18676
rect 45892 18620 47068 18676
rect 47954 18620 47964 18676
rect 48020 18620 48300 18676
rect 48356 18620 48366 18676
rect 51314 18620 51324 18676
rect 51380 18620 53004 18676
rect 53060 18620 53070 18676
rect 53638 18620 53676 18676
rect 53732 18620 53742 18676
rect 55412 18620 57456 18676
rect 354 18508 364 18564
rect 420 18508 3388 18564
rect 3444 18508 3454 18564
rect 4162 18508 4172 18564
rect 4228 18508 5852 18564
rect 5908 18508 6412 18564
rect 6468 18508 6478 18564
rect 8194 18508 8204 18564
rect 8260 18508 11340 18564
rect 11396 18508 11406 18564
rect 12674 18508 12684 18564
rect 12740 18508 14924 18564
rect 14980 18508 14990 18564
rect 16258 18508 16268 18564
rect 16324 18508 20412 18564
rect 20468 18508 20478 18564
rect 23492 18508 24388 18564
rect 25442 18508 25452 18564
rect 25508 18508 27188 18564
rect 27346 18508 27356 18564
rect 27412 18508 27692 18564
rect 27748 18508 27758 18564
rect 28690 18508 28700 18564
rect 28756 18508 29708 18564
rect 29764 18508 30044 18564
rect 30100 18508 30110 18564
rect 33170 18508 33180 18564
rect 33236 18508 34300 18564
rect 34356 18508 34366 18564
rect 34514 18508 34524 18564
rect 34580 18508 35980 18564
rect 36036 18508 36046 18564
rect 36530 18508 36540 18564
rect 36596 18508 36988 18564
rect 37044 18508 37054 18564
rect 38612 18508 42644 18564
rect 43026 18508 43036 18564
rect 43092 18508 43708 18564
rect 43764 18508 43774 18564
rect 27132 18452 27188 18508
rect 44604 18452 44660 18620
rect 47012 18564 47068 18620
rect 57344 18592 57456 18620
rect 44818 18508 44828 18564
rect 44884 18508 46732 18564
rect 46788 18508 46798 18564
rect 47012 18508 49084 18564
rect 49140 18508 49150 18564
rect 50866 18508 50876 18564
rect 50932 18508 51212 18564
rect 51268 18508 51278 18564
rect 52098 18508 52108 18564
rect 52164 18508 52174 18564
rect 53106 18508 53116 18564
rect 53172 18508 53564 18564
rect 53620 18508 53630 18564
rect 52108 18452 52164 18508
rect 1250 18396 1260 18452
rect 1316 18396 2604 18452
rect 2660 18396 2670 18452
rect 4274 18396 4284 18452
rect 4340 18396 6188 18452
rect 6244 18396 6524 18452
rect 6580 18396 6590 18452
rect 7298 18396 7308 18452
rect 7364 18396 7420 18452
rect 7476 18396 7486 18452
rect 7970 18396 7980 18452
rect 8036 18396 9100 18452
rect 9156 18396 9166 18452
rect 9314 18396 9324 18452
rect 9380 18396 10556 18452
rect 10612 18396 11228 18452
rect 11284 18396 11294 18452
rect 11732 18396 12236 18452
rect 12292 18396 12908 18452
rect 12964 18396 12974 18452
rect 13234 18396 13244 18452
rect 13300 18396 14812 18452
rect 14868 18396 14878 18452
rect 14998 18396 15036 18452
rect 15092 18396 15102 18452
rect 17126 18396 17164 18452
rect 17220 18396 17230 18452
rect 18022 18396 18060 18452
rect 18116 18396 18126 18452
rect 20290 18396 20300 18452
rect 20356 18396 24892 18452
rect 24948 18396 26236 18452
rect 26292 18396 26302 18452
rect 27132 18396 29372 18452
rect 29428 18396 29438 18452
rect 30258 18396 30268 18452
rect 30324 18396 32732 18452
rect 32788 18396 33516 18452
rect 33572 18396 34412 18452
rect 34468 18396 34478 18452
rect 35084 18396 35308 18452
rect 37090 18396 37100 18452
rect 37156 18396 38780 18452
rect 38836 18396 38846 18452
rect 40450 18396 40460 18452
rect 40516 18396 40908 18452
rect 40964 18396 41580 18452
rect 41636 18396 41646 18452
rect 42242 18396 42252 18452
rect 42308 18396 43260 18452
rect 43316 18396 43326 18452
rect 44258 18396 44268 18452
rect 44324 18396 44660 18452
rect 45378 18396 45388 18452
rect 45444 18396 49420 18452
rect 49476 18396 49486 18452
rect 49634 18396 49644 18452
rect 49700 18396 50204 18452
rect 50260 18396 50270 18452
rect 51314 18396 51324 18452
rect 51380 18396 52164 18452
rect 52406 18396 52444 18452
rect 52500 18396 52510 18452
rect 52658 18396 52668 18452
rect 52724 18396 54684 18452
rect 54740 18396 54750 18452
rect 11732 18340 11788 18396
rect 35084 18340 35140 18396
rect 3126 18284 3164 18340
rect 3220 18284 3230 18340
rect 4274 18284 4284 18340
rect 4340 18284 6916 18340
rect 7074 18284 7084 18340
rect 7140 18284 9436 18340
rect 9492 18284 9502 18340
rect 9986 18284 9996 18340
rect 10052 18284 10668 18340
rect 10724 18284 10734 18340
rect 10994 18284 11004 18340
rect 11060 18284 11788 18340
rect 12002 18284 12012 18340
rect 12068 18284 14252 18340
rect 14308 18284 14318 18340
rect 17042 18284 17052 18340
rect 17108 18284 21308 18340
rect 21364 18284 21374 18340
rect 23090 18284 23100 18340
rect 23156 18284 26124 18340
rect 26180 18284 26190 18340
rect 28354 18284 28364 18340
rect 28420 18284 31276 18340
rect 31332 18284 31342 18340
rect 31490 18284 31500 18340
rect 31556 18284 35140 18340
rect 35252 18340 35308 18396
rect 35252 18284 35420 18340
rect 35476 18284 35486 18340
rect 35746 18284 35756 18340
rect 35812 18284 36316 18340
rect 36372 18284 36382 18340
rect 37090 18284 37100 18340
rect 37156 18284 37324 18340
rect 37380 18284 37390 18340
rect 37538 18284 37548 18340
rect 37604 18284 45668 18340
rect 46946 18284 46956 18340
rect 47012 18284 47180 18340
rect 47236 18284 47246 18340
rect 50866 18284 50876 18340
rect 50932 18284 51772 18340
rect 51828 18284 51838 18340
rect 52098 18284 52108 18340
rect 52164 18284 52332 18340
rect 52388 18284 52398 18340
rect 54786 18284 54796 18340
rect 54852 18284 56364 18340
rect 56420 18284 56430 18340
rect 0 18228 112 18256
rect 0 18172 924 18228
rect 980 18172 990 18228
rect 1362 18172 1372 18228
rect 1428 18172 1708 18228
rect 1764 18172 1774 18228
rect 4284 18172 6636 18228
rect 6692 18172 6702 18228
rect 0 18144 112 18172
rect 4284 18116 4340 18172
rect 242 18060 252 18116
rect 308 18060 4340 18116
rect 5506 18060 5516 18116
rect 5572 18060 5628 18116
rect 5684 18060 5694 18116
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 6860 18004 6916 18284
rect 9762 18172 9772 18228
rect 9828 18172 12348 18228
rect 12404 18172 12414 18228
rect 12898 18172 12908 18228
rect 12964 18172 13020 18228
rect 13076 18172 13086 18228
rect 16258 18172 16268 18228
rect 16324 18172 17948 18228
rect 18004 18172 18014 18228
rect 21522 18172 21532 18228
rect 21588 18172 26796 18228
rect 26852 18172 26862 18228
rect 27234 18172 27244 18228
rect 27300 18172 30828 18228
rect 30884 18172 30894 18228
rect 31378 18172 31388 18228
rect 31444 18172 36988 18228
rect 37044 18172 37054 18228
rect 37762 18172 37772 18228
rect 37828 18172 41020 18228
rect 41076 18172 41086 18228
rect 41906 18172 41916 18228
rect 41972 18172 44828 18228
rect 44884 18172 44894 18228
rect 7746 18060 7756 18116
rect 7812 18060 7868 18116
rect 7924 18060 8988 18116
rect 9044 18060 9054 18116
rect 9538 18060 9548 18116
rect 9604 18060 10892 18116
rect 10948 18060 10958 18116
rect 11442 18060 11452 18116
rect 11508 18060 16044 18116
rect 16100 18060 16110 18116
rect 19394 18060 19404 18116
rect 19460 18060 22764 18116
rect 22820 18060 22830 18116
rect 24882 18060 24892 18116
rect 24948 18060 25452 18116
rect 25508 18060 25518 18116
rect 27346 18060 27356 18116
rect 27412 18060 31724 18116
rect 31780 18060 31790 18116
rect 31892 18060 33740 18116
rect 33796 18060 34412 18116
rect 34468 18060 34478 18116
rect 34972 18060 36204 18116
rect 36260 18060 36270 18116
rect 40114 18060 40124 18116
rect 40180 18060 42140 18116
rect 42196 18060 42206 18116
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 30828 18004 30884 18060
rect 31892 18004 31948 18060
rect 1474 17948 1484 18004
rect 1540 17948 4284 18004
rect 4340 17948 4350 18004
rect 5058 17948 5068 18004
rect 5124 17948 5404 18004
rect 5460 17948 5470 18004
rect 6860 17948 12460 18004
rect 12516 17948 12526 18004
rect 14690 17948 14700 18004
rect 14756 17948 14924 18004
rect 14980 17948 14990 18004
rect 15932 17948 23548 18004
rect 23604 17948 23614 18004
rect 30818 17948 30828 18004
rect 30884 17948 30894 18004
rect 31490 17948 31500 18004
rect 31556 17948 31948 18004
rect 33058 17948 33068 18004
rect 33124 17948 33292 18004
rect 33348 17948 33358 18004
rect 15932 17892 15988 17948
rect 34972 17892 35028 18060
rect 44454 18004 44464 18060
rect 44520 18004 44568 18060
rect 44624 18004 44672 18060
rect 44728 18004 44738 18060
rect 45612 18004 45668 18284
rect 57344 18228 57456 18256
rect 45826 18172 45836 18228
rect 45892 18172 50092 18228
rect 50148 18172 50158 18228
rect 51538 18172 51548 18228
rect 51604 18172 52892 18228
rect 52948 18172 54012 18228
rect 54068 18172 54078 18228
rect 54450 18172 54460 18228
rect 54516 18172 55244 18228
rect 55300 18172 55310 18228
rect 55458 18172 55468 18228
rect 55524 18172 57456 18228
rect 57344 18144 57456 18172
rect 48850 18060 48860 18116
rect 48916 18060 53676 18116
rect 53732 18060 53742 18116
rect 35186 17948 35196 18004
rect 35252 17948 38444 18004
rect 38500 17948 38510 18004
rect 40786 17948 40796 18004
rect 40852 17948 43148 18004
rect 43204 17948 43214 18004
rect 45612 17948 47852 18004
rect 47908 17948 52276 18004
rect 52434 17948 52444 18004
rect 52500 17948 52668 18004
rect 52724 17948 52734 18004
rect 53414 17948 53452 18004
rect 53508 17948 53518 18004
rect 53676 17948 55692 18004
rect 55748 17948 55758 18004
rect 52220 17892 52276 17948
rect 53676 17892 53732 17948
rect 3602 17836 3612 17892
rect 3668 17836 5740 17892
rect 5796 17836 5806 17892
rect 6178 17836 6188 17892
rect 6244 17836 8540 17892
rect 8596 17836 8606 17892
rect 8866 17836 8876 17892
rect 8932 17836 11452 17892
rect 11508 17836 11518 17892
rect 14802 17836 14812 17892
rect 14868 17836 15932 17892
rect 15988 17836 15998 17892
rect 16146 17836 16156 17892
rect 16212 17836 18956 17892
rect 19012 17836 19022 17892
rect 19170 17836 19180 17892
rect 19236 17836 20188 17892
rect 20244 17836 20254 17892
rect 20402 17836 20412 17892
rect 20468 17836 31052 17892
rect 31108 17836 31118 17892
rect 31724 17836 34188 17892
rect 34244 17836 34254 17892
rect 34972 17836 35084 17892
rect 35140 17836 35150 17892
rect 35298 17836 35308 17892
rect 35364 17836 37100 17892
rect 37156 17836 37166 17892
rect 37314 17836 37324 17892
rect 37380 17836 37884 17892
rect 37940 17836 37950 17892
rect 38108 17836 48244 17892
rect 48738 17836 48748 17892
rect 48804 17836 50652 17892
rect 50708 17836 51996 17892
rect 52052 17836 52062 17892
rect 52220 17836 53732 17892
rect 54684 17836 55356 17892
rect 55412 17836 55422 17892
rect 56354 17836 56364 17892
rect 56420 17836 57036 17892
rect 57092 17836 57102 17892
rect 0 17780 112 17808
rect 0 17724 5628 17780
rect 5684 17724 5694 17780
rect 6290 17724 6300 17780
rect 6356 17724 12012 17780
rect 12068 17724 12796 17780
rect 12852 17724 12862 17780
rect 13010 17724 13020 17780
rect 13076 17724 16940 17780
rect 16996 17724 17006 17780
rect 17154 17724 17164 17780
rect 17220 17724 29484 17780
rect 29540 17724 29550 17780
rect 0 17696 112 17724
rect 31724 17668 31780 17836
rect 38108 17780 38164 17836
rect 32946 17724 32956 17780
rect 33012 17724 34636 17780
rect 34692 17724 34702 17780
rect 34860 17724 38164 17780
rect 38434 17724 38444 17780
rect 38500 17724 41468 17780
rect 41524 17724 41534 17780
rect 41682 17724 41692 17780
rect 41748 17724 45388 17780
rect 45444 17724 45454 17780
rect 47030 17724 47068 17780
rect 47124 17724 47134 17780
rect 34860 17668 34916 17724
rect 45388 17668 45444 17724
rect 48188 17668 48244 17836
rect 50082 17724 50092 17780
rect 50148 17724 50204 17780
rect 50260 17724 50270 17780
rect 51762 17724 51772 17780
rect 51828 17724 52332 17780
rect 52388 17724 52398 17780
rect 54684 17668 54740 17836
rect 57344 17780 57456 17808
rect 54898 17724 54908 17780
rect 54964 17724 55804 17780
rect 55860 17724 55870 17780
rect 57138 17724 57148 17780
rect 57204 17724 57456 17780
rect 57344 17696 57456 17724
rect 2118 17612 2156 17668
rect 2212 17612 2222 17668
rect 3378 17612 3388 17668
rect 3444 17612 3948 17668
rect 4004 17612 4014 17668
rect 5842 17612 5852 17668
rect 5908 17612 6972 17668
rect 7028 17612 7532 17668
rect 7588 17612 7598 17668
rect 8754 17612 8764 17668
rect 8820 17612 9100 17668
rect 9156 17612 12236 17668
rect 12292 17612 13356 17668
rect 13412 17612 13916 17668
rect 13972 17612 14476 17668
rect 14532 17612 15876 17668
rect 16034 17612 16044 17668
rect 16100 17612 20748 17668
rect 20804 17612 20814 17668
rect 21298 17612 21308 17668
rect 21364 17612 22428 17668
rect 22484 17612 22494 17668
rect 25078 17612 25116 17668
rect 25172 17612 25182 17668
rect 26226 17612 26236 17668
rect 26292 17612 27356 17668
rect 27412 17612 27422 17668
rect 30146 17612 30156 17668
rect 30212 17612 30380 17668
rect 30436 17612 30446 17668
rect 31014 17612 31052 17668
rect 31108 17612 31118 17668
rect 31714 17612 31724 17668
rect 31780 17612 31790 17668
rect 32274 17612 32284 17668
rect 32340 17612 34916 17668
rect 41010 17612 41020 17668
rect 41076 17612 44044 17668
rect 44100 17612 44110 17668
rect 45388 17612 47628 17668
rect 47684 17612 47694 17668
rect 48188 17612 51100 17668
rect 51156 17612 51166 17668
rect 52098 17612 52108 17668
rect 52164 17612 55020 17668
rect 55076 17612 55086 17668
rect 15820 17556 15876 17612
rect 1362 17500 1372 17556
rect 1428 17500 1708 17556
rect 1764 17500 1774 17556
rect 2706 17500 2716 17556
rect 2772 17500 3612 17556
rect 3668 17500 15540 17556
rect 15820 17500 16156 17556
rect 16212 17500 16222 17556
rect 21186 17500 21196 17556
rect 21252 17500 27748 17556
rect 27906 17500 27916 17556
rect 27972 17500 28028 17556
rect 28084 17500 33404 17556
rect 33460 17500 33470 17556
rect 33954 17500 33964 17556
rect 34020 17500 34412 17556
rect 34468 17500 34478 17556
rect 38994 17500 39004 17556
rect 39060 17500 47292 17556
rect 47348 17500 47358 17556
rect 47618 17500 47628 17556
rect 47684 17500 48076 17556
rect 48132 17500 48142 17556
rect 48290 17500 48300 17556
rect 48356 17500 49980 17556
rect 50036 17500 50046 17556
rect 50194 17500 50204 17556
rect 50260 17500 54684 17556
rect 54740 17500 54750 17556
rect 15484 17444 15540 17500
rect 27692 17444 27748 17500
rect 3490 17388 3500 17444
rect 3556 17388 4396 17444
rect 4452 17388 4462 17444
rect 4722 17388 4732 17444
rect 4788 17388 5068 17444
rect 5124 17388 5292 17444
rect 5348 17388 5358 17444
rect 5730 17388 5740 17444
rect 5796 17388 6188 17444
rect 6244 17388 6254 17444
rect 6748 17388 9156 17444
rect 9314 17388 9324 17444
rect 9380 17388 10668 17444
rect 10724 17388 10734 17444
rect 11004 17388 12796 17444
rect 12852 17388 15260 17444
rect 15316 17388 15326 17444
rect 15484 17388 24220 17444
rect 24276 17388 27468 17444
rect 27524 17388 27534 17444
rect 27692 17388 31500 17444
rect 31556 17388 31566 17444
rect 36306 17388 36316 17444
rect 36372 17388 37772 17444
rect 37828 17388 37838 17444
rect 38070 17388 38108 17444
rect 38164 17388 38174 17444
rect 41234 17388 41244 17444
rect 41300 17388 51436 17444
rect 51492 17388 51502 17444
rect 0 17332 112 17360
rect 6748 17332 6804 17388
rect 9100 17332 9156 17388
rect 11004 17332 11060 17388
rect 57344 17332 57456 17360
rect 0 17276 3388 17332
rect 4946 17276 4956 17332
rect 5012 17276 6804 17332
rect 6962 17276 6972 17332
rect 7028 17276 8764 17332
rect 8820 17276 8830 17332
rect 9100 17276 11060 17332
rect 11218 17276 11228 17332
rect 11284 17276 16604 17332
rect 16660 17276 18732 17332
rect 18788 17276 18798 17332
rect 18956 17276 20916 17332
rect 24770 17276 24780 17332
rect 24836 17276 43260 17332
rect 43316 17276 43326 17332
rect 45490 17276 45500 17332
rect 45556 17276 45948 17332
rect 46004 17276 47516 17332
rect 47572 17276 47582 17332
rect 48178 17276 48188 17332
rect 48244 17276 50092 17332
rect 50148 17276 50428 17332
rect 50484 17276 51548 17332
rect 51604 17276 54124 17332
rect 54180 17276 55188 17332
rect 55794 17276 55804 17332
rect 55860 17276 57456 17332
rect 0 17248 112 17276
rect 3332 17108 3388 17276
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 18956 17220 19012 17276
rect 20860 17220 20916 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 43794 17220 43804 17276
rect 43860 17220 43908 17276
rect 43964 17220 44012 17276
rect 44068 17220 44078 17276
rect 53004 17220 53060 17276
rect 55132 17220 55188 17276
rect 57344 17248 57456 17276
rect 4274 17164 4284 17220
rect 4340 17164 5964 17220
rect 6020 17164 6030 17220
rect 6514 17164 6524 17220
rect 6580 17164 7980 17220
rect 8036 17164 8046 17220
rect 10322 17164 10332 17220
rect 10388 17164 13244 17220
rect 13300 17164 13310 17220
rect 13570 17164 13580 17220
rect 13636 17164 14924 17220
rect 14980 17164 16828 17220
rect 16884 17164 16894 17220
rect 18386 17164 18396 17220
rect 18452 17164 19012 17220
rect 19282 17164 19292 17220
rect 19348 17164 20076 17220
rect 20132 17164 20142 17220
rect 20850 17164 20860 17220
rect 20916 17164 21756 17220
rect 21812 17164 21822 17220
rect 24210 17164 24220 17220
rect 24276 17164 26460 17220
rect 26516 17164 26526 17220
rect 29026 17164 29036 17220
rect 29092 17164 41020 17220
rect 41076 17164 41086 17220
rect 41458 17164 41468 17220
rect 41524 17164 42868 17220
rect 44146 17164 44156 17220
rect 44212 17164 45836 17220
rect 45892 17164 45902 17220
rect 46498 17164 46508 17220
rect 46564 17164 47404 17220
rect 47460 17164 47470 17220
rect 47618 17164 47628 17220
rect 47684 17164 52444 17220
rect 52500 17164 52510 17220
rect 52994 17164 53004 17220
rect 53060 17164 53070 17220
rect 55122 17164 55132 17220
rect 55188 17164 55198 17220
rect 20076 17108 20132 17164
rect 42812 17108 42868 17164
rect 1026 17052 1036 17108
rect 1092 17052 3220 17108
rect 3332 17052 7084 17108
rect 7140 17052 7150 17108
rect 8530 17052 8540 17108
rect 8596 17052 9716 17108
rect 3164 16996 3220 17052
rect 9660 16996 9716 17052
rect 10780 17052 15148 17108
rect 15474 17052 15484 17108
rect 15540 17052 17164 17108
rect 17220 17052 17230 17108
rect 17714 17052 17724 17108
rect 17780 17052 19516 17108
rect 19572 17052 19582 17108
rect 20076 17052 23772 17108
rect 23828 17052 28140 17108
rect 28196 17052 28206 17108
rect 29698 17052 29708 17108
rect 29764 17052 30268 17108
rect 30324 17052 30334 17108
rect 30930 17052 30940 17108
rect 30996 17052 33852 17108
rect 33908 17052 33918 17108
rect 34066 17052 34076 17108
rect 34132 17052 34412 17108
rect 34468 17052 34478 17108
rect 34850 17052 34860 17108
rect 34916 17052 35308 17108
rect 37202 17052 37212 17108
rect 37268 17052 41748 17108
rect 41906 17052 41916 17108
rect 41972 17052 42588 17108
rect 42644 17052 42654 17108
rect 42812 17052 49084 17108
rect 49140 17052 49150 17108
rect 51314 17052 51324 17108
rect 51380 17052 52444 17108
rect 52500 17052 52510 17108
rect 53554 17052 53564 17108
rect 53620 17052 54012 17108
rect 54068 17052 54078 17108
rect 242 16940 252 16996
rect 308 16940 1372 16996
rect 1428 16940 1438 16996
rect 1810 16940 1820 16996
rect 1876 16940 2716 16996
rect 2772 16940 2782 16996
rect 3164 16940 5180 16996
rect 5236 16940 5246 16996
rect 5394 16940 5404 16996
rect 5460 16940 5964 16996
rect 6020 16940 6030 16996
rect 7970 16940 7980 16996
rect 8036 16940 8988 16996
rect 9044 16940 9054 16996
rect 9650 16940 9660 16996
rect 9716 16940 10556 16996
rect 10612 16940 10622 16996
rect 0 16884 112 16912
rect 0 16828 588 16884
rect 644 16828 654 16884
rect 3154 16828 3164 16884
rect 3220 16828 7756 16884
rect 7812 16828 7822 16884
rect 8866 16828 8876 16884
rect 8932 16828 9996 16884
rect 10052 16828 10062 16884
rect 0 16800 112 16828
rect 10780 16772 10836 17052
rect 15092 16996 15148 17052
rect 35252 16996 35308 17052
rect 41692 16996 41748 17052
rect 13906 16940 13916 16996
rect 13972 16940 14980 16996
rect 15092 16940 21028 16996
rect 21298 16940 21308 16996
rect 21364 16940 24220 16996
rect 24276 16940 24286 16996
rect 25106 16940 25116 16996
rect 25172 16940 28812 16996
rect 28868 16940 28878 16996
rect 32834 16940 32844 16996
rect 32900 16940 34524 16996
rect 34580 16940 34590 16996
rect 34934 16940 34972 16996
rect 35028 16940 35038 16996
rect 35252 16940 35532 16996
rect 35588 16940 37380 16996
rect 41692 16940 44940 16996
rect 44996 16940 45006 16996
rect 45154 16940 45164 16996
rect 45220 16940 45836 16996
rect 45892 16940 45902 16996
rect 47394 16940 47404 16996
rect 47460 16940 49196 16996
rect 49252 16940 49980 16996
rect 50036 16940 50046 16996
rect 51762 16940 51772 16996
rect 51828 16940 54684 16996
rect 54740 16940 54908 16996
rect 54964 16940 54974 16996
rect 14924 16884 14980 16940
rect 14924 16828 15372 16884
rect 15428 16828 16716 16884
rect 16772 16828 16782 16884
rect 18946 16828 18956 16884
rect 19012 16828 19964 16884
rect 20020 16828 20030 16884
rect 20972 16772 21028 16940
rect 21298 16828 21308 16884
rect 21364 16828 22428 16884
rect 22484 16828 22988 16884
rect 23044 16828 23054 16884
rect 23314 16828 23324 16884
rect 23380 16828 24108 16884
rect 24164 16828 24174 16884
rect 24658 16828 24668 16884
rect 24724 16828 25228 16884
rect 25284 16828 25294 16884
rect 25750 16828 25788 16884
rect 25844 16828 28588 16884
rect 28644 16828 28654 16884
rect 31826 16828 31836 16884
rect 31892 16828 32508 16884
rect 32564 16828 32574 16884
rect 33282 16828 33292 16884
rect 33348 16828 34188 16884
rect 34244 16828 34254 16884
rect 34412 16828 35140 16884
rect 35410 16828 35420 16884
rect 35476 16828 37268 16884
rect 34412 16772 34468 16828
rect 466 16716 476 16772
rect 532 16716 588 16772
rect 644 16716 654 16772
rect 1036 16716 1260 16772
rect 1316 16716 1326 16772
rect 2258 16716 2268 16772
rect 2324 16716 2940 16772
rect 2996 16716 3006 16772
rect 3378 16716 3388 16772
rect 3444 16716 4172 16772
rect 4228 16716 4900 16772
rect 5170 16716 5180 16772
rect 5236 16716 6748 16772
rect 6804 16716 6814 16772
rect 7522 16716 7532 16772
rect 7588 16716 10836 16772
rect 11106 16716 11116 16772
rect 11172 16716 13244 16772
rect 13300 16716 13310 16772
rect 13458 16716 13468 16772
rect 13524 16716 13804 16772
rect 13860 16716 14140 16772
rect 14196 16716 14206 16772
rect 15586 16716 15596 16772
rect 15652 16716 16492 16772
rect 16548 16716 16604 16772
rect 16660 16716 16670 16772
rect 17042 16716 17052 16772
rect 17108 16716 19124 16772
rect 20972 16716 32844 16772
rect 32900 16716 32910 16772
rect 33058 16716 33068 16772
rect 33124 16716 34468 16772
rect 35084 16772 35140 16828
rect 35084 16716 36036 16772
rect 36194 16716 36204 16772
rect 36260 16716 36988 16772
rect 37044 16716 37054 16772
rect 1036 16660 1092 16716
rect 1026 16604 1036 16660
rect 1092 16604 1102 16660
rect 2146 16604 2156 16660
rect 2212 16604 4172 16660
rect 4228 16604 4238 16660
rect 4844 16548 4900 16716
rect 19068 16660 19124 16716
rect 5954 16604 5964 16660
rect 6020 16604 7084 16660
rect 7140 16604 7150 16660
rect 7410 16604 7420 16660
rect 7476 16604 7644 16660
rect 7700 16604 7710 16660
rect 11778 16604 11788 16660
rect 11844 16604 13916 16660
rect 13972 16604 13982 16660
rect 15250 16604 15260 16660
rect 15316 16604 17836 16660
rect 17892 16604 17902 16660
rect 19068 16604 21252 16660
rect 22194 16604 22204 16660
rect 22260 16604 29148 16660
rect 29204 16604 34300 16660
rect 34356 16604 34366 16660
rect 35074 16604 35084 16660
rect 35140 16604 35420 16660
rect 35476 16604 35486 16660
rect 3154 16492 3164 16548
rect 3220 16492 3724 16548
rect 3780 16492 3790 16548
rect 4050 16492 4060 16548
rect 4116 16492 4172 16548
rect 4228 16492 4238 16548
rect 4844 16492 9772 16548
rect 9828 16492 9838 16548
rect 9986 16492 9996 16548
rect 10052 16492 10668 16548
rect 10724 16492 10734 16548
rect 11330 16492 11340 16548
rect 11396 16492 13692 16548
rect 13748 16492 13758 16548
rect 20150 16492 20188 16548
rect 20244 16492 20254 16548
rect 0 16436 112 16464
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 21196 16436 21252 16604
rect 35980 16548 36036 16716
rect 37212 16660 37268 16828
rect 37324 16772 37380 16940
rect 57344 16884 57456 16912
rect 38770 16828 38780 16884
rect 38836 16828 40908 16884
rect 40964 16828 40974 16884
rect 41916 16828 45052 16884
rect 45108 16828 45118 16884
rect 45938 16828 45948 16884
rect 46004 16828 46284 16884
rect 46340 16828 46350 16884
rect 46946 16828 46956 16884
rect 47012 16828 47292 16884
rect 47348 16828 50988 16884
rect 51044 16828 51054 16884
rect 51324 16828 57456 16884
rect 41916 16772 41972 16828
rect 51324 16772 51380 16828
rect 57344 16800 57456 16828
rect 37324 16716 41972 16772
rect 42130 16716 42140 16772
rect 42196 16716 42364 16772
rect 42420 16716 42430 16772
rect 42578 16716 42588 16772
rect 42644 16716 43036 16772
rect 43092 16716 48300 16772
rect 48356 16716 48366 16772
rect 48514 16716 48524 16772
rect 48580 16716 48636 16772
rect 48692 16716 48702 16772
rect 49410 16716 49420 16772
rect 49476 16716 49532 16772
rect 49588 16716 49598 16772
rect 50194 16716 50204 16772
rect 50260 16716 51380 16772
rect 53106 16716 53116 16772
rect 53172 16716 54236 16772
rect 54292 16716 54908 16772
rect 54964 16716 54974 16772
rect 37212 16604 39228 16660
rect 39284 16604 42364 16660
rect 42420 16604 42430 16660
rect 43362 16604 43372 16660
rect 43428 16604 46620 16660
rect 46676 16604 46686 16660
rect 47394 16604 47404 16660
rect 47460 16604 50764 16660
rect 50820 16604 50830 16660
rect 52994 16604 53004 16660
rect 53060 16604 55132 16660
rect 55188 16604 55198 16660
rect 47404 16548 47460 16604
rect 21522 16492 21532 16548
rect 21588 16492 23324 16548
rect 23380 16492 23390 16548
rect 26114 16492 26124 16548
rect 26180 16492 27244 16548
rect 27300 16492 27310 16548
rect 28914 16492 28924 16548
rect 28980 16492 29484 16548
rect 29540 16492 29550 16548
rect 29698 16492 29708 16548
rect 29764 16492 31388 16548
rect 31444 16492 31454 16548
rect 31938 16492 31948 16548
rect 32004 16492 33180 16548
rect 33236 16492 33246 16548
rect 34850 16492 34860 16548
rect 34916 16492 35308 16548
rect 35364 16492 35374 16548
rect 35980 16492 39564 16548
rect 39620 16492 39630 16548
rect 39788 16492 44268 16548
rect 44324 16492 44334 16548
rect 45490 16492 45500 16548
rect 45556 16492 47460 16548
rect 47740 16492 52892 16548
rect 52948 16492 53676 16548
rect 53732 16492 53742 16548
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 39788 16436 39844 16492
rect 44454 16436 44464 16492
rect 44520 16436 44568 16492
rect 44624 16436 44672 16492
rect 44728 16436 44738 16492
rect 47740 16436 47796 16492
rect 57344 16436 57456 16464
rect 0 16380 588 16436
rect 644 16380 654 16436
rect 2930 16380 2940 16436
rect 2996 16380 3388 16436
rect 3444 16380 3454 16436
rect 3602 16380 3612 16436
rect 3668 16380 4172 16436
rect 4228 16380 4238 16436
rect 5506 16380 5516 16436
rect 5572 16380 6300 16436
rect 6356 16380 6366 16436
rect 8978 16380 8988 16436
rect 9044 16380 11004 16436
rect 11060 16380 11070 16436
rect 13794 16380 13804 16436
rect 13860 16380 14476 16436
rect 14532 16380 14542 16436
rect 14690 16380 14700 16436
rect 14756 16380 20972 16436
rect 21028 16380 21038 16436
rect 21196 16380 24108 16436
rect 24164 16380 24174 16436
rect 27010 16380 27020 16436
rect 27076 16380 30380 16436
rect 30436 16380 30446 16436
rect 31378 16380 31388 16436
rect 31444 16380 32508 16436
rect 32564 16380 32574 16436
rect 33058 16380 33068 16436
rect 33124 16380 37548 16436
rect 37604 16380 37614 16436
rect 38994 16380 39004 16436
rect 39060 16380 39844 16436
rect 41430 16380 41468 16436
rect 41524 16380 41534 16436
rect 44930 16380 44940 16436
rect 44996 16380 45612 16436
rect 45668 16380 45678 16436
rect 47170 16380 47180 16436
rect 47236 16380 47796 16436
rect 48850 16380 48860 16436
rect 48916 16380 50316 16436
rect 50372 16380 50382 16436
rect 51538 16380 51548 16436
rect 51604 16380 52108 16436
rect 52164 16380 53340 16436
rect 53396 16380 53406 16436
rect 55122 16380 55132 16436
rect 55188 16380 57456 16436
rect 0 16352 112 16380
rect 57344 16352 57456 16380
rect 1362 16268 1372 16324
rect 1428 16268 6524 16324
rect 6580 16268 6590 16324
rect 6850 16268 6860 16324
rect 6916 16268 7420 16324
rect 7476 16268 7486 16324
rect 9426 16268 9436 16324
rect 9492 16268 10332 16324
rect 10388 16268 10398 16324
rect 10546 16268 10556 16324
rect 10612 16268 17388 16324
rect 17444 16268 17454 16324
rect 19618 16268 19628 16324
rect 19684 16268 21196 16324
rect 21252 16268 21756 16324
rect 21812 16268 21822 16324
rect 22866 16268 22876 16324
rect 22932 16268 25900 16324
rect 25956 16268 26124 16324
rect 26180 16268 26190 16324
rect 26674 16268 26684 16324
rect 26740 16268 28700 16324
rect 28756 16268 28766 16324
rect 29586 16268 29596 16324
rect 29652 16268 29820 16324
rect 29876 16268 29886 16324
rect 30566 16268 30604 16324
rect 30660 16268 30670 16324
rect 32834 16268 32844 16324
rect 32900 16268 51996 16324
rect 52052 16268 52062 16324
rect 52322 16268 52332 16324
rect 52388 16268 53452 16324
rect 53508 16268 53518 16324
rect 55010 16268 55020 16324
rect 55076 16268 56028 16324
rect 56084 16268 56094 16324
rect 56354 16268 56364 16324
rect 56420 16268 56700 16324
rect 56756 16268 56766 16324
rect 1922 16156 1932 16212
rect 1988 16156 7196 16212
rect 7252 16156 7262 16212
rect 11106 16156 11116 16212
rect 11172 16156 11900 16212
rect 11956 16156 11966 16212
rect 13122 16156 13132 16212
rect 13188 16156 14700 16212
rect 14756 16156 14766 16212
rect 16034 16156 16044 16212
rect 16100 16156 16492 16212
rect 16548 16156 16558 16212
rect 18470 16156 18508 16212
rect 18564 16156 18574 16212
rect 18732 16156 23100 16212
rect 23156 16156 23166 16212
rect 23538 16156 23548 16212
rect 23604 16156 24892 16212
rect 24948 16156 24958 16212
rect 26786 16156 26796 16212
rect 18732 16100 18788 16156
rect 26852 16100 26908 16212
rect 27234 16156 27244 16212
rect 27300 16156 29932 16212
rect 29988 16156 29998 16212
rect 32386 16156 32396 16212
rect 32452 16156 32956 16212
rect 33012 16156 33022 16212
rect 33170 16156 33180 16212
rect 33236 16156 33852 16212
rect 33908 16156 33918 16212
rect 34290 16156 34300 16212
rect 34356 16156 35084 16212
rect 35140 16156 35150 16212
rect 37762 16156 37772 16212
rect 37828 16156 38332 16212
rect 38388 16156 38398 16212
rect 41346 16156 41356 16212
rect 41412 16156 45052 16212
rect 45108 16156 45118 16212
rect 45378 16156 45388 16212
rect 45444 16156 45454 16212
rect 47506 16156 47516 16212
rect 47572 16156 48972 16212
rect 49028 16156 49038 16212
rect 50194 16156 50204 16212
rect 50260 16156 50876 16212
rect 50932 16156 50942 16212
rect 51202 16156 51212 16212
rect 51268 16156 54740 16212
rect 1250 16044 1260 16100
rect 1316 16044 1820 16100
rect 1876 16044 1886 16100
rect 3602 16044 3612 16100
rect 3668 16044 4060 16100
rect 4116 16044 4126 16100
rect 4946 16044 4956 16100
rect 5012 16044 6076 16100
rect 6132 16044 6142 16100
rect 6290 16044 6300 16100
rect 6356 16044 6972 16100
rect 7028 16044 7038 16100
rect 7298 16044 7308 16100
rect 7364 16044 10108 16100
rect 10164 16044 10174 16100
rect 14018 16044 14028 16100
rect 14084 16044 16940 16100
rect 16996 16044 17006 16100
rect 17826 16044 17836 16100
rect 17892 16044 18788 16100
rect 19730 16044 19740 16100
rect 19796 16044 20524 16100
rect 20580 16044 20590 16100
rect 20962 16044 20972 16100
rect 21028 16044 21644 16100
rect 21700 16044 21710 16100
rect 22306 16044 22316 16100
rect 22372 16044 24220 16100
rect 24276 16044 24286 16100
rect 26852 16044 30604 16100
rect 30660 16044 30670 16100
rect 31042 16044 31052 16100
rect 31108 16044 32284 16100
rect 32340 16044 32350 16100
rect 32834 16044 32844 16100
rect 32900 16044 35980 16100
rect 36036 16044 36876 16100
rect 36932 16044 36942 16100
rect 37314 16044 37324 16100
rect 37380 16044 37884 16100
rect 37940 16044 37950 16100
rect 38882 16044 38892 16100
rect 38948 16044 41916 16100
rect 41972 16044 42812 16100
rect 42868 16044 44828 16100
rect 44884 16044 45164 16100
rect 45220 16044 45230 16100
rect 0 15988 112 16016
rect 10108 15988 10164 16044
rect 45388 15988 45444 16156
rect 54684 16100 54740 16156
rect 56028 16156 56252 16212
rect 56308 16156 56318 16212
rect 56028 16100 56084 16156
rect 46498 16044 46508 16100
rect 46564 16044 49196 16100
rect 49252 16044 49262 16100
rect 51426 16044 51436 16100
rect 51492 16044 52332 16100
rect 52388 16044 52398 16100
rect 54674 16044 54684 16100
rect 54740 16044 54750 16100
rect 56018 16044 56028 16100
rect 56084 16044 56094 16100
rect 57344 15988 57456 16016
rect 0 15932 9212 15988
rect 9268 15932 9278 15988
rect 10108 15932 16716 15988
rect 16772 15932 16782 15988
rect 18162 15932 18172 15988
rect 18228 15932 20412 15988
rect 20468 15932 20478 15988
rect 21298 15932 21308 15988
rect 21364 15932 23660 15988
rect 23716 15932 23726 15988
rect 24098 15932 24108 15988
rect 24164 15932 26684 15988
rect 26740 15932 26750 15988
rect 26898 15932 26908 15988
rect 26964 15932 31164 15988
rect 31220 15932 31230 15988
rect 31602 15932 31612 15988
rect 31668 15932 40236 15988
rect 40292 15932 40460 15988
rect 40516 15932 40526 15988
rect 41570 15932 41580 15988
rect 41636 15932 44380 15988
rect 44436 15932 44940 15988
rect 44996 15932 45006 15988
rect 45378 15932 45388 15988
rect 45444 15932 45454 15988
rect 45602 15932 45612 15988
rect 45668 15932 46620 15988
rect 46676 15932 46686 15988
rect 47058 15932 47068 15988
rect 47124 15932 48748 15988
rect 48804 15932 48814 15988
rect 49410 15932 49420 15988
rect 49476 15932 50092 15988
rect 50148 15932 50158 15988
rect 50642 15932 50652 15988
rect 50708 15932 57456 15988
rect 0 15904 112 15932
rect 57344 15904 57456 15932
rect 2818 15820 2828 15876
rect 2884 15820 3164 15876
rect 3220 15820 3276 15876
rect 3332 15820 3342 15876
rect 3602 15820 3612 15876
rect 3668 15820 4788 15876
rect 4946 15820 4956 15876
rect 5012 15820 10556 15876
rect 10612 15820 10622 15876
rect 12002 15820 12012 15876
rect 12068 15820 15260 15876
rect 15316 15820 15326 15876
rect 15586 15820 15596 15876
rect 15652 15820 23436 15876
rect 23492 15820 23502 15876
rect 23660 15820 25116 15876
rect 25172 15820 25182 15876
rect 27794 15820 27804 15876
rect 27860 15820 31052 15876
rect 31108 15820 31118 15876
rect 31378 15820 31388 15876
rect 31444 15820 32284 15876
rect 32340 15820 32732 15876
rect 32788 15820 32798 15876
rect 33618 15820 33628 15876
rect 33684 15820 34188 15876
rect 34244 15820 34254 15876
rect 34402 15820 34412 15876
rect 34468 15820 34972 15876
rect 35028 15820 35038 15876
rect 35746 15820 35756 15876
rect 35812 15820 50428 15876
rect 50484 15820 50494 15876
rect 50866 15820 50876 15876
rect 50932 15820 54348 15876
rect 54404 15820 54572 15876
rect 54628 15820 54638 15876
rect 4732 15764 4788 15820
rect 23660 15764 23716 15820
rect 1250 15708 1260 15764
rect 1316 15708 1932 15764
rect 1988 15708 1998 15764
rect 2258 15708 2268 15764
rect 2324 15708 3500 15764
rect 3556 15708 3566 15764
rect 4732 15708 13244 15764
rect 13300 15708 13310 15764
rect 13570 15708 13580 15764
rect 13636 15708 14252 15764
rect 14308 15708 19852 15764
rect 19908 15708 22876 15764
rect 22932 15708 22942 15764
rect 23090 15708 23100 15764
rect 23156 15708 23548 15764
rect 23604 15708 23716 15764
rect 30594 15708 30604 15764
rect 30660 15708 37100 15764
rect 37156 15708 37166 15764
rect 45052 15708 45388 15764
rect 48962 15708 48972 15764
rect 49028 15708 50764 15764
rect 50820 15708 51548 15764
rect 51604 15708 51614 15764
rect 51986 15708 51996 15764
rect 52052 15708 55244 15764
rect 55300 15708 55310 15764
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 43794 15652 43804 15708
rect 43860 15652 43908 15708
rect 43964 15652 44012 15708
rect 44068 15652 44078 15708
rect 45052 15652 45108 15708
rect 3042 15596 3052 15652
rect 3108 15596 3612 15652
rect 3668 15596 3678 15652
rect 5730 15596 5740 15652
rect 5796 15596 5964 15652
rect 6020 15596 6030 15652
rect 7074 15596 7084 15652
rect 7140 15596 7644 15652
rect 7700 15596 7710 15652
rect 8082 15596 8092 15652
rect 8148 15596 9100 15652
rect 9156 15596 9166 15652
rect 9538 15596 9548 15652
rect 9604 15596 11452 15652
rect 11508 15596 11518 15652
rect 13458 15596 13468 15652
rect 13524 15596 19292 15652
rect 19348 15596 19358 15652
rect 20860 15596 21532 15652
rect 21588 15596 21598 15652
rect 21746 15596 21756 15652
rect 21812 15596 22708 15652
rect 22978 15596 22988 15652
rect 23044 15596 23660 15652
rect 23716 15596 23726 15652
rect 29810 15596 29820 15652
rect 29876 15596 31948 15652
rect 32004 15596 32014 15652
rect 32274 15596 32284 15652
rect 32340 15596 34020 15652
rect 34178 15596 34188 15652
rect 34244 15596 37436 15652
rect 37492 15596 37502 15652
rect 40226 15596 40236 15652
rect 40292 15596 43372 15652
rect 43428 15596 43438 15652
rect 44930 15596 44940 15652
rect 44996 15596 45108 15652
rect 45332 15652 45388 15708
rect 45332 15596 48188 15652
rect 48244 15596 48916 15652
rect 0 15540 112 15568
rect 20860 15540 20916 15596
rect 22652 15540 22708 15596
rect 33964 15540 34020 15596
rect 48860 15540 48916 15596
rect 57344 15540 57456 15568
rect 0 15484 4004 15540
rect 4134 15484 4172 15540
rect 4228 15484 4238 15540
rect 5292 15484 8652 15540
rect 8708 15484 8718 15540
rect 9314 15484 9324 15540
rect 9380 15484 10108 15540
rect 10164 15484 13580 15540
rect 13636 15484 13646 15540
rect 14354 15484 14364 15540
rect 14420 15484 17052 15540
rect 17108 15484 17118 15540
rect 17724 15484 20916 15540
rect 21270 15484 21308 15540
rect 21364 15484 21374 15540
rect 21858 15484 21868 15540
rect 21924 15484 22428 15540
rect 22484 15484 22494 15540
rect 22652 15484 33180 15540
rect 33236 15484 33246 15540
rect 33964 15484 37548 15540
rect 37604 15484 37614 15540
rect 37986 15484 37996 15540
rect 38052 15484 38108 15540
rect 38164 15484 38174 15540
rect 41122 15484 41132 15540
rect 41188 15484 43708 15540
rect 43764 15484 45388 15540
rect 45444 15484 45454 15540
rect 46834 15484 46844 15540
rect 46900 15484 48300 15540
rect 48356 15484 48636 15540
rect 48692 15484 48702 15540
rect 48860 15484 49644 15540
rect 49700 15484 49710 15540
rect 50530 15484 50540 15540
rect 50596 15484 52108 15540
rect 52164 15484 52174 15540
rect 52994 15484 53004 15540
rect 53060 15484 53676 15540
rect 53732 15484 54572 15540
rect 54628 15484 54638 15540
rect 55346 15484 55356 15540
rect 55412 15484 56140 15540
rect 56196 15484 56206 15540
rect 56588 15484 57456 15540
rect 0 15456 112 15484
rect 3948 15428 4004 15484
rect 5292 15428 5348 15484
rect 2706 15372 2716 15428
rect 2772 15372 3052 15428
rect 3108 15372 3118 15428
rect 3948 15372 5348 15428
rect 5506 15372 5516 15428
rect 5572 15372 6524 15428
rect 6580 15372 6590 15428
rect 7196 15372 9996 15428
rect 10052 15372 10062 15428
rect 10210 15372 10220 15428
rect 10276 15372 10556 15428
rect 10612 15372 10622 15428
rect 12338 15372 12348 15428
rect 12404 15372 13636 15428
rect 7196 15316 7252 15372
rect 13580 15316 13636 15372
rect 1922 15260 1932 15316
rect 1988 15260 2492 15316
rect 2548 15260 2558 15316
rect 3154 15260 3164 15316
rect 3220 15260 3612 15316
rect 3668 15260 3678 15316
rect 5142 15260 5180 15316
rect 5236 15260 5246 15316
rect 6626 15260 6636 15316
rect 6692 15260 7252 15316
rect 8978 15260 8988 15316
rect 9044 15260 12908 15316
rect 12964 15260 12974 15316
rect 13570 15260 13580 15316
rect 13636 15260 13646 15316
rect 16482 15260 16492 15316
rect 16548 15260 17164 15316
rect 17220 15260 17230 15316
rect 17724 15204 17780 15484
rect 37548 15428 37604 15484
rect 56588 15428 56644 15484
rect 57344 15456 57456 15484
rect 18946 15372 18956 15428
rect 19012 15372 36540 15428
rect 36596 15372 36606 15428
rect 37548 15372 38444 15428
rect 38500 15372 38510 15428
rect 41794 15372 41804 15428
rect 41860 15372 43148 15428
rect 43204 15372 43214 15428
rect 43586 15372 43596 15428
rect 43652 15372 44268 15428
rect 44324 15372 46508 15428
rect 46564 15372 46574 15428
rect 46722 15372 46732 15428
rect 46788 15372 46956 15428
rect 47012 15372 47022 15428
rect 47730 15372 47740 15428
rect 47796 15372 48692 15428
rect 48850 15372 48860 15428
rect 48916 15372 53676 15428
rect 53732 15372 53742 15428
rect 55346 15372 55356 15428
rect 55412 15372 56644 15428
rect 48636 15316 48692 15372
rect 17948 15260 18172 15316
rect 18228 15260 18238 15316
rect 19282 15260 19292 15316
rect 19348 15260 31500 15316
rect 31556 15260 31566 15316
rect 31714 15260 31724 15316
rect 31780 15260 32284 15316
rect 32340 15260 32350 15316
rect 32834 15260 32844 15316
rect 32900 15260 33516 15316
rect 33572 15260 37548 15316
rect 37604 15260 37614 15316
rect 38210 15260 38220 15316
rect 38276 15260 38286 15316
rect 38434 15260 38444 15316
rect 38500 15260 40460 15316
rect 40516 15260 40526 15316
rect 40674 15260 40684 15316
rect 40740 15260 41916 15316
rect 41972 15260 41982 15316
rect 42354 15260 42364 15316
rect 42420 15260 44156 15316
rect 44212 15260 44222 15316
rect 44930 15260 44940 15316
rect 44996 15260 45164 15316
rect 45220 15260 45230 15316
rect 45378 15260 45388 15316
rect 45444 15260 45482 15316
rect 47170 15260 47180 15316
rect 47236 15260 48188 15316
rect 48244 15260 48254 15316
rect 48636 15260 48972 15316
rect 49028 15260 49038 15316
rect 49382 15260 49420 15316
rect 49476 15260 49486 15316
rect 49634 15260 49644 15316
rect 49700 15260 53340 15316
rect 53396 15260 53406 15316
rect 17948 15204 18004 15260
rect 38220 15204 38276 15260
rect 1474 15148 1484 15204
rect 1540 15148 3948 15204
rect 4004 15148 4014 15204
rect 4274 15148 4284 15204
rect 4340 15148 4956 15204
rect 5012 15148 5022 15204
rect 5282 15148 5292 15204
rect 5348 15148 9660 15204
rect 9716 15148 9726 15204
rect 9986 15148 9996 15204
rect 10052 15148 10892 15204
rect 10948 15148 10958 15204
rect 12114 15148 12124 15204
rect 12180 15148 14364 15204
rect 14420 15148 14430 15204
rect 14914 15148 14924 15204
rect 14980 15148 15372 15204
rect 15428 15148 15438 15204
rect 16146 15148 16156 15204
rect 16212 15148 16604 15204
rect 16660 15148 17780 15204
rect 17938 15148 17948 15204
rect 18004 15148 21084 15204
rect 21140 15148 23212 15204
rect 23268 15148 23278 15204
rect 24210 15148 24220 15204
rect 24276 15148 27244 15204
rect 27300 15148 27310 15204
rect 30258 15148 30268 15204
rect 30324 15148 31612 15204
rect 31668 15148 31678 15204
rect 33730 15148 33740 15204
rect 33796 15148 34748 15204
rect 34804 15148 34814 15204
rect 37090 15148 37100 15204
rect 37156 15148 38276 15204
rect 38434 15148 38444 15204
rect 38500 15148 38780 15204
rect 38836 15148 38846 15204
rect 39554 15148 39564 15204
rect 39620 15148 43036 15204
rect 43092 15148 43102 15204
rect 43820 15148 46172 15204
rect 46228 15148 46238 15204
rect 46946 15148 46956 15204
rect 47012 15148 50204 15204
rect 50260 15148 50270 15204
rect 53554 15148 53564 15204
rect 53620 15148 54908 15204
rect 54964 15148 54974 15204
rect 0 15092 112 15120
rect 43820 15092 43876 15148
rect 57344 15092 57456 15120
rect 0 15036 5012 15092
rect 5618 15036 5628 15092
rect 5684 15036 6748 15092
rect 6804 15036 6814 15092
rect 6962 15036 6972 15092
rect 7028 15036 9436 15092
rect 9492 15036 9502 15092
rect 9762 15036 9772 15092
rect 9828 15036 35756 15092
rect 35812 15036 35822 15092
rect 35970 15036 35980 15092
rect 36036 15036 41188 15092
rect 41346 15036 41356 15092
rect 41412 15036 43876 15092
rect 44034 15036 44044 15092
rect 44100 15036 44268 15092
rect 44324 15036 44334 15092
rect 44706 15036 44716 15092
rect 44772 15036 44940 15092
rect 44996 15036 45006 15092
rect 47506 15036 47516 15092
rect 47572 15036 48860 15092
rect 48916 15036 48926 15092
rect 49858 15036 49868 15092
rect 49924 15036 57456 15092
rect 0 15008 112 15036
rect 4956 14980 5012 15036
rect 41132 14980 41188 15036
rect 57344 15008 57456 15036
rect 2930 14924 2940 14980
rect 2996 14924 4060 14980
rect 4116 14924 4126 14980
rect 4946 14924 4956 14980
rect 5012 14924 5022 14980
rect 5282 14924 5292 14980
rect 5348 14924 6076 14980
rect 6132 14924 6142 14980
rect 6822 14924 6860 14980
rect 6916 14924 6926 14980
rect 7074 14924 7084 14980
rect 7140 14924 12348 14980
rect 12404 14924 12740 14980
rect 12898 14924 12908 14980
rect 12964 14924 14924 14980
rect 14980 14924 17164 14980
rect 17220 14924 17230 14980
rect 17490 14924 17500 14980
rect 17556 14924 22428 14980
rect 22484 14924 22494 14980
rect 29362 14924 29372 14980
rect 29428 14924 32844 14980
rect 32900 14924 32910 14980
rect 37538 14924 37548 14980
rect 37604 14924 39340 14980
rect 39396 14924 39406 14980
rect 41132 14924 44324 14980
rect 44930 14924 44940 14980
rect 44996 14924 46620 14980
rect 46676 14924 46686 14980
rect 47618 14924 47628 14980
rect 47684 14924 47852 14980
rect 47908 14924 47918 14980
rect 48626 14924 48636 14980
rect 48692 14924 49532 14980
rect 49588 14924 49598 14980
rect 52770 14924 52780 14980
rect 52836 14924 52846 14980
rect 52994 14924 53004 14980
rect 53060 14924 53676 14980
rect 53732 14924 53742 14980
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 12684 14868 12740 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 5058 14812 5068 14868
rect 5124 14812 8092 14868
rect 8148 14812 12124 14868
rect 12180 14812 12190 14868
rect 12684 14812 13244 14868
rect 13300 14812 13310 14868
rect 14130 14812 14140 14868
rect 14196 14812 15372 14868
rect 15428 14812 15438 14868
rect 15596 14812 18956 14868
rect 19012 14812 19022 14868
rect 19730 14812 19740 14868
rect 19796 14812 20076 14868
rect 20132 14812 20142 14868
rect 20962 14812 20972 14868
rect 21028 14812 21756 14868
rect 21812 14812 21822 14868
rect 24892 14812 30268 14868
rect 30324 14812 30334 14868
rect 30930 14812 30940 14868
rect 30996 14812 31164 14868
rect 31220 14812 31230 14868
rect 32722 14812 32732 14868
rect 32788 14812 36092 14868
rect 36148 14812 36158 14868
rect 38770 14812 38780 14868
rect 38836 14812 41020 14868
rect 41076 14812 41086 14868
rect 42466 14812 42476 14868
rect 42532 14812 42700 14868
rect 42756 14812 42766 14868
rect 15596 14756 15652 14812
rect 24892 14756 24948 14812
rect 44268 14756 44324 14924
rect 44454 14868 44464 14924
rect 44520 14868 44568 14924
rect 44624 14868 44672 14924
rect 44728 14868 44738 14924
rect 52780 14868 52836 14924
rect 45154 14812 45164 14868
rect 45220 14812 45948 14868
rect 46004 14812 46014 14868
rect 46162 14812 46172 14868
rect 46228 14812 47180 14868
rect 47236 14812 47246 14868
rect 47618 14812 47628 14868
rect 47684 14812 48748 14868
rect 48804 14812 48814 14868
rect 49522 14812 49532 14868
rect 49588 14812 50204 14868
rect 50260 14812 50270 14868
rect 51426 14812 51436 14868
rect 51492 14812 52556 14868
rect 52612 14812 52622 14868
rect 52780 14812 55580 14868
rect 55636 14812 55646 14868
rect 2370 14700 2380 14756
rect 2436 14700 3276 14756
rect 3332 14700 3342 14756
rect 4610 14700 4620 14756
rect 4676 14700 5180 14756
rect 5236 14700 5246 14756
rect 5730 14700 5740 14756
rect 5796 14700 6748 14756
rect 6804 14700 6814 14756
rect 8642 14700 8652 14756
rect 8708 14700 8876 14756
rect 8932 14700 8942 14756
rect 12786 14700 12796 14756
rect 12852 14700 15036 14756
rect 15092 14700 15652 14756
rect 15810 14700 15820 14756
rect 15876 14700 24948 14756
rect 29334 14700 29372 14756
rect 29428 14700 29438 14756
rect 29586 14700 29596 14756
rect 29652 14700 41356 14756
rect 41412 14700 41422 14756
rect 41906 14700 41916 14756
rect 41972 14700 44044 14756
rect 44100 14700 44110 14756
rect 44268 14700 47516 14756
rect 47572 14700 47582 14756
rect 48066 14700 48076 14756
rect 48132 14700 48188 14756
rect 48244 14700 48254 14756
rect 48486 14700 48524 14756
rect 48580 14700 48590 14756
rect 48962 14700 48972 14756
rect 49028 14700 50876 14756
rect 50932 14700 51660 14756
rect 51716 14700 51726 14756
rect 51986 14700 51996 14756
rect 52052 14700 53340 14756
rect 53396 14700 53406 14756
rect 56018 14700 56028 14756
rect 56084 14700 56588 14756
rect 56644 14700 56654 14756
rect 0 14644 112 14672
rect 57344 14644 57456 14672
rect 0 14588 700 14644
rect 756 14588 766 14644
rect 1810 14588 1820 14644
rect 1876 14588 2268 14644
rect 2324 14588 2334 14644
rect 2482 14588 2492 14644
rect 2548 14588 6076 14644
rect 6132 14588 6142 14644
rect 6626 14588 6636 14644
rect 6692 14588 7196 14644
rect 7252 14588 7262 14644
rect 7858 14588 7868 14644
rect 7924 14588 8428 14644
rect 8484 14588 9884 14644
rect 9940 14588 12572 14644
rect 12628 14588 12638 14644
rect 13794 14588 13804 14644
rect 13860 14588 49532 14644
rect 49588 14588 49598 14644
rect 49756 14588 54124 14644
rect 54180 14588 54460 14644
rect 54516 14588 54526 14644
rect 57026 14588 57036 14644
rect 57092 14588 57456 14644
rect 0 14560 112 14588
rect 49756 14532 49812 14588
rect 57344 14560 57456 14588
rect 1138 14476 1148 14532
rect 1204 14476 1596 14532
rect 1652 14476 4956 14532
rect 5012 14476 5022 14532
rect 5394 14476 5404 14532
rect 5460 14476 5628 14532
rect 5684 14476 5694 14532
rect 5842 14476 5852 14532
rect 5908 14476 6300 14532
rect 6356 14476 6366 14532
rect 6738 14476 6748 14532
rect 6804 14476 11004 14532
rect 11060 14476 11788 14532
rect 12114 14476 12124 14532
rect 12180 14476 12236 14532
rect 12292 14476 12302 14532
rect 12562 14476 12572 14532
rect 12628 14476 12908 14532
rect 12964 14476 13692 14532
rect 13748 14476 13758 14532
rect 17714 14476 17724 14532
rect 17780 14476 17836 14532
rect 17892 14476 17902 14532
rect 18162 14476 18172 14532
rect 18228 14476 18396 14532
rect 18452 14476 18462 14532
rect 18946 14476 18956 14532
rect 19012 14476 20636 14532
rect 20692 14476 20702 14532
rect 21298 14476 21308 14532
rect 21364 14476 22316 14532
rect 22372 14476 22382 14532
rect 24108 14476 24220 14532
rect 24276 14476 24286 14532
rect 25106 14476 25116 14532
rect 25172 14476 25676 14532
rect 25732 14476 25742 14532
rect 27234 14476 27244 14532
rect 27300 14476 31164 14532
rect 31220 14476 31612 14532
rect 31668 14476 31678 14532
rect 33954 14476 33964 14532
rect 34020 14476 34860 14532
rect 34916 14476 34926 14532
rect 35522 14476 35532 14532
rect 35588 14476 41580 14532
rect 41636 14476 41646 14532
rect 43026 14476 43036 14532
rect 43092 14476 43148 14532
rect 43204 14476 43932 14532
rect 43988 14476 43998 14532
rect 44930 14476 44940 14532
rect 44996 14476 45724 14532
rect 45780 14476 45790 14532
rect 46134 14476 46172 14532
rect 46228 14476 49812 14532
rect 52658 14476 52668 14532
rect 52724 14476 52892 14532
rect 52948 14476 52958 14532
rect 56364 14476 56588 14532
rect 56644 14476 56654 14532
rect 11732 14420 11788 14476
rect 24108 14420 24164 14476
rect 56364 14420 56420 14476
rect 354 14364 364 14420
rect 420 14364 1036 14420
rect 1092 14364 2156 14420
rect 2212 14364 2222 14420
rect 3612 14364 9548 14420
rect 9604 14364 9614 14420
rect 11732 14364 12964 14420
rect 13234 14364 13244 14420
rect 13300 14364 14364 14420
rect 14420 14364 15708 14420
rect 15764 14364 15774 14420
rect 17714 14364 17724 14420
rect 17780 14364 22092 14420
rect 22148 14364 24164 14420
rect 24322 14364 24332 14420
rect 24388 14364 25900 14420
rect 25956 14364 25966 14420
rect 26124 14364 27244 14420
rect 27300 14364 27310 14420
rect 28578 14364 28588 14420
rect 28644 14364 29036 14420
rect 29092 14364 29102 14420
rect 30258 14364 30268 14420
rect 30324 14364 38668 14420
rect 39330 14364 39340 14420
rect 39396 14364 42028 14420
rect 42084 14364 42094 14420
rect 43586 14364 43596 14420
rect 43652 14364 46060 14420
rect 46116 14364 46126 14420
rect 47394 14364 47404 14420
rect 47460 14364 47964 14420
rect 48020 14364 48030 14420
rect 48402 14364 48412 14420
rect 48468 14364 48972 14420
rect 49028 14364 49038 14420
rect 50082 14364 50092 14420
rect 50148 14364 50428 14420
rect 50484 14364 50494 14420
rect 51772 14364 53788 14420
rect 53844 14364 53854 14420
rect 56354 14364 56364 14420
rect 56420 14364 56430 14420
rect 0 14196 112 14224
rect 3612 14196 3668 14364
rect 12908 14308 12964 14364
rect 3826 14252 3836 14308
rect 3892 14252 4844 14308
rect 4900 14252 4910 14308
rect 5170 14252 5180 14308
rect 5236 14252 6076 14308
rect 6132 14252 7084 14308
rect 7140 14252 7150 14308
rect 7308 14252 12572 14308
rect 12628 14252 12638 14308
rect 12908 14252 16380 14308
rect 16436 14252 16446 14308
rect 16604 14252 18956 14308
rect 19012 14252 19022 14308
rect 19842 14252 19852 14308
rect 19908 14252 25228 14308
rect 25284 14252 25294 14308
rect 7308 14196 7364 14252
rect 16604 14196 16660 14252
rect 26124 14196 26180 14364
rect 38612 14308 38668 14364
rect 29138 14252 29148 14308
rect 29204 14252 29484 14308
rect 29540 14252 29550 14308
rect 30034 14252 30044 14308
rect 30100 14252 32844 14308
rect 32900 14252 32910 14308
rect 33842 14252 33852 14308
rect 33908 14252 34972 14308
rect 35028 14252 35420 14308
rect 35476 14252 35486 14308
rect 37090 14252 37100 14308
rect 37156 14252 37996 14308
rect 38052 14252 38062 14308
rect 38612 14252 39788 14308
rect 39844 14252 39854 14308
rect 40012 14252 51436 14308
rect 51492 14252 51502 14308
rect 40012 14196 40068 14252
rect 0 14140 3668 14196
rect 4722 14140 4732 14196
rect 4788 14140 7364 14196
rect 13570 14140 13580 14196
rect 13636 14140 15036 14196
rect 15092 14140 16660 14196
rect 17490 14140 17500 14196
rect 17556 14140 21532 14196
rect 21588 14140 21598 14196
rect 24210 14140 24220 14196
rect 24276 14140 26180 14196
rect 26236 14140 27020 14196
rect 27076 14140 27086 14196
rect 27346 14140 27356 14196
rect 27412 14140 28924 14196
rect 28980 14140 28990 14196
rect 31826 14140 31836 14196
rect 31892 14140 40068 14196
rect 40562 14140 40572 14196
rect 40628 14140 41804 14196
rect 41860 14140 41870 14196
rect 43026 14140 43036 14196
rect 43092 14140 43484 14196
rect 43540 14140 43550 14196
rect 44818 14140 44828 14196
rect 44884 14140 47404 14196
rect 47460 14140 47470 14196
rect 47954 14140 47964 14196
rect 48020 14140 49196 14196
rect 49252 14140 49262 14196
rect 0 14112 112 14140
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 26236 14084 26292 14140
rect 43794 14084 43804 14140
rect 43860 14084 43908 14140
rect 43964 14084 44012 14140
rect 44068 14084 44078 14140
rect 51772 14084 51828 14364
rect 56130 14252 56140 14308
rect 56196 14252 56812 14308
rect 56868 14252 56878 14308
rect 57344 14196 57456 14224
rect 52098 14140 52108 14196
rect 52164 14140 54572 14196
rect 54628 14140 54638 14196
rect 57250 14140 57260 14196
rect 57316 14140 57456 14196
rect 57344 14112 57456 14140
rect 2146 14028 2156 14084
rect 2212 14028 2716 14084
rect 2772 14028 3052 14084
rect 3108 14028 3118 14084
rect 4162 14028 4172 14084
rect 4228 14028 5180 14084
rect 5236 14028 5246 14084
rect 5394 14028 5404 14084
rect 5460 14028 8316 14084
rect 8372 14028 8382 14084
rect 9212 14028 17780 14084
rect 19506 14028 19516 14084
rect 19572 14028 20972 14084
rect 21028 14028 21038 14084
rect 24882 14028 24892 14084
rect 24948 14028 26292 14084
rect 26450 14028 26460 14084
rect 26516 14028 29260 14084
rect 29316 14028 29326 14084
rect 30258 14028 30268 14084
rect 30324 14028 32844 14084
rect 32900 14028 33292 14084
rect 33348 14028 33358 14084
rect 35298 14028 35308 14084
rect 35364 14028 38220 14084
rect 38276 14028 38286 14084
rect 38658 14028 38668 14084
rect 38724 14028 43596 14084
rect 43652 14028 43662 14084
rect 44146 14028 44156 14084
rect 44212 14028 44940 14084
rect 44996 14028 45006 14084
rect 46386 14028 46396 14084
rect 46452 14028 51828 14084
rect 53106 14028 53116 14084
rect 53172 14028 53676 14084
rect 53732 14028 53742 14084
rect 130 13916 140 13972
rect 196 13916 3164 13972
rect 3220 13916 3500 13972
rect 3556 13916 3566 13972
rect 4946 13916 4956 13972
rect 5012 13916 7868 13972
rect 7924 13916 7934 13972
rect 9212 13860 9268 14028
rect 17724 13972 17780 14028
rect 9650 13916 9660 13972
rect 9716 13916 9996 13972
rect 10052 13916 10062 13972
rect 10210 13916 10220 13972
rect 10276 13916 11228 13972
rect 11284 13916 11294 13972
rect 12114 13916 12124 13972
rect 12180 13916 13020 13972
rect 13076 13916 13086 13972
rect 13542 13916 13580 13972
rect 13636 13916 13646 13972
rect 14924 13916 15596 13972
rect 15652 13916 15662 13972
rect 16818 13916 16828 13972
rect 16884 13916 17388 13972
rect 17444 13916 17454 13972
rect 17724 13916 39620 13972
rect 39778 13916 39788 13972
rect 39844 13916 42924 13972
rect 42980 13916 42990 13972
rect 43138 13916 43148 13972
rect 43204 13916 45500 13972
rect 45556 13916 45566 13972
rect 47954 13916 47964 13972
rect 48020 13916 48524 13972
rect 48580 13916 48590 13972
rect 48850 13916 48860 13972
rect 48916 13916 49532 13972
rect 49588 13916 49598 13972
rect 51874 13916 51884 13972
rect 51940 13916 55692 13972
rect 55748 13916 55758 13972
rect 14924 13860 14980 13916
rect 39564 13860 39620 13916
rect 1698 13804 1708 13860
rect 1764 13804 9268 13860
rect 10108 13804 11228 13860
rect 11284 13804 14980 13860
rect 15092 13804 31836 13860
rect 31892 13804 31902 13860
rect 32162 13804 32172 13860
rect 32228 13804 32284 13860
rect 32340 13804 32350 13860
rect 32946 13804 32956 13860
rect 33012 13804 33180 13860
rect 33236 13804 33246 13860
rect 37538 13804 37548 13860
rect 37604 13804 38892 13860
rect 38948 13804 38958 13860
rect 39564 13804 43372 13860
rect 43428 13804 43438 13860
rect 43698 13804 43708 13860
rect 43764 13804 46172 13860
rect 46228 13804 46238 13860
rect 46396 13804 48860 13860
rect 48916 13804 48926 13860
rect 51986 13804 51996 13860
rect 52052 13804 53116 13860
rect 53172 13804 53182 13860
rect 0 13748 112 13776
rect 10108 13748 10164 13804
rect 0 13692 3388 13748
rect 3490 13692 3500 13748
rect 3556 13692 6188 13748
rect 6244 13692 6254 13748
rect 6738 13692 6748 13748
rect 6804 13692 6916 13748
rect 7074 13692 7084 13748
rect 7140 13692 7420 13748
rect 7476 13692 7486 13748
rect 8194 13692 8204 13748
rect 8260 13692 10164 13748
rect 10406 13692 10444 13748
rect 10500 13692 10510 13748
rect 10966 13692 11004 13748
rect 11060 13692 11070 13748
rect 11218 13692 11228 13748
rect 11284 13692 13356 13748
rect 13412 13692 13422 13748
rect 13570 13692 13580 13748
rect 13636 13692 14700 13748
rect 14756 13692 14766 13748
rect 0 13664 112 13692
rect 3332 13636 3388 13692
rect 6860 13636 6916 13692
rect 15092 13636 15148 13804
rect 46396 13748 46452 13804
rect 57344 13748 57456 13776
rect 17602 13692 17612 13748
rect 17668 13692 19740 13748
rect 19796 13692 19806 13748
rect 20850 13692 20860 13748
rect 20916 13692 21420 13748
rect 21476 13692 21486 13748
rect 21858 13692 21868 13748
rect 21924 13692 24892 13748
rect 24948 13692 24958 13748
rect 25218 13692 25228 13748
rect 25284 13692 33068 13748
rect 33124 13692 33134 13748
rect 33282 13692 33292 13748
rect 33348 13692 39564 13748
rect 39620 13692 39630 13748
rect 40898 13692 40908 13748
rect 40964 13692 41580 13748
rect 41636 13692 41646 13748
rect 43138 13692 43148 13748
rect 43204 13692 44492 13748
rect 44548 13692 44558 13748
rect 44706 13692 44716 13748
rect 44772 13692 46452 13748
rect 47170 13692 47180 13748
rect 47236 13692 49308 13748
rect 49364 13692 49374 13748
rect 49746 13692 49756 13748
rect 49812 13692 57456 13748
rect 57344 13664 57456 13692
rect 3332 13580 4732 13636
rect 4788 13580 4798 13636
rect 5068 13580 6636 13636
rect 6692 13580 6702 13636
rect 6860 13580 15148 13636
rect 15362 13580 15372 13636
rect 15428 13580 17948 13636
rect 18004 13580 18014 13636
rect 19282 13580 19292 13636
rect 19348 13580 23100 13636
rect 23156 13580 23166 13636
rect 23650 13580 23660 13636
rect 23716 13580 25732 13636
rect 25890 13580 25900 13636
rect 25956 13580 26236 13636
rect 26292 13580 26302 13636
rect 29250 13580 29260 13636
rect 29316 13580 29484 13636
rect 29540 13580 29550 13636
rect 32050 13580 32060 13636
rect 32116 13580 33292 13636
rect 33348 13580 34244 13636
rect 34374 13580 34412 13636
rect 34468 13580 34478 13636
rect 34626 13580 34636 13636
rect 34692 13580 36316 13636
rect 36372 13580 36382 13636
rect 36754 13580 36764 13636
rect 36820 13580 37380 13636
rect 37958 13580 37996 13636
rect 38052 13580 38556 13636
rect 38612 13580 38622 13636
rect 41458 13580 41468 13636
rect 41524 13580 43372 13636
rect 43428 13580 44940 13636
rect 44996 13580 45006 13636
rect 47282 13580 47292 13636
rect 47348 13580 47852 13636
rect 47908 13580 47918 13636
rect 48514 13580 48524 13636
rect 48580 13580 50764 13636
rect 50820 13580 50830 13636
rect 52518 13580 52556 13636
rect 52612 13580 52622 13636
rect 52994 13580 53004 13636
rect 53060 13580 54348 13636
rect 54404 13580 54414 13636
rect 5068 13524 5124 13580
rect 25676 13524 25732 13580
rect 34188 13524 34244 13580
rect 37324 13524 37380 13580
rect 1362 13468 1372 13524
rect 1428 13468 2604 13524
rect 2660 13468 2670 13524
rect 3014 13468 3052 13524
rect 3108 13468 5124 13524
rect 5282 13468 5292 13524
rect 5348 13468 5516 13524
rect 5572 13468 5582 13524
rect 6150 13468 6188 13524
rect 6244 13468 6254 13524
rect 6402 13468 6412 13524
rect 6468 13468 8428 13524
rect 8484 13468 8494 13524
rect 9538 13468 9548 13524
rect 9604 13468 11116 13524
rect 11172 13468 11182 13524
rect 15138 13468 15148 13524
rect 15204 13468 16156 13524
rect 16212 13468 16222 13524
rect 18498 13468 18508 13524
rect 18564 13468 19068 13524
rect 19124 13468 19134 13524
rect 19730 13468 19740 13524
rect 19796 13468 20748 13524
rect 20804 13468 20814 13524
rect 21074 13468 21084 13524
rect 21140 13468 22092 13524
rect 22148 13468 22158 13524
rect 22418 13468 22428 13524
rect 22484 13468 25452 13524
rect 25508 13468 25518 13524
rect 25676 13468 26124 13524
rect 26180 13468 26190 13524
rect 28242 13468 28252 13524
rect 28308 13468 32172 13524
rect 32228 13468 32238 13524
rect 34188 13468 37100 13524
rect 37156 13468 37166 13524
rect 37324 13468 40460 13524
rect 40516 13468 40526 13524
rect 42354 13468 42364 13524
rect 42420 13468 43596 13524
rect 43652 13468 43662 13524
rect 43820 13468 44044 13524
rect 44100 13468 44110 13524
rect 44268 13468 44884 13524
rect 45154 13468 45164 13524
rect 45220 13468 48412 13524
rect 48468 13468 48478 13524
rect 49606 13468 49644 13524
rect 49700 13468 49710 13524
rect 50876 13468 53452 13524
rect 53508 13468 53518 13524
rect 55122 13468 55132 13524
rect 55188 13468 56140 13524
rect 56196 13468 56206 13524
rect 5068 13412 5124 13468
rect 43820 13412 43876 13468
rect 5058 13356 5068 13412
rect 5124 13356 5134 13412
rect 5618 13356 5628 13412
rect 5684 13356 6748 13412
rect 6804 13356 6814 13412
rect 7186 13356 7196 13412
rect 7252 13356 24388 13412
rect 24892 13356 25788 13412
rect 25844 13356 28140 13412
rect 28196 13356 34860 13412
rect 34916 13356 34926 13412
rect 36530 13356 36540 13412
rect 36596 13356 39116 13412
rect 39172 13356 39182 13412
rect 43362 13356 43372 13412
rect 43428 13356 43876 13412
rect 0 13300 112 13328
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 0 13244 2380 13300
rect 2436 13244 2446 13300
rect 4956 13244 6412 13300
rect 6468 13244 6478 13300
rect 6626 13244 6636 13300
rect 6692 13244 8316 13300
rect 8372 13244 8382 13300
rect 9426 13244 9436 13300
rect 9492 13244 11004 13300
rect 11060 13244 11564 13300
rect 11620 13244 11630 13300
rect 14914 13244 14924 13300
rect 14980 13244 15372 13300
rect 15428 13244 15438 13300
rect 16594 13244 16604 13300
rect 16660 13244 17836 13300
rect 17892 13244 18060 13300
rect 18116 13244 23548 13300
rect 23604 13244 23660 13300
rect 23716 13244 23726 13300
rect 0 13216 112 13244
rect 4956 13188 5012 13244
rect 24332 13188 24388 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 24892 13188 24948 13356
rect 44268 13300 44324 13468
rect 44828 13412 44884 13468
rect 50876 13412 50932 13468
rect 44828 13356 50204 13412
rect 50260 13356 50270 13412
rect 50866 13356 50876 13412
rect 50932 13356 50942 13412
rect 52098 13356 52108 13412
rect 52164 13356 52220 13412
rect 52276 13356 52286 13412
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 57344 13300 57456 13328
rect 29922 13244 29932 13300
rect 29988 13244 35532 13300
rect 35588 13244 35598 13300
rect 37314 13244 37324 13300
rect 37380 13244 37548 13300
rect 37604 13244 44324 13300
rect 44930 13244 44940 13300
rect 44996 13244 48300 13300
rect 48356 13244 48366 13300
rect 48514 13244 48524 13300
rect 48580 13244 48972 13300
rect 49028 13244 49038 13300
rect 49186 13244 49196 13300
rect 49252 13244 54124 13300
rect 54180 13244 54190 13300
rect 54898 13244 54908 13300
rect 54964 13244 57456 13300
rect 57344 13216 57456 13244
rect 2258 13132 2268 13188
rect 2324 13132 3052 13188
rect 3108 13132 3276 13188
rect 3332 13132 3342 13188
rect 3938 13132 3948 13188
rect 4004 13132 5012 13188
rect 5068 13132 6972 13188
rect 7028 13132 7038 13188
rect 7718 13132 7756 13188
rect 7812 13132 10220 13188
rect 10276 13132 10286 13188
rect 10546 13132 10556 13188
rect 10612 13132 11340 13188
rect 11396 13132 11406 13188
rect 12450 13132 12460 13188
rect 12516 13132 12908 13188
rect 12964 13132 12974 13188
rect 13906 13132 13916 13188
rect 13972 13132 14476 13188
rect 14532 13132 14542 13188
rect 15250 13132 15260 13188
rect 15316 13132 15484 13188
rect 15540 13132 15550 13188
rect 20178 13132 20188 13188
rect 20244 13132 22988 13188
rect 23044 13132 23054 13188
rect 23650 13132 23660 13188
rect 23716 13132 23772 13188
rect 23828 13132 23838 13188
rect 24332 13132 24948 13188
rect 25666 13132 25676 13188
rect 25732 13132 25788 13188
rect 25844 13132 25854 13188
rect 26852 13132 43484 13188
rect 43540 13132 43550 13188
rect 43932 13132 47516 13188
rect 47572 13132 47582 13188
rect 48066 13132 48076 13188
rect 48132 13132 48636 13188
rect 48692 13132 48702 13188
rect 48850 13132 48860 13188
rect 48916 13132 52668 13188
rect 52724 13132 52734 13188
rect 54646 13132 54684 13188
rect 54740 13132 54750 13188
rect 5068 13076 5124 13132
rect 26852 13076 26908 13132
rect 43932 13076 43988 13132
rect 1698 13020 1708 13076
rect 1764 13020 3500 13076
rect 3556 13020 3566 13076
rect 4610 13020 4620 13076
rect 4676 13020 4686 13076
rect 4946 13020 4956 13076
rect 5012 13020 5124 13076
rect 5506 13020 5516 13076
rect 5572 13020 5740 13076
rect 5796 13020 5806 13076
rect 6178 13020 6188 13076
rect 6244 13020 6300 13076
rect 6356 13020 6366 13076
rect 8082 13020 8092 13076
rect 8148 13020 8988 13076
rect 9044 13020 9054 13076
rect 9650 13020 9660 13076
rect 9716 13020 13804 13076
rect 13860 13020 14476 13076
rect 14532 13020 14542 13076
rect 18610 13020 18620 13076
rect 18676 13020 19404 13076
rect 19460 13020 19470 13076
rect 20962 13020 20972 13076
rect 21028 13020 23212 13076
rect 23268 13020 23278 13076
rect 23426 13020 23436 13076
rect 23492 13020 26908 13076
rect 27010 13020 27020 13076
rect 27076 13020 27692 13076
rect 27748 13020 27758 13076
rect 28690 13020 28700 13076
rect 28756 13020 30156 13076
rect 30212 13020 31164 13076
rect 31220 13020 32620 13076
rect 32676 13020 32686 13076
rect 38882 13020 38892 13076
rect 38948 13020 40908 13076
rect 40964 13020 43988 13076
rect 44594 13020 44604 13076
rect 44660 13020 44940 13076
rect 44996 13020 45006 13076
rect 45126 13020 45164 13076
rect 45220 13020 45230 13076
rect 46162 13020 46172 13076
rect 46228 13020 46844 13076
rect 46900 13020 46910 13076
rect 47394 13020 47404 13076
rect 47460 13020 56588 13076
rect 56644 13020 56654 13076
rect 4620 12964 4676 13020
rect 2482 12908 2492 12964
rect 2548 12908 4564 12964
rect 4620 12908 5292 12964
rect 5348 12908 6748 12964
rect 6804 12908 6814 12964
rect 7522 12908 7532 12964
rect 7588 12908 9100 12964
rect 9156 12908 9166 12964
rect 10546 12908 10556 12964
rect 10612 12908 10892 12964
rect 10948 12908 10958 12964
rect 12114 12908 12124 12964
rect 12180 12908 13132 12964
rect 13188 12908 13198 12964
rect 13682 12908 13692 12964
rect 13748 12908 17500 12964
rect 17556 12908 17566 12964
rect 20178 12908 20188 12964
rect 20244 12908 21308 12964
rect 21364 12908 21374 12964
rect 21522 12908 21532 12964
rect 21588 12908 22428 12964
rect 22484 12908 22494 12964
rect 22642 12908 22652 12964
rect 22708 12908 29148 12964
rect 29204 12908 33068 12964
rect 33124 12908 33134 12964
rect 36866 12908 36876 12964
rect 36932 12908 37324 12964
rect 37380 12908 38108 12964
rect 38164 12908 40516 12964
rect 41010 12908 41020 12964
rect 41076 12908 41244 12964
rect 41300 12908 41310 12964
rect 41794 12908 41804 12964
rect 41860 12908 43260 12964
rect 43316 12908 43326 12964
rect 43474 12908 43484 12964
rect 43540 12908 44380 12964
rect 44436 12908 44446 12964
rect 44604 12908 48972 12964
rect 49028 12908 49038 12964
rect 50418 12908 50428 12964
rect 50484 12908 52332 12964
rect 52388 12908 52556 12964
rect 52612 12908 52622 12964
rect 0 12852 112 12880
rect 4508 12852 4564 12908
rect 40460 12852 40516 12908
rect 44604 12852 44660 12908
rect 57344 12852 57456 12880
rect 0 12796 140 12852
rect 196 12796 206 12852
rect 2146 12796 2156 12852
rect 2212 12796 4452 12852
rect 4508 12796 6412 12852
rect 6468 12796 6478 12852
rect 7186 12796 7196 12852
rect 7252 12796 8652 12852
rect 8708 12796 8718 12852
rect 16268 12796 16828 12852
rect 16884 12796 17276 12852
rect 17332 12796 17342 12852
rect 18946 12796 18956 12852
rect 19012 12796 20860 12852
rect 20916 12796 20926 12852
rect 21410 12796 21420 12852
rect 21476 12796 26236 12852
rect 26292 12796 26302 12852
rect 27010 12796 27020 12852
rect 27076 12796 31836 12852
rect 31892 12796 31902 12852
rect 33068 12796 36204 12852
rect 36260 12796 36270 12852
rect 39218 12796 39228 12852
rect 39284 12796 40236 12852
rect 40292 12796 40302 12852
rect 40460 12796 44660 12852
rect 44716 12796 51772 12852
rect 51828 12796 51838 12852
rect 53330 12796 53340 12852
rect 53396 12796 57456 12852
rect 0 12768 112 12796
rect 4396 12740 4452 12796
rect 16268 12740 16324 12796
rect 33068 12740 33124 12796
rect 39228 12740 39284 12796
rect 44716 12740 44772 12796
rect 57344 12768 57456 12796
rect 2818 12684 2828 12740
rect 2884 12684 4340 12740
rect 4396 12684 5292 12740
rect 5348 12684 8204 12740
rect 8260 12684 8270 12740
rect 8530 12684 8540 12740
rect 8596 12684 16324 12740
rect 16482 12684 16492 12740
rect 16548 12684 30044 12740
rect 30100 12684 30110 12740
rect 33058 12684 33068 12740
rect 33124 12684 33134 12740
rect 33394 12684 33404 12740
rect 33460 12684 39284 12740
rect 39442 12684 39452 12740
rect 39508 12684 39788 12740
rect 39844 12684 40572 12740
rect 40628 12684 43260 12740
rect 43316 12684 43326 12740
rect 43474 12684 43484 12740
rect 43540 12684 44212 12740
rect 44594 12684 44604 12740
rect 44660 12684 44772 12740
rect 44930 12684 44940 12740
rect 44996 12684 49756 12740
rect 49812 12684 49822 12740
rect 50978 12684 50988 12740
rect 51044 12684 51436 12740
rect 51492 12684 51502 12740
rect 2258 12572 2268 12628
rect 2324 12572 3612 12628
rect 3668 12572 3678 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 4284 12516 4340 12684
rect 44156 12628 44212 12684
rect 4498 12572 4508 12628
rect 4564 12572 9268 12628
rect 11106 12572 11116 12628
rect 11172 12572 13020 12628
rect 13076 12572 13086 12628
rect 13234 12572 13244 12628
rect 13300 12572 23660 12628
rect 23716 12572 23726 12628
rect 24210 12572 24220 12628
rect 24276 12572 24444 12628
rect 24500 12572 24510 12628
rect 25890 12572 25900 12628
rect 25956 12572 26124 12628
rect 26180 12572 26190 12628
rect 30706 12572 30716 12628
rect 30772 12572 35084 12628
rect 35140 12572 35150 12628
rect 36194 12572 36204 12628
rect 36260 12572 42252 12628
rect 42308 12572 42318 12628
rect 43026 12572 43036 12628
rect 43092 12572 43148 12628
rect 43204 12572 43214 12628
rect 44156 12572 44940 12628
rect 44996 12572 45006 12628
rect 46470 12572 46508 12628
rect 46564 12572 46574 12628
rect 47282 12572 47292 12628
rect 47348 12572 49196 12628
rect 49252 12572 49262 12628
rect 9212 12516 9268 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 354 12460 364 12516
rect 420 12460 2940 12516
rect 2996 12460 3006 12516
rect 3378 12460 3388 12516
rect 3444 12460 3482 12516
rect 4284 12460 4396 12516
rect 4452 12460 4462 12516
rect 5730 12460 5740 12516
rect 5796 12460 5806 12516
rect 5964 12460 6300 12516
rect 6356 12460 7196 12516
rect 7252 12460 7262 12516
rect 8642 12460 8652 12516
rect 8708 12460 8988 12516
rect 9044 12460 9054 12516
rect 9212 12460 14924 12516
rect 14980 12460 14990 12516
rect 15092 12460 21028 12516
rect 21522 12460 21532 12516
rect 21588 12460 22652 12516
rect 22708 12460 22718 12516
rect 25218 12460 25228 12516
rect 25284 12460 25564 12516
rect 25620 12460 25630 12516
rect 26114 12460 26124 12516
rect 26180 12460 27804 12516
rect 27860 12460 28924 12516
rect 28980 12460 28990 12516
rect 29138 12460 29148 12516
rect 29204 12460 40796 12516
rect 40852 12460 41804 12516
rect 41860 12460 41870 12516
rect 42130 12460 42140 12516
rect 42196 12460 43484 12516
rect 43540 12460 43550 12516
rect 45602 12460 45612 12516
rect 45668 12460 46844 12516
rect 46900 12460 47852 12516
rect 47908 12460 47918 12516
rect 48290 12460 48300 12516
rect 48356 12460 48972 12516
rect 49028 12460 49038 12516
rect 0 12404 112 12432
rect 5740 12404 5796 12460
rect 5964 12404 6020 12460
rect 15092 12404 15148 12460
rect 20972 12404 21028 12460
rect 57344 12404 57456 12432
rect 0 12348 140 12404
rect 196 12348 206 12404
rect 2146 12348 2156 12404
rect 2212 12348 5292 12404
rect 5740 12348 6020 12404
rect 6738 12348 6748 12404
rect 6804 12348 7420 12404
rect 7476 12348 7486 12404
rect 8194 12348 8204 12404
rect 8260 12348 11564 12404
rect 11620 12348 11630 12404
rect 11778 12348 11788 12404
rect 11844 12348 12236 12404
rect 12292 12348 12302 12404
rect 12460 12348 15148 12404
rect 15362 12348 15372 12404
rect 15428 12348 17836 12404
rect 17892 12348 18508 12404
rect 18564 12348 18574 12404
rect 20972 12348 49420 12404
rect 49476 12348 49486 12404
rect 50642 12348 50652 12404
rect 50708 12348 51100 12404
rect 51156 12348 51996 12404
rect 52052 12348 52556 12404
rect 52612 12348 52622 12404
rect 55682 12348 55692 12404
rect 55748 12348 57456 12404
rect 0 12320 112 12348
rect 5236 12292 5292 12348
rect 1138 12236 1148 12292
rect 1204 12236 2380 12292
rect 2436 12236 2446 12292
rect 3266 12236 3276 12292
rect 3332 12236 4508 12292
rect 4564 12236 4574 12292
rect 4918 12236 4956 12292
rect 5012 12236 5022 12292
rect 5236 12236 11788 12292
rect 11844 12236 11854 12292
rect 12460 12180 12516 12348
rect 57344 12320 57456 12348
rect 14130 12236 14140 12292
rect 14196 12236 15428 12292
rect 17938 12236 17948 12292
rect 18004 12236 24164 12292
rect 25218 12236 25228 12292
rect 25284 12236 28700 12292
rect 28756 12236 28766 12292
rect 28914 12236 28924 12292
rect 28980 12236 31836 12292
rect 31892 12236 33852 12292
rect 33908 12236 33918 12292
rect 34626 12236 34636 12292
rect 34692 12236 34972 12292
rect 35028 12236 35038 12292
rect 37090 12236 37100 12292
rect 37156 12236 55916 12292
rect 55972 12236 55982 12292
rect 15372 12180 15428 12236
rect 24108 12180 24164 12236
rect 18 12124 28 12180
rect 84 12124 140 12180
rect 196 12124 206 12180
rect 1894 12124 1932 12180
rect 1988 12124 1998 12180
rect 3266 12124 3276 12180
rect 3332 12124 3500 12180
rect 3556 12124 3566 12180
rect 3714 12124 3724 12180
rect 3780 12124 5180 12180
rect 5236 12124 5246 12180
rect 5618 12124 5628 12180
rect 5684 12124 6972 12180
rect 7028 12124 7038 12180
rect 7410 12124 7420 12180
rect 7476 12124 12516 12180
rect 13010 12124 13020 12180
rect 13076 12124 14140 12180
rect 14196 12124 14700 12180
rect 14756 12124 14766 12180
rect 15372 12124 15932 12180
rect 15988 12124 18396 12180
rect 18452 12124 18462 12180
rect 19058 12124 19068 12180
rect 19124 12124 19852 12180
rect 19908 12124 19918 12180
rect 20066 12124 20076 12180
rect 20132 12124 21644 12180
rect 21700 12124 21710 12180
rect 23090 12124 23100 12180
rect 23156 12124 23884 12180
rect 23940 12124 23950 12180
rect 24108 12124 25452 12180
rect 25508 12124 25518 12180
rect 26338 12124 26348 12180
rect 26404 12124 26684 12180
rect 26740 12124 26750 12180
rect 31266 12124 31276 12180
rect 31332 12124 31724 12180
rect 31780 12124 31790 12180
rect 32946 12124 32956 12180
rect 33012 12124 33852 12180
rect 33908 12124 33964 12180
rect 34020 12124 34030 12180
rect 38882 12124 38892 12180
rect 38948 12124 40796 12180
rect 40852 12124 40862 12180
rect 42914 12124 42924 12180
rect 42980 12124 45388 12180
rect 45444 12124 45454 12180
rect 46386 12124 46396 12180
rect 46452 12124 46620 12180
rect 46676 12124 46686 12180
rect 46946 12124 46956 12180
rect 47012 12124 49028 12180
rect 49186 12124 49196 12180
rect 49252 12124 52668 12180
rect 52724 12124 52734 12180
rect 53442 12124 53452 12180
rect 53508 12124 54012 12180
rect 54068 12124 55132 12180
rect 55188 12124 55198 12180
rect 2818 12012 2828 12068
rect 2884 12012 4172 12068
rect 4228 12012 4238 12068
rect 4834 12012 4844 12068
rect 4900 12012 5572 12068
rect 5842 12012 5852 12068
rect 5908 12012 6300 12068
rect 6356 12012 6366 12068
rect 6514 12012 6524 12068
rect 6580 12012 7644 12068
rect 7700 12012 7710 12068
rect 7858 12012 7868 12068
rect 7924 12012 11116 12068
rect 11172 12012 11182 12068
rect 11330 12012 11340 12068
rect 11396 12012 17612 12068
rect 17668 12012 17678 12068
rect 19170 12012 19180 12068
rect 19236 12012 20300 12068
rect 20356 12012 20972 12068
rect 21028 12012 21038 12068
rect 21942 12012 21980 12068
rect 22036 12012 22046 12068
rect 22530 12012 22540 12068
rect 22596 12012 23324 12068
rect 23380 12012 23390 12068
rect 23538 12012 23548 12068
rect 23604 12012 23614 12068
rect 23986 12012 23996 12068
rect 24052 12012 28476 12068
rect 28532 12012 28542 12068
rect 31574 12012 31612 12068
rect 31668 12012 31678 12068
rect 31938 12012 31948 12068
rect 32004 12012 34524 12068
rect 34580 12012 34590 12068
rect 35756 12012 39004 12068
rect 39060 12012 39070 12068
rect 39330 12012 39340 12068
rect 39396 12012 39676 12068
rect 39732 12012 47348 12068
rect 47842 12012 47852 12068
rect 47908 12012 48300 12068
rect 48356 12012 48366 12068
rect 48514 12012 48524 12068
rect 48580 12012 48618 12068
rect 0 11956 112 11984
rect 5516 11956 5572 12012
rect 23548 11956 23604 12012
rect 0 11900 1148 11956
rect 1204 11900 1214 11956
rect 3266 11900 3276 11956
rect 3332 11900 3612 11956
rect 3668 11900 3678 11956
rect 5516 11900 6020 11956
rect 6290 11900 6300 11956
rect 6356 11900 6748 11956
rect 6804 11900 6814 11956
rect 7298 11900 7308 11956
rect 7364 11900 9660 11956
rect 9716 11900 9726 11956
rect 12338 11900 12348 11956
rect 12404 11900 14308 11956
rect 14466 11900 14476 11956
rect 14532 11900 23100 11956
rect 23156 11900 23166 11956
rect 23548 11900 23660 11956
rect 23716 11900 29148 11956
rect 29204 11900 29214 11956
rect 30370 11900 30380 11956
rect 30436 11900 34972 11956
rect 35028 11900 35038 11956
rect 0 11872 112 11900
rect 5964 11844 6020 11900
rect 14252 11844 14308 11900
rect 1222 11788 1260 11844
rect 1316 11788 1326 11844
rect 2034 11788 2044 11844
rect 2100 11788 3500 11844
rect 3556 11788 3566 11844
rect 5964 11788 8204 11844
rect 8260 11788 8270 11844
rect 9538 11788 9548 11844
rect 9604 11788 9996 11844
rect 10052 11788 10062 11844
rect 11106 11788 11116 11844
rect 11172 11788 12012 11844
rect 12068 11788 12078 11844
rect 13804 11788 13916 11844
rect 13972 11788 13982 11844
rect 14252 11788 15372 11844
rect 15428 11788 15438 11844
rect 15586 11788 15596 11844
rect 15652 11788 16156 11844
rect 16212 11788 16222 11844
rect 21970 11788 21980 11844
rect 22036 11788 22764 11844
rect 22820 11788 22830 11844
rect 23538 11788 23548 11844
rect 23604 11788 23772 11844
rect 23828 11788 23838 11844
rect 25554 11788 25564 11844
rect 25620 11788 26684 11844
rect 26740 11788 26750 11844
rect 26852 11788 27692 11844
rect 27748 11788 30156 11844
rect 30212 11788 30222 11844
rect 31826 11788 31836 11844
rect 31892 11788 32564 11844
rect 34178 11788 34188 11844
rect 34244 11788 35532 11844
rect 35588 11788 35598 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 13804 11732 13860 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 26852 11732 26908 11788
rect 32508 11732 32564 11788
rect 35756 11732 35812 12012
rect 47292 11956 47348 12012
rect 48972 11956 49028 12124
rect 50306 12012 50316 12068
rect 50372 12012 53564 12068
rect 53620 12012 53630 12068
rect 54422 12012 54460 12068
rect 54516 12012 54526 12068
rect 57344 11956 57456 11984
rect 36306 11900 36316 11956
rect 36372 11900 37548 11956
rect 37604 11900 37614 11956
rect 40348 11900 44828 11956
rect 44884 11900 44894 11956
rect 45826 11900 45836 11956
rect 45892 11900 47068 11956
rect 47124 11900 47134 11956
rect 47282 11900 47292 11956
rect 47348 11900 47358 11956
rect 47842 11900 47852 11956
rect 47908 11900 48748 11956
rect 48804 11900 48814 11956
rect 48972 11900 50428 11956
rect 50484 11900 50494 11956
rect 52658 11900 52668 11956
rect 52724 11900 53788 11956
rect 53844 11900 54124 11956
rect 54180 11900 54190 11956
rect 55122 11900 55132 11956
rect 55188 11900 55580 11956
rect 55636 11900 55646 11956
rect 56242 11900 56252 11956
rect 56308 11900 57456 11956
rect 40348 11844 40404 11900
rect 57344 11872 57456 11900
rect 37650 11788 37660 11844
rect 37716 11788 37996 11844
rect 38052 11788 40404 11844
rect 42802 11788 42812 11844
rect 42868 11788 42924 11844
rect 42980 11788 42990 11844
rect 43250 11788 43260 11844
rect 43316 11788 44268 11844
rect 44324 11788 44334 11844
rect 46694 11788 46732 11844
rect 46788 11788 46798 11844
rect 47282 11788 47292 11844
rect 47348 11788 48300 11844
rect 48356 11788 48366 11844
rect 48626 11788 48636 11844
rect 48692 11788 49084 11844
rect 49140 11788 49150 11844
rect 50194 11788 50204 11844
rect 50260 11788 51324 11844
rect 51380 11788 51390 11844
rect 52070 11788 52108 11844
rect 52164 11788 52174 11844
rect 52434 11788 52444 11844
rect 52500 11788 53004 11844
rect 53060 11788 53070 11844
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 5954 11676 5964 11732
rect 6020 11676 12964 11732
rect 13122 11676 13132 11732
rect 13188 11676 13860 11732
rect 14476 11676 15260 11732
rect 15316 11676 15326 11732
rect 15698 11676 15708 11732
rect 15764 11676 16604 11732
rect 16660 11676 16670 11732
rect 18834 11676 18844 11732
rect 18900 11676 19516 11732
rect 19572 11676 19740 11732
rect 19796 11676 19806 11732
rect 21298 11676 21308 11732
rect 21364 11676 22204 11732
rect 22260 11676 22270 11732
rect 22428 11676 24220 11732
rect 24276 11676 24286 11732
rect 26562 11676 26572 11732
rect 26628 11676 26908 11732
rect 27010 11676 27020 11732
rect 27076 11676 28252 11732
rect 28308 11676 28318 11732
rect 29026 11676 29036 11732
rect 29092 11676 32284 11732
rect 32340 11676 32350 11732
rect 32508 11676 35812 11732
rect 36642 11676 36652 11732
rect 36708 11676 37100 11732
rect 37156 11676 37166 11732
rect 38098 11676 38108 11732
rect 38164 11676 38332 11732
rect 38388 11676 38398 11732
rect 38882 11676 38892 11732
rect 38948 11676 41020 11732
rect 41076 11676 41086 11732
rect 45490 11676 45500 11732
rect 45556 11676 55020 11732
rect 55076 11676 55086 11732
rect 1250 11564 1260 11620
rect 1316 11564 1820 11620
rect 1876 11564 4956 11620
rect 5012 11564 5022 11620
rect 5170 11564 5180 11620
rect 5236 11564 5628 11620
rect 5684 11564 5694 11620
rect 6626 11564 6636 11620
rect 6692 11564 8036 11620
rect 8194 11564 8204 11620
rect 8260 11564 9324 11620
rect 9380 11564 9492 11620
rect 9622 11564 9660 11620
rect 9716 11564 9726 11620
rect 9986 11564 9996 11620
rect 10052 11564 11564 11620
rect 11620 11564 11630 11620
rect 0 11508 112 11536
rect 7980 11508 8036 11564
rect 9436 11508 9492 11564
rect 12908 11508 12964 11676
rect 14476 11620 14532 11676
rect 13570 11564 13580 11620
rect 13636 11564 14532 11620
rect 14690 11564 14700 11620
rect 14756 11564 15036 11620
rect 15092 11564 15102 11620
rect 15334 11564 15372 11620
rect 15428 11564 15438 11620
rect 15586 11564 15596 11620
rect 15652 11564 15690 11620
rect 16146 11564 16156 11620
rect 16212 11564 17836 11620
rect 17892 11564 17902 11620
rect 18722 11564 18732 11620
rect 18788 11564 20188 11620
rect 20244 11564 20254 11620
rect 16156 11508 16212 11564
rect 22428 11508 22484 11676
rect 22866 11564 22876 11620
rect 22932 11564 24332 11620
rect 24388 11564 24398 11620
rect 25442 11564 25452 11620
rect 25508 11564 35308 11620
rect 35364 11564 35644 11620
rect 35700 11564 35710 11620
rect 35858 11564 35868 11620
rect 35924 11564 36540 11620
rect 36596 11564 36606 11620
rect 38612 11564 40348 11620
rect 40404 11564 40414 11620
rect 42242 11564 42252 11620
rect 42308 11564 42476 11620
rect 42532 11564 42542 11620
rect 43026 11564 43036 11620
rect 43092 11564 49084 11620
rect 49140 11564 49150 11620
rect 49522 11564 49532 11620
rect 49588 11564 50092 11620
rect 50148 11564 50158 11620
rect 50726 11564 50764 11620
rect 50820 11564 50830 11620
rect 51874 11564 51884 11620
rect 51940 11564 52332 11620
rect 52388 11564 52398 11620
rect 52546 11564 52556 11620
rect 52612 11564 53564 11620
rect 53620 11564 53630 11620
rect 56354 11564 56364 11620
rect 56420 11564 56476 11620
rect 56532 11564 56542 11620
rect 38612 11508 38668 11564
rect 57344 11508 57456 11536
rect 0 11452 644 11508
rect 802 11452 812 11508
rect 868 11452 1596 11508
rect 1652 11452 1662 11508
rect 4946 11452 4956 11508
rect 5012 11452 5404 11508
rect 5460 11452 5470 11508
rect 5842 11452 5852 11508
rect 5908 11452 6300 11508
rect 6356 11452 6366 11508
rect 6738 11452 6748 11508
rect 6804 11452 6972 11508
rect 7028 11452 7084 11508
rect 7140 11452 7150 11508
rect 7980 11452 9212 11508
rect 9268 11452 9278 11508
rect 9436 11452 10332 11508
rect 10388 11452 11676 11508
rect 11732 11452 11900 11508
rect 11956 11452 11966 11508
rect 12908 11458 15316 11508
rect 15484 11458 15764 11508
rect 15932 11458 16212 11508
rect 12908 11452 16212 11458
rect 16482 11452 16492 11508
rect 16548 11452 19460 11508
rect 19618 11452 19628 11508
rect 19684 11452 20748 11508
rect 20804 11452 20814 11508
rect 22194 11452 22204 11508
rect 22260 11452 22484 11508
rect 23426 11452 23436 11508
rect 23492 11452 29316 11508
rect 29922 11452 29932 11508
rect 29988 11452 30268 11508
rect 30324 11452 30334 11508
rect 34738 11452 34748 11508
rect 34804 11452 38668 11508
rect 38994 11452 39004 11508
rect 39060 11452 40908 11508
rect 40964 11452 40974 11508
rect 41122 11452 41132 11508
rect 41188 11452 42028 11508
rect 42084 11452 42588 11508
rect 42644 11452 42654 11508
rect 44034 11452 44044 11508
rect 44100 11452 45612 11508
rect 45668 11452 45678 11508
rect 47394 11452 47404 11508
rect 47460 11452 48748 11508
rect 48804 11452 48814 11508
rect 48962 11452 48972 11508
rect 49028 11452 52892 11508
rect 52948 11452 52958 11508
rect 53116 11452 57456 11508
rect 0 11424 112 11452
rect 588 11396 644 11452
rect 15260 11402 15540 11452
rect 15708 11402 15988 11452
rect 19404 11396 19460 11452
rect 588 11340 2492 11396
rect 2548 11340 2558 11396
rect 5170 11340 5180 11396
rect 5236 11340 6972 11396
rect 7028 11340 7038 11396
rect 9426 11340 9436 11396
rect 9492 11340 9996 11396
rect 10052 11340 10062 11396
rect 11106 11340 11116 11396
rect 11172 11340 15036 11396
rect 15092 11340 15102 11396
rect 16370 11340 16380 11396
rect 16436 11340 17388 11396
rect 17444 11340 19180 11396
rect 19236 11340 19246 11396
rect 19404 11340 25452 11396
rect 25508 11340 25518 11396
rect 26786 11340 26796 11396
rect 26852 11340 27580 11396
rect 27636 11340 27646 11396
rect 28018 11340 28028 11396
rect 28084 11340 28812 11396
rect 28868 11340 28878 11396
rect 29260 11284 29316 11452
rect 29474 11340 29484 11396
rect 29540 11340 30156 11396
rect 30212 11340 30222 11396
rect 33170 11340 33180 11396
rect 33236 11340 36652 11396
rect 36708 11340 38668 11396
rect 39106 11340 39116 11396
rect 39172 11340 43372 11396
rect 43428 11340 43438 11396
rect 44118 11340 44156 11396
rect 44212 11340 44222 11396
rect 47842 11340 47852 11396
rect 47908 11340 48524 11396
rect 48580 11340 48636 11396
rect 48692 11340 48702 11396
rect 38612 11284 38668 11340
rect 53116 11284 53172 11452
rect 57344 11424 57456 11452
rect 3266 11228 3276 11284
rect 3332 11228 3724 11284
rect 3780 11228 3790 11284
rect 4162 11228 4172 11284
rect 4228 11228 5292 11284
rect 5348 11228 5358 11284
rect 5618 11228 5628 11284
rect 5684 11228 7868 11284
rect 7924 11228 7934 11284
rect 8194 11228 8204 11284
rect 8260 11228 8428 11284
rect 8484 11228 8494 11284
rect 8876 11228 8988 11284
rect 9044 11228 9054 11284
rect 11666 11228 11676 11284
rect 11732 11228 12236 11284
rect 12292 11228 12302 11284
rect 13346 11228 13356 11284
rect 13412 11228 14364 11284
rect 14420 11228 14430 11284
rect 14578 11228 14588 11284
rect 14644 11228 17948 11284
rect 18004 11228 18014 11284
rect 21298 11228 21308 11284
rect 21364 11228 26572 11284
rect 26628 11228 26638 11284
rect 29260 11228 37100 11284
rect 37156 11228 37166 11284
rect 38612 11228 39340 11284
rect 39396 11228 39406 11284
rect 39554 11228 39564 11284
rect 39620 11228 40236 11284
rect 40292 11228 40302 11284
rect 44034 11228 44044 11284
rect 44100 11228 44940 11284
rect 44996 11228 45006 11284
rect 46274 11228 46284 11284
rect 46340 11228 51772 11284
rect 51828 11228 51838 11284
rect 53106 11228 53116 11284
rect 53172 11228 53182 11284
rect 8876 11172 8932 11228
rect 690 11116 700 11172
rect 756 11116 1596 11172
rect 1652 11116 1662 11172
rect 3612 11116 8932 11172
rect 9090 11116 9100 11172
rect 9156 11116 12124 11172
rect 12180 11116 12190 11172
rect 13906 11116 13916 11172
rect 13972 11116 16156 11172
rect 16212 11116 16604 11172
rect 16660 11116 16670 11172
rect 16930 11116 16940 11172
rect 16996 11116 17724 11172
rect 17780 11116 17790 11172
rect 18470 11116 18508 11172
rect 18564 11116 18574 11172
rect 19170 11116 19180 11172
rect 19236 11116 20860 11172
rect 20916 11116 21756 11172
rect 21812 11116 21822 11172
rect 23762 11116 23772 11172
rect 23828 11116 25788 11172
rect 25844 11116 25854 11172
rect 26124 11116 27244 11172
rect 27300 11116 28700 11172
rect 28756 11116 28766 11172
rect 32162 11116 32172 11172
rect 32228 11116 34524 11172
rect 34580 11116 34590 11172
rect 37314 11116 37324 11172
rect 37380 11116 40124 11172
rect 40180 11116 40908 11172
rect 40964 11116 40974 11172
rect 43596 11116 46732 11172
rect 46788 11116 46798 11172
rect 46946 11116 46956 11172
rect 47012 11116 56028 11172
rect 56084 11116 56094 11172
rect 0 11060 112 11088
rect 3612 11060 3668 11116
rect 17724 11060 17780 11116
rect 26124 11060 26180 11116
rect 37324 11060 37380 11116
rect 0 11004 812 11060
rect 868 11004 878 11060
rect 2930 11004 2940 11060
rect 2996 11004 3668 11060
rect 4386 11004 4396 11060
rect 4452 11004 5628 11060
rect 5684 11004 5694 11060
rect 5954 11004 5964 11060
rect 6020 11004 9436 11060
rect 9492 11004 9660 11060
rect 9716 11004 9726 11060
rect 10210 11004 10220 11060
rect 10276 11004 15036 11060
rect 15092 11004 16268 11060
rect 16324 11004 16334 11060
rect 17724 11004 22428 11060
rect 22484 11004 22494 11060
rect 24210 11004 24220 11060
rect 24276 11004 26180 11060
rect 26338 11004 26348 11060
rect 26404 11004 29932 11060
rect 29988 11004 29998 11060
rect 32610 11004 32620 11060
rect 32676 11004 37380 11060
rect 38612 11004 40348 11060
rect 40404 11004 42812 11060
rect 42868 11004 42878 11060
rect 0 10976 112 11004
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 38612 10948 38668 11004
rect 43596 10948 43652 11116
rect 57344 11060 57456 11088
rect 44258 11004 44268 11060
rect 44324 11004 46956 11060
rect 47012 11004 47022 11060
rect 47590 11004 47628 11060
rect 47684 11004 47694 11060
rect 48402 11004 48412 11060
rect 48468 11004 48524 11060
rect 48580 11004 48590 11060
rect 52994 11004 53004 11060
rect 53060 11004 57456 11060
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 57344 10976 57456 11004
rect 1362 10892 1372 10948
rect 1428 10892 3668 10948
rect 4162 10892 4172 10948
rect 4228 10892 8428 10948
rect 8484 10892 8494 10948
rect 9090 10892 9100 10948
rect 9156 10892 12348 10948
rect 12404 10892 12414 10948
rect 14354 10892 14364 10948
rect 14420 10892 17500 10948
rect 17556 10892 20076 10948
rect 20132 10892 20142 10948
rect 21858 10892 21868 10948
rect 21924 10892 22204 10948
rect 22260 10892 22270 10948
rect 22530 10892 22540 10948
rect 22596 10892 23324 10948
rect 23380 10892 23390 10948
rect 26002 10892 26012 10948
rect 26068 10892 30380 10948
rect 30436 10892 30446 10948
rect 32732 10892 38668 10948
rect 38994 10892 39004 10948
rect 39060 10892 43652 10948
rect 44482 10892 44492 10948
rect 44548 10892 53564 10948
rect 53620 10892 53630 10948
rect 53778 10892 53788 10948
rect 53844 10892 53882 10948
rect 3612 10836 3668 10892
rect 32732 10836 32788 10892
rect 3612 10780 5180 10836
rect 5236 10780 5404 10836
rect 5460 10780 5470 10836
rect 5618 10780 5628 10836
rect 5684 10780 5964 10836
rect 6020 10780 6030 10836
rect 6178 10780 6188 10836
rect 6244 10780 6300 10836
rect 6356 10780 7084 10836
rect 7140 10780 7150 10836
rect 10546 10780 10556 10836
rect 10612 10780 10892 10836
rect 10948 10780 10958 10836
rect 11106 10780 11116 10836
rect 11172 10780 13636 10836
rect 13794 10780 13804 10836
rect 13860 10780 14924 10836
rect 14980 10780 15260 10836
rect 15316 10780 15326 10836
rect 15474 10780 15484 10836
rect 15540 10780 16268 10836
rect 16324 10780 16334 10836
rect 16594 10780 16604 10836
rect 16660 10780 16716 10836
rect 16772 10780 16782 10836
rect 17266 10780 17276 10836
rect 17332 10780 19964 10836
rect 20020 10780 26348 10836
rect 26404 10780 26414 10836
rect 26562 10780 26572 10836
rect 26628 10780 32788 10836
rect 32844 10780 56308 10836
rect 13580 10724 13636 10780
rect 17276 10724 17332 10780
rect 32844 10724 32900 10780
rect 3332 10668 8876 10724
rect 8932 10668 8942 10724
rect 9762 10668 9772 10724
rect 9828 10668 11452 10724
rect 11508 10668 11518 10724
rect 12450 10668 12460 10724
rect 12516 10668 12908 10724
rect 12964 10668 12974 10724
rect 13580 10668 14700 10724
rect 14756 10668 17332 10724
rect 20962 10668 20972 10724
rect 21028 10668 21420 10724
rect 21476 10668 22204 10724
rect 22260 10668 22270 10724
rect 22418 10668 22428 10724
rect 22484 10668 25284 10724
rect 25442 10668 25452 10724
rect 25508 10668 28028 10724
rect 28084 10668 28094 10724
rect 29222 10668 29260 10724
rect 29316 10668 29326 10724
rect 31052 10668 32900 10724
rect 37202 10668 37212 10724
rect 37268 10668 44492 10724
rect 44548 10668 44558 10724
rect 44706 10668 44716 10724
rect 44772 10668 48188 10724
rect 48244 10668 48254 10724
rect 49382 10668 49420 10724
rect 49476 10668 49486 10724
rect 49634 10668 49644 10724
rect 49700 10668 53788 10724
rect 53844 10668 53854 10724
rect 0 10612 112 10640
rect 3332 10612 3388 10668
rect 25228 10612 25284 10668
rect 31052 10612 31108 10668
rect 56252 10612 56308 10780
rect 57344 10612 57456 10640
rect 0 10556 3388 10612
rect 3602 10556 3612 10612
rect 3668 10556 4844 10612
rect 4900 10556 4910 10612
rect 5058 10556 5068 10612
rect 5124 10556 5134 10612
rect 5282 10556 5292 10612
rect 5348 10556 5516 10612
rect 5572 10556 5582 10612
rect 5954 10556 5964 10612
rect 6020 10556 6860 10612
rect 6916 10556 6926 10612
rect 7634 10556 7644 10612
rect 7700 10556 8316 10612
rect 8372 10556 8382 10612
rect 8530 10556 8540 10612
rect 8596 10556 10332 10612
rect 10388 10556 11004 10612
rect 11060 10556 11172 10612
rect 11554 10556 11564 10612
rect 11620 10556 12348 10612
rect 12404 10556 12414 10612
rect 12684 10556 13244 10612
rect 13300 10556 13310 10612
rect 14578 10556 14588 10612
rect 14644 10556 14924 10612
rect 14980 10556 15092 10612
rect 15670 10556 15708 10612
rect 15764 10556 16828 10612
rect 16884 10556 17836 10612
rect 17892 10556 17902 10612
rect 18498 10556 18508 10612
rect 18564 10556 18956 10612
rect 19012 10556 21196 10612
rect 21252 10556 21262 10612
rect 21420 10556 23716 10612
rect 23874 10556 23884 10612
rect 23940 10556 24444 10612
rect 24500 10556 24510 10612
rect 24966 10556 25004 10612
rect 25060 10556 25070 10612
rect 25228 10556 25452 10612
rect 25508 10556 25518 10612
rect 25666 10556 25676 10612
rect 25732 10556 26460 10612
rect 26516 10556 31108 10612
rect 31238 10556 31276 10612
rect 31332 10556 31342 10612
rect 35746 10556 35756 10612
rect 35812 10556 36764 10612
rect 36820 10556 36830 10612
rect 38612 10556 39732 10612
rect 40450 10556 40460 10612
rect 40516 10556 41020 10612
rect 41076 10556 41086 10612
rect 42242 10556 42252 10612
rect 42308 10556 45276 10612
rect 45332 10556 45342 10612
rect 47730 10556 47740 10612
rect 47796 10556 48412 10612
rect 48468 10556 48478 10612
rect 49298 10556 49308 10612
rect 49364 10556 49756 10612
rect 49812 10556 49822 10612
rect 51986 10556 51996 10612
rect 52052 10556 52062 10612
rect 52770 10556 52780 10612
rect 52836 10556 52892 10612
rect 52948 10556 53676 10612
rect 53732 10556 53742 10612
rect 55346 10556 55356 10612
rect 55412 10556 56028 10612
rect 56084 10556 56094 10612
rect 56252 10556 57456 10612
rect 0 10528 112 10556
rect 5068 10500 5124 10556
rect 7644 10500 7700 10556
rect 1922 10444 1932 10500
rect 1988 10444 5124 10500
rect 5954 10444 5964 10500
rect 6020 10444 6076 10500
rect 6132 10444 6142 10500
rect 6626 10444 6636 10500
rect 6692 10444 7700 10500
rect 11116 10500 11172 10556
rect 12684 10500 12740 10556
rect 15036 10500 15092 10556
rect 11116 10444 12740 10500
rect 12898 10444 12908 10500
rect 12964 10444 14476 10500
rect 14532 10444 14542 10500
rect 15036 10444 15484 10500
rect 15540 10444 16716 10500
rect 16772 10444 16782 10500
rect 21420 10388 21476 10556
rect 23660 10500 23716 10556
rect 38612 10500 38668 10556
rect 22306 10444 22316 10500
rect 22372 10444 22540 10500
rect 22596 10444 22606 10500
rect 22764 10444 22988 10500
rect 23044 10444 23436 10500
rect 23492 10444 23502 10500
rect 23660 10444 26572 10500
rect 26628 10444 26638 10500
rect 30146 10444 30156 10500
rect 30212 10444 38668 10500
rect 3378 10332 3388 10388
rect 3444 10332 3500 10388
rect 3556 10332 3566 10388
rect 4162 10332 4172 10388
rect 4228 10332 4844 10388
rect 4900 10332 4910 10388
rect 5058 10332 5068 10388
rect 5124 10332 5134 10388
rect 5282 10332 5292 10388
rect 5348 10332 7644 10388
rect 7700 10332 7710 10388
rect 9426 10332 9436 10388
rect 9492 10332 9772 10388
rect 9828 10332 9838 10388
rect 9986 10332 9996 10388
rect 10052 10332 11788 10388
rect 11844 10332 11854 10388
rect 12562 10332 12572 10388
rect 12628 10332 13468 10388
rect 13524 10332 13534 10388
rect 15362 10332 15372 10388
rect 15428 10332 15596 10388
rect 15652 10332 15662 10388
rect 15810 10332 15820 10388
rect 15876 10332 21476 10388
rect 5068 10276 5124 10332
rect 22764 10276 22820 10444
rect 39676 10388 39732 10556
rect 51996 10500 52052 10556
rect 57344 10528 57456 10556
rect 39890 10444 39900 10500
rect 39956 10444 40124 10500
rect 40180 10444 42028 10500
rect 42084 10444 42094 10500
rect 44370 10444 44380 10500
rect 44436 10444 45948 10500
rect 46004 10444 46014 10500
rect 46722 10444 46732 10500
rect 46788 10444 47964 10500
rect 48020 10444 52668 10500
rect 52724 10444 52734 10500
rect 56242 10444 56252 10500
rect 56308 10444 56364 10500
rect 56420 10444 56430 10500
rect 22988 10332 23996 10388
rect 24052 10332 24062 10388
rect 24332 10332 25620 10388
rect 25778 10332 25788 10388
rect 25844 10332 26012 10388
rect 26068 10332 26078 10388
rect 29026 10332 29036 10388
rect 29092 10332 29596 10388
rect 29652 10332 29662 10388
rect 30258 10332 30268 10388
rect 30324 10332 33292 10388
rect 33348 10332 33358 10388
rect 33506 10332 33516 10388
rect 33572 10332 39340 10388
rect 39396 10332 39406 10388
rect 39676 10332 44156 10388
rect 44212 10332 44222 10388
rect 44594 10332 44604 10388
rect 44660 10332 46060 10388
rect 46116 10332 46126 10388
rect 47852 10332 49532 10388
rect 49588 10332 49598 10388
rect 49746 10332 49756 10388
rect 49812 10332 52220 10388
rect 52276 10332 52286 10388
rect 54450 10332 54460 10388
rect 54516 10332 55020 10388
rect 55076 10332 55086 10388
rect 56102 10332 56140 10388
rect 56196 10332 56206 10388
rect 22988 10276 23044 10332
rect 24332 10276 24388 10332
rect 242 10220 252 10276
rect 308 10220 1820 10276
rect 1876 10220 1886 10276
rect 2370 10220 2380 10276
rect 2436 10220 4172 10276
rect 4228 10220 4238 10276
rect 5068 10220 6076 10276
rect 6132 10220 6142 10276
rect 6262 10220 6300 10276
rect 6356 10220 6366 10276
rect 6636 10220 7196 10276
rect 7252 10220 7262 10276
rect 7970 10220 7980 10276
rect 8036 10220 8092 10276
rect 8148 10220 8158 10276
rect 9650 10220 9660 10276
rect 9716 10220 22820 10276
rect 22978 10220 22988 10276
rect 23044 10220 23054 10276
rect 23650 10220 23660 10276
rect 23716 10220 24388 10276
rect 25564 10276 25620 10332
rect 33516 10276 33572 10332
rect 25564 10220 26348 10276
rect 26404 10220 26414 10276
rect 28466 10220 28476 10276
rect 28532 10220 31948 10276
rect 32050 10220 32060 10276
rect 32116 10220 33572 10276
rect 35410 10220 35420 10276
rect 35476 10220 41132 10276
rect 41188 10220 41198 10276
rect 41916 10220 44268 10276
rect 44324 10220 44334 10276
rect 0 10164 112 10192
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 6636 10164 6692 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 0 10108 3388 10164
rect 5282 10108 5292 10164
rect 5348 10108 6692 10164
rect 6850 10108 6860 10164
rect 6916 10108 8876 10164
rect 8932 10108 8942 10164
rect 9538 10108 9548 10164
rect 9604 10108 11564 10164
rect 11620 10108 11630 10164
rect 11788 10108 13356 10164
rect 13412 10108 13422 10164
rect 14018 10108 14028 10164
rect 14084 10108 18676 10164
rect 19058 10108 19068 10164
rect 19124 10108 23212 10164
rect 23268 10108 23278 10164
rect 0 10080 112 10108
rect 3332 10052 3388 10108
rect 11788 10052 11844 10108
rect 3332 9996 8204 10052
rect 8260 9996 8270 10052
rect 9202 9996 9212 10052
rect 9268 9996 9436 10052
rect 9492 9996 9660 10052
rect 9716 9996 9726 10052
rect 10098 9996 10108 10052
rect 10164 9996 11004 10052
rect 11060 9996 11070 10052
rect 11442 9996 11452 10052
rect 11508 9996 11844 10052
rect 14690 9996 14700 10052
rect 14756 9996 15260 10052
rect 15316 9996 15326 10052
rect 15586 9996 15596 10052
rect 15652 9996 15876 10052
rect 16034 9996 16044 10052
rect 16100 9996 16492 10052
rect 16548 9996 18060 10052
rect 18116 9996 18126 10052
rect 15820 9940 15876 9996
rect 18620 9940 18676 10108
rect 31892 10052 31948 10220
rect 41916 10164 41972 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 33170 10108 33180 10164
rect 33236 10108 34300 10164
rect 34356 10108 34366 10164
rect 34514 10108 34524 10164
rect 34580 10108 35980 10164
rect 36036 10108 37212 10164
rect 37268 10108 37278 10164
rect 37538 10108 37548 10164
rect 37604 10108 41972 10164
rect 42102 10108 42140 10164
rect 42196 10108 42206 10164
rect 46386 10108 46396 10164
rect 46452 10108 47404 10164
rect 47460 10108 47470 10164
rect 47852 10052 47908 10332
rect 48850 10220 48860 10276
rect 48916 10220 50764 10276
rect 50820 10220 50830 10276
rect 57344 10164 57456 10192
rect 48066 10108 48076 10164
rect 48132 10108 48142 10164
rect 48514 10108 48524 10164
rect 48580 10108 49308 10164
rect 49364 10108 49374 10164
rect 49634 10108 49644 10164
rect 49700 10108 51660 10164
rect 51716 10108 51726 10164
rect 51874 10108 51884 10164
rect 51940 10108 53900 10164
rect 53956 10108 53966 10164
rect 54786 10108 54796 10164
rect 54852 10108 57456 10164
rect 19394 9996 19404 10052
rect 19460 9996 20188 10052
rect 20244 9996 21868 10052
rect 21924 9996 21934 10052
rect 22726 9996 22764 10052
rect 22820 9996 22830 10052
rect 26114 9996 26124 10052
rect 26180 9996 27356 10052
rect 27412 9996 27422 10052
rect 31892 9996 33964 10052
rect 34020 9996 34030 10052
rect 34402 9996 34412 10052
rect 34468 9996 35868 10052
rect 35924 9996 35934 10052
rect 41430 9996 41468 10052
rect 41524 9996 41534 10052
rect 43586 9996 43596 10052
rect 43652 9996 44492 10052
rect 44548 9996 45724 10052
rect 45780 9996 47908 10052
rect 48076 10052 48132 10108
rect 57344 10080 57456 10108
rect 48076 9996 50204 10052
rect 50260 9996 50270 10052
rect 51426 9996 51436 10052
rect 51492 9996 51996 10052
rect 52052 9996 52062 10052
rect 53442 9996 53452 10052
rect 53508 9996 53676 10052
rect 53732 9996 53742 10052
rect 56326 9996 56364 10052
rect 56420 9996 56430 10052
rect 3378 9884 3388 9940
rect 3444 9884 4732 9940
rect 4788 9884 8652 9940
rect 8708 9884 8718 9940
rect 9314 9884 9324 9940
rect 9380 9884 9884 9940
rect 9940 9884 9950 9940
rect 10770 9884 10780 9940
rect 10836 9884 11340 9940
rect 11396 9884 11406 9940
rect 12226 9884 12236 9940
rect 12292 9884 12796 9940
rect 12852 9884 12862 9940
rect 15820 9884 15988 9940
rect 16146 9884 16156 9940
rect 16212 9884 17724 9940
rect 17780 9884 17790 9940
rect 18620 9884 19404 9940
rect 19460 9884 21532 9940
rect 21588 9884 21598 9940
rect 21746 9884 21756 9940
rect 21812 9884 22092 9940
rect 22148 9884 27916 9940
rect 27972 9884 27982 9940
rect 28242 9884 28252 9940
rect 28308 9884 37212 9940
rect 37268 9884 37278 9940
rect 41794 9884 41804 9940
rect 41860 9884 44044 9940
rect 44100 9884 44110 9940
rect 44258 9884 44268 9940
rect 44324 9884 48972 9940
rect 49028 9884 49038 9940
rect 49382 9884 49420 9940
rect 49476 9884 49486 9940
rect 49746 9884 49756 9940
rect 49812 9884 54012 9940
rect 54068 9884 54078 9940
rect 15932 9828 15988 9884
rect 1484 9772 2156 9828
rect 2212 9772 2222 9828
rect 2454 9772 2492 9828
rect 2548 9772 2558 9828
rect 3938 9772 3948 9828
rect 4004 9772 4284 9828
rect 4340 9772 4350 9828
rect 5282 9772 5292 9828
rect 5348 9772 6412 9828
rect 6468 9772 6478 9828
rect 6738 9772 6748 9828
rect 6804 9772 7420 9828
rect 7476 9772 7486 9828
rect 7858 9772 7868 9828
rect 7924 9772 13580 9828
rect 13636 9772 13804 9828
rect 13860 9772 14588 9828
rect 14644 9772 14654 9828
rect 15932 9772 16828 9828
rect 16884 9772 16894 9828
rect 17266 9772 17276 9828
rect 17332 9772 18116 9828
rect 0 9716 112 9744
rect 1484 9716 1540 9772
rect 18060 9716 18116 9772
rect 20860 9772 21196 9828
rect 21252 9772 26684 9828
rect 26740 9772 26750 9828
rect 27458 9772 27468 9828
rect 27524 9772 29596 9828
rect 29652 9772 29662 9828
rect 31378 9772 31388 9828
rect 31444 9772 33404 9828
rect 33460 9772 33470 9828
rect 34626 9772 34636 9828
rect 34692 9772 34748 9828
rect 34804 9772 34814 9828
rect 35074 9772 35084 9828
rect 35140 9772 36876 9828
rect 36932 9772 36942 9828
rect 43026 9772 43036 9828
rect 43092 9772 43932 9828
rect 43988 9772 43998 9828
rect 44146 9772 44156 9828
rect 44212 9772 47068 9828
rect 47124 9772 47134 9828
rect 47842 9772 47852 9828
rect 47908 9772 48412 9828
rect 48468 9772 48478 9828
rect 49298 9772 49308 9828
rect 49364 9772 50764 9828
rect 50820 9772 52220 9828
rect 52276 9772 52286 9828
rect 20860 9716 20916 9772
rect 57344 9716 57456 9744
rect 0 9660 1540 9716
rect 1596 9660 9324 9716
rect 9380 9660 9390 9716
rect 9650 9660 9660 9716
rect 9716 9660 11452 9716
rect 11508 9660 11518 9716
rect 11676 9660 13132 9716
rect 13188 9660 13198 9716
rect 14476 9660 15316 9716
rect 16034 9660 16044 9716
rect 16100 9660 16940 9716
rect 16996 9660 17836 9716
rect 17892 9660 17902 9716
rect 18060 9660 18732 9716
rect 18788 9660 18798 9716
rect 19170 9660 19180 9716
rect 19236 9660 20916 9716
rect 24322 9660 24332 9716
rect 24388 9660 34412 9716
rect 34468 9660 34478 9716
rect 35634 9660 35644 9716
rect 35700 9660 47180 9716
rect 47236 9660 47246 9716
rect 47394 9660 47404 9716
rect 47460 9660 48188 9716
rect 48244 9660 48254 9716
rect 49186 9660 49196 9716
rect 49252 9660 55916 9716
rect 55972 9660 55982 9716
rect 56364 9660 57456 9716
rect 0 9632 112 9660
rect 0 9268 112 9296
rect 1596 9268 1652 9660
rect 11676 9604 11732 9660
rect 14476 9604 14532 9660
rect 2482 9548 2492 9604
rect 2548 9548 2716 9604
rect 2772 9548 2782 9604
rect 4274 9548 4284 9604
rect 4340 9548 6972 9604
rect 7028 9548 7868 9604
rect 7924 9548 7934 9604
rect 8306 9548 8316 9604
rect 8372 9548 8652 9604
rect 8708 9548 8718 9604
rect 9100 9548 11732 9604
rect 11890 9548 11900 9604
rect 11956 9548 12572 9604
rect 12628 9548 12638 9604
rect 13010 9548 13020 9604
rect 13076 9548 14532 9604
rect 15260 9604 15316 9660
rect 15260 9548 16100 9604
rect 16258 9548 16268 9604
rect 16324 9548 17500 9604
rect 17556 9548 26908 9604
rect 27682 9548 27692 9604
rect 27748 9548 31388 9604
rect 31444 9548 31454 9604
rect 31714 9548 31724 9604
rect 31780 9548 32396 9604
rect 32452 9548 36428 9604
rect 36484 9548 37212 9604
rect 37268 9548 37278 9604
rect 39442 9548 39452 9604
rect 39508 9548 45388 9604
rect 45444 9548 45454 9604
rect 47170 9548 47180 9604
rect 47236 9548 47964 9604
rect 48020 9548 48030 9604
rect 51762 9548 51772 9604
rect 51828 9548 52556 9604
rect 52612 9548 52622 9604
rect 9100 9492 9156 9548
rect 16044 9492 16100 9548
rect 26852 9492 26908 9548
rect 56364 9492 56420 9660
rect 57344 9632 57456 9660
rect 2482 9436 2492 9492
rect 2548 9436 3388 9492
rect 3444 9436 3454 9492
rect 4274 9436 4284 9492
rect 4340 9436 9156 9492
rect 9314 9436 9324 9492
rect 9380 9436 13804 9492
rect 13860 9436 13870 9492
rect 15250 9436 15260 9492
rect 15316 9436 15652 9492
rect 15782 9436 15820 9492
rect 15876 9436 15886 9492
rect 16044 9436 16492 9492
rect 16548 9436 16558 9492
rect 17826 9436 17836 9492
rect 17892 9436 22876 9492
rect 22932 9436 22942 9492
rect 26852 9436 32844 9492
rect 32900 9436 32910 9492
rect 33058 9436 33068 9492
rect 33124 9436 33134 9492
rect 33282 9436 33292 9492
rect 33348 9436 37268 9492
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 15596 9380 15652 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 4386 9324 4396 9380
rect 4452 9324 9660 9380
rect 9716 9324 9726 9380
rect 10994 9324 11004 9380
rect 11060 9324 11788 9380
rect 11844 9324 11854 9380
rect 13234 9324 13244 9380
rect 13300 9324 14644 9380
rect 15596 9324 16044 9380
rect 16100 9324 16110 9380
rect 16258 9324 16268 9380
rect 16324 9324 16604 9380
rect 16660 9324 16670 9380
rect 16930 9324 16940 9380
rect 16996 9324 19068 9380
rect 19124 9324 19134 9380
rect 20962 9324 20972 9380
rect 21028 9324 23660 9380
rect 23716 9324 23726 9380
rect 24322 9324 24332 9380
rect 24388 9324 26572 9380
rect 26628 9324 26638 9380
rect 26786 9324 26796 9380
rect 26852 9324 30044 9380
rect 30100 9324 30110 9380
rect 14588 9268 14644 9324
rect 33068 9268 33124 9436
rect 37212 9380 37268 9436
rect 38780 9436 40348 9492
rect 40404 9436 40414 9492
rect 44594 9436 44604 9492
rect 44660 9436 45052 9492
rect 45108 9436 45118 9492
rect 45378 9436 45388 9492
rect 45444 9436 56420 9492
rect 38780 9380 38836 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 35970 9324 35980 9380
rect 36036 9324 36316 9380
rect 36372 9324 36382 9380
rect 37212 9324 38780 9380
rect 38836 9324 38846 9380
rect 38994 9324 39004 9380
rect 39060 9324 41020 9380
rect 41076 9324 41086 9380
rect 42690 9324 42700 9380
rect 42756 9324 43484 9380
rect 43540 9324 43550 9380
rect 44146 9324 44156 9380
rect 44212 9324 52892 9380
rect 52948 9324 52958 9380
rect 57344 9268 57456 9296
rect 0 9212 476 9268
rect 532 9212 542 9268
rect 1484 9212 1652 9268
rect 2146 9212 2156 9268
rect 2212 9212 5068 9268
rect 5124 9212 5134 9268
rect 5506 9212 5516 9268
rect 5572 9212 6188 9268
rect 6244 9212 6254 9268
rect 6962 9212 6972 9268
rect 7028 9212 9100 9268
rect 9156 9212 9166 9268
rect 9426 9212 9436 9268
rect 9492 9212 9548 9268
rect 9604 9212 9614 9268
rect 9846 9212 9884 9268
rect 9940 9212 9950 9268
rect 10098 9212 10108 9268
rect 10164 9212 14364 9268
rect 14420 9212 14430 9268
rect 14588 9212 18396 9268
rect 18452 9212 18462 9268
rect 20738 9212 20748 9268
rect 20804 9212 21756 9268
rect 21812 9212 21822 9268
rect 23090 9212 23100 9268
rect 23156 9212 24220 9268
rect 24276 9212 26908 9268
rect 26964 9212 26974 9268
rect 28802 9212 28812 9268
rect 28868 9212 33124 9268
rect 33394 9212 33404 9268
rect 33460 9212 36764 9268
rect 36820 9212 36830 9268
rect 36978 9212 36988 9268
rect 37044 9212 39452 9268
rect 39508 9212 39518 9268
rect 43362 9212 43372 9268
rect 43428 9212 49308 9268
rect 49364 9212 49374 9268
rect 49970 9212 49980 9268
rect 50036 9212 50540 9268
rect 50596 9212 50606 9268
rect 50754 9212 50764 9268
rect 50820 9212 52332 9268
rect 52388 9212 53564 9268
rect 53620 9212 53630 9268
rect 54114 9212 54124 9268
rect 54180 9212 57456 9268
rect 0 9184 112 9212
rect 1222 8988 1260 9044
rect 1316 8988 1326 9044
rect 0 8820 112 8848
rect 1484 8820 1540 9212
rect 57344 9184 57456 9212
rect 1698 9100 1708 9156
rect 1764 9100 6636 9156
rect 6692 9100 6702 9156
rect 7746 9100 7756 9156
rect 7812 9100 52332 9156
rect 52388 9100 52398 9156
rect 53442 9100 53452 9156
rect 53508 9100 56028 9156
rect 56084 9100 56094 9156
rect 3332 8988 6748 9044
rect 6804 8988 6814 9044
rect 7298 8988 7308 9044
rect 7364 8988 7980 9044
rect 8036 8988 8046 9044
rect 8204 8988 14140 9044
rect 14196 8988 14206 9044
rect 14690 8988 14700 9044
rect 14756 8988 15596 9044
rect 15652 8988 16716 9044
rect 16772 8988 16782 9044
rect 17490 8988 17500 9044
rect 17556 8988 18620 9044
rect 18676 8988 18686 9044
rect 18834 8988 18844 9044
rect 18900 8988 22316 9044
rect 22372 8988 23436 9044
rect 23492 8988 23502 9044
rect 23650 8988 23660 9044
rect 23716 8988 27692 9044
rect 27748 8988 27758 9044
rect 27906 8988 27916 9044
rect 27972 8988 29036 9044
rect 29092 8988 29102 9044
rect 32806 8988 32844 9044
rect 32900 8988 32910 9044
rect 38434 8988 38444 9044
rect 38500 8988 38668 9044
rect 38724 8988 38734 9044
rect 39890 8988 39900 9044
rect 39956 8988 42588 9044
rect 42644 8988 46900 9044
rect 48178 8988 48188 9044
rect 48244 8988 50764 9044
rect 50820 8988 50830 9044
rect 52658 8988 52668 9044
rect 52724 8988 53340 9044
rect 53396 8988 53406 9044
rect 56354 8988 56364 9044
rect 56420 8988 57372 9044
rect 57428 8988 57438 9044
rect 3332 8932 3388 8988
rect 3042 8876 3052 8932
rect 3108 8876 3388 8932
rect 3490 8876 3500 8932
rect 3556 8876 3948 8932
rect 4004 8876 4014 8932
rect 4274 8876 4284 8932
rect 4340 8876 5180 8932
rect 5236 8876 5246 8932
rect 5842 8876 5852 8932
rect 5908 8876 6748 8932
rect 6804 8876 7868 8932
rect 7924 8876 7934 8932
rect 0 8764 1540 8820
rect 3602 8764 3612 8820
rect 3668 8764 5572 8820
rect 5730 8764 5740 8820
rect 5796 8764 6076 8820
rect 6132 8764 7420 8820
rect 7476 8764 7486 8820
rect 0 8736 112 8764
rect 5516 8708 5572 8764
rect 8204 8708 8260 8988
rect 8642 8876 8652 8932
rect 8708 8876 43036 8932
rect 43092 8876 43102 8932
rect 44034 8876 44044 8932
rect 44100 8876 44828 8932
rect 44884 8876 44894 8932
rect 46844 8820 46900 8988
rect 47170 8876 47180 8932
rect 47236 8876 48076 8932
rect 48132 8876 48142 8932
rect 53330 8876 53340 8932
rect 53396 8876 53564 8932
rect 53620 8876 53630 8932
rect 57344 8820 57456 8848
rect 8418 8764 8428 8820
rect 8484 8764 11004 8820
rect 11060 8764 11070 8820
rect 11554 8764 11564 8820
rect 11620 8764 15708 8820
rect 15764 8764 15774 8820
rect 18844 8764 43372 8820
rect 43428 8764 43438 8820
rect 43596 8764 45164 8820
rect 45220 8764 45230 8820
rect 46834 8764 46844 8820
rect 46900 8764 46910 8820
rect 49522 8764 49532 8820
rect 49588 8764 50316 8820
rect 50372 8764 50382 8820
rect 52210 8764 52220 8820
rect 52276 8764 52668 8820
rect 52724 8764 52734 8820
rect 53218 8764 53228 8820
rect 53284 8764 53788 8820
rect 53844 8764 54348 8820
rect 54404 8764 54414 8820
rect 54572 8764 57456 8820
rect 18844 8708 18900 8764
rect 43596 8708 43652 8764
rect 54572 8708 54628 8764
rect 57344 8736 57456 8764
rect 5058 8652 5068 8708
rect 5124 8652 5292 8708
rect 5348 8652 5358 8708
rect 5516 8652 8260 8708
rect 9314 8652 9324 8708
rect 9380 8652 18900 8708
rect 19842 8652 19852 8708
rect 19908 8652 23660 8708
rect 23716 8652 23726 8708
rect 26646 8652 26684 8708
rect 26740 8652 26750 8708
rect 30370 8652 30380 8708
rect 30436 8652 38668 8708
rect 38724 8652 40236 8708
rect 40292 8652 40302 8708
rect 41010 8652 41020 8708
rect 41076 8652 43652 8708
rect 44930 8652 44940 8708
rect 44996 8652 49980 8708
rect 50036 8652 50046 8708
rect 50530 8652 50540 8708
rect 50596 8652 54628 8708
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 2706 8540 2716 8596
rect 2772 8540 4284 8596
rect 4340 8540 4350 8596
rect 4946 8540 4956 8596
rect 5012 8540 13356 8596
rect 13412 8540 13422 8596
rect 13570 8540 13580 8596
rect 13636 8540 18060 8596
rect 18116 8540 18126 8596
rect 18610 8540 18620 8596
rect 18676 8540 24332 8596
rect 24388 8540 24398 8596
rect 26562 8540 26572 8596
rect 26628 8540 30604 8596
rect 30660 8540 32172 8596
rect 32228 8540 32238 8596
rect 33394 8540 33404 8596
rect 33460 8540 34636 8596
rect 34692 8540 34702 8596
rect 35644 8540 40908 8596
rect 40964 8540 40974 8596
rect 41122 8540 41132 8596
rect 41188 8540 44268 8596
rect 44324 8540 44334 8596
rect 48626 8540 48636 8596
rect 48692 8540 48972 8596
rect 49028 8540 49038 8596
rect 50372 8540 55468 8596
rect 55524 8540 55534 8596
rect 35644 8484 35700 8540
rect 50372 8484 50428 8540
rect 2034 8428 2044 8484
rect 2100 8428 3052 8484
rect 3108 8428 3118 8484
rect 4060 8428 5628 8484
rect 5684 8428 5694 8484
rect 6290 8428 6300 8484
rect 6356 8428 6636 8484
rect 6692 8428 6702 8484
rect 8092 8428 12796 8484
rect 12852 8428 12862 8484
rect 13234 8428 13244 8484
rect 13300 8428 14252 8484
rect 14308 8428 14318 8484
rect 14466 8428 14476 8484
rect 14532 8428 18060 8484
rect 18116 8428 18126 8484
rect 18386 8428 18396 8484
rect 18452 8428 19180 8484
rect 19236 8428 19246 8484
rect 19740 8428 20804 8484
rect 21298 8428 21308 8484
rect 21364 8428 23100 8484
rect 23156 8428 28588 8484
rect 28644 8428 28654 8484
rect 30482 8428 30492 8484
rect 30548 8428 32620 8484
rect 32676 8428 32686 8484
rect 33506 8428 33516 8484
rect 33572 8428 35700 8484
rect 35756 8428 50428 8484
rect 52770 8428 52780 8484
rect 52836 8428 53900 8484
rect 53956 8428 53966 8484
rect 0 8372 112 8400
rect 0 8316 812 8372
rect 868 8316 878 8372
rect 1586 8316 1596 8372
rect 1652 8316 3612 8372
rect 3668 8316 3678 8372
rect 0 8288 112 8316
rect 4060 8260 4116 8428
rect 5282 8316 5292 8372
rect 5348 8316 6524 8372
rect 6580 8316 6590 8372
rect 2034 8204 2044 8260
rect 2100 8204 3164 8260
rect 3220 8204 4116 8260
rect 4274 8204 4284 8260
rect 4340 8204 4508 8260
rect 4564 8204 4574 8260
rect 5170 8204 5180 8260
rect 5236 8204 5516 8260
rect 5572 8204 5582 8260
rect 5954 8204 5964 8260
rect 6020 8204 6972 8260
rect 7028 8204 7038 8260
rect 8092 8148 8148 8428
rect 19740 8372 19796 8428
rect 20748 8372 20804 8428
rect 12562 8316 12572 8372
rect 12628 8316 13468 8372
rect 13524 8316 13534 8372
rect 14914 8316 14924 8372
rect 14980 8316 16940 8372
rect 16996 8316 17006 8372
rect 17164 8316 18452 8372
rect 18610 8316 18620 8372
rect 18676 8316 19796 8372
rect 19954 8316 19964 8372
rect 20020 8316 20524 8372
rect 20580 8316 20590 8372
rect 20748 8316 21196 8372
rect 21252 8316 21262 8372
rect 23314 8316 23324 8372
rect 23380 8316 23548 8372
rect 23604 8316 23614 8372
rect 25442 8316 25452 8372
rect 25508 8316 26124 8372
rect 26180 8316 26190 8372
rect 26338 8316 26348 8372
rect 26404 8316 31612 8372
rect 31668 8316 31678 8372
rect 31826 8316 31836 8372
rect 31892 8316 32396 8372
rect 32452 8316 34188 8372
rect 34244 8316 34254 8372
rect 17164 8260 17220 8316
rect 8642 8204 8652 8260
rect 8708 8204 9548 8260
rect 9604 8204 9614 8260
rect 10294 8204 10332 8260
rect 10388 8204 10398 8260
rect 10882 8204 10892 8260
rect 10948 8204 11900 8260
rect 11956 8204 11966 8260
rect 14690 8204 14700 8260
rect 14756 8204 15596 8260
rect 15652 8204 16268 8260
rect 16324 8204 16334 8260
rect 16818 8204 16828 8260
rect 16884 8204 17220 8260
rect 17350 8204 17388 8260
rect 17444 8204 17454 8260
rect 17938 8204 17948 8260
rect 18004 8204 18060 8260
rect 18116 8204 18126 8260
rect 18396 8148 18452 8316
rect 32732 8260 32788 8316
rect 19058 8204 19068 8260
rect 19124 8204 20972 8260
rect 21028 8204 22316 8260
rect 22372 8204 22382 8260
rect 23436 8204 23884 8260
rect 23940 8204 24332 8260
rect 24388 8204 24398 8260
rect 24994 8204 25004 8260
rect 25060 8204 26012 8260
rect 26068 8204 26078 8260
rect 26674 8204 26684 8260
rect 26740 8204 27468 8260
rect 27524 8204 27534 8260
rect 27906 8204 27916 8260
rect 27972 8204 29820 8260
rect 29876 8204 29886 8260
rect 30370 8204 30380 8260
rect 30436 8204 31388 8260
rect 31444 8204 31454 8260
rect 31724 8204 32284 8260
rect 32340 8204 32508 8260
rect 32564 8204 32574 8260
rect 32722 8204 32732 8260
rect 32788 8204 32798 8260
rect 33730 8204 33740 8260
rect 33796 8204 34412 8260
rect 34468 8204 34478 8260
rect 23436 8148 23492 8204
rect 31724 8148 31780 8204
rect 1698 8092 1708 8148
rect 1764 8092 8148 8148
rect 8204 8092 9884 8148
rect 9940 8092 9950 8148
rect 10658 8092 10668 8148
rect 10724 8092 11564 8148
rect 11620 8092 11630 8148
rect 14578 8092 14588 8148
rect 14644 8092 14700 8148
rect 14756 8092 17612 8148
rect 17668 8092 18060 8148
rect 18116 8092 18126 8148
rect 18396 8092 19852 8148
rect 19908 8092 19918 8148
rect 20066 8092 20076 8148
rect 20132 8092 22764 8148
rect 22820 8092 23492 8148
rect 23548 8092 25452 8148
rect 25508 8092 25518 8148
rect 25676 8092 27356 8148
rect 27412 8092 31780 8148
rect 31938 8092 31948 8148
rect 32004 8092 33180 8148
rect 33236 8092 33246 8148
rect 34402 8092 34412 8148
rect 34468 8092 35420 8148
rect 35476 8092 35486 8148
rect 8204 8036 8260 8092
rect 23548 8036 23604 8092
rect 25676 8036 25732 8092
rect 1474 7980 1484 8036
rect 1540 7980 1596 8036
rect 1652 7980 1662 8036
rect 1810 7980 1820 8036
rect 1876 7980 3388 8036
rect 3444 7980 3454 8036
rect 3602 7980 3612 8036
rect 3668 7980 6300 8036
rect 6356 7980 6366 8036
rect 6738 7980 6748 8036
rect 6804 7980 8260 8036
rect 11778 7980 11788 8036
rect 11844 7980 23604 8036
rect 23660 7980 25676 8036
rect 25732 7980 25742 8036
rect 25890 7980 25900 8036
rect 25956 7980 26908 8036
rect 28578 7980 28588 8036
rect 28644 7980 30772 8036
rect 31714 7980 31724 8036
rect 31780 7980 32844 8036
rect 32900 7980 33852 8036
rect 33908 7980 33918 8036
rect 0 7924 112 7952
rect 23660 7924 23716 7980
rect 0 7868 3388 7924
rect 4162 7868 4172 7924
rect 4228 7868 7532 7924
rect 7588 7868 7598 7924
rect 7746 7868 7756 7924
rect 7812 7868 9100 7924
rect 9156 7868 10556 7924
rect 10612 7868 12068 7924
rect 12226 7868 12236 7924
rect 12292 7868 23716 7924
rect 26852 7924 26908 7980
rect 30716 7924 30772 7980
rect 35756 7924 35812 8428
rect 57344 8372 57456 8400
rect 37650 8316 37660 8372
rect 37716 8316 38332 8372
rect 38388 8316 38398 8372
rect 38612 8316 39900 8372
rect 39956 8316 39966 8372
rect 41570 8316 41580 8372
rect 41636 8316 41804 8372
rect 41860 8316 41870 8372
rect 42438 8316 42476 8372
rect 42532 8316 42542 8372
rect 43026 8316 43036 8372
rect 43092 8316 47516 8372
rect 47572 8316 47582 8372
rect 50978 8316 50988 8372
rect 51044 8316 54124 8372
rect 54180 8316 54190 8372
rect 55692 8316 57456 8372
rect 36306 8204 36316 8260
rect 36372 8204 37772 8260
rect 37828 8204 37838 8260
rect 38612 8148 38668 8316
rect 41010 8204 41020 8260
rect 41076 8204 43820 8260
rect 43876 8204 43886 8260
rect 47926 8204 47964 8260
rect 48020 8204 48030 8260
rect 50978 8204 50988 8260
rect 51044 8204 52892 8260
rect 52948 8204 52958 8260
rect 55692 8148 55748 8316
rect 57344 8288 57456 8316
rect 56354 8204 56364 8260
rect 56420 8204 57148 8260
rect 57204 8204 57214 8260
rect 36866 8092 36876 8148
rect 36932 8092 38668 8148
rect 43138 8092 43148 8148
rect 43204 8092 43932 8148
rect 43988 8092 43998 8148
rect 46956 8092 50652 8148
rect 50708 8092 51996 8148
rect 52052 8092 52062 8148
rect 52322 8092 52332 8148
rect 52388 8092 55748 8148
rect 40786 7980 40796 8036
rect 40852 7980 41356 8036
rect 41412 7980 44044 8036
rect 44100 7980 44110 8036
rect 46956 7924 47012 8092
rect 47730 7980 47740 8036
rect 47796 7980 48188 8036
rect 48244 7980 48254 8036
rect 49858 7980 49868 8036
rect 49924 7980 50316 8036
rect 50372 7980 51156 8036
rect 51874 7980 51884 8036
rect 51940 7980 54796 8036
rect 54852 7980 54862 8036
rect 51100 7924 51156 7980
rect 57344 7924 57456 7952
rect 26852 7868 30156 7924
rect 30212 7868 30222 7924
rect 30706 7868 30716 7924
rect 30772 7868 32060 7924
rect 32116 7868 32126 7924
rect 32274 7868 32284 7924
rect 32340 7868 35812 7924
rect 41682 7868 41692 7924
rect 41748 7868 43596 7924
rect 43652 7868 43662 7924
rect 45826 7868 45836 7924
rect 45892 7868 46956 7924
rect 47012 7868 47022 7924
rect 47170 7868 47180 7924
rect 47236 7868 50764 7924
rect 50820 7868 50830 7924
rect 51090 7868 51100 7924
rect 51156 7868 52220 7924
rect 52276 7868 53340 7924
rect 53396 7868 53406 7924
rect 53666 7868 53676 7924
rect 53732 7868 57456 7924
rect 0 7840 112 7868
rect 2594 7756 2604 7812
rect 2660 7756 2670 7812
rect 2604 7588 2660 7756
rect 3332 7700 3388 7868
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 12012 7812 12068 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 57344 7840 57456 7868
rect 6402 7756 6412 7812
rect 6468 7756 11788 7812
rect 11844 7756 11854 7812
rect 12012 7756 14364 7812
rect 14420 7756 14430 7812
rect 14914 7756 14924 7812
rect 14980 7756 15372 7812
rect 15428 7756 15438 7812
rect 16034 7756 16044 7812
rect 16100 7756 16828 7812
rect 16884 7756 16894 7812
rect 17042 7756 17052 7812
rect 17108 7756 17612 7812
rect 17668 7756 17678 7812
rect 19282 7756 19292 7812
rect 19348 7756 20636 7812
rect 20692 7756 20702 7812
rect 25442 7756 25452 7812
rect 25508 7756 27020 7812
rect 27076 7756 27086 7812
rect 27794 7756 27804 7812
rect 27860 7756 30380 7812
rect 30436 7756 30446 7812
rect 32050 7756 32060 7812
rect 32116 7756 33740 7812
rect 33796 7756 33806 7812
rect 34076 7756 40460 7812
rect 40516 7756 40526 7812
rect 44146 7756 44156 7812
rect 44212 7756 44828 7812
rect 44884 7756 45612 7812
rect 45668 7756 46508 7812
rect 46564 7756 48300 7812
rect 48356 7756 48366 7812
rect 48850 7756 48860 7812
rect 48916 7756 56028 7812
rect 56084 7756 56094 7812
rect 34076 7700 34132 7756
rect 2818 7644 2828 7700
rect 2884 7644 3164 7700
rect 3220 7644 3230 7700
rect 3332 7644 6300 7700
rect 6356 7644 6366 7700
rect 8418 7644 8428 7700
rect 8484 7644 13132 7700
rect 13188 7644 13198 7700
rect 13458 7644 13468 7700
rect 13524 7644 24668 7700
rect 24724 7644 24734 7700
rect 26114 7644 26124 7700
rect 26180 7644 26684 7700
rect 26740 7644 27132 7700
rect 27188 7644 27198 7700
rect 30034 7644 30044 7700
rect 30100 7644 34132 7700
rect 37090 7644 37100 7700
rect 37156 7644 40236 7700
rect 40292 7644 40302 7700
rect 40450 7644 40460 7700
rect 40516 7644 44268 7700
rect 44324 7644 45836 7700
rect 45892 7644 45902 7700
rect 48290 7644 48300 7700
rect 48356 7644 49868 7700
rect 49924 7644 49934 7700
rect 51426 7644 51436 7700
rect 51492 7644 53004 7700
rect 53060 7644 53070 7700
rect 53330 7644 53340 7700
rect 53396 7644 56588 7700
rect 56644 7644 56654 7700
rect 466 7532 476 7588
rect 532 7532 5684 7588
rect 6374 7532 6412 7588
rect 6468 7532 6478 7588
rect 8194 7532 8204 7588
rect 8260 7532 8652 7588
rect 8708 7532 8718 7588
rect 10098 7532 10108 7588
rect 10164 7532 12012 7588
rect 12068 7532 14812 7588
rect 14868 7532 14878 7588
rect 15026 7532 15036 7588
rect 15092 7532 16492 7588
rect 16548 7532 16558 7588
rect 16706 7532 16716 7588
rect 16772 7532 22204 7588
rect 22260 7532 22270 7588
rect 23314 7532 23324 7588
rect 23380 7532 25116 7588
rect 25172 7532 25182 7588
rect 25340 7532 26684 7588
rect 26740 7532 26750 7588
rect 26852 7532 27804 7588
rect 27860 7532 27870 7588
rect 32498 7532 32508 7588
rect 32564 7532 33516 7588
rect 33572 7532 33582 7588
rect 33740 7532 53564 7588
rect 53620 7532 53630 7588
rect 0 7476 112 7504
rect 5628 7476 5684 7532
rect 25340 7476 25396 7532
rect 26852 7476 26908 7532
rect 33740 7476 33796 7532
rect 57344 7476 57456 7504
rect 0 7420 2268 7476
rect 2324 7420 2334 7476
rect 3938 7420 3948 7476
rect 4004 7420 4956 7476
rect 5012 7420 5022 7476
rect 5618 7420 5628 7476
rect 5684 7420 6524 7476
rect 6580 7420 6590 7476
rect 8530 7420 8540 7476
rect 8596 7420 9660 7476
rect 9716 7420 9726 7476
rect 9986 7420 9996 7476
rect 10052 7420 10108 7476
rect 10164 7420 10174 7476
rect 10546 7420 10556 7476
rect 10612 7420 11676 7476
rect 11732 7420 11742 7476
rect 11890 7420 11900 7476
rect 11956 7420 12348 7476
rect 12404 7420 12414 7476
rect 13542 7420 13580 7476
rect 13636 7420 16156 7476
rect 16212 7420 19292 7476
rect 19348 7420 19358 7476
rect 19842 7420 19852 7476
rect 19908 7420 20972 7476
rect 21028 7420 21038 7476
rect 21186 7420 21196 7476
rect 21252 7420 25396 7476
rect 25890 7420 25900 7476
rect 25956 7420 26908 7476
rect 29148 7420 30940 7476
rect 30996 7420 31006 7476
rect 31378 7420 31388 7476
rect 31444 7420 33796 7476
rect 34850 7420 34860 7476
rect 34916 7420 35868 7476
rect 35924 7420 35934 7476
rect 38434 7420 38444 7476
rect 38500 7420 39340 7476
rect 39396 7420 39406 7476
rect 39862 7420 39900 7476
rect 39956 7420 39966 7476
rect 40226 7420 40236 7476
rect 40292 7420 47180 7476
rect 47236 7420 47246 7476
rect 48290 7420 48300 7476
rect 48356 7420 51548 7476
rect 51604 7420 51614 7476
rect 53004 7420 57456 7476
rect 0 7392 112 7420
rect 29148 7364 29204 7420
rect 242 7308 252 7364
rect 308 7308 3612 7364
rect 3668 7308 3678 7364
rect 4162 7308 4172 7364
rect 4228 7308 4396 7364
rect 4452 7308 14252 7364
rect 14308 7308 14318 7364
rect 14466 7308 14476 7364
rect 14532 7308 14924 7364
rect 14980 7308 14990 7364
rect 15810 7308 15820 7364
rect 15876 7308 16492 7364
rect 16548 7308 17388 7364
rect 17444 7308 17454 7364
rect 19852 7308 20188 7364
rect 20244 7308 20254 7364
rect 24658 7308 24668 7364
rect 24724 7308 29204 7364
rect 30258 7308 30268 7364
rect 30324 7308 31948 7364
rect 32004 7308 32014 7364
rect 33170 7308 33180 7364
rect 33236 7308 41244 7364
rect 41300 7308 41580 7364
rect 41636 7308 41646 7364
rect 42018 7308 42028 7364
rect 42084 7308 42140 7364
rect 42196 7308 42206 7364
rect 42354 7308 42364 7364
rect 42420 7308 44828 7364
rect 44884 7308 48860 7364
rect 48916 7308 48926 7364
rect 51090 7308 51100 7364
rect 51156 7308 52556 7364
rect 52612 7308 52622 7364
rect 19852 7252 19908 7308
rect 354 7196 364 7252
rect 420 7196 1260 7252
rect 1316 7196 1326 7252
rect 4834 7196 4844 7252
rect 4900 7196 7644 7252
rect 7700 7196 7710 7252
rect 8306 7196 8316 7252
rect 8372 7196 8652 7252
rect 8708 7196 8718 7252
rect 8978 7196 8988 7252
rect 9044 7196 9054 7252
rect 9314 7196 9324 7252
rect 9380 7196 14028 7252
rect 14084 7196 14094 7252
rect 14354 7196 14364 7252
rect 14420 7196 16268 7252
rect 16324 7196 19908 7252
rect 20066 7196 20076 7252
rect 20132 7196 21644 7252
rect 21700 7196 21710 7252
rect 21868 7196 44884 7252
rect 8988 7140 9044 7196
rect 21868 7140 21924 7196
rect 1474 7084 1484 7140
rect 1540 7084 4116 7140
rect 4274 7084 4284 7140
rect 4340 7084 4350 7140
rect 4946 7084 4956 7140
rect 5012 7084 5404 7140
rect 5460 7084 5470 7140
rect 5618 7084 5628 7140
rect 5684 7084 9044 7140
rect 9314 7084 9324 7140
rect 9380 7084 11116 7140
rect 11172 7084 11182 7140
rect 12450 7084 12460 7140
rect 12516 7084 13244 7140
rect 13300 7084 14476 7140
rect 14532 7084 14542 7140
rect 17938 7084 17948 7140
rect 18004 7084 20860 7140
rect 20916 7084 21924 7140
rect 26450 7084 26460 7140
rect 26516 7084 32508 7140
rect 32564 7084 32574 7140
rect 32722 7084 32732 7140
rect 32788 7084 37548 7140
rect 37604 7084 37614 7140
rect 38210 7084 38220 7140
rect 38276 7084 41580 7140
rect 41636 7084 41646 7140
rect 41794 7084 41804 7140
rect 41860 7084 42924 7140
rect 42980 7084 44156 7140
rect 44212 7084 44222 7140
rect 0 7028 112 7056
rect 0 6972 700 7028
rect 756 6972 766 7028
rect 3350 6972 3388 7028
rect 3444 6972 3454 7028
rect 0 6944 112 6972
rect 1138 6860 1148 6916
rect 1204 6860 1484 6916
rect 1540 6860 1550 6916
rect 4060 6804 4116 7084
rect 4284 6916 4340 7084
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 41804 7028 41860 7084
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 44828 7028 44884 7196
rect 46610 7084 46620 7140
rect 46676 7084 51324 7140
rect 51380 7084 51390 7140
rect 53004 7028 53060 7420
rect 57344 7392 57456 7420
rect 53218 7196 53228 7252
rect 53284 7196 53788 7252
rect 53844 7196 53854 7252
rect 56242 7084 56252 7140
rect 56308 7084 56318 7140
rect 5282 6972 5292 7028
rect 5348 6972 5404 7028
rect 5460 6972 5470 7028
rect 7186 6972 7196 7028
rect 7252 6972 14364 7028
rect 14420 6972 14430 7028
rect 15922 6972 15932 7028
rect 15988 6972 22876 7028
rect 22932 6972 22942 7028
rect 25106 6972 25116 7028
rect 25172 6972 30268 7028
rect 30324 6972 30334 7028
rect 33506 6972 33516 7028
rect 33572 6972 34356 7028
rect 34514 6972 34524 7028
rect 34580 6972 36316 7028
rect 36372 6972 36382 7028
rect 36540 6972 36652 7028
rect 36708 6972 41860 7028
rect 44828 6972 53060 7028
rect 56252 7028 56308 7084
rect 57344 7028 57456 7056
rect 56252 6972 57456 7028
rect 34300 6916 34356 6972
rect 36540 6916 36596 6972
rect 57344 6944 57456 6972
rect 4284 6860 6412 6916
rect 6468 6860 6478 6916
rect 6636 6860 7980 6916
rect 8036 6860 8046 6916
rect 8194 6860 8204 6916
rect 8260 6860 8876 6916
rect 8932 6860 8942 6916
rect 10770 6860 10780 6916
rect 10836 6860 13580 6916
rect 13636 6860 13646 6916
rect 13794 6860 13804 6916
rect 13860 6860 31836 6916
rect 31892 6860 31902 6916
rect 33058 6860 33068 6916
rect 33124 6860 33628 6916
rect 33684 6860 33694 6916
rect 34300 6860 35420 6916
rect 35476 6860 35486 6916
rect 35858 6860 35868 6916
rect 35924 6860 36596 6916
rect 37314 6860 37324 6916
rect 37380 6860 42252 6916
rect 42308 6860 42924 6916
rect 42980 6860 45724 6916
rect 45780 6860 45790 6916
rect 45938 6860 45948 6916
rect 46004 6860 46620 6916
rect 46676 6860 46686 6916
rect 54086 6860 54124 6916
rect 54180 6860 54190 6916
rect 6636 6804 6692 6860
rect 1362 6748 1372 6804
rect 1428 6748 1932 6804
rect 1988 6748 3388 6804
rect 4060 6748 6692 6804
rect 7074 6748 7084 6804
rect 7140 6748 9100 6804
rect 9156 6748 9166 6804
rect 11218 6748 11228 6804
rect 11284 6748 14588 6804
rect 14644 6748 14654 6804
rect 15250 6748 15260 6804
rect 15316 6748 15932 6804
rect 15988 6748 15998 6804
rect 18050 6748 18060 6804
rect 18116 6748 20076 6804
rect 20132 6748 20142 6804
rect 21970 6748 21980 6804
rect 22036 6748 22204 6804
rect 22260 6748 22270 6804
rect 23538 6748 23548 6804
rect 23604 6748 25116 6804
rect 25172 6748 25182 6804
rect 26898 6748 26908 6804
rect 26964 6748 30492 6804
rect 30548 6748 30558 6804
rect 33058 6748 33068 6804
rect 33124 6748 34748 6804
rect 34804 6748 35028 6804
rect 35186 6748 35196 6804
rect 35252 6748 35644 6804
rect 35700 6748 35710 6804
rect 36306 6748 36316 6804
rect 36372 6748 38220 6804
rect 38276 6748 38286 6804
rect 38434 6748 38444 6804
rect 38500 6748 41356 6804
rect 41412 6748 41422 6804
rect 41570 6748 41580 6804
rect 41636 6748 42364 6804
rect 42420 6748 45444 6804
rect 45602 6748 45612 6804
rect 45668 6748 46284 6804
rect 46340 6748 46350 6804
rect 3332 6692 3388 6748
rect 34972 6692 35028 6748
rect 40796 6692 40852 6748
rect 3332 6636 4452 6692
rect 4610 6636 4620 6692
rect 4676 6636 8876 6692
rect 8932 6636 8942 6692
rect 9090 6636 9100 6692
rect 9156 6636 9212 6692
rect 9268 6636 9996 6692
rect 10052 6636 10062 6692
rect 11778 6636 11788 6692
rect 11844 6636 15372 6692
rect 15428 6636 15438 6692
rect 15698 6636 15708 6692
rect 15764 6636 16604 6692
rect 16660 6636 16670 6692
rect 17042 6636 17052 6692
rect 17108 6636 18284 6692
rect 18340 6636 18620 6692
rect 18676 6636 18686 6692
rect 19170 6636 19180 6692
rect 19236 6636 19852 6692
rect 19908 6636 20188 6692
rect 20244 6636 20254 6692
rect 20626 6636 20636 6692
rect 20692 6636 24332 6692
rect 24388 6636 24398 6692
rect 24854 6636 24892 6692
rect 24948 6636 24958 6692
rect 25218 6636 25228 6692
rect 25284 6636 25900 6692
rect 25956 6636 25966 6692
rect 27122 6636 27132 6692
rect 27188 6636 27692 6692
rect 27748 6636 27758 6692
rect 28326 6636 28364 6692
rect 28420 6636 28430 6692
rect 29362 6636 29372 6692
rect 29428 6636 31388 6692
rect 31444 6636 31454 6692
rect 31612 6636 33404 6692
rect 33460 6636 33470 6692
rect 33618 6636 33628 6692
rect 33684 6636 34916 6692
rect 34972 6636 35532 6692
rect 35588 6636 35598 6692
rect 39554 6636 39564 6692
rect 39620 6636 40572 6692
rect 40628 6636 40638 6692
rect 40786 6636 40796 6692
rect 40852 6636 40862 6692
rect 41570 6636 41580 6692
rect 41636 6636 43036 6692
rect 43092 6636 44380 6692
rect 44436 6636 44446 6692
rect 0 6580 112 6608
rect 4396 6580 4452 6636
rect 31612 6580 31668 6636
rect 34860 6580 34916 6636
rect 0 6524 2828 6580
rect 2884 6524 2894 6580
rect 4396 6524 5516 6580
rect 5572 6524 5582 6580
rect 6626 6524 6636 6580
rect 6692 6524 6972 6580
rect 7028 6524 7868 6580
rect 7924 6524 9100 6580
rect 9156 6524 9166 6580
rect 10322 6524 10332 6580
rect 10388 6524 11452 6580
rect 11508 6524 11518 6580
rect 11890 6524 11900 6580
rect 11956 6524 14700 6580
rect 14756 6524 14766 6580
rect 15586 6524 15596 6580
rect 15652 6524 16940 6580
rect 16996 6524 17006 6580
rect 17154 6524 17164 6580
rect 17220 6524 19516 6580
rect 19572 6524 19582 6580
rect 19730 6524 19740 6580
rect 19796 6524 21756 6580
rect 21812 6524 21822 6580
rect 23426 6524 23436 6580
rect 23492 6524 23996 6580
rect 24052 6524 29484 6580
rect 29540 6524 31668 6580
rect 33142 6524 33180 6580
rect 33236 6524 33246 6580
rect 33506 6524 33516 6580
rect 33572 6524 34188 6580
rect 34244 6524 34636 6580
rect 34692 6524 34702 6580
rect 34860 6524 39788 6580
rect 39844 6524 39854 6580
rect 40114 6524 40124 6580
rect 40180 6524 40236 6580
rect 40292 6524 40302 6580
rect 40450 6524 40460 6580
rect 40516 6524 44268 6580
rect 44324 6524 44334 6580
rect 0 6496 112 6524
rect 45388 6468 45444 6748
rect 45714 6636 45724 6692
rect 45780 6636 50540 6692
rect 50596 6636 50652 6692
rect 50708 6636 50718 6692
rect 53554 6636 53564 6692
rect 53620 6636 55916 6692
rect 55972 6636 55982 6692
rect 57344 6580 57456 6608
rect 47170 6524 47180 6580
rect 47236 6524 53340 6580
rect 53396 6524 53406 6580
rect 53666 6524 53676 6580
rect 53732 6524 53742 6580
rect 55458 6524 55468 6580
rect 55524 6524 57456 6580
rect 53676 6468 53732 6524
rect 57344 6496 57456 6524
rect 2370 6412 2380 6468
rect 2436 6412 4172 6468
rect 4228 6412 4238 6468
rect 5142 6412 5180 6468
rect 5236 6412 5852 6468
rect 5908 6412 5918 6468
rect 6402 6412 6412 6468
rect 6468 6412 7308 6468
rect 7364 6412 7374 6468
rect 8642 6412 8652 6468
rect 8708 6412 9716 6468
rect 10658 6412 10668 6468
rect 10724 6412 11116 6468
rect 11172 6412 11182 6468
rect 11666 6412 11676 6468
rect 11732 6412 14252 6468
rect 14308 6412 14318 6468
rect 15036 6412 18732 6468
rect 18788 6412 18798 6468
rect 23660 6412 25452 6468
rect 25508 6412 25518 6468
rect 26226 6412 26236 6468
rect 26292 6412 26460 6468
rect 26516 6412 26526 6468
rect 31714 6412 31724 6468
rect 31780 6412 32508 6468
rect 32564 6412 35084 6468
rect 35140 6412 35196 6468
rect 35252 6412 35262 6468
rect 36530 6412 36540 6468
rect 36596 6412 41020 6468
rect 41076 6412 41086 6468
rect 42130 6412 42140 6468
rect 42196 6412 44324 6468
rect 44482 6412 44492 6468
rect 44548 6412 44940 6468
rect 44996 6412 45006 6468
rect 45388 6412 52780 6468
rect 52836 6412 52846 6468
rect 53676 6412 54460 6468
rect 54516 6412 56252 6468
rect 56308 6412 56318 6468
rect 1362 6300 1372 6356
rect 1428 6300 3388 6356
rect 3444 6300 3454 6356
rect 4274 6300 4284 6356
rect 4340 6300 5292 6356
rect 5348 6300 5628 6356
rect 5684 6300 5694 6356
rect 6178 6300 6188 6356
rect 6244 6300 6636 6356
rect 6692 6300 6702 6356
rect 6962 6300 6972 6356
rect 7028 6300 7084 6356
rect 7140 6300 8148 6356
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 8092 6244 8148 6300
rect 9660 6244 9716 6412
rect 9874 6300 9884 6356
rect 9940 6300 12236 6356
rect 12292 6300 12302 6356
rect 15036 6244 15092 6412
rect 23660 6356 23716 6412
rect 26236 6356 26292 6412
rect 44268 6356 44324 6412
rect 15250 6300 15260 6356
rect 15316 6300 15596 6356
rect 15652 6300 15662 6356
rect 15922 6300 15932 6356
rect 15988 6300 18508 6356
rect 18564 6300 18574 6356
rect 18946 6300 18956 6356
rect 19012 6300 23716 6356
rect 24322 6300 24332 6356
rect 24388 6300 26292 6356
rect 26348 6300 33068 6356
rect 33124 6300 33134 6356
rect 33282 6300 33292 6356
rect 33348 6300 34748 6356
rect 34804 6300 34814 6356
rect 34962 6300 34972 6356
rect 35028 6300 36428 6356
rect 36484 6300 36494 6356
rect 37986 6300 37996 6356
rect 38052 6300 39676 6356
rect 39732 6300 39742 6356
rect 44268 6300 45836 6356
rect 45892 6300 45902 6356
rect 50754 6300 50764 6356
rect 50820 6300 54348 6356
rect 54404 6300 54414 6356
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 26348 6244 26404 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 242 6188 252 6244
rect 308 6188 3500 6244
rect 3556 6188 3566 6244
rect 4274 6188 4284 6244
rect 4340 6188 6860 6244
rect 6916 6188 6926 6244
rect 8092 6188 9100 6244
rect 9156 6188 9166 6244
rect 9660 6188 10780 6244
rect 10836 6188 10846 6244
rect 11106 6188 11116 6244
rect 11172 6188 12124 6244
rect 12180 6188 12190 6244
rect 13346 6188 13356 6244
rect 13412 6188 15092 6244
rect 16482 6188 16492 6244
rect 16548 6188 23716 6244
rect 24434 6188 24444 6244
rect 24500 6188 26404 6244
rect 32956 6188 36540 6244
rect 36596 6188 36606 6244
rect 44146 6188 44156 6244
rect 44212 6188 44940 6244
rect 44996 6188 45006 6244
rect 45154 6188 45164 6244
rect 45220 6188 48412 6244
rect 48468 6188 48478 6244
rect 51202 6188 51212 6244
rect 51268 6188 52108 6244
rect 52164 6188 52174 6244
rect 52770 6188 52780 6244
rect 52836 6188 55132 6244
rect 55188 6188 55198 6244
rect 0 6132 112 6160
rect 23660 6132 23716 6188
rect 32956 6132 33012 6188
rect 57344 6132 57456 6160
rect 0 6076 700 6132
rect 756 6076 766 6132
rect 1362 6076 1372 6132
rect 1428 6076 6244 6132
rect 6402 6076 6412 6132
rect 6468 6076 16716 6132
rect 16772 6076 16782 6132
rect 17714 6076 17724 6132
rect 17780 6076 17948 6132
rect 18004 6076 18014 6132
rect 18946 6076 18956 6132
rect 19012 6076 23100 6132
rect 23156 6076 23166 6132
rect 23660 6076 25228 6132
rect 25284 6076 25294 6132
rect 27234 6076 27244 6132
rect 27300 6076 28476 6132
rect 28532 6076 28542 6132
rect 32946 6076 32956 6132
rect 33012 6076 33022 6132
rect 34178 6076 34188 6132
rect 34244 6076 34524 6132
rect 34580 6076 35980 6132
rect 36036 6076 36046 6132
rect 36204 6076 47068 6132
rect 47124 6076 47134 6132
rect 51762 6076 51772 6132
rect 51828 6076 52444 6132
rect 52500 6076 52510 6132
rect 52658 6076 52668 6132
rect 52724 6076 57456 6132
rect 0 6048 112 6076
rect 6188 6020 6244 6076
rect 36204 6020 36260 6076
rect 57344 6048 57456 6076
rect 1586 5964 1596 6020
rect 1652 5964 2828 6020
rect 2884 5964 4844 6020
rect 4900 5964 4910 6020
rect 6188 5964 11564 6020
rect 11620 5964 11630 6020
rect 11778 5964 11788 6020
rect 11844 5964 11882 6020
rect 11974 5964 12012 6020
rect 12068 5964 12078 6020
rect 12226 5964 12236 6020
rect 12292 5964 12908 6020
rect 12964 5964 12974 6020
rect 14466 5964 14476 6020
rect 14532 5964 15484 6020
rect 15540 5964 15550 6020
rect 15810 5964 15820 6020
rect 15876 5964 16268 6020
rect 16324 5964 16334 6020
rect 20402 5964 20412 6020
rect 20468 5964 24668 6020
rect 24724 5964 24734 6020
rect 26338 5964 26348 6020
rect 26404 5964 26684 6020
rect 26740 5964 26750 6020
rect 27458 5964 27468 6020
rect 27524 5964 36260 6020
rect 36418 5964 36428 6020
rect 36484 5964 53564 6020
rect 53620 5964 53630 6020
rect 2370 5852 2380 5908
rect 2436 5852 3052 5908
rect 3108 5852 3388 5908
rect 4050 5852 4060 5908
rect 4116 5852 5964 5908
rect 6020 5852 6030 5908
rect 6290 5852 6300 5908
rect 6356 5852 7980 5908
rect 8036 5852 8046 5908
rect 8530 5852 8540 5908
rect 8596 5852 9324 5908
rect 9380 5852 9390 5908
rect 10098 5852 10108 5908
rect 10164 5852 10892 5908
rect 10948 5852 15596 5908
rect 15652 5852 15662 5908
rect 15810 5852 15820 5908
rect 15876 5852 18396 5908
rect 18452 5852 18462 5908
rect 21074 5852 21084 5908
rect 21140 5852 21868 5908
rect 21924 5852 21934 5908
rect 24210 5852 24220 5908
rect 24276 5852 25004 5908
rect 25060 5852 27804 5908
rect 27860 5852 27870 5908
rect 29148 5852 33180 5908
rect 33236 5852 33246 5908
rect 33394 5852 33404 5908
rect 33460 5852 34860 5908
rect 34916 5852 34926 5908
rect 35074 5852 35084 5908
rect 35140 5852 35178 5908
rect 35410 5852 35420 5908
rect 35476 5852 36540 5908
rect 36596 5852 36606 5908
rect 38098 5852 38108 5908
rect 38164 5852 48748 5908
rect 48804 5852 48814 5908
rect 3332 5796 3388 5852
rect 29148 5796 29204 5852
rect 3332 5740 5180 5796
rect 5236 5740 5246 5796
rect 5842 5740 5852 5796
rect 5908 5740 7196 5796
rect 7252 5740 7262 5796
rect 7410 5740 7420 5796
rect 7476 5740 8764 5796
rect 8820 5740 8830 5796
rect 9650 5740 9660 5796
rect 9716 5740 10332 5796
rect 10388 5740 10398 5796
rect 14578 5740 14588 5796
rect 14644 5740 15932 5796
rect 15988 5740 15998 5796
rect 19058 5740 19068 5796
rect 19124 5740 21420 5796
rect 21476 5740 21486 5796
rect 22866 5740 22876 5796
rect 22932 5740 24556 5796
rect 24612 5740 24622 5796
rect 27570 5740 27580 5796
rect 27636 5740 29204 5796
rect 29362 5740 29372 5796
rect 29428 5740 29932 5796
rect 29988 5740 29998 5796
rect 30146 5740 30156 5796
rect 30212 5740 32620 5796
rect 32676 5740 39900 5796
rect 39956 5740 39966 5796
rect 40114 5740 40124 5796
rect 40180 5740 40348 5796
rect 40404 5740 40414 5796
rect 41458 5740 41468 5796
rect 41524 5740 44156 5796
rect 44212 5740 44222 5796
rect 44930 5740 44940 5796
rect 44996 5740 48972 5796
rect 49028 5740 50876 5796
rect 50932 5740 50942 5796
rect 54898 5740 54908 5796
rect 54964 5740 56140 5796
rect 56196 5740 56206 5796
rect 0 5684 112 5712
rect 57344 5684 57456 5712
rect 0 5628 420 5684
rect 3826 5628 3836 5684
rect 3892 5628 15148 5684
rect 0 5600 112 5628
rect 364 5572 420 5628
rect 15092 5572 15148 5628
rect 18172 5628 27860 5684
rect 28018 5628 28028 5684
rect 28084 5628 28700 5684
rect 28756 5628 28766 5684
rect 29250 5628 29260 5684
rect 29316 5628 32732 5684
rect 32788 5628 33068 5684
rect 33124 5628 33134 5684
rect 34290 5628 34300 5684
rect 34356 5628 35084 5684
rect 35140 5628 35150 5684
rect 36754 5628 36764 5684
rect 36820 5628 38444 5684
rect 38500 5628 39340 5684
rect 39396 5628 39406 5684
rect 41356 5628 48636 5684
rect 48692 5628 48702 5684
rect 50372 5628 57456 5684
rect 18172 5572 18228 5628
rect 27804 5572 27860 5628
rect 41356 5572 41412 5628
rect 50372 5572 50428 5628
rect 57344 5600 57456 5628
rect 364 5516 3164 5572
rect 3220 5516 3230 5572
rect 5170 5516 5180 5572
rect 5236 5516 6748 5572
rect 6804 5516 6814 5572
rect 7634 5516 7644 5572
rect 7700 5516 11340 5572
rect 11396 5516 11406 5572
rect 14578 5516 14588 5572
rect 14644 5516 14700 5572
rect 14756 5516 14766 5572
rect 14914 5516 14924 5572
rect 14980 5516 15018 5572
rect 15092 5516 18228 5572
rect 18386 5516 18396 5572
rect 18452 5516 19628 5572
rect 19684 5516 19694 5572
rect 19954 5516 19964 5572
rect 20020 5516 20030 5572
rect 20962 5516 20972 5572
rect 21028 5516 21756 5572
rect 21812 5516 21822 5572
rect 25218 5516 25228 5572
rect 25284 5516 25564 5572
rect 25620 5516 27580 5572
rect 27636 5516 27646 5572
rect 27804 5516 41412 5572
rect 43586 5516 43596 5572
rect 43652 5516 44268 5572
rect 44324 5516 44334 5572
rect 47058 5516 47068 5572
rect 47124 5516 50428 5572
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 19964 5460 20020 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 690 5404 700 5460
rect 756 5404 3388 5460
rect 3490 5404 3500 5460
rect 3556 5404 4284 5460
rect 4340 5404 4350 5460
rect 6626 5404 6636 5460
rect 6692 5404 6860 5460
rect 6916 5404 8092 5460
rect 8148 5404 8158 5460
rect 9202 5404 9212 5460
rect 9268 5404 19460 5460
rect 19964 5404 20860 5460
rect 20916 5404 21644 5460
rect 21700 5404 21710 5460
rect 23650 5404 23660 5460
rect 23716 5404 23726 5460
rect 24892 5404 25900 5460
rect 25956 5404 27692 5460
rect 27748 5404 27758 5460
rect 33058 5404 33068 5460
rect 33124 5404 33292 5460
rect 33348 5404 33358 5460
rect 33964 5404 43540 5460
rect 44818 5404 44828 5460
rect 44884 5404 44922 5460
rect 3332 5348 3388 5404
rect 19404 5348 19460 5404
rect 23660 5348 23716 5404
rect 2482 5292 2492 5348
rect 2548 5292 2558 5348
rect 3332 5292 7812 5348
rect 7970 5292 7980 5348
rect 8036 5292 9436 5348
rect 9492 5292 9502 5348
rect 9884 5292 10892 5348
rect 10948 5292 10958 5348
rect 12450 5292 12460 5348
rect 12516 5292 19068 5348
rect 19124 5292 19134 5348
rect 19404 5292 23716 5348
rect 0 5236 112 5264
rect 0 5180 1708 5236
rect 1764 5180 1774 5236
rect 0 5152 112 5180
rect 2492 5012 2548 5292
rect 7756 5236 7812 5292
rect 9884 5236 9940 5292
rect 3490 5180 3500 5236
rect 3556 5180 7084 5236
rect 7140 5180 7150 5236
rect 7756 5180 9940 5236
rect 10098 5180 10108 5236
rect 10164 5180 12236 5236
rect 12292 5180 12302 5236
rect 12898 5180 12908 5236
rect 12964 5180 14140 5236
rect 14196 5180 14476 5236
rect 14532 5180 14542 5236
rect 15250 5180 15260 5236
rect 15316 5180 18620 5236
rect 18676 5180 18686 5236
rect 19180 5180 20972 5236
rect 21028 5180 21038 5236
rect 19180 5124 19236 5180
rect 24892 5124 24948 5404
rect 26002 5292 26012 5348
rect 26068 5292 26796 5348
rect 26852 5292 26862 5348
rect 27234 5292 27244 5348
rect 27300 5292 28588 5348
rect 28644 5292 28654 5348
rect 32834 5292 32844 5348
rect 32900 5292 33740 5348
rect 33796 5292 33806 5348
rect 33964 5236 34020 5404
rect 43484 5348 43540 5404
rect 34626 5292 34636 5348
rect 34692 5292 34748 5348
rect 34804 5292 34814 5348
rect 35298 5292 35308 5348
rect 35364 5292 43428 5348
rect 43484 5292 55468 5348
rect 55524 5292 55534 5348
rect 43372 5236 43428 5292
rect 57344 5236 57456 5264
rect 25106 5180 25116 5236
rect 25172 5180 28028 5236
rect 28084 5180 28094 5236
rect 28242 5180 28252 5236
rect 28308 5180 34020 5236
rect 40338 5180 40348 5236
rect 40404 5180 41020 5236
rect 41076 5180 41356 5236
rect 41412 5180 41422 5236
rect 42578 5180 42588 5236
rect 42644 5180 43204 5236
rect 43372 5180 49420 5236
rect 49476 5180 52556 5236
rect 52612 5180 52622 5236
rect 56130 5180 56140 5236
rect 56196 5180 57456 5236
rect 43148 5124 43204 5180
rect 57344 5152 57456 5180
rect 2678 5068 2716 5124
rect 2772 5068 2782 5124
rect 3602 5068 3612 5124
rect 3668 5068 5516 5124
rect 5572 5068 5582 5124
rect 5730 5068 5740 5124
rect 5796 5068 7308 5124
rect 7364 5068 7980 5124
rect 8036 5068 8046 5124
rect 8530 5068 8540 5124
rect 8596 5068 9772 5124
rect 9828 5068 9838 5124
rect 10770 5068 10780 5124
rect 10836 5068 11116 5124
rect 11172 5068 11900 5124
rect 11956 5068 11966 5124
rect 12338 5068 12348 5124
rect 12404 5068 12414 5124
rect 12646 5068 12684 5124
rect 12740 5068 12750 5124
rect 13122 5068 13132 5124
rect 13188 5068 13198 5124
rect 13906 5068 13916 5124
rect 13972 5068 15820 5124
rect 15876 5068 15886 5124
rect 16146 5068 16156 5124
rect 16212 5068 16996 5124
rect 12348 5012 12404 5068
rect 13132 5012 13188 5068
rect 16940 5012 16996 5068
rect 18396 5068 18956 5124
rect 19012 5068 19022 5124
rect 19170 5068 19180 5124
rect 19236 5068 19246 5124
rect 19730 5068 19740 5124
rect 19796 5068 20300 5124
rect 20356 5068 20366 5124
rect 20514 5068 20524 5124
rect 20580 5068 20618 5124
rect 21410 5068 21420 5124
rect 21476 5068 22316 5124
rect 22372 5068 22382 5124
rect 22754 5068 22764 5124
rect 22820 5068 24948 5124
rect 25890 5068 25900 5124
rect 25956 5068 27020 5124
rect 27076 5068 27916 5124
rect 27972 5068 27982 5124
rect 32274 5068 32284 5124
rect 32340 5068 37548 5124
rect 37604 5068 37614 5124
rect 37874 5068 37884 5124
rect 37940 5068 40460 5124
rect 40516 5068 41244 5124
rect 41300 5068 42140 5124
rect 42196 5068 42206 5124
rect 42588 5068 43092 5124
rect 43148 5068 43484 5124
rect 43540 5068 43596 5124
rect 43652 5068 43662 5124
rect 44258 5068 44268 5124
rect 44324 5068 44380 5124
rect 44436 5068 44446 5124
rect 44594 5068 44604 5124
rect 44660 5068 44940 5124
rect 44996 5068 45006 5124
rect 46610 5068 46620 5124
rect 46676 5068 49756 5124
rect 49812 5068 49822 5124
rect 53106 5068 53116 5124
rect 53172 5068 54908 5124
rect 54964 5068 54974 5124
rect 56242 5068 56252 5124
rect 56308 5068 57036 5124
rect 57092 5068 57102 5124
rect 18396 5012 18452 5068
rect 42588 5012 42644 5068
rect 43036 5012 43092 5068
rect 2380 4956 2548 5012
rect 2930 4956 2940 5012
rect 2996 4956 8988 5012
rect 9044 4956 9054 5012
rect 10546 4956 10556 5012
rect 10612 4956 13188 5012
rect 13570 4956 13580 5012
rect 13636 4956 15148 5012
rect 15204 4956 15214 5012
rect 16930 4956 16940 5012
rect 16996 4956 17006 5012
rect 18386 4956 18396 5012
rect 18452 4956 18462 5012
rect 18722 4956 18732 5012
rect 18788 4956 35532 5012
rect 35588 4956 35598 5012
rect 36978 4956 36988 5012
rect 37044 4956 37996 5012
rect 38052 4956 38062 5012
rect 38546 4956 38556 5012
rect 38612 4956 42644 5012
rect 42774 4956 42812 5012
rect 42868 4956 42878 5012
rect 43036 4956 46676 5012
rect 46806 4956 46844 5012
rect 46900 4956 46910 5012
rect 49298 4956 49308 5012
rect 49364 4956 55916 5012
rect 55972 4956 55982 5012
rect 2380 4900 2436 4956
rect 46620 4900 46676 4956
rect 2370 4844 2380 4900
rect 2436 4844 2446 4900
rect 4172 4844 5628 4900
rect 5684 4844 5694 4900
rect 6290 4844 6300 4900
rect 6356 4844 8876 4900
rect 8932 4844 8942 4900
rect 9090 4844 9100 4900
rect 9156 4844 12124 4900
rect 12180 4844 12190 4900
rect 12338 4844 12348 4900
rect 12404 4844 13468 4900
rect 13524 4844 13534 4900
rect 14578 4844 14588 4900
rect 14644 4844 14700 4900
rect 14756 4844 14766 4900
rect 15092 4844 31724 4900
rect 31780 4844 31790 4900
rect 31938 4844 31948 4900
rect 32004 4844 35308 4900
rect 35364 4844 35374 4900
rect 38658 4844 38668 4900
rect 38724 4844 39116 4900
rect 39172 4844 39182 4900
rect 41122 4844 41132 4900
rect 41188 4844 44156 4900
rect 44212 4844 44222 4900
rect 44818 4844 44828 4900
rect 44884 4844 44940 4900
rect 44996 4844 45006 4900
rect 46620 4844 47964 4900
rect 48020 4844 48030 4900
rect 50306 4844 50316 4900
rect 50372 4844 53956 4900
rect 0 4788 112 4816
rect 0 4732 3612 4788
rect 3668 4732 3678 4788
rect 0 4704 112 4732
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 4172 4618 4228 4844
rect 15092 4788 15148 4844
rect 53900 4788 53956 4844
rect 57344 4788 57456 4816
rect 5282 4732 5292 4788
rect 5348 4732 5628 4788
rect 5684 4732 5694 4788
rect 7298 4732 7308 4788
rect 7364 4732 15148 4788
rect 15250 4732 15260 4788
rect 15316 4732 16604 4788
rect 16660 4732 16670 4788
rect 17490 4732 17500 4788
rect 17556 4732 18956 4788
rect 19012 4732 19022 4788
rect 21074 4732 21084 4788
rect 21140 4732 21756 4788
rect 21812 4732 21822 4788
rect 26982 4732 27020 4788
rect 27076 4732 27086 4788
rect 29026 4732 29036 4788
rect 29092 4732 29372 4788
rect 29428 4732 29438 4788
rect 30370 4732 30380 4788
rect 30436 4732 31948 4788
rect 32004 4732 32014 4788
rect 32162 4732 32172 4788
rect 32228 4732 35756 4788
rect 35812 4732 35822 4788
rect 35970 4732 35980 4788
rect 36036 4732 43596 4788
rect 43652 4732 43662 4788
rect 44156 4732 50428 4788
rect 51538 4732 51548 4788
rect 51604 4732 52556 4788
rect 52612 4732 52622 4788
rect 53900 4732 57456 4788
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 4386 4620 4396 4676
rect 4452 4620 7756 4676
rect 7812 4620 17892 4676
rect 18050 4620 18060 4676
rect 18116 4620 20300 4676
rect 20356 4620 20366 4676
rect 20738 4620 20748 4676
rect 20804 4620 21532 4676
rect 21588 4620 21598 4676
rect 24210 4620 24220 4676
rect 24276 4620 29148 4676
rect 29204 4620 29214 4676
rect 31826 4620 31836 4676
rect 31892 4620 43652 4676
rect 4060 4564 4228 4618
rect 17836 4564 17892 4620
rect 43596 4564 43652 4620
rect 44156 4564 44212 4732
rect 50372 4676 50428 4732
rect 57344 4704 57456 4732
rect 50372 4620 55020 4676
rect 55076 4620 55086 4676
rect 2594 4508 2604 4564
rect 2660 4508 2940 4564
rect 2996 4508 3006 4564
rect 3938 4508 3948 4564
rect 4004 4562 4228 4564
rect 4004 4508 4116 4562
rect 4284 4508 7420 4564
rect 7476 4508 7486 4564
rect 7970 4508 7980 4564
rect 8036 4508 8652 4564
rect 8708 4508 8718 4564
rect 8866 4508 8876 4564
rect 8932 4508 9436 4564
rect 9492 4508 9502 4564
rect 10434 4508 10444 4564
rect 10500 4508 13020 4564
rect 13076 4508 13086 4564
rect 14578 4508 14588 4564
rect 14644 4508 16268 4564
rect 16324 4508 16828 4564
rect 16884 4508 16894 4564
rect 17836 4508 20972 4564
rect 21028 4508 21038 4564
rect 43596 4508 44212 4564
rect 44818 4508 44828 4564
rect 44884 4508 45500 4564
rect 45556 4508 45566 4564
rect 48738 4508 48748 4564
rect 48804 4508 52668 4564
rect 52724 4508 52734 4564
rect 0 4340 112 4368
rect 4284 4340 4340 4508
rect 4610 4396 4620 4452
rect 4676 4396 11564 4452
rect 11620 4396 11630 4452
rect 12114 4396 12124 4452
rect 12180 4396 12908 4452
rect 12964 4396 12974 4452
rect 14018 4396 14028 4452
rect 14084 4396 18284 4452
rect 18340 4396 18350 4452
rect 18498 4396 18508 4452
rect 18564 4396 21084 4452
rect 21140 4396 21150 4452
rect 21522 4396 21532 4452
rect 21588 4396 28252 4452
rect 28308 4396 28318 4452
rect 28578 4396 28588 4452
rect 28644 4396 30604 4452
rect 30660 4396 31276 4452
rect 31332 4396 31342 4452
rect 31948 4396 38108 4452
rect 38164 4396 38174 4452
rect 38322 4396 38332 4452
rect 38388 4396 38780 4452
rect 38836 4396 38846 4452
rect 39890 4396 39900 4452
rect 39956 4396 44604 4452
rect 44660 4396 44670 4452
rect 31948 4340 32004 4396
rect 57344 4340 57456 4368
rect 0 4284 3276 4340
rect 3332 4284 3342 4340
rect 3714 4284 3724 4340
rect 3780 4284 4340 4340
rect 4498 4284 4508 4340
rect 4564 4284 9548 4340
rect 9604 4284 9614 4340
rect 10098 4284 10108 4340
rect 10164 4284 13468 4340
rect 13524 4284 15148 4340
rect 15922 4284 15932 4340
rect 15988 4284 18396 4340
rect 18452 4284 18462 4340
rect 19954 4284 19964 4340
rect 20020 4284 20636 4340
rect 20692 4284 20702 4340
rect 22082 4284 22092 4340
rect 22148 4284 23660 4340
rect 23716 4284 23726 4340
rect 23874 4284 23884 4340
rect 23940 4284 27916 4340
rect 27972 4284 27982 4340
rect 30818 4284 30828 4340
rect 30884 4284 32004 4340
rect 32582 4284 32620 4340
rect 32676 4284 32686 4340
rect 33730 4284 33740 4340
rect 33796 4284 34076 4340
rect 34132 4284 34142 4340
rect 35718 4284 35756 4340
rect 35812 4284 35822 4340
rect 36418 4284 36428 4340
rect 36484 4284 36876 4340
rect 36932 4284 36942 4340
rect 37538 4284 37548 4340
rect 37604 4284 38556 4340
rect 38612 4284 38622 4340
rect 44482 4284 44492 4340
rect 44548 4284 46508 4340
rect 46564 4284 46574 4340
rect 53554 4284 53564 4340
rect 53620 4284 57456 4340
rect 0 4256 112 4284
rect 15092 4228 15148 4284
rect 57344 4256 57456 4284
rect 1782 4172 1820 4228
rect 1876 4172 1886 4228
rect 2258 4172 2268 4228
rect 2324 4172 6300 4228
rect 6356 4172 6366 4228
rect 6962 4172 6972 4228
rect 7028 4172 7308 4228
rect 7364 4172 7374 4228
rect 7522 4172 7532 4228
rect 7588 4172 8092 4228
rect 8148 4172 8158 4228
rect 9426 4172 9436 4228
rect 9492 4172 10668 4228
rect 10724 4172 10734 4228
rect 13346 4172 13356 4228
rect 13412 4172 13580 4228
rect 13636 4172 13916 4228
rect 13972 4172 13982 4228
rect 15092 4172 18956 4228
rect 19012 4172 19022 4228
rect 19964 4172 32284 4228
rect 32340 4172 32350 4228
rect 32722 4172 32732 4228
rect 32788 4172 37212 4228
rect 37268 4172 37278 4228
rect 44034 4172 44044 4228
rect 44100 4172 55916 4228
rect 55972 4172 55982 4228
rect 1362 4060 1372 4116
rect 1428 4060 2380 4116
rect 2436 4060 2716 4116
rect 2772 4060 2782 4116
rect 3602 4060 3612 4116
rect 3668 4060 7588 4116
rect 8306 4060 8316 4116
rect 8372 4060 11900 4116
rect 11956 4060 11966 4116
rect 13804 4060 14924 4116
rect 14980 4060 14990 4116
rect 16258 4060 16268 4116
rect 16324 4060 17052 4116
rect 17108 4060 17118 4116
rect 7532 4004 7588 4060
rect 13804 4004 13860 4060
rect 466 3948 476 4004
rect 532 3948 3500 4004
rect 3556 3948 3566 4004
rect 4134 3948 4172 4004
rect 4228 3948 4238 4004
rect 5954 3948 5964 4004
rect 6020 3948 6524 4004
rect 6580 3948 6590 4004
rect 7522 3948 7532 4004
rect 7588 3948 7598 4004
rect 8082 3948 8092 4004
rect 8148 3948 13860 4004
rect 14018 3948 14028 4004
rect 14084 3948 16828 4004
rect 16884 3948 16894 4004
rect 0 3892 112 3920
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 19964 3892 20020 4172
rect 20178 4060 20188 4116
rect 20244 4060 22652 4116
rect 22708 4060 22718 4116
rect 23986 4060 23996 4116
rect 24052 4060 24220 4116
rect 24276 4060 24286 4116
rect 31602 4060 31612 4116
rect 31668 4060 32508 4116
rect 32564 4060 32574 4116
rect 32732 4060 35980 4116
rect 36036 4060 36046 4116
rect 43586 4060 43596 4116
rect 43652 4060 52332 4116
rect 52388 4060 52398 4116
rect 52882 4060 52892 4116
rect 52948 4060 53564 4116
rect 53620 4060 53630 4116
rect 32732 4004 32788 4060
rect 22754 3948 22764 4004
rect 22820 3948 23884 4004
rect 23940 3948 23950 4004
rect 31490 3948 31500 4004
rect 31556 3948 32788 4004
rect 33618 3948 33628 4004
rect 33684 3948 44268 4004
rect 44324 3948 44334 4004
rect 45378 3948 45388 4004
rect 45444 3948 50204 4004
rect 50260 3948 50270 4004
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 57344 3892 57456 3920
rect 0 3836 3500 3892
rect 3556 3836 3566 3892
rect 5618 3836 5628 3892
rect 5684 3836 9660 3892
rect 9716 3836 9726 3892
rect 11218 3836 11228 3892
rect 11284 3836 20020 3892
rect 20178 3836 20188 3892
rect 20244 3836 22652 3892
rect 22708 3836 22718 3892
rect 29148 3836 44156 3892
rect 44212 3836 44222 3892
rect 46050 3836 46060 3892
rect 46116 3836 46172 3892
rect 46228 3836 46508 3892
rect 46564 3836 46574 3892
rect 47058 3836 47068 3892
rect 47124 3836 57456 3892
rect 0 3808 112 3836
rect 29148 3780 29204 3836
rect 57344 3808 57456 3836
rect 802 3724 812 3780
rect 868 3724 1372 3780
rect 1428 3724 1438 3780
rect 3332 3724 7868 3780
rect 7924 3724 7934 3780
rect 9734 3724 9772 3780
rect 9828 3724 9838 3780
rect 11078 3724 11116 3780
rect 11172 3724 11182 3780
rect 12982 3724 13020 3780
rect 13076 3724 13086 3780
rect 14242 3724 14252 3780
rect 14308 3724 15932 3780
rect 15988 3724 16716 3780
rect 16772 3724 16782 3780
rect 19618 3724 19628 3780
rect 19684 3724 21644 3780
rect 21700 3724 21710 3780
rect 23538 3724 23548 3780
rect 23604 3724 26012 3780
rect 26068 3724 26078 3780
rect 26562 3724 26572 3780
rect 26628 3724 26796 3780
rect 26852 3724 26862 3780
rect 27682 3724 27692 3780
rect 27748 3724 28476 3780
rect 28532 3724 28542 3780
rect 29138 3724 29148 3780
rect 29204 3724 29214 3780
rect 32050 3724 32060 3780
rect 32116 3724 32172 3780
rect 32228 3724 32238 3780
rect 33842 3724 33852 3780
rect 33908 3724 36652 3780
rect 36708 3724 36718 3780
rect 37986 3724 37996 3780
rect 38052 3724 38668 3780
rect 38724 3724 38734 3780
rect 40002 3724 40012 3780
rect 40068 3724 50764 3780
rect 50820 3724 50830 3780
rect 53778 3724 53788 3780
rect 53844 3724 54012 3780
rect 54068 3724 54078 3780
rect 55318 3724 55356 3780
rect 55412 3724 55422 3780
rect 3332 3668 3388 3724
rect 802 3612 812 3668
rect 868 3612 3388 3668
rect 3490 3612 3500 3668
rect 3556 3612 7476 3668
rect 7634 3612 7644 3668
rect 7700 3612 12684 3668
rect 12740 3612 12750 3668
rect 14130 3612 14140 3668
rect 14196 3612 14924 3668
rect 14980 3612 18732 3668
rect 18788 3612 19628 3668
rect 19684 3612 19694 3668
rect 19842 3612 19852 3668
rect 19908 3612 21756 3668
rect 21812 3612 21822 3668
rect 28102 3612 28140 3668
rect 28196 3612 32284 3668
rect 32340 3612 32350 3668
rect 32722 3612 32732 3668
rect 32788 3612 34412 3668
rect 34468 3612 34478 3668
rect 35634 3612 35644 3668
rect 35700 3612 35868 3668
rect 35924 3612 35934 3668
rect 36306 3612 36316 3668
rect 36372 3612 36764 3668
rect 36820 3612 36830 3668
rect 40870 3612 40908 3668
rect 40964 3612 40974 3668
rect 44146 3612 44156 3668
rect 44212 3612 44492 3668
rect 44548 3612 45052 3668
rect 45108 3612 45118 3668
rect 46386 3612 46396 3668
rect 46452 3612 47068 3668
rect 47124 3612 47134 3668
rect 47842 3612 47852 3668
rect 47908 3612 54908 3668
rect 54964 3612 54974 3668
rect 7420 3556 7476 3612
rect 1474 3500 1484 3556
rect 1540 3500 1596 3556
rect 1652 3500 1662 3556
rect 2370 3500 2380 3556
rect 2436 3500 7196 3556
rect 7252 3500 7262 3556
rect 7420 3500 9492 3556
rect 10098 3500 10108 3556
rect 10164 3500 15148 3556
rect 16146 3500 16156 3556
rect 16212 3500 16604 3556
rect 16660 3500 16670 3556
rect 17602 3500 17612 3556
rect 17668 3500 18172 3556
rect 18228 3500 18238 3556
rect 18498 3500 18508 3556
rect 18564 3500 24220 3556
rect 24276 3500 24286 3556
rect 26086 3500 26124 3556
rect 26180 3500 28700 3556
rect 28756 3500 28766 3556
rect 29362 3500 29372 3556
rect 29428 3500 30156 3556
rect 30212 3500 30222 3556
rect 31126 3500 31164 3556
rect 31220 3500 31230 3556
rect 35522 3500 35532 3556
rect 35588 3500 40404 3556
rect 45154 3500 45164 3556
rect 45220 3500 46732 3556
rect 46788 3500 46798 3556
rect 47394 3500 47404 3556
rect 47460 3500 48748 3556
rect 48804 3500 48814 3556
rect 0 3444 112 3472
rect 9436 3444 9492 3500
rect 15092 3444 15148 3500
rect 0 3388 476 3444
rect 532 3388 542 3444
rect 2940 3388 3332 3444
rect 3388 3388 3398 3444
rect 3490 3388 3500 3444
rect 3556 3388 5068 3444
rect 5124 3388 5134 3444
rect 8372 3388 9212 3444
rect 9268 3388 9278 3444
rect 9436 3388 14028 3444
rect 14084 3388 14094 3444
rect 15092 3388 16492 3444
rect 16548 3388 16558 3444
rect 18834 3388 18844 3444
rect 18900 3388 20860 3444
rect 20916 3388 20926 3444
rect 21074 3388 21084 3444
rect 21140 3388 26460 3444
rect 26516 3388 26526 3444
rect 31892 3388 35420 3444
rect 35476 3388 36092 3444
rect 36148 3388 36158 3444
rect 36866 3388 36876 3444
rect 36932 3388 37884 3444
rect 37940 3388 37950 3444
rect 0 3360 112 3388
rect 2940 3332 2996 3388
rect 8372 3332 8428 3388
rect 31892 3332 31948 3388
rect 40348 3332 40404 3500
rect 57344 3444 57456 3472
rect 40562 3388 40572 3444
rect 40628 3388 41692 3444
rect 41748 3388 41758 3444
rect 43260 3388 44044 3444
rect 44100 3388 44110 3444
rect 44258 3388 44268 3444
rect 44324 3388 49084 3444
rect 49140 3388 49150 3444
rect 49308 3388 51100 3444
rect 51156 3388 51166 3444
rect 53788 3388 57456 3444
rect 43260 3332 43316 3388
rect 49308 3332 49364 3388
rect 53788 3332 53844 3388
rect 57344 3360 57456 3388
rect 2930 3276 2940 3332
rect 2996 3276 3006 3332
rect 3266 3276 3276 3332
rect 3332 3276 6692 3332
rect 6850 3276 6860 3332
rect 6916 3276 8428 3332
rect 14130 3276 14140 3332
rect 14196 3276 14252 3332
rect 14308 3276 14318 3332
rect 14924 3276 15820 3332
rect 15876 3276 15886 3332
rect 18498 3276 18508 3332
rect 18564 3276 21532 3332
rect 21588 3276 21598 3332
rect 22194 3276 22204 3332
rect 22260 3276 31948 3332
rect 33954 3276 33964 3332
rect 34020 3276 35308 3332
rect 37426 3276 37436 3332
rect 37492 3276 39228 3332
rect 39284 3276 39294 3332
rect 40348 3276 43316 3332
rect 43474 3276 43484 3332
rect 43540 3276 44828 3332
rect 44884 3276 44894 3332
rect 45500 3276 49364 3332
rect 49522 3276 49532 3332
rect 49588 3276 53844 3332
rect 6636 3220 6692 3276
rect 6636 3164 7980 3220
rect 8036 3164 8046 3220
rect 9314 3164 9324 3220
rect 9380 3164 14700 3220
rect 14756 3164 14766 3220
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 14924 3108 14980 3276
rect 35252 3220 35308 3276
rect 5954 3052 5964 3108
rect 6020 3052 13020 3108
rect 13076 3052 13086 3108
rect 13794 3052 13804 3108
rect 13860 3052 14980 3108
rect 15092 3164 22876 3220
rect 22932 3164 22942 3220
rect 23314 3164 23324 3220
rect 23380 3164 23436 3220
rect 23492 3164 23502 3220
rect 24322 3164 24332 3220
rect 24388 3164 25452 3220
rect 25508 3164 25518 3220
rect 25666 3164 25676 3220
rect 25732 3164 28028 3220
rect 28084 3164 28094 3220
rect 28354 3164 28364 3220
rect 28420 3164 29260 3220
rect 29316 3164 29326 3220
rect 30482 3164 30492 3220
rect 30548 3164 34412 3220
rect 34468 3164 34478 3220
rect 35252 3164 36204 3220
rect 36260 3164 42364 3220
rect 42420 3164 42430 3220
rect 0 2996 112 3024
rect 15092 2996 15148 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 18946 3052 18956 3108
rect 19012 3052 23548 3108
rect 23604 3052 23614 3108
rect 24210 3052 24220 3108
rect 24276 3052 26460 3108
rect 26516 3052 26526 3108
rect 27122 3052 27132 3108
rect 27188 3052 28588 3108
rect 28644 3052 28654 3108
rect 29922 3052 29932 3108
rect 29988 3052 35980 3108
rect 36036 3052 36046 3108
rect 36194 3052 36204 3108
rect 36260 3052 43484 3108
rect 43540 3052 43550 3108
rect 45500 2996 45556 3276
rect 47506 3164 47516 3220
rect 47572 3164 55804 3220
rect 55860 3164 55870 3220
rect 46946 3052 46956 3108
rect 47012 3052 52220 3108
rect 52276 3052 53116 3108
rect 53172 3052 53182 3108
rect 56242 3052 56252 3108
rect 56308 3052 56924 3108
rect 56980 3052 56990 3108
rect 57344 2996 57456 3024
rect 0 2940 4340 2996
rect 4498 2940 4508 2996
rect 4564 2940 15148 2996
rect 16146 2940 16156 2996
rect 16212 2940 32956 2996
rect 33012 2940 33022 2996
rect 35074 2940 35084 2996
rect 35140 2940 37660 2996
rect 37716 2940 37726 2996
rect 40002 2940 40012 2996
rect 40068 2940 40684 2996
rect 40740 2940 40750 2996
rect 40898 2940 40908 2996
rect 40964 2940 45556 2996
rect 45714 2940 45724 2996
rect 45780 2940 46564 2996
rect 48402 2940 48412 2996
rect 48468 2940 52108 2996
rect 52164 2940 52174 2996
rect 56364 2940 57456 2996
rect 0 2912 112 2940
rect 4284 2884 4340 2940
rect 46508 2884 46564 2940
rect 690 2828 700 2884
rect 756 2828 3388 2884
rect 3444 2828 3454 2884
rect 4284 2828 7756 2884
rect 7812 2828 7822 2884
rect 8316 2828 13020 2884
rect 13076 2828 13086 2884
rect 13794 2828 13804 2884
rect 13860 2828 14476 2884
rect 14532 2828 14542 2884
rect 17266 2828 17276 2884
rect 17332 2828 17500 2884
rect 17556 2828 17948 2884
rect 18004 2828 18014 2884
rect 18610 2828 18620 2884
rect 18676 2828 20300 2884
rect 20356 2828 25676 2884
rect 25732 2828 25742 2884
rect 26422 2828 26460 2884
rect 26516 2828 26526 2884
rect 31714 2828 31724 2884
rect 31780 2828 46284 2884
rect 46340 2828 46350 2884
rect 46508 2828 48412 2884
rect 48468 2828 48478 2884
rect 48626 2828 48636 2884
rect 48692 2828 55916 2884
rect 55972 2828 55982 2884
rect 914 2716 924 2772
rect 980 2716 2268 2772
rect 2324 2716 2334 2772
rect 3714 2716 3724 2772
rect 3780 2716 4508 2772
rect 4564 2716 4574 2772
rect 5058 2716 5068 2772
rect 5124 2716 6636 2772
rect 6692 2716 6702 2772
rect 8054 2716 8092 2772
rect 8148 2716 8158 2772
rect 8316 2660 8372 2828
rect 56364 2772 56420 2940
rect 57344 2912 57456 2940
rect 8642 2716 8652 2772
rect 8708 2716 8876 2772
rect 8932 2716 8942 2772
rect 9212 2716 11228 2772
rect 11284 2716 11294 2772
rect 12226 2716 12236 2772
rect 12292 2716 13580 2772
rect 13636 2716 13646 2772
rect 13804 2716 15596 2772
rect 15652 2716 15662 2772
rect 18498 2716 18508 2772
rect 18564 2716 19068 2772
rect 19124 2716 19134 2772
rect 19506 2716 19516 2772
rect 19572 2716 21196 2772
rect 21252 2716 21262 2772
rect 21410 2716 21420 2772
rect 21476 2716 22428 2772
rect 22484 2716 22494 2772
rect 23874 2716 23884 2772
rect 23940 2716 24220 2772
rect 24276 2716 24286 2772
rect 25330 2716 25340 2772
rect 25396 2716 27804 2772
rect 27860 2716 27870 2772
rect 31938 2716 31948 2772
rect 32004 2716 32172 2772
rect 32228 2716 32238 2772
rect 32946 2716 32956 2772
rect 33012 2716 33292 2772
rect 33348 2716 33358 2772
rect 33702 2716 33740 2772
rect 33796 2716 33806 2772
rect 34178 2716 34188 2772
rect 34244 2716 34300 2772
rect 34356 2716 34366 2772
rect 35158 2716 35196 2772
rect 35252 2716 35262 2772
rect 35746 2716 35756 2772
rect 35812 2716 36316 2772
rect 36372 2716 36382 2772
rect 36614 2716 36652 2772
rect 36708 2716 36718 2772
rect 37286 2716 37324 2772
rect 37380 2716 37390 2772
rect 38546 2716 38556 2772
rect 38612 2716 39116 2772
rect 39172 2716 39182 2772
rect 39330 2716 39340 2772
rect 39396 2716 39564 2772
rect 39620 2716 39630 2772
rect 42102 2716 42140 2772
rect 42196 2716 42206 2772
rect 43586 2716 43596 2772
rect 43652 2716 45500 2772
rect 45556 2716 45566 2772
rect 45714 2716 45724 2772
rect 45780 2716 48860 2772
rect 48916 2716 48926 2772
rect 49084 2716 56420 2772
rect 9212 2660 9268 2716
rect 13804 2660 13860 2716
rect 49084 2660 49140 2716
rect 466 2604 476 2660
rect 532 2604 6692 2660
rect 6822 2604 6860 2660
rect 6916 2604 6926 2660
rect 7298 2604 7308 2660
rect 7364 2604 8372 2660
rect 8642 2604 8652 2660
rect 8708 2604 9268 2660
rect 9650 2604 9660 2660
rect 9716 2604 13860 2660
rect 14690 2604 14700 2660
rect 14756 2604 16548 2660
rect 16706 2604 16716 2660
rect 16772 2604 17164 2660
rect 17220 2604 17230 2660
rect 18050 2604 18060 2660
rect 18116 2604 19180 2660
rect 19236 2604 19246 2660
rect 19954 2604 19964 2660
rect 20020 2604 23100 2660
rect 23156 2604 23166 2660
rect 23398 2604 23436 2660
rect 23492 2604 23502 2660
rect 28998 2604 29036 2660
rect 29092 2604 29102 2660
rect 32050 2604 32060 2660
rect 32116 2604 38892 2660
rect 38948 2604 38958 2660
rect 40338 2604 40348 2660
rect 40404 2604 41132 2660
rect 41188 2604 41198 2660
rect 43362 2604 43372 2660
rect 43428 2604 44156 2660
rect 44212 2604 44222 2660
rect 45378 2604 45388 2660
rect 45444 2604 48244 2660
rect 48738 2604 48748 2660
rect 48804 2604 49140 2660
rect 49298 2604 49308 2660
rect 49364 2604 55244 2660
rect 55300 2604 55310 2660
rect 0 2548 112 2576
rect 6636 2548 6692 2604
rect 16492 2548 16548 2604
rect 48188 2548 48244 2604
rect 57344 2548 57456 2576
rect 0 2492 6580 2548
rect 6636 2492 12796 2548
rect 12852 2492 12862 2548
rect 13010 2492 13020 2548
rect 13076 2492 16436 2548
rect 16492 2492 17724 2548
rect 17780 2492 17790 2548
rect 18274 2492 18284 2548
rect 18340 2492 20076 2548
rect 20132 2492 20142 2548
rect 21186 2492 21196 2548
rect 21252 2492 24108 2548
rect 24164 2492 24174 2548
rect 24434 2492 24444 2548
rect 24500 2492 27916 2548
rect 27972 2492 30716 2548
rect 30772 2492 30782 2548
rect 31714 2492 31724 2548
rect 31780 2492 33292 2548
rect 33348 2492 33358 2548
rect 35746 2492 35756 2548
rect 35812 2492 36988 2548
rect 37044 2492 37054 2548
rect 37986 2492 37996 2548
rect 38052 2492 41468 2548
rect 41524 2492 41534 2548
rect 43138 2492 43148 2548
rect 43204 2492 43932 2548
rect 43988 2492 43998 2548
rect 44258 2492 44268 2548
rect 44324 2492 45276 2548
rect 45332 2492 45342 2548
rect 45826 2492 45836 2548
rect 45892 2492 47852 2548
rect 47908 2492 47918 2548
rect 48178 2492 48188 2548
rect 48244 2492 48254 2548
rect 48402 2492 48412 2548
rect 48468 2492 57456 2548
rect 0 2464 112 2492
rect 6524 2436 6580 2492
rect 16380 2436 16436 2492
rect 57344 2464 57456 2492
rect 2706 2380 2716 2436
rect 2772 2380 4284 2436
rect 4340 2380 4350 2436
rect 6524 2380 13916 2436
rect 13972 2380 13982 2436
rect 14242 2380 14252 2436
rect 14308 2380 15540 2436
rect 16380 2380 18620 2436
rect 18676 2380 18686 2436
rect 18834 2380 18844 2436
rect 18900 2380 19852 2436
rect 19908 2380 20748 2436
rect 20804 2380 20814 2436
rect 21410 2380 21420 2436
rect 21476 2380 23772 2436
rect 23828 2380 23838 2436
rect 30258 2380 30268 2436
rect 30324 2380 32060 2436
rect 32116 2380 32126 2436
rect 32274 2380 32284 2436
rect 32340 2380 38164 2436
rect 40562 2380 40572 2436
rect 40628 2380 44324 2436
rect 45938 2380 45948 2436
rect 46004 2380 47516 2436
rect 47572 2380 47582 2436
rect 48402 2380 48412 2436
rect 48468 2380 48478 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 2818 2268 2828 2324
rect 2884 2268 4060 2324
rect 4116 2268 4126 2324
rect 5058 2268 5068 2324
rect 5124 2268 8540 2324
rect 8596 2268 8606 2324
rect 8764 2268 15260 2324
rect 15316 2268 15326 2324
rect 8764 2212 8820 2268
rect 15484 2212 15540 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 38108 2324 38164 2380
rect 17602 2268 17612 2324
rect 17668 2268 21308 2324
rect 21364 2268 21374 2324
rect 23538 2268 23548 2324
rect 23604 2268 24220 2324
rect 24276 2268 24286 2324
rect 24882 2268 24892 2324
rect 24948 2268 25340 2324
rect 25396 2268 25406 2324
rect 28914 2268 28924 2324
rect 28980 2268 33964 2324
rect 34020 2268 34030 2324
rect 34860 2268 37884 2324
rect 37940 2268 37950 2324
rect 38108 2268 43708 2324
rect 24892 2212 24948 2268
rect 34860 2212 34916 2268
rect 3154 2156 3164 2212
rect 3220 2156 5180 2212
rect 5236 2156 5246 2212
rect 6178 2156 6188 2212
rect 6244 2156 6412 2212
rect 6468 2156 6478 2212
rect 7298 2156 7308 2212
rect 7364 2156 8820 2212
rect 9622 2156 9660 2212
rect 9716 2156 9726 2212
rect 12226 2156 12236 2212
rect 12292 2156 14924 2212
rect 14980 2156 14990 2212
rect 15484 2156 19012 2212
rect 19282 2156 19292 2212
rect 19348 2156 19516 2212
rect 19572 2156 19582 2212
rect 19740 2156 20076 2212
rect 20132 2156 22652 2212
rect 22708 2156 22718 2212
rect 22866 2156 22876 2212
rect 22932 2156 24948 2212
rect 25190 2156 25228 2212
rect 25284 2156 25294 2212
rect 26226 2156 26236 2212
rect 26292 2156 26572 2212
rect 26628 2156 26638 2212
rect 27020 2156 34916 2212
rect 35074 2156 35084 2212
rect 35140 2156 35644 2212
rect 35700 2156 35710 2212
rect 36082 2156 36092 2212
rect 36148 2156 37548 2212
rect 37604 2156 37614 2212
rect 38210 2156 38220 2212
rect 38276 2156 38332 2212
rect 38388 2156 38398 2212
rect 40674 2156 40684 2212
rect 40740 2156 40796 2212
rect 40852 2156 40862 2212
rect 42914 2156 42924 2212
rect 42980 2156 43260 2212
rect 43316 2156 43326 2212
rect 0 2100 112 2128
rect 18956 2100 19012 2156
rect 19740 2100 19796 2156
rect 27020 2100 27076 2156
rect 43652 2100 43708 2268
rect 44268 2212 44324 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 48412 2324 48468 2380
rect 45154 2268 45164 2324
rect 45220 2268 47292 2324
rect 47348 2268 47358 2324
rect 47516 2268 48468 2324
rect 47516 2212 47572 2268
rect 44268 2156 45612 2212
rect 45668 2156 45678 2212
rect 46246 2156 46284 2212
rect 46340 2156 46350 2212
rect 47170 2156 47180 2212
rect 47236 2156 47572 2212
rect 48038 2156 48076 2212
rect 48132 2156 48142 2212
rect 48402 2156 48412 2212
rect 48468 2156 49196 2212
rect 49252 2156 49262 2212
rect 57344 2100 57456 2128
rect 0 2044 3276 2100
rect 3332 2044 3342 2100
rect 4722 2044 4732 2100
rect 4788 2044 6188 2100
rect 6244 2044 6254 2100
rect 6626 2044 6636 2100
rect 6692 2044 8428 2100
rect 8530 2044 8540 2100
rect 8596 2044 14588 2100
rect 14644 2044 14654 2100
rect 16828 2044 17724 2100
rect 17780 2044 18060 2100
rect 18116 2044 18126 2100
rect 18246 2044 18284 2100
rect 18340 2044 18350 2100
rect 18956 2044 19796 2100
rect 22530 2044 22540 2100
rect 22596 2044 27076 2100
rect 29586 2044 29596 2100
rect 29652 2044 31948 2100
rect 32946 2044 32956 2100
rect 33012 2044 34188 2100
rect 34244 2044 34254 2100
rect 36082 2044 36092 2100
rect 36148 2044 37884 2100
rect 37940 2044 37950 2100
rect 39554 2044 39564 2100
rect 39620 2044 43484 2100
rect 43540 2044 43550 2100
rect 43652 2044 57456 2100
rect 0 2016 112 2044
rect 8372 1988 8428 2044
rect 16828 1988 16884 2044
rect 31892 1988 31948 2044
rect 57344 2016 57456 2044
rect 2034 1932 2044 1988
rect 2100 1932 8204 1988
rect 8260 1932 8270 1988
rect 8372 1932 9324 1988
rect 9380 1932 9390 1988
rect 9650 1932 9660 1988
rect 9716 1932 10220 1988
rect 10276 1932 10286 1988
rect 10546 1932 10556 1988
rect 10612 1932 12348 1988
rect 12404 1932 12414 1988
rect 12870 1932 12908 1988
rect 12964 1932 14252 1988
rect 14308 1932 14318 1988
rect 15026 1932 15036 1988
rect 15092 1932 16884 1988
rect 17938 1932 17948 1988
rect 18004 1932 18732 1988
rect 18788 1932 18798 1988
rect 19170 1932 19180 1988
rect 19236 1932 19516 1988
rect 19572 1932 19852 1988
rect 19908 1932 19918 1988
rect 23090 1932 23100 1988
rect 23156 1932 25116 1988
rect 25172 1932 25182 1988
rect 25330 1932 25340 1988
rect 25396 1932 30380 1988
rect 30436 1932 30446 1988
rect 31892 1932 36428 1988
rect 36484 1932 36494 1988
rect 42466 1932 42476 1988
rect 42532 1932 45836 1988
rect 45892 1932 45902 1988
rect 46610 1932 46620 1988
rect 46676 1932 49196 1988
rect 49252 1932 49262 1988
rect 2930 1820 2940 1876
rect 2996 1820 3612 1876
rect 3668 1820 3678 1876
rect 4498 1820 4508 1876
rect 4564 1820 11564 1876
rect 11620 1820 11630 1876
rect 33842 1820 33852 1876
rect 33908 1820 36316 1876
rect 36372 1820 36382 1876
rect 43362 1820 43372 1876
rect 43428 1820 46956 1876
rect 47012 1820 47022 1876
rect 48150 1820 48188 1876
rect 48244 1820 48254 1876
rect 1362 1708 1372 1764
rect 1428 1708 1932 1764
rect 1988 1708 13468 1764
rect 13524 1708 13534 1764
rect 14354 1708 14364 1764
rect 14420 1708 16044 1764
rect 16100 1708 16110 1764
rect 18050 1708 18060 1764
rect 18116 1708 18620 1764
rect 18676 1708 18686 1764
rect 19170 1708 19180 1764
rect 19236 1708 21420 1764
rect 21476 1708 21486 1764
rect 21970 1708 21980 1764
rect 22036 1708 25676 1764
rect 25732 1708 25742 1764
rect 31154 1708 31164 1764
rect 31220 1708 34076 1764
rect 34132 1708 34142 1764
rect 35970 1708 35980 1764
rect 36036 1708 40908 1764
rect 40964 1708 40974 1764
rect 41906 1708 41916 1764
rect 41972 1708 47404 1764
rect 47460 1708 47470 1764
rect 0 1652 112 1680
rect 57344 1652 57456 1680
rect 0 1596 3388 1652
rect 3444 1596 3454 1652
rect 6038 1596 6076 1652
rect 6132 1596 6142 1652
rect 6300 1596 7196 1652
rect 7252 1596 7262 1652
rect 7410 1596 7420 1652
rect 7476 1596 7980 1652
rect 8036 1596 8046 1652
rect 8278 1596 8316 1652
rect 8372 1596 8382 1652
rect 9174 1596 9212 1652
rect 9268 1596 9278 1652
rect 11414 1596 11452 1652
rect 11508 1596 11518 1652
rect 11666 1596 11676 1652
rect 11732 1596 11956 1652
rect 12310 1596 12348 1652
rect 12404 1596 12414 1652
rect 13206 1596 13244 1652
rect 13300 1596 13310 1652
rect 14242 1596 14252 1652
rect 14308 1596 14588 1652
rect 14644 1596 14654 1652
rect 14802 1596 14812 1652
rect 14868 1596 15036 1652
rect 15092 1596 15102 1652
rect 15894 1596 15932 1652
rect 15988 1596 15998 1652
rect 16342 1596 16380 1652
rect 16436 1596 16446 1652
rect 16790 1596 16828 1652
rect 16884 1596 16894 1652
rect 17238 1596 17276 1652
rect 17332 1596 17342 1652
rect 18134 1596 18172 1652
rect 18228 1596 18238 1652
rect 20374 1596 20412 1652
rect 20468 1596 20478 1652
rect 20738 1596 20748 1652
rect 20804 1596 21756 1652
rect 21812 1596 21822 1652
rect 23510 1596 23548 1652
rect 23604 1596 23614 1652
rect 24210 1596 24220 1652
rect 24276 1596 30268 1652
rect 30324 1596 30334 1652
rect 31602 1596 31612 1652
rect 31668 1596 35308 1652
rect 35364 1596 35374 1652
rect 38770 1596 38780 1652
rect 38836 1596 40012 1652
rect 40068 1596 40078 1652
rect 44594 1596 44604 1652
rect 44660 1596 47628 1652
rect 47684 1596 47694 1652
rect 50092 1596 57456 1652
rect 0 1568 112 1596
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 6300 1540 6356 1596
rect 11900 1540 11956 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 1110 1484 1148 1540
rect 1204 1484 1214 1540
rect 1558 1484 1596 1540
rect 1652 1484 1662 1540
rect 4386 1484 4396 1540
rect 4452 1484 6356 1540
rect 6962 1484 6972 1540
rect 7028 1484 8204 1540
rect 8260 1484 8270 1540
rect 8754 1484 8764 1540
rect 8820 1484 8988 1540
rect 9044 1484 9054 1540
rect 10994 1484 11004 1540
rect 11060 1484 11676 1540
rect 11732 1484 11742 1540
rect 11900 1484 15036 1540
rect 15092 1484 15102 1540
rect 19954 1484 19964 1540
rect 20020 1484 20860 1540
rect 20916 1484 20926 1540
rect 24322 1484 24332 1540
rect 24388 1484 29932 1540
rect 29988 1484 29998 1540
rect 39442 1484 39452 1540
rect 39508 1484 43708 1540
rect 45154 1484 45164 1540
rect 45220 1484 48636 1540
rect 48692 1484 48702 1540
rect 43652 1428 43708 1484
rect 578 1372 588 1428
rect 644 1372 2940 1428
rect 2996 1372 3006 1428
rect 3332 1372 16380 1428
rect 16436 1372 16446 1428
rect 16594 1372 16604 1428
rect 16660 1372 19516 1428
rect 19572 1372 19582 1428
rect 21634 1372 21644 1428
rect 21700 1372 25004 1428
rect 25060 1372 25070 1428
rect 25778 1372 25788 1428
rect 25844 1372 28812 1428
rect 28868 1372 28878 1428
rect 29138 1372 29148 1428
rect 29204 1372 30044 1428
rect 30100 1372 31724 1428
rect 31780 1372 31790 1428
rect 33954 1372 33964 1428
rect 34020 1372 35532 1428
rect 35588 1372 35598 1428
rect 38770 1372 38780 1428
rect 38836 1372 41132 1428
rect 41188 1372 41198 1428
rect 43652 1372 45276 1428
rect 45332 1372 45342 1428
rect 46722 1372 46732 1428
rect 46788 1372 49868 1428
rect 49924 1372 49934 1428
rect 3332 1316 3388 1372
rect 50092 1316 50148 1596
rect 57344 1568 57456 1596
rect 54338 1484 54348 1540
rect 54404 1484 55804 1540
rect 55860 1484 55870 1540
rect 51874 1372 51884 1428
rect 51940 1372 54460 1428
rect 54516 1372 54526 1428
rect 2594 1260 2604 1316
rect 2660 1260 3388 1316
rect 4274 1260 4284 1316
rect 4340 1260 8148 1316
rect 8418 1260 8428 1316
rect 8484 1260 9884 1316
rect 9940 1260 9950 1316
rect 10220 1260 12796 1316
rect 12852 1260 12862 1316
rect 13010 1260 13020 1316
rect 13076 1260 28028 1316
rect 28084 1260 28094 1316
rect 28690 1260 28700 1316
rect 28756 1260 30156 1316
rect 30212 1260 30222 1316
rect 31892 1260 50148 1316
rect 50866 1260 50876 1316
rect 50932 1260 55356 1316
rect 55412 1260 55422 1316
rect 0 1204 112 1232
rect 8092 1204 8148 1260
rect 10220 1204 10276 1260
rect 31892 1204 31948 1260
rect 57344 1204 57456 1232
rect 0 1148 868 1204
rect 998 1148 1036 1204
rect 1092 1148 1102 1204
rect 1810 1148 1820 1204
rect 1876 1148 2268 1204
rect 2324 1148 2334 1204
rect 3378 1148 3388 1204
rect 3444 1148 4172 1204
rect 4228 1148 4238 1204
rect 4806 1148 4844 1204
rect 4900 1148 4910 1204
rect 5618 1148 5628 1204
rect 5684 1148 5852 1204
rect 5908 1148 5918 1204
rect 6850 1148 6860 1204
rect 6916 1148 7868 1204
rect 7924 1148 7934 1204
rect 8092 1148 8540 1204
rect 8596 1148 8606 1204
rect 8726 1148 8764 1204
rect 8820 1148 8830 1204
rect 9874 1148 9884 1204
rect 9940 1148 10276 1204
rect 10434 1148 10444 1204
rect 10500 1148 12572 1204
rect 12628 1148 12638 1204
rect 15474 1148 15484 1204
rect 15540 1148 16716 1204
rect 16772 1148 16782 1204
rect 18722 1148 18732 1204
rect 18788 1148 24668 1204
rect 24724 1148 24734 1204
rect 24882 1148 24892 1204
rect 24948 1148 26236 1204
rect 26292 1148 26302 1204
rect 30146 1148 30156 1204
rect 30212 1148 31052 1204
rect 31108 1148 31118 1204
rect 31266 1148 31276 1204
rect 31332 1148 31948 1204
rect 34626 1148 34636 1204
rect 34692 1148 36876 1204
rect 36932 1148 36942 1204
rect 37622 1148 37660 1204
rect 37716 1148 37726 1204
rect 39414 1148 39452 1204
rect 39508 1148 39518 1204
rect 43250 1148 43260 1204
rect 43316 1148 46956 1204
rect 47012 1148 47022 1204
rect 55412 1148 57456 1204
rect 0 1120 112 1148
rect 812 980 868 1148
rect 55412 1092 55468 1148
rect 57344 1120 57456 1148
rect 1362 1036 1372 1092
rect 1428 1036 11228 1092
rect 11284 1036 11294 1092
rect 11554 1036 11564 1092
rect 11620 1036 15764 1092
rect 16370 1036 16380 1092
rect 16436 1036 22316 1092
rect 22372 1036 22382 1092
rect 24434 1036 24444 1092
rect 24500 1036 27020 1092
rect 27076 1036 27086 1092
rect 29026 1036 29036 1092
rect 29092 1036 34748 1092
rect 34804 1036 34814 1092
rect 41458 1036 41468 1092
rect 41524 1036 43596 1092
rect 43652 1036 43662 1092
rect 44034 1036 44044 1092
rect 44100 1036 45332 1092
rect 47282 1036 47292 1092
rect 47348 1036 49420 1092
rect 49476 1036 49486 1092
rect 50866 1036 50876 1092
rect 50932 1036 52332 1092
rect 52388 1036 52398 1092
rect 52658 1036 52668 1092
rect 52724 1036 55468 1092
rect 15708 980 15764 1036
rect 812 924 3388 980
rect 3490 924 3500 980
rect 3556 924 5012 980
rect 5170 924 5180 980
rect 5236 924 8092 980
rect 8148 924 8158 980
rect 9986 924 9996 980
rect 10052 924 12516 980
rect 13906 924 13916 980
rect 13972 924 14140 980
rect 14196 924 14206 980
rect 15708 924 18508 980
rect 18564 924 18574 980
rect 21634 924 21644 980
rect 21700 924 23100 980
rect 23156 924 23166 980
rect 23314 924 23324 980
rect 23380 924 26684 980
rect 26740 924 26750 980
rect 27122 924 27132 980
rect 27188 924 28924 980
rect 28980 924 28990 980
rect 30370 924 30380 980
rect 30436 924 34076 980
rect 34132 924 34142 980
rect 37426 924 37436 980
rect 37492 924 39788 980
rect 39844 924 39854 980
rect 40226 924 40236 980
rect 40292 924 45052 980
rect 45108 924 45118 980
rect 3332 868 3388 924
rect 4956 868 5012 924
rect 3332 812 4284 868
rect 4340 812 4350 868
rect 4956 812 11564 868
rect 11620 812 11630 868
rect 0 756 112 784
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 12460 756 12516 924
rect 45276 868 45332 1036
rect 46834 924 46844 980
rect 46900 924 50540 980
rect 50596 924 50606 980
rect 13654 812 13692 868
rect 13748 812 13758 868
rect 13916 812 23324 868
rect 23380 812 23390 868
rect 33394 812 33404 868
rect 33460 812 37324 868
rect 37380 812 37390 868
rect 42354 812 42364 868
rect 42420 812 44324 868
rect 45276 812 52780 868
rect 52836 812 52846 868
rect 13916 756 13972 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 0 700 3388 756
rect 5170 700 5180 756
rect 5236 700 6636 756
rect 6692 700 6702 756
rect 7522 700 7532 756
rect 7588 700 10892 756
rect 10948 700 10958 756
rect 11862 700 11900 756
rect 11956 700 11966 756
rect 12460 700 13972 756
rect 0 672 112 700
rect 3332 644 3388 700
rect 15092 644 15148 756
rect 15204 700 15214 756
rect 15446 700 15484 756
rect 15540 700 15550 756
rect 20626 700 20636 756
rect 20692 700 21308 756
rect 21364 700 21374 756
rect 22614 700 22652 756
rect 22708 700 22718 756
rect 22866 700 22876 756
rect 22932 700 24332 756
rect 24388 700 24398 756
rect 24882 700 24892 756
rect 24948 700 26908 756
rect 30706 700 30716 756
rect 30772 700 34412 756
rect 34468 700 34478 756
rect 38322 700 38332 756
rect 38388 700 40460 756
rect 40516 700 40526 756
rect 26852 644 26908 700
rect 44268 644 44324 812
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 57344 756 57456 784
rect 47702 700 47740 756
rect 47796 700 47806 756
rect 50082 700 50092 756
rect 50148 700 51772 756
rect 51828 700 51838 756
rect 52098 700 52108 756
rect 52164 700 57456 756
rect 57344 672 57456 700
rect 2034 588 2044 644
rect 2100 588 2156 644
rect 2212 588 2222 644
rect 2454 588 2492 644
rect 2548 588 2558 644
rect 3332 588 15148 644
rect 21410 588 21420 644
rect 21476 588 25340 644
rect 25396 588 25406 644
rect 26852 588 44044 644
rect 44100 588 44110 644
rect 44268 588 48300 644
rect 48356 588 48366 644
rect 49970 588 49980 644
rect 50036 588 54012 644
rect 54068 588 54078 644
rect 3266 476 3276 532
rect 3332 476 16268 532
rect 16324 476 16334 532
rect 20626 476 20636 532
rect 20692 476 24892 532
rect 24948 476 24958 532
rect 25106 476 25116 532
rect 25172 476 27580 532
rect 27636 476 27646 532
rect 28354 476 28364 532
rect 28420 476 29372 532
rect 29428 476 29438 532
rect 32050 476 32060 532
rect 32116 476 35980 532
rect 36036 476 36046 532
rect 36530 476 36540 532
rect 36596 476 39116 532
rect 39172 476 39182 532
rect 41010 476 41020 532
rect 41076 476 46732 532
rect 46788 476 46798 532
rect 5394 364 5404 420
rect 5460 364 13020 420
rect 13076 364 13086 420
rect 15138 364 15148 420
rect 15204 364 19068 420
rect 19124 364 19134 420
rect 22754 364 22764 420
rect 22820 364 26236 420
rect 26292 364 26302 420
rect 34738 364 34748 420
rect 34804 364 37212 420
rect 37268 364 37278 420
rect 39218 364 39228 420
rect 39284 364 43148 420
rect 43204 364 43214 420
rect 44146 364 44156 420
rect 44212 364 49644 420
rect 49700 364 49710 420
rect 0 308 112 336
rect 57344 308 57456 336
rect 0 252 7308 308
rect 7364 252 7374 308
rect 7718 252 7756 308
rect 7812 252 7822 308
rect 7970 252 7980 308
rect 8036 252 15148 308
rect 23202 252 23212 308
rect 23268 252 24444 308
rect 24500 252 24510 308
rect 26450 252 26460 308
rect 26516 252 28476 308
rect 28532 252 28542 308
rect 30258 252 30268 308
rect 30324 252 33516 308
rect 33572 252 33582 308
rect 34290 252 34300 308
rect 34356 252 37996 308
rect 38052 252 38062 308
rect 43810 252 43820 308
rect 43876 252 48972 308
rect 49028 252 49038 308
rect 50306 252 50316 308
rect 50372 252 57456 308
rect 0 224 112 252
rect 15092 196 15148 252
rect 57344 224 57456 252
rect 7186 140 7196 196
rect 7252 140 10332 196
rect 10388 140 12908 196
rect 12964 140 12974 196
rect 15092 140 30492 196
rect 30548 140 30558 196
rect 32498 140 32508 196
rect 32564 140 36764 196
rect 36820 140 36830 196
rect 39778 140 39788 196
rect 39844 140 49980 196
rect 50036 140 50046 196
rect 54226 140 54236 196
rect 54292 140 54302 196
rect 54236 84 54292 140
rect 7634 28 7644 84
rect 7700 28 10780 84
rect 10836 28 10846 84
rect 13458 28 13468 84
rect 13524 28 22876 84
rect 22932 28 22942 84
rect 24266 28 24276 84
rect 24332 28 32732 84
rect 32788 28 32798 84
rect 36754 28 36764 84
rect 36820 28 54292 84
<< via3 >>
rect 46844 57372 46900 57428
rect 48524 57372 48580 57428
rect 45276 57260 45332 57316
rect 6188 57148 6244 57204
rect 22764 57148 22820 57204
rect 21308 57036 21364 57092
rect 38444 57036 38500 57092
rect 46844 57036 46900 57092
rect 16492 56924 16548 56980
rect 27804 56812 27860 56868
rect 44268 56812 44324 56868
rect 476 56700 532 56756
rect 55804 56700 55860 56756
rect 44828 56588 44884 56644
rect 48636 56476 48692 56532
rect 52444 56476 52500 56532
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 43804 56420 43860 56476
rect 43908 56420 43964 56476
rect 44012 56420 44068 56476
rect 3388 56364 3444 56420
rect 34972 56364 35028 56420
rect 42812 56364 42868 56420
rect 252 56252 308 56308
rect 5068 56252 5124 56308
rect 44156 56252 44212 56308
rect 46284 56140 46340 56196
rect 2940 56028 2996 56084
rect 27132 56028 27188 56084
rect 31724 56028 31780 56084
rect 32508 56028 32564 56084
rect 33404 56028 33460 56084
rect 34748 56028 34804 56084
rect 42364 56028 42420 56084
rect 812 55804 868 55860
rect 21980 55916 22036 55972
rect 25900 55916 25956 55972
rect 43036 55916 43092 55972
rect 45948 55916 46004 55972
rect 26460 55804 26516 55860
rect 29596 55804 29652 55860
rect 30044 55804 30100 55860
rect 32284 55804 32340 55860
rect 34300 55804 34356 55860
rect 35756 55804 35812 55860
rect 37324 55804 37380 55860
rect 38556 55804 38612 55860
rect 39116 55804 39172 55860
rect 44940 55804 44996 55860
rect 47404 55804 47460 55860
rect 52108 55804 52164 55860
rect 54348 55804 54404 55860
rect 55580 55804 55636 55860
rect 13356 55692 13412 55748
rect 28812 55692 28868 55748
rect 35196 55692 35252 55748
rect 44156 55692 44212 55748
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 44464 55636 44520 55692
rect 44568 55636 44624 55692
rect 44672 55636 44728 55692
rect 4956 55580 5012 55636
rect 14812 55580 14868 55636
rect 41468 55580 41524 55636
rect 43260 55580 43316 55636
rect 45052 55580 45108 55636
rect 45500 55580 45556 55636
rect 9436 55468 9492 55524
rect 9660 55468 9716 55524
rect 25788 55468 25844 55524
rect 27580 55468 27636 55524
rect 28028 55468 28084 55524
rect 29372 55468 29428 55524
rect 30716 55468 30772 55524
rect 34524 55468 34580 55524
rect 35420 55468 35476 55524
rect 38332 55468 38388 55524
rect 40236 55468 40292 55524
rect 46060 55468 46116 55524
rect 46844 55468 46900 55524
rect 47292 55468 47348 55524
rect 48972 55468 49028 55524
rect 49420 55468 49476 55524
rect 49980 55468 50036 55524
rect 50876 55468 50932 55524
rect 1708 55356 1764 55412
rect 6860 55356 6916 55412
rect 30156 55356 30212 55412
rect 30492 55356 30548 55412
rect 30828 55356 30884 55412
rect 33852 55356 33908 55412
rect 34188 55356 34244 55412
rect 36316 55356 36372 55412
rect 37884 55356 37940 55412
rect 39452 55356 39508 55412
rect 40684 55356 40740 55412
rect 52444 55356 52500 55412
rect 3052 55244 3108 55300
rect 3276 55244 3332 55300
rect 8204 55244 8260 55300
rect 8540 55244 8596 55300
rect 10444 55244 10500 55300
rect 14812 55244 14868 55300
rect 15596 55244 15652 55300
rect 19740 55244 19796 55300
rect 21644 55244 21700 55300
rect 22540 55244 22596 55300
rect 26908 55244 26964 55300
rect 32172 55244 32228 55300
rect 32732 55244 32788 55300
rect 44156 55244 44212 55300
rect 46396 55244 46452 55300
rect 54012 55244 54068 55300
rect 33180 55132 33236 55188
rect 51436 55132 51492 55188
rect 4284 55020 4340 55076
rect 13132 55020 13188 55076
rect 13468 55020 13524 55076
rect 15372 55020 15428 55076
rect 18284 55020 18340 55076
rect 41356 55020 41412 55076
rect 140 54908 196 54964
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 3388 54796 3444 54852
rect 20636 54796 20692 54852
rect 33292 54908 33348 54964
rect 48188 54908 48244 54964
rect 43804 54852 43860 54908
rect 43908 54852 43964 54908
rect 44012 54852 44068 54908
rect 30380 54796 30436 54852
rect 32396 54796 32452 54852
rect 37772 54796 37828 54852
rect 43484 54796 43540 54852
rect 45388 54796 45444 54852
rect 12796 54684 12852 54740
rect 48524 54684 48580 54740
rect 51996 54684 52052 54740
rect 13356 54572 13412 54628
rect 32844 54572 32900 54628
rect 36540 54572 36596 54628
rect 38780 54572 38836 54628
rect 39900 54572 39956 54628
rect 1372 54460 1428 54516
rect 40908 54460 40964 54516
rect 46172 54460 46228 54516
rect 50092 54460 50148 54516
rect 54684 54460 54740 54516
rect 2492 54348 2548 54404
rect 5964 54348 6020 54404
rect 8988 54348 9044 54404
rect 18620 54348 18676 54404
rect 26684 54348 26740 54404
rect 9772 54236 9828 54292
rect 14476 54236 14532 54292
rect 15148 54236 15204 54292
rect 15372 54236 15428 54292
rect 23436 54236 23492 54292
rect 27244 54236 27300 54292
rect 27916 54236 27972 54292
rect 32396 54236 32452 54292
rect 33068 54236 33124 54292
rect 36876 54236 36932 54292
rect 40460 54236 40516 54292
rect 55468 54236 55524 54292
rect 55692 54236 55748 54292
rect 7644 54124 7700 54180
rect 7868 54124 7924 54180
rect 14028 54124 14084 54180
rect 20860 54124 20916 54180
rect 1260 54012 1316 54068
rect 3612 54012 3668 54068
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 44464 54068 44520 54124
rect 44568 54068 44624 54124
rect 44672 54068 44728 54124
rect 18732 54012 18788 54068
rect 19964 54012 20020 54068
rect 20188 54012 20244 54068
rect 36652 54012 36708 54068
rect 36876 54012 36932 54068
rect 43372 54012 43428 54068
rect 48524 54012 48580 54068
rect 48860 54012 48916 54068
rect 6412 53900 6468 53956
rect 8428 53900 8484 53956
rect 35084 53900 35140 53956
rect 43484 53900 43540 53956
rect 53788 53900 53844 53956
rect 3388 53788 3444 53844
rect 7308 53788 7364 53844
rect 25564 53788 25620 53844
rect 26796 53788 26852 53844
rect 35532 53788 35588 53844
rect 36764 53788 36820 53844
rect 43596 53788 43652 53844
rect 12460 53676 12516 53732
rect 13804 53676 13860 53732
rect 14252 53676 14308 53732
rect 22092 53676 22148 53732
rect 22988 53676 23044 53732
rect 6636 53564 6692 53620
rect 11564 53564 11620 53620
rect 20188 53564 20244 53620
rect 21084 53564 21140 53620
rect 25228 53564 25284 53620
rect 3388 53452 3444 53508
rect 6972 53452 7028 53508
rect 11676 53452 11732 53508
rect 23324 53452 23380 53508
rect 31500 53676 31556 53732
rect 47516 53676 47572 53732
rect 50764 53676 50820 53732
rect 51548 53676 51604 53732
rect 52556 53676 52612 53732
rect 53900 53676 53956 53732
rect 48524 53564 48580 53620
rect 3500 53340 3556 53396
rect 7420 53340 7476 53396
rect 9996 53340 10052 53396
rect 20300 53340 20356 53396
rect 30604 53452 30660 53508
rect 31164 53452 31220 53508
rect 51100 53452 51156 53508
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 26796 53340 26852 53396
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 4172 53228 4228 53284
rect 6076 53228 6132 53284
rect 8652 53228 8708 53284
rect 10668 53228 10724 53284
rect 14252 53228 14308 53284
rect 24220 53228 24276 53284
rect 43372 53228 43428 53284
rect 43804 53284 43860 53340
rect 43908 53284 43964 53340
rect 44012 53284 44068 53340
rect 53452 53228 53508 53284
rect 8428 53116 8484 53172
rect 13244 53116 13300 53172
rect 15596 53116 15652 53172
rect 17724 53116 17780 53172
rect 19852 53116 19908 53172
rect 31836 53116 31892 53172
rect 45164 53116 45220 53172
rect 3164 53004 3220 53060
rect 7308 53004 7364 53060
rect 13580 53004 13636 53060
rect 42700 53004 42756 53060
rect 45724 53004 45780 53060
rect 45948 53004 46004 53060
rect 50092 53004 50148 53060
rect 51324 53004 51380 53060
rect 1932 52892 1988 52948
rect 2828 52892 2884 52948
rect 4172 52892 4228 52948
rect 6972 52892 7028 52948
rect 16268 52892 16324 52948
rect 17724 52892 17780 52948
rect 35868 52892 35924 52948
rect 55244 52892 55300 52948
rect 2604 52780 2660 52836
rect 3276 52780 3332 52836
rect 6748 52780 6804 52836
rect 15708 52780 15764 52836
rect 31164 52780 31220 52836
rect 5852 52668 5908 52724
rect 6076 52668 6132 52724
rect 7868 52668 7924 52724
rect 19628 52668 19684 52724
rect 19852 52668 19908 52724
rect 22316 52668 22372 52724
rect 29036 52668 29092 52724
rect 37436 52668 37492 52724
rect 41804 52668 41860 52724
rect 43372 52668 43428 52724
rect 16380 52556 16436 52612
rect 18172 52556 18228 52612
rect 19964 52556 20020 52612
rect 24220 52556 24276 52612
rect 26124 52556 26180 52612
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 44464 52500 44520 52556
rect 44568 52500 44624 52556
rect 44672 52500 44728 52556
rect 50988 52780 51044 52836
rect 48300 52668 48356 52724
rect 49196 52668 49252 52724
rect 56924 52668 56980 52724
rect 48636 52556 48692 52612
rect 33292 52444 33348 52500
rect 35084 52444 35140 52500
rect 41356 52444 41412 52500
rect 48412 52444 48468 52500
rect 48860 52444 48916 52500
rect 53116 52444 53172 52500
rect 3500 52332 3556 52388
rect 8092 52332 8148 52388
rect 8988 52332 9044 52388
rect 12124 52332 12180 52388
rect 16716 52332 16772 52388
rect 16940 52332 16996 52388
rect 25004 52332 25060 52388
rect 25900 52332 25956 52388
rect 26572 52332 26628 52388
rect 29708 52332 29764 52388
rect 43036 52332 43092 52388
rect 6636 52220 6692 52276
rect 10668 52220 10724 52276
rect 17052 52220 17108 52276
rect 32620 52220 32676 52276
rect 34636 52220 34692 52276
rect 35868 52220 35924 52276
rect 37436 52220 37492 52276
rect 40348 52220 40404 52276
rect 40572 52220 40628 52276
rect 50988 52220 51044 52276
rect 51884 52220 51940 52276
rect 2604 52108 2660 52164
rect 14252 52108 14308 52164
rect 14924 52108 14980 52164
rect 19180 52108 19236 52164
rect 21532 52108 21588 52164
rect 25900 52108 25956 52164
rect 4172 51996 4228 52052
rect 5964 51996 6020 52052
rect 7308 51996 7364 52052
rect 29708 52108 29764 52164
rect 30828 52108 30884 52164
rect 32956 52108 33012 52164
rect 34412 52108 34468 52164
rect 45612 52108 45668 52164
rect 54124 52108 54180 52164
rect 20972 51996 21028 52052
rect 29484 51996 29540 52052
rect 40796 51996 40852 52052
rect 49644 51996 49700 52052
rect 52668 51996 52724 52052
rect 3388 51884 3444 51940
rect 10108 51884 10164 51940
rect 1932 51772 1988 51828
rect 14252 51772 14308 51828
rect 14924 51772 14980 51828
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 4172 51660 4228 51716
rect 13580 51660 13636 51716
rect 23100 51660 23156 51716
rect 43804 51716 43860 51772
rect 43908 51716 43964 51772
rect 44012 51716 44068 51772
rect 54236 51660 54292 51716
rect 55132 51660 55188 51716
rect 1596 51548 1652 51604
rect 12124 51548 12180 51604
rect 49868 51548 49924 51604
rect 50092 51548 50148 51604
rect 55356 51548 55412 51604
rect 57260 51548 57316 51604
rect 3388 51436 3444 51492
rect 7420 51436 7476 51492
rect 3612 51324 3668 51380
rect 8428 51324 8484 51380
rect 15484 51324 15540 51380
rect 45164 51436 45220 51492
rect 50204 51436 50260 51492
rect 30044 51324 30100 51380
rect 30268 51324 30324 51380
rect 31164 51324 31220 51380
rect 32732 51324 32788 51380
rect 33964 51324 34020 51380
rect 45948 51324 46004 51380
rect 50316 51324 50372 51380
rect 51660 51324 51716 51380
rect 10668 51212 10724 51268
rect 12684 51212 12740 51268
rect 15036 51212 15092 51268
rect 29820 51212 29876 51268
rect 32620 51212 32676 51268
rect 38220 51212 38276 51268
rect 52780 51436 52836 51492
rect 54460 51324 54516 51380
rect 40348 51212 40404 51268
rect 41916 51212 41972 51268
rect 2380 51100 2436 51156
rect 3388 51100 3444 51156
rect 6524 51100 6580 51156
rect 23212 51100 23268 51156
rect 30044 51100 30100 51156
rect 33516 51100 33572 51156
rect 34860 51100 34916 51156
rect 40124 51100 40180 51156
rect 43372 51100 43428 51156
rect 50204 51100 50260 51156
rect 53676 51100 53732 51156
rect 54236 51100 54292 51156
rect 57148 51100 57204 51156
rect 7084 50988 7140 51044
rect 23660 50988 23716 51044
rect 28588 50988 28644 51044
rect 41580 50988 41636 51044
rect 43484 50988 43540 51044
rect 44268 50988 44324 51044
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 44464 50932 44520 50988
rect 44568 50932 44624 50988
rect 44672 50932 44728 50988
rect 2716 50876 2772 50932
rect 3500 50876 3556 50932
rect 23548 50876 23604 50932
rect 33292 50876 33348 50932
rect 50092 50876 50148 50932
rect 50428 50876 50484 50932
rect 51212 50876 51268 50932
rect 52444 50876 52500 50932
rect 52668 50876 52724 50932
rect 55356 50876 55412 50932
rect 5404 50764 5460 50820
rect 30268 50764 30324 50820
rect 32732 50764 32788 50820
rect 50204 50764 50260 50820
rect 50540 50764 50596 50820
rect 53564 50764 53620 50820
rect 5292 50652 5348 50708
rect 12348 50652 12404 50708
rect 15036 50652 15092 50708
rect 25340 50652 25396 50708
rect 30940 50652 30996 50708
rect 50764 50652 50820 50708
rect 54796 50764 54852 50820
rect 55020 50764 55076 50820
rect 54236 50652 54292 50708
rect 7868 50540 7924 50596
rect 15260 50540 15316 50596
rect 24220 50540 24276 50596
rect 25004 50540 25060 50596
rect 29260 50540 29316 50596
rect 32396 50540 32452 50596
rect 43596 50540 43652 50596
rect 44268 50540 44324 50596
rect 48524 50540 48580 50596
rect 51212 50540 51268 50596
rect 52332 50540 52388 50596
rect 54796 50540 54852 50596
rect 1820 50428 1876 50484
rect 3276 50428 3332 50484
rect 12348 50428 12404 50484
rect 12684 50428 12740 50484
rect 1148 50316 1204 50372
rect 6076 50316 6132 50372
rect 8764 50316 8820 50372
rect 26460 50428 26516 50484
rect 29932 50428 29988 50484
rect 38892 50428 38948 50484
rect 43372 50428 43428 50484
rect 45948 50428 46004 50484
rect 49532 50428 49588 50484
rect 51996 50428 52052 50484
rect 52780 50428 52836 50484
rect 53004 50428 53060 50484
rect 12460 50316 12516 50372
rect 23100 50316 23156 50372
rect 26796 50316 26852 50372
rect 29484 50316 29540 50372
rect 37548 50316 37604 50372
rect 37772 50316 37828 50372
rect 43148 50316 43204 50372
rect 49644 50316 49700 50372
rect 50652 50316 50708 50372
rect 51436 50316 51492 50372
rect 52220 50316 52276 50372
rect 16828 50204 16884 50260
rect 20860 50204 20916 50260
rect 22652 50204 22708 50260
rect 23660 50204 23716 50260
rect 41804 50204 41860 50260
rect 44156 50204 44212 50260
rect 45164 50204 45220 50260
rect 48748 50204 48804 50260
rect 52556 50204 52612 50260
rect 52892 50204 52948 50260
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 43804 50148 43860 50204
rect 43908 50148 43964 50204
rect 44012 50148 44068 50204
rect 19740 50092 19796 50148
rect 28140 50092 28196 50148
rect 30044 50092 30100 50148
rect 31612 50092 31668 50148
rect 36540 50092 36596 50148
rect 54460 50092 54516 50148
rect 700 49980 756 50036
rect 12012 49980 12068 50036
rect 24220 49980 24276 50036
rect 34972 49980 35028 50036
rect 2044 49868 2100 49924
rect 10892 49868 10948 49924
rect 2268 49756 2324 49812
rect 8428 49756 8484 49812
rect 9100 49756 9156 49812
rect 10220 49756 10276 49812
rect 12012 49756 12068 49812
rect 16940 49756 16996 49812
rect 18844 49756 18900 49812
rect 23660 49756 23716 49812
rect 29036 49756 29092 49812
rect 38444 49756 38500 49812
rect 41356 49756 41412 49812
rect 1596 49644 1652 49700
rect 4956 49644 5012 49700
rect 16492 49644 16548 49700
rect 17052 49644 17108 49700
rect 25228 49644 25284 49700
rect 34636 49644 34692 49700
rect 41804 49644 41860 49700
rect 42140 49644 42196 49700
rect 43148 49644 43204 49700
rect 51212 49644 51268 49700
rect 55804 49644 55860 49700
rect 13580 49532 13636 49588
rect 18172 49532 18228 49588
rect 18956 49532 19012 49588
rect 22428 49532 22484 49588
rect 23212 49532 23268 49588
rect 24220 49532 24276 49588
rect 29708 49532 29764 49588
rect 30604 49532 30660 49588
rect 37100 49532 37156 49588
rect 38892 49532 38948 49588
rect 52332 49532 52388 49588
rect 52556 49532 52612 49588
rect 56588 49532 56644 49588
rect 2380 49420 2436 49476
rect 7980 49420 8036 49476
rect 18508 49420 18564 49476
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 2716 49308 2772 49364
rect 3612 49308 3668 49364
rect 6188 49308 6244 49364
rect 38220 49420 38276 49476
rect 38444 49420 38500 49476
rect 42028 49420 42084 49476
rect 51772 49420 51828 49476
rect 56028 49420 56084 49476
rect 44464 49364 44520 49420
rect 44568 49364 44624 49420
rect 44672 49364 44728 49420
rect 28140 49308 28196 49364
rect 30940 49308 30996 49364
rect 31388 49308 31444 49364
rect 32172 49308 32228 49364
rect 34076 49308 34132 49364
rect 34300 49308 34356 49364
rect 3388 49196 3444 49252
rect 6076 49196 6132 49252
rect 11340 49196 11396 49252
rect 14588 49196 14644 49252
rect 19852 49196 19908 49252
rect 30604 49196 30660 49252
rect 34188 49196 34244 49252
rect 45724 49196 45780 49252
rect 49980 49196 50036 49252
rect 1596 49084 1652 49140
rect 1932 49084 1988 49140
rect 2716 49084 2772 49140
rect 5068 49084 5124 49140
rect 6748 49084 6804 49140
rect 10668 49084 10724 49140
rect 15484 49084 15540 49140
rect 17052 49084 17108 49140
rect 22204 49084 22260 49140
rect 30380 49084 30436 49140
rect 34636 49084 34692 49140
rect 2268 48972 2324 49028
rect 3500 48972 3556 49028
rect 12460 48972 12516 49028
rect 15036 48972 15092 49028
rect 16044 48972 16100 49028
rect 45388 48972 45444 49028
rect 4284 48860 4340 48916
rect 5180 48860 5236 48916
rect 19180 48860 19236 48916
rect 20748 48860 20804 48916
rect 22204 48860 22260 48916
rect 26796 48860 26852 48916
rect 41580 48860 41636 48916
rect 44156 48860 44212 48916
rect 45836 48860 45892 48916
rect 46620 48860 46676 48916
rect 48636 48860 48692 48916
rect 51100 48860 51156 48916
rect 53676 48860 53732 48916
rect 812 48748 868 48804
rect 3164 48748 3220 48804
rect 5516 48748 5572 48804
rect 35084 48748 35140 48804
rect 45724 48748 45780 48804
rect 11004 48636 11060 48692
rect 12796 48636 12852 48692
rect 15484 48636 15540 48692
rect 16492 48636 16548 48692
rect 26572 48636 26628 48692
rect 27692 48636 27748 48692
rect 40796 48636 40852 48692
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 43804 48580 43860 48636
rect 43908 48580 43964 48636
rect 44012 48580 44068 48636
rect 11228 48524 11284 48580
rect 17500 48524 17556 48580
rect 20972 48524 21028 48580
rect 24220 48524 24276 48580
rect 28364 48524 28420 48580
rect 30604 48524 30660 48580
rect 31500 48524 31556 48580
rect 33964 48524 34020 48580
rect 44156 48524 44212 48580
rect 53340 48524 53396 48580
rect 1708 48412 1764 48468
rect 2044 48412 2100 48468
rect 3164 48412 3220 48468
rect 5068 48412 5124 48468
rect 19852 48412 19908 48468
rect 23548 48412 23604 48468
rect 25340 48412 25396 48468
rect 30044 48412 30100 48468
rect 32284 48412 32340 48468
rect 49196 48412 49252 48468
rect 7980 48300 8036 48356
rect 12348 48300 12404 48356
rect 21980 48300 22036 48356
rect 34860 48300 34916 48356
rect 35308 48300 35364 48356
rect 48748 48300 48804 48356
rect 53116 48300 53172 48356
rect 54908 48300 54964 48356
rect 2380 48188 2436 48244
rect 10892 48188 10948 48244
rect 11452 48188 11508 48244
rect 20972 48188 21028 48244
rect 29484 48188 29540 48244
rect 31388 48188 31444 48244
rect 41916 48188 41972 48244
rect 48300 48188 48356 48244
rect 49308 48188 49364 48244
rect 51212 48188 51268 48244
rect 16828 48076 16884 48132
rect 25676 48076 25732 48132
rect 26124 48076 26180 48132
rect 35308 48076 35364 48132
rect 53788 48188 53844 48244
rect 7756 47964 7812 48020
rect 10332 47964 10388 48020
rect 13468 47964 13524 48020
rect 13692 47964 13748 48020
rect 19180 47964 19236 48020
rect 20076 47964 20132 48020
rect 21420 47964 21476 48020
rect 30380 47964 30436 48020
rect 31276 47964 31332 48020
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 38220 47852 38276 47908
rect 43148 47852 43204 47908
rect 43596 47852 43652 47908
rect 44464 47796 44520 47852
rect 44568 47796 44624 47852
rect 44672 47796 44728 47852
rect 1708 47740 1764 47796
rect 3612 47740 3668 47796
rect 13468 47740 13524 47796
rect 15036 47740 15092 47796
rect 29596 47740 29652 47796
rect 32396 47740 32452 47796
rect 32844 47740 32900 47796
rect 50092 47740 50148 47796
rect 51324 47740 51380 47796
rect 55020 47740 55076 47796
rect 4172 47628 4228 47684
rect 6076 47628 6132 47684
rect 9212 47628 9268 47684
rect 11228 47628 11284 47684
rect 18060 47628 18116 47684
rect 28364 47628 28420 47684
rect 34076 47628 34132 47684
rect 43596 47628 43652 47684
rect 17164 47516 17220 47572
rect 53004 47628 53060 47684
rect 53676 47628 53732 47684
rect 44268 47516 44324 47572
rect 49980 47516 50036 47572
rect 20636 47404 20692 47460
rect 26460 47404 26516 47460
rect 28476 47404 28532 47460
rect 29260 47404 29316 47460
rect 29484 47404 29540 47460
rect 43596 47404 43652 47460
rect 52444 47404 52500 47460
rect 3388 47292 3444 47348
rect 5180 47292 5236 47348
rect 16492 47292 16548 47348
rect 30268 47292 30324 47348
rect 33180 47292 33236 47348
rect 34860 47292 34916 47348
rect 47964 47292 48020 47348
rect 48188 47292 48244 47348
rect 51436 47292 51492 47348
rect 7756 47180 7812 47236
rect 18508 47180 18564 47236
rect 29596 47180 29652 47236
rect 6748 47068 6804 47124
rect 7420 47068 7476 47124
rect 7868 47068 7924 47124
rect 10332 47068 10388 47124
rect 13020 47068 13076 47124
rect 22764 47068 22820 47124
rect 26460 47068 26516 47124
rect 49084 47068 49140 47124
rect 50204 47068 50260 47124
rect 52668 47068 52724 47124
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 43804 47012 43860 47068
rect 43908 47012 43964 47068
rect 44012 47012 44068 47068
rect 1932 46956 1988 47012
rect 3612 46956 3668 47012
rect 14252 46956 14308 47012
rect 14812 46956 14868 47012
rect 28252 46956 28308 47012
rect 34972 46956 35028 47012
rect 37100 46956 37156 47012
rect 40012 46956 40068 47012
rect 41020 46956 41076 47012
rect 43372 46956 43428 47012
rect 44156 46956 44212 47012
rect 48300 46956 48356 47012
rect 22764 46844 22820 46900
rect 3388 46732 3444 46788
rect 3612 46732 3668 46788
rect 5740 46732 5796 46788
rect 14588 46732 14644 46788
rect 15036 46732 15092 46788
rect 27020 46732 27076 46788
rect 7756 46620 7812 46676
rect 10220 46620 10276 46676
rect 12908 46620 12964 46676
rect 14252 46620 14308 46676
rect 25116 46620 25172 46676
rect 924 46508 980 46564
rect 13804 46508 13860 46564
rect 14924 46508 14980 46564
rect 21980 46508 22036 46564
rect 25004 46508 25060 46564
rect 31612 46844 31668 46900
rect 34636 46844 34692 46900
rect 49196 46844 49252 46900
rect 49644 46844 49700 46900
rect 50652 46956 50708 47012
rect 55020 46956 55076 47012
rect 55804 46844 55860 46900
rect 29036 46732 29092 46788
rect 30156 46732 30212 46788
rect 31948 46732 32004 46788
rect 49420 46732 49476 46788
rect 50316 46732 50372 46788
rect 53004 46732 53060 46788
rect 30828 46620 30884 46676
rect 32844 46620 32900 46676
rect 36764 46620 36820 46676
rect 41804 46620 41860 46676
rect 53116 46620 53172 46676
rect 56252 46620 56308 46676
rect 28140 46508 28196 46564
rect 40124 46508 40180 46564
rect 40572 46508 40628 46564
rect 45164 46508 45220 46564
rect 364 46396 420 46452
rect 3388 46396 3444 46452
rect 5740 46396 5796 46452
rect 10892 46396 10948 46452
rect 14588 46396 14644 46452
rect 15932 46396 15988 46452
rect 17276 46396 17332 46452
rect 18172 46396 18228 46452
rect 28924 46396 28980 46452
rect 35644 46396 35700 46452
rect 36092 46396 36148 46452
rect 41692 46396 41748 46452
rect 42476 46396 42532 46452
rect 46956 46396 47012 46452
rect 48300 46396 48356 46452
rect 49644 46396 49700 46452
rect 5180 46284 5236 46340
rect 11340 46284 11396 46340
rect 16828 46284 16884 46340
rect 29036 46284 29092 46340
rect 31388 46284 31444 46340
rect 36764 46284 36820 46340
rect 41580 46284 41636 46340
rect 44156 46284 44212 46340
rect 47180 46284 47236 46340
rect 48748 46284 48804 46340
rect 49868 46284 49924 46340
rect 51212 46284 51268 46340
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 44464 46228 44520 46284
rect 44568 46228 44624 46284
rect 44672 46228 44728 46284
rect 17500 46172 17556 46228
rect 49084 46172 49140 46228
rect 51884 46172 51940 46228
rect 9996 46060 10052 46116
rect 12236 46060 12292 46116
rect 12908 46060 12964 46116
rect 14252 46060 14308 46116
rect 14812 46060 14868 46116
rect 23212 46060 23268 46116
rect 27468 46060 27524 46116
rect 28924 46060 28980 46116
rect 30828 46060 30884 46116
rect 32844 46060 32900 46116
rect 34636 46060 34692 46116
rect 35532 46060 35588 46116
rect 35980 46060 36036 46116
rect 39228 46060 39284 46116
rect 55804 46060 55860 46116
rect 1148 45948 1204 46004
rect 2044 45948 2100 46004
rect 3500 45948 3556 46004
rect 5628 45948 5684 46004
rect 7420 45948 7476 46004
rect 14924 45948 14980 46004
rect 21196 45948 21252 46004
rect 21532 45948 21588 46004
rect 28364 45948 28420 46004
rect 37772 45948 37828 46004
rect 42476 45948 42532 46004
rect 49084 45948 49140 46004
rect 49532 45948 49588 46004
rect 49868 45948 49924 46004
rect 50540 45948 50596 46004
rect 54908 45948 54964 46004
rect 3388 45836 3444 45892
rect 9884 45836 9940 45892
rect 11788 45836 11844 45892
rect 22092 45836 22148 45892
rect 23100 45836 23156 45892
rect 24892 45836 24948 45892
rect 30828 45836 30884 45892
rect 37660 45836 37716 45892
rect 39564 45836 39620 45892
rect 41916 45836 41972 45892
rect 49196 45836 49252 45892
rect 25564 45724 25620 45780
rect 54908 45724 54964 45780
rect 3276 45612 3332 45668
rect 7532 45612 7588 45668
rect 8988 45612 9044 45668
rect 11452 45612 11508 45668
rect 21196 45612 21252 45668
rect 22764 45612 22820 45668
rect 29820 45612 29876 45668
rect 48860 45612 48916 45668
rect 53116 45612 53172 45668
rect 5068 45500 5124 45556
rect 6972 45500 7028 45556
rect 11116 45500 11172 45556
rect 25228 45500 25284 45556
rect 39788 45500 39844 45556
rect 48748 45500 48804 45556
rect 49756 45500 49812 45556
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 43804 45444 43860 45500
rect 43908 45444 43964 45500
rect 44012 45444 44068 45500
rect 6636 45388 6692 45444
rect 25452 45388 25508 45444
rect 27916 45388 27972 45444
rect 31948 45388 32004 45444
rect 33740 45388 33796 45444
rect 34860 45388 34916 45444
rect 35532 45388 35588 45444
rect 42252 45388 42308 45444
rect 45612 45388 45668 45444
rect 51996 45388 52052 45444
rect 4284 45276 4340 45332
rect 5628 45276 5684 45332
rect 6300 45276 6356 45332
rect 53788 45500 53844 45556
rect 55356 45388 55412 45444
rect 31052 45276 31108 45332
rect 41020 45276 41076 45332
rect 42588 45276 42644 45332
rect 47628 45276 47684 45332
rect 50428 45276 50484 45332
rect 53116 45276 53172 45332
rect 56140 45276 56196 45332
rect 3612 45164 3668 45220
rect 4172 45164 4228 45220
rect 4844 45164 4900 45220
rect 6188 45164 6244 45220
rect 8316 45164 8372 45220
rect 13916 45164 13972 45220
rect 17612 45164 17668 45220
rect 21980 45164 22036 45220
rect 22540 45164 22596 45220
rect 23548 45164 23604 45220
rect 38668 45164 38724 45220
rect 39564 45164 39620 45220
rect 56476 45164 56532 45220
rect 3276 45052 3332 45108
rect 3388 45052 3444 45108
rect 14700 45052 14756 45108
rect 16044 45052 16100 45108
rect 21196 45052 21252 45108
rect 33628 45052 33684 45108
rect 41804 45052 41860 45108
rect 42252 45052 42308 45108
rect 1036 44940 1092 44996
rect 5628 44940 5684 44996
rect 16268 44940 16324 44996
rect 18620 44940 18676 44996
rect 22540 44940 22596 44996
rect 27356 44940 27412 44996
rect 30156 44940 30212 44996
rect 40012 44940 40068 44996
rect 48524 44940 48580 44996
rect 49196 44940 49252 44996
rect 50316 44940 50372 44996
rect 51436 44940 51492 44996
rect 4844 44828 4900 44884
rect 10780 44828 10836 44884
rect 22204 44828 22260 44884
rect 39228 44828 39284 44884
rect 42028 44828 42084 44884
rect 2044 44716 2100 44772
rect 6300 44716 6356 44772
rect 11004 44716 11060 44772
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 25900 44716 25956 44772
rect 5180 44604 5236 44660
rect 11116 44604 11172 44660
rect 13580 44604 13636 44660
rect 18956 44604 19012 44660
rect 18172 44492 18228 44548
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 49756 44828 49812 44884
rect 53788 44828 53844 44884
rect 54124 44828 54180 44884
rect 54908 44828 54964 44884
rect 53564 44716 53620 44772
rect 54460 44716 54516 44772
rect 44464 44660 44520 44716
rect 44568 44660 44624 44716
rect 44672 44660 44728 44716
rect 21196 44604 21252 44660
rect 26684 44604 26740 44660
rect 28140 44604 28196 44660
rect 40348 44604 40404 44660
rect 42700 44604 42756 44660
rect 42924 44604 42980 44660
rect 30604 44492 30660 44548
rect 1932 44380 1988 44436
rect 2604 44380 2660 44436
rect 4284 44380 4340 44436
rect 6188 44380 6244 44436
rect 13356 44380 13412 44436
rect 16940 44380 16996 44436
rect 41244 44380 41300 44436
rect 41804 44380 41860 44436
rect 45836 44380 45892 44436
rect 48748 44380 48804 44436
rect 53900 44380 53956 44436
rect 3276 44268 3332 44324
rect 8764 44268 8820 44324
rect 11228 44268 11284 44324
rect 13468 44268 13524 44324
rect 20860 44268 20916 44324
rect 28924 44268 28980 44324
rect 30716 44268 30772 44324
rect 50988 44268 51044 44324
rect 51436 44268 51492 44324
rect 54124 44268 54180 44324
rect 4284 44156 4340 44212
rect 5068 44156 5124 44212
rect 6636 44156 6692 44212
rect 7532 44156 7588 44212
rect 27020 44156 27076 44212
rect 29372 44156 29428 44212
rect 44156 44156 44212 44212
rect 53900 44156 53956 44212
rect 54796 44156 54852 44212
rect 7980 44044 8036 44100
rect 20972 44044 21028 44100
rect 26684 44044 26740 44100
rect 26908 44044 26964 44100
rect 31500 44044 31556 44100
rect 34076 44044 34132 44100
rect 38668 44044 38724 44100
rect 812 43932 868 43988
rect 1596 43932 1652 43988
rect 6972 43932 7028 43988
rect 7868 43932 7924 43988
rect 18508 43932 18564 43988
rect 21308 43932 21364 43988
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 54348 44044 54404 44100
rect 55020 44044 55076 44100
rect 48524 43932 48580 43988
rect 48748 43932 48804 43988
rect 43804 43876 43860 43932
rect 43908 43876 43964 43932
rect 44012 43876 44068 43932
rect 8764 43820 8820 43876
rect 10556 43820 10612 43876
rect 25004 43820 25060 43876
rect 38220 43820 38276 43876
rect 39340 43820 39396 43876
rect 39788 43820 39844 43876
rect 44156 43820 44212 43876
rect 53004 43820 53060 43876
rect 53228 43820 53284 43876
rect 56140 43820 56196 43876
rect 12684 43708 12740 43764
rect 12908 43708 12964 43764
rect 20076 43708 20132 43764
rect 29708 43708 29764 43764
rect 37212 43708 37268 43764
rect 38444 43708 38500 43764
rect 50092 43708 50148 43764
rect 54796 43708 54852 43764
rect 13468 43596 13524 43652
rect 31276 43596 31332 43652
rect 54684 43596 54740 43652
rect 55020 43596 55076 43652
rect 3276 43484 3332 43540
rect 3612 43484 3668 43540
rect 4844 43484 4900 43540
rect 5740 43484 5796 43540
rect 7084 43484 7140 43540
rect 15820 43484 15876 43540
rect 16940 43484 16996 43540
rect 19852 43484 19908 43540
rect 25004 43484 25060 43540
rect 52668 43484 52724 43540
rect 53564 43484 53620 43540
rect 56140 43484 56196 43540
rect 57372 43484 57428 43540
rect 1596 43372 1652 43428
rect 32956 43372 33012 43428
rect 33180 43372 33236 43428
rect 47852 43372 47908 43428
rect 50988 43372 51044 43428
rect 51324 43372 51380 43428
rect 6636 43260 6692 43316
rect 6972 43260 7028 43316
rect 19292 43260 19348 43316
rect 37772 43260 37828 43316
rect 53564 43260 53620 43316
rect 1148 43148 1204 43204
rect 4284 43148 4340 43204
rect 6748 43148 6804 43204
rect 20972 43148 21028 43204
rect 27244 43148 27300 43204
rect 41020 43148 41076 43204
rect 43148 43148 43204 43204
rect 50372 43148 50428 43204
rect 55020 43148 55076 43204
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 3388 43036 3444 43092
rect 9548 43036 9604 43092
rect 28364 43036 28420 43092
rect 40460 43036 40516 43092
rect 42252 43036 42308 43092
rect 44464 43092 44520 43148
rect 44568 43092 44624 43148
rect 44672 43092 44728 43148
rect 52444 43036 52500 43092
rect 54796 43036 54852 43092
rect 700 42924 756 42980
rect 16716 42924 16772 42980
rect 17164 42924 17220 42980
rect 34860 42924 34916 42980
rect 37660 42924 37716 42980
rect 45164 42924 45220 42980
rect 48524 42924 48580 42980
rect 50988 42924 51044 42980
rect 54572 42924 54628 42980
rect 3612 42812 3668 42868
rect 8988 42812 9044 42868
rect 11900 42812 11956 42868
rect 13356 42812 13412 42868
rect 17612 42812 17668 42868
rect 20076 42812 20132 42868
rect 28364 42812 28420 42868
rect 34412 42812 34468 42868
rect 40348 42812 40404 42868
rect 41244 42812 41300 42868
rect 41580 42812 41636 42868
rect 46620 42812 46676 42868
rect 50204 42812 50260 42868
rect 53676 42812 53732 42868
rect 56028 42812 56084 42868
rect 3500 42700 3556 42756
rect 7308 42700 7364 42756
rect 23100 42700 23156 42756
rect 39340 42700 39396 42756
rect 50540 42700 50596 42756
rect 52108 42700 52164 42756
rect 52444 42700 52500 42756
rect 12460 42588 12516 42644
rect 20972 42588 21028 42644
rect 35420 42588 35476 42644
rect 41132 42588 41188 42644
rect 45836 42588 45892 42644
rect 49196 42588 49252 42644
rect 52892 42588 52948 42644
rect 54796 42588 54852 42644
rect 2268 42476 2324 42532
rect 3388 42476 3444 42532
rect 18956 42476 19012 42532
rect 25228 42476 25284 42532
rect 29148 42476 29204 42532
rect 32956 42476 33012 42532
rect 35084 42476 35140 42532
rect 35980 42476 36036 42532
rect 38668 42476 38724 42532
rect 41356 42476 41412 42532
rect 50428 42476 50484 42532
rect 3500 42364 3556 42420
rect 4844 42364 4900 42420
rect 12572 42364 12628 42420
rect 14700 42364 14756 42420
rect 15820 42364 15876 42420
rect 20300 42364 20356 42420
rect 21308 42364 21364 42420
rect 55580 42364 55636 42420
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 43804 42308 43860 42364
rect 43908 42308 43964 42364
rect 44012 42308 44068 42364
rect 9324 42252 9380 42308
rect 22764 42252 22820 42308
rect 27468 42252 27524 42308
rect 28364 42252 28420 42308
rect 38220 42252 38276 42308
rect 44156 42252 44212 42308
rect 45388 42252 45444 42308
rect 2940 42140 2996 42196
rect 48076 42252 48132 42308
rect 51772 42252 51828 42308
rect 52668 42252 52724 42308
rect 52892 42252 52948 42308
rect 53788 42252 53844 42308
rect 10556 42140 10612 42196
rect 13020 42140 13076 42196
rect 14812 42140 14868 42196
rect 47628 42140 47684 42196
rect 50204 42140 50260 42196
rect 50428 42140 50484 42196
rect 52108 42140 52164 42196
rect 12012 42028 12068 42084
rect 13580 42028 13636 42084
rect 25452 42028 25508 42084
rect 31388 42028 31444 42084
rect 53788 42028 53844 42084
rect 55356 42028 55412 42084
rect 55580 42028 55636 42084
rect 56140 42028 56196 42084
rect 56812 42028 56868 42084
rect 19516 41916 19572 41972
rect 24220 41916 24276 41972
rect 31164 41916 31220 41972
rect 32060 41916 32116 41972
rect 32396 41916 32452 41972
rect 32620 41916 32676 41972
rect 34076 41916 34132 41972
rect 41020 41916 41076 41972
rect 46508 41916 46564 41972
rect 46956 41916 47012 41972
rect 1596 41804 1652 41860
rect 4172 41804 4228 41860
rect 5068 41804 5124 41860
rect 5516 41804 5572 41860
rect 8764 41804 8820 41860
rect 29148 41804 29204 41860
rect 37436 41804 37492 41860
rect 2492 41692 2548 41748
rect 18508 41692 18564 41748
rect 22876 41692 22932 41748
rect 30604 41692 30660 41748
rect 47964 41692 48020 41748
rect 49196 41692 49252 41748
rect 53676 41692 53732 41748
rect 55468 41692 55524 41748
rect 812 41580 868 41636
rect 8876 41580 8932 41636
rect 10892 41580 10948 41636
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 41244 41580 41300 41636
rect 44156 41580 44212 41636
rect 49868 41580 49924 41636
rect 53116 41580 53172 41636
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 44464 41524 44520 41580
rect 44568 41524 44624 41580
rect 44672 41524 44728 41580
rect 2380 41468 2436 41524
rect 3052 41468 3108 41524
rect 3612 41468 3668 41524
rect 4172 41468 4228 41524
rect 9548 41468 9604 41524
rect 23212 41468 23268 41524
rect 34748 41468 34804 41524
rect 36764 41468 36820 41524
rect 48860 41468 48916 41524
rect 51548 41468 51604 41524
rect 700 41356 756 41412
rect 6972 41356 7028 41412
rect 19292 41356 19348 41412
rect 40908 41356 40964 41412
rect 55356 41356 55412 41412
rect 56364 41356 56420 41412
rect 13580 41244 13636 41300
rect 13804 41244 13860 41300
rect 14364 41244 14420 41300
rect 1708 41132 1764 41188
rect 2044 41132 2100 41188
rect 39004 41244 39060 41300
rect 41916 41244 41972 41300
rect 49868 41244 49924 41300
rect 52668 41244 52724 41300
rect 54348 41244 54404 41300
rect 5628 41132 5684 41188
rect 8428 41132 8484 41188
rect 9996 41132 10052 41188
rect 12012 41132 12068 41188
rect 13468 41132 13524 41188
rect 26572 41132 26628 41188
rect 28140 41132 28196 41188
rect 29036 41132 29092 41188
rect 29484 41132 29540 41188
rect 30940 41132 30996 41188
rect 36540 41132 36596 41188
rect 43596 41132 43652 41188
rect 44156 41132 44212 41188
rect 45164 41132 45220 41188
rect 46956 41132 47012 41188
rect 55804 41132 55860 41188
rect 57036 41132 57092 41188
rect 4284 41020 4340 41076
rect 23436 41020 23492 41076
rect 24220 41020 24276 41076
rect 31388 41020 31444 41076
rect 33628 41020 33684 41076
rect 33964 41020 34020 41076
rect 35196 41020 35252 41076
rect 50204 41020 50260 41076
rect 3612 40908 3668 40964
rect 8876 40908 8932 40964
rect 9548 40908 9604 40964
rect 14140 40908 14196 40964
rect 16828 40908 16884 40964
rect 22316 40908 22372 40964
rect 29820 40908 29876 40964
rect 3388 40796 3444 40852
rect 6972 40796 7028 40852
rect 35084 40796 35140 40852
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 47964 40908 48020 40964
rect 50316 40908 50372 40964
rect 50428 40908 50484 40964
rect 52444 40908 52500 40964
rect 54348 40908 54404 40964
rect 53340 40796 53396 40852
rect 43804 40740 43860 40796
rect 43908 40740 43964 40796
rect 44012 40740 44068 40796
rect 4172 40684 4228 40740
rect 5180 40684 5236 40740
rect 12460 40684 12516 40740
rect 16268 40684 16324 40740
rect 22316 40684 22372 40740
rect 33964 40684 34020 40740
rect 34300 40684 34356 40740
rect 35644 40684 35700 40740
rect 20972 40572 21028 40628
rect 49868 40572 49924 40628
rect 50540 40572 50596 40628
rect 5740 40460 5796 40516
rect 23212 40460 23268 40516
rect 29036 40460 29092 40516
rect 31388 40460 31444 40516
rect 32060 40460 32116 40516
rect 36092 40460 36148 40516
rect 37548 40460 37604 40516
rect 42588 40460 42644 40516
rect 48524 40460 48580 40516
rect 50204 40460 50260 40516
rect 53340 40460 53396 40516
rect 3052 40348 3108 40404
rect 10556 40348 10612 40404
rect 11900 40348 11956 40404
rect 12236 40348 12292 40404
rect 1148 40236 1204 40292
rect 12460 40236 12516 40292
rect 13020 40236 13076 40292
rect 16940 40348 16996 40404
rect 27020 40348 27076 40404
rect 48076 40348 48132 40404
rect 50988 40348 51044 40404
rect 16604 40236 16660 40292
rect 18172 40236 18228 40292
rect 19852 40236 19908 40292
rect 24892 40236 24948 40292
rect 34972 40236 35028 40292
rect 49308 40236 49364 40292
rect 10668 40124 10724 40180
rect 11452 40124 11508 40180
rect 26908 40124 26964 40180
rect 35980 40124 36036 40180
rect 41580 40124 41636 40180
rect 53452 40124 53508 40180
rect 4172 40012 4228 40068
rect 22764 40012 22820 40068
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 2268 39900 2324 39956
rect 7308 39900 7364 39956
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 34748 40012 34804 40068
rect 40012 40012 40068 40068
rect 45164 40012 45220 40068
rect 50428 40012 50484 40068
rect 51660 40012 51716 40068
rect 44464 39956 44520 40012
rect 44568 39956 44624 40012
rect 44672 39956 44728 40012
rect 22316 39900 22372 39956
rect 45388 39900 45444 39956
rect 47068 39900 47124 39956
rect 55692 39900 55748 39956
rect 8876 39788 8932 39844
rect 9212 39788 9268 39844
rect 9548 39788 9604 39844
rect 10668 39788 10724 39844
rect 13020 39788 13076 39844
rect 35196 39788 35252 39844
rect 41580 39788 41636 39844
rect 47180 39788 47236 39844
rect 52892 39788 52948 39844
rect 9884 39676 9940 39732
rect 11788 39676 11844 39732
rect 14588 39676 14644 39732
rect 16716 39676 16772 39732
rect 23212 39676 23268 39732
rect 26796 39676 26852 39732
rect 35420 39676 35476 39732
rect 42588 39676 42644 39732
rect 45164 39676 45220 39732
rect 1148 39564 1204 39620
rect 3052 39564 3108 39620
rect 5740 39564 5796 39620
rect 26124 39564 26180 39620
rect 26684 39564 26740 39620
rect 53340 39564 53396 39620
rect 56140 39564 56196 39620
rect 9548 39452 9604 39508
rect 12572 39452 12628 39508
rect 13020 39452 13076 39508
rect 13356 39452 13412 39508
rect 14140 39452 14196 39508
rect 26348 39452 26404 39508
rect 40124 39452 40180 39508
rect 45948 39452 46004 39508
rect 25228 39340 25284 39396
rect 28588 39340 28644 39396
rect 47068 39340 47124 39396
rect 48524 39340 48580 39396
rect 52444 39340 52500 39396
rect 53788 39340 53844 39396
rect 4172 39228 4228 39284
rect 10892 39228 10948 39284
rect 13132 39228 13188 39284
rect 15932 39228 15988 39284
rect 30716 39228 30772 39284
rect 34860 39228 34916 39284
rect 38892 39228 38948 39284
rect 39676 39228 39732 39284
rect 40124 39228 40180 39284
rect 50428 39228 50484 39284
rect 50652 39228 50708 39284
rect 54348 39228 54404 39284
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 43804 39172 43860 39228
rect 43908 39172 43964 39228
rect 44012 39172 44068 39228
rect 1036 39116 1092 39172
rect 4844 39116 4900 39172
rect 27020 39116 27076 39172
rect 33292 39116 33348 39172
rect 49308 39116 49364 39172
rect 49868 39116 49924 39172
rect 1820 39004 1876 39060
rect 2044 39004 2100 39060
rect 3500 39004 3556 39060
rect 6188 39004 6244 39060
rect 12460 39004 12516 39060
rect 25228 39004 25284 39060
rect 2492 38892 2548 38948
rect 25452 38892 25508 38948
rect 35532 38892 35588 38948
rect 36764 38892 36820 38948
rect 700 38780 756 38836
rect 4956 38780 5012 38836
rect 5292 38780 5348 38836
rect 7980 38780 8036 38836
rect 8428 38780 8484 38836
rect 10332 38780 10388 38836
rect 10780 38780 10836 38836
rect 13132 38780 13188 38836
rect 25116 38780 25172 38836
rect 40348 39004 40404 39060
rect 50092 39004 50148 39060
rect 50428 39004 50484 39060
rect 45948 38780 46004 38836
rect 50204 38780 50260 38836
rect 2940 38668 2996 38724
rect 5180 38668 5236 38724
rect 9548 38668 9604 38724
rect 14588 38668 14644 38724
rect 18172 38668 18228 38724
rect 26908 38668 26964 38724
rect 29260 38668 29316 38724
rect 33516 38668 33572 38724
rect 45164 38668 45220 38724
rect 47292 38668 47348 38724
rect 48076 38668 48132 38724
rect 50652 38668 50708 38724
rect 56700 38668 56756 38724
rect 7756 38556 7812 38612
rect 10892 38556 10948 38612
rect 15372 38556 15428 38612
rect 15596 38556 15652 38612
rect 25452 38556 25508 38612
rect 30828 38556 30884 38612
rect 31500 38556 31556 38612
rect 31948 38556 32004 38612
rect 14588 38444 14644 38500
rect 33516 38444 33572 38500
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 39676 38556 39732 38612
rect 54684 38556 54740 38612
rect 35196 38444 35252 38500
rect 41356 38444 41412 38500
rect 41916 38444 41972 38500
rect 44940 38444 44996 38500
rect 47852 38444 47908 38500
rect 44464 38388 44520 38444
rect 44568 38388 44624 38444
rect 44672 38388 44728 38444
rect 5068 38332 5124 38388
rect 11340 38332 11396 38388
rect 12684 38332 12740 38388
rect 15372 38332 15428 38388
rect 20972 38332 21028 38388
rect 24220 38332 24276 38388
rect 25116 38332 25172 38388
rect 29372 38332 29428 38388
rect 33740 38332 33796 38388
rect 35868 38332 35924 38388
rect 42140 38332 42196 38388
rect 54572 38332 54628 38388
rect 56364 38332 56420 38388
rect 56812 38332 56868 38388
rect 2268 38220 2324 38276
rect 7868 38220 7924 38276
rect 27692 38220 27748 38276
rect 39564 38220 39620 38276
rect 41804 38220 41860 38276
rect 49308 38220 49364 38276
rect 53900 38220 53956 38276
rect 56700 38220 56756 38276
rect 1596 38108 1652 38164
rect 9884 38108 9940 38164
rect 14252 38108 14308 38164
rect 18956 38108 19012 38164
rect 30828 38108 30884 38164
rect 41356 38108 41412 38164
rect 48412 38108 48468 38164
rect 5628 37996 5684 38052
rect 13132 37996 13188 38052
rect 14700 37996 14756 38052
rect 29036 37996 29092 38052
rect 31052 37996 31108 38052
rect 53340 37996 53396 38052
rect 2044 37884 2100 37940
rect 2940 37884 2996 37940
rect 5516 37884 5572 37940
rect 45836 37884 45892 37940
rect 14588 37772 14644 37828
rect 49308 37772 49364 37828
rect 55356 37772 55412 37828
rect 4284 37660 4340 37716
rect 5292 37660 5348 37716
rect 8428 37660 8484 37716
rect 12012 37660 12068 37716
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 12684 37660 12740 37716
rect 41804 37660 41860 37716
rect 42140 37660 42196 37716
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 43804 37604 43860 37660
rect 43908 37604 43964 37660
rect 44012 37604 44068 37660
rect 3500 37548 3556 37604
rect 4172 37548 4228 37604
rect 4956 37548 5012 37604
rect 7868 37548 7924 37604
rect 25116 37548 25172 37604
rect 26908 37548 26964 37604
rect 31836 37548 31892 37604
rect 54348 37548 54404 37604
rect 55356 37548 55412 37604
rect 33628 37436 33684 37492
rect 54124 37436 54180 37492
rect 55244 37436 55300 37492
rect 2156 37324 2212 37380
rect 36092 37324 36148 37380
rect 41244 37324 41300 37380
rect 42700 37324 42756 37380
rect 50092 37324 50148 37380
rect 53228 37324 53284 37380
rect 55132 37324 55188 37380
rect 1484 37212 1540 37268
rect 5068 37212 5124 37268
rect 17724 37212 17780 37268
rect 24892 37212 24948 37268
rect 27244 37212 27300 37268
rect 31948 37212 32004 37268
rect 39564 37212 39620 37268
rect 39788 37212 39844 37268
rect 41916 37212 41972 37268
rect 50540 37212 50596 37268
rect 4172 37100 4228 37156
rect 4844 37100 4900 37156
rect 5516 37100 5572 37156
rect 10332 37100 10388 37156
rect 23436 37100 23492 37156
rect 28252 37100 28308 37156
rect 29932 37100 29988 37156
rect 50652 37100 50708 37156
rect 51548 37100 51604 37156
rect 55132 37100 55188 37156
rect 7980 36988 8036 37044
rect 9436 36988 9492 37044
rect 15708 36988 15764 37044
rect 43596 36988 43652 37044
rect 49196 36988 49252 37044
rect 50540 36988 50596 37044
rect 50764 36988 50820 37044
rect 52892 36988 52948 37044
rect 53788 36988 53844 37044
rect 54460 36988 54516 37044
rect 4284 36876 4340 36932
rect 4844 36876 4900 36932
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 17388 36876 17444 36932
rect 26796 36876 26852 36932
rect 29932 36876 29988 36932
rect 40572 36876 40628 36932
rect 41356 36876 41412 36932
rect 41692 36876 41748 36932
rect 44156 36876 44212 36932
rect 51660 36876 51716 36932
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 44464 36820 44520 36876
rect 44568 36820 44624 36876
rect 44672 36820 44728 36876
rect 588 36764 644 36820
rect 5068 36764 5124 36820
rect 6300 36764 6356 36820
rect 13132 36764 13188 36820
rect 22204 36764 22260 36820
rect 24220 36764 24276 36820
rect 24892 36764 24948 36820
rect 34860 36764 34916 36820
rect 41244 36764 41300 36820
rect 46508 36764 46564 36820
rect 46732 36764 46788 36820
rect 47404 36764 47460 36820
rect 56252 36764 56308 36820
rect 57036 36764 57092 36820
rect 2044 36652 2100 36708
rect 6860 36652 6916 36708
rect 13580 36652 13636 36708
rect 37436 36652 37492 36708
rect 42476 36652 42532 36708
rect 9660 36540 9716 36596
rect 14924 36540 14980 36596
rect 38220 36540 38276 36596
rect 42700 36540 42756 36596
rect 51772 36540 51828 36596
rect 52780 36540 52836 36596
rect 56924 36540 56980 36596
rect 20860 36428 20916 36484
rect 37548 36428 37604 36484
rect 48748 36428 48804 36484
rect 53340 36428 53396 36484
rect 3052 36316 3108 36372
rect 5964 36316 6020 36372
rect 8652 36316 8708 36372
rect 27132 36316 27188 36372
rect 29932 36316 29988 36372
rect 30380 36316 30436 36372
rect 41132 36316 41188 36372
rect 49084 36316 49140 36372
rect 50764 36316 50820 36372
rect 54796 36316 54852 36372
rect 46508 36204 46564 36260
rect 46956 36204 47012 36260
rect 52108 36204 52164 36260
rect 5740 36092 5796 36148
rect 13580 36092 13636 36148
rect 15372 36092 15428 36148
rect 31612 36092 31668 36148
rect 35196 36092 35252 36148
rect 47516 36092 47572 36148
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 43804 36036 43860 36092
rect 43908 36036 43964 36092
rect 44012 36036 44068 36092
rect 22428 35980 22484 36036
rect 24220 35980 24276 36036
rect 25228 35980 25284 36036
rect 27356 35980 27412 36036
rect 40124 35980 40180 36036
rect 43596 35980 43652 36036
rect 46732 35980 46788 36036
rect 6076 35868 6132 35924
rect 7868 35868 7924 35924
rect 8876 35868 8932 35924
rect 3388 35756 3444 35812
rect 5740 35756 5796 35812
rect 8428 35756 8484 35812
rect 52444 35868 52500 35924
rect 9436 35756 9492 35812
rect 11788 35756 11844 35812
rect 54796 35756 54852 35812
rect 56476 35756 56532 35812
rect 17388 35644 17444 35700
rect 30044 35644 30100 35700
rect 33292 35644 33348 35700
rect 33628 35644 33684 35700
rect 40908 35644 40964 35700
rect 50428 35644 50484 35700
rect 55356 35644 55412 35700
rect 55580 35644 55636 35700
rect 8428 35532 8484 35588
rect 9436 35532 9492 35588
rect 14364 35532 14420 35588
rect 17612 35532 17668 35588
rect 19740 35532 19796 35588
rect 39676 35532 39732 35588
rect 43036 35532 43092 35588
rect 6300 35420 6356 35476
rect 6636 35420 6692 35476
rect 7980 35420 8036 35476
rect 22876 35420 22932 35476
rect 23660 35420 23716 35476
rect 24220 35420 24276 35476
rect 25116 35420 25172 35476
rect 29148 35420 29204 35476
rect 29820 35420 29876 35476
rect 34188 35420 34244 35476
rect 35980 35420 36036 35476
rect 37212 35420 37268 35476
rect 42252 35420 42308 35476
rect 46396 35420 46452 35476
rect 47292 35420 47348 35476
rect 5292 35308 5348 35364
rect 6972 35308 7028 35364
rect 11340 35308 11396 35364
rect 35420 35308 35476 35364
rect 37100 35308 37156 35364
rect 48524 35308 48580 35364
rect 51548 35308 51604 35364
rect 51884 35308 51940 35364
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 3052 35196 3108 35252
rect 5964 35196 6020 35252
rect 22764 35196 22820 35252
rect 6076 35084 6132 35140
rect 7196 35084 7252 35140
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 44464 35252 44520 35308
rect 44568 35252 44624 35308
rect 44672 35252 44728 35308
rect 28700 35196 28756 35252
rect 38444 35196 38500 35252
rect 39004 35196 39060 35252
rect 46172 35196 46228 35252
rect 47740 35196 47796 35252
rect 20636 35084 20692 35140
rect 25564 35084 25620 35140
rect 38668 35084 38724 35140
rect 51100 35196 51156 35252
rect 51772 35196 51828 35252
rect 53452 35196 53508 35252
rect 57260 35196 57316 35252
rect 50988 35084 51044 35140
rect 13580 34972 13636 35028
rect 17724 34972 17780 35028
rect 22428 34972 22484 35028
rect 31836 34972 31892 35028
rect 36988 34972 37044 35028
rect 37660 34972 37716 35028
rect 8428 34860 8484 34916
rect 25676 34860 25732 34916
rect 27692 34860 27748 34916
rect 30940 34860 30996 34916
rect 31500 34860 31556 34916
rect 39900 34860 39956 34916
rect 8764 34748 8820 34804
rect 9996 34748 10052 34804
rect 14812 34748 14868 34804
rect 21532 34748 21588 34804
rect 25452 34748 25508 34804
rect 39676 34748 39732 34804
rect 15596 34636 15652 34692
rect 27132 34636 27188 34692
rect 31948 34636 32004 34692
rect 40348 34636 40404 34692
rect 6412 34524 6468 34580
rect 7756 34524 7812 34580
rect 21420 34524 21476 34580
rect 39564 34524 39620 34580
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 8988 34412 9044 34468
rect 14252 34412 14308 34468
rect 16156 34412 16212 34468
rect 19740 34412 19796 34468
rect 23436 34412 23492 34468
rect 23660 34412 23716 34468
rect 24892 34412 24948 34468
rect 34300 34412 34356 34468
rect 46732 34748 46788 34804
rect 47292 34748 47348 34804
rect 50204 34748 50260 34804
rect 46956 34636 47012 34692
rect 52780 34748 52836 34804
rect 57148 34748 57204 34804
rect 50316 34524 50372 34580
rect 52108 34524 52164 34580
rect 52892 34524 52948 34580
rect 43804 34468 43860 34524
rect 43908 34468 43964 34524
rect 44012 34468 44068 34524
rect 50652 34412 50708 34468
rect 47180 34300 47236 34356
rect 5516 34188 5572 34244
rect 9996 34188 10052 34244
rect 12460 34188 12516 34244
rect 15372 34188 15428 34244
rect 18284 34188 18340 34244
rect 24892 34188 24948 34244
rect 46956 34188 47012 34244
rect 47292 34188 47348 34244
rect 50652 34188 50708 34244
rect 4284 34076 4340 34132
rect 13692 34076 13748 34132
rect 14252 34076 14308 34132
rect 14588 34076 14644 34132
rect 17052 34076 17108 34132
rect 22876 34076 22932 34132
rect 40348 34076 40404 34132
rect 46396 34076 46452 34132
rect 51884 34076 51940 34132
rect 54124 34076 54180 34132
rect 2492 33964 2548 34020
rect 5292 33964 5348 34020
rect 9100 33964 9156 34020
rect 17388 33964 17444 34020
rect 24892 33964 24948 34020
rect 32508 33964 32564 34020
rect 33852 33964 33908 34020
rect 48636 33964 48692 34020
rect 55020 33964 55076 34020
rect 1932 33852 1988 33908
rect 7196 33852 7252 33908
rect 11004 33852 11060 33908
rect 11788 33852 11844 33908
rect 13356 33852 13412 33908
rect 22876 33852 22932 33908
rect 27356 33852 27412 33908
rect 35308 33852 35364 33908
rect 38108 33852 38164 33908
rect 40460 33852 40516 33908
rect 47180 33852 47236 33908
rect 2268 33740 2324 33796
rect 4284 33740 4340 33796
rect 4844 33740 4900 33796
rect 14252 33740 14308 33796
rect 15372 33740 15428 33796
rect 15596 33740 15652 33796
rect 16828 33740 16884 33796
rect 18956 33740 19012 33796
rect 24892 33740 24948 33796
rect 25116 33740 25172 33796
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 2716 33516 2772 33572
rect 5628 33516 5684 33572
rect 2044 33404 2100 33460
rect 7980 33292 8036 33348
rect 11452 33292 11508 33348
rect 51100 33740 51156 33796
rect 44464 33684 44520 33740
rect 44568 33684 44624 33740
rect 44672 33684 44728 33740
rect 39676 33628 39732 33684
rect 47292 33628 47348 33684
rect 47964 33628 48020 33684
rect 52780 33628 52836 33684
rect 53340 33628 53396 33684
rect 47628 33572 47684 33628
rect 13916 33516 13972 33572
rect 30380 33516 30436 33572
rect 31164 33516 31220 33572
rect 45948 33516 46004 33572
rect 46732 33516 46788 33572
rect 48412 33516 48468 33572
rect 49308 33516 49364 33572
rect 51100 33516 51156 33572
rect 16492 33404 16548 33460
rect 21420 33404 21476 33460
rect 23212 33404 23268 33460
rect 30716 33404 30772 33460
rect 38444 33404 38500 33460
rect 40124 33404 40180 33460
rect 52892 33404 52948 33460
rect 54236 33404 54292 33460
rect 13468 33292 13524 33348
rect 17388 33292 17444 33348
rect 37100 33292 37156 33348
rect 38108 33292 38164 33348
rect 39676 33292 39732 33348
rect 43596 33292 43652 33348
rect 31836 33180 31892 33236
rect 49084 33292 49140 33348
rect 50092 33292 50148 33348
rect 53900 33292 53956 33348
rect 42700 33180 42756 33236
rect 49980 33180 50036 33236
rect 50204 33180 50260 33236
rect 50652 33180 50708 33236
rect 55916 33180 55972 33236
rect 5964 33068 6020 33124
rect 18508 33068 18564 33124
rect 22988 33068 23044 33124
rect 23660 33068 23716 33124
rect 25900 33068 25956 33124
rect 26572 33068 26628 33124
rect 27916 33068 27972 33124
rect 33068 33068 33124 33124
rect 33516 33068 33572 33124
rect 38892 33068 38948 33124
rect 53004 33068 53060 33124
rect 53340 33068 53396 33124
rect 7084 32956 7140 33012
rect 8428 32956 8484 33012
rect 41580 32956 41636 33012
rect 41916 32956 41972 33012
rect 42700 32956 42756 33012
rect 50652 32956 50708 33012
rect 51100 32956 51156 33012
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 4284 32844 4340 32900
rect 11340 32844 11396 32900
rect 20636 32844 20692 32900
rect 22876 32844 22932 32900
rect 3612 32732 3668 32788
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 43804 32900 43860 32956
rect 43908 32900 43964 32956
rect 44012 32900 44068 32956
rect 24892 32844 24948 32900
rect 52444 32844 52500 32900
rect 15708 32732 15764 32788
rect 16940 32732 16996 32788
rect 18956 32732 19012 32788
rect 21868 32732 21924 32788
rect 25900 32732 25956 32788
rect 32396 32732 32452 32788
rect 36204 32732 36260 32788
rect 44940 32732 44996 32788
rect 49420 32732 49476 32788
rect 54684 32732 54740 32788
rect 18284 32620 18340 32676
rect 35868 32620 35924 32676
rect 38220 32620 38276 32676
rect 49980 32620 50036 32676
rect 52892 32620 52948 32676
rect 7196 32508 7252 32564
rect 11452 32508 11508 32564
rect 12236 32508 12292 32564
rect 13916 32508 13972 32564
rect 16268 32508 16324 32564
rect 16828 32508 16884 32564
rect 24892 32508 24948 32564
rect 31724 32508 31780 32564
rect 32508 32508 32564 32564
rect 41468 32508 41524 32564
rect 45612 32508 45668 32564
rect 47292 32508 47348 32564
rect 51772 32508 51828 32564
rect 1260 32396 1316 32452
rect 1708 32396 1764 32452
rect 3612 32396 3668 32452
rect 7532 32396 7588 32452
rect 7980 32396 8036 32452
rect 17388 32396 17444 32452
rect 21308 32396 21364 32452
rect 25676 32396 25732 32452
rect 29372 32396 29428 32452
rect 35308 32396 35364 32452
rect 39228 32396 39284 32452
rect 43596 32396 43652 32452
rect 44940 32396 44996 32452
rect 7084 32284 7140 32340
rect 8428 32284 8484 32340
rect 13692 32284 13748 32340
rect 14140 32284 14196 32340
rect 14700 32284 14756 32340
rect 29708 32284 29764 32340
rect 37100 32284 37156 32340
rect 37436 32284 37492 32340
rect 37996 32284 38052 32340
rect 49196 32284 49252 32340
rect 2716 32172 2772 32228
rect 9548 32172 9604 32228
rect 23660 32172 23716 32228
rect 35308 32172 35364 32228
rect 39004 32172 39060 32228
rect 44156 32172 44212 32228
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 44464 32116 44520 32172
rect 44568 32116 44624 32172
rect 44672 32116 44728 32172
rect 47964 32172 48020 32228
rect 50988 32172 51044 32228
rect 6412 32060 6468 32116
rect 7980 32060 8036 32116
rect 17500 32060 17556 32116
rect 22876 32060 22932 32116
rect 39228 32060 39284 32116
rect 51884 32060 51940 32116
rect 52556 32060 52612 32116
rect 12236 31948 12292 32004
rect 21196 31948 21252 32004
rect 25900 31948 25956 32004
rect 39676 31948 39732 32004
rect 47628 31948 47684 32004
rect 51772 31948 51828 32004
rect 2156 31836 2212 31892
rect 3388 31836 3444 31892
rect 3612 31836 3668 31892
rect 16716 31836 16772 31892
rect 26236 31836 26292 31892
rect 26572 31836 26628 31892
rect 32956 31836 33012 31892
rect 36540 31836 36596 31892
rect 36876 31836 36932 31892
rect 39340 31836 39396 31892
rect 40908 31836 40964 31892
rect 47068 31836 47124 31892
rect 54124 31836 54180 31892
rect 4284 31724 4340 31780
rect 5180 31724 5236 31780
rect 9884 31724 9940 31780
rect 12908 31724 12964 31780
rect 17836 31724 17892 31780
rect 18284 31724 18340 31780
rect 23100 31724 23156 31780
rect 37660 31724 37716 31780
rect 38668 31724 38724 31780
rect 41692 31724 41748 31780
rect 45836 31724 45892 31780
rect 53452 31724 53508 31780
rect 10332 31612 10388 31668
rect 23548 31612 23604 31668
rect 27916 31612 27972 31668
rect 28700 31612 28756 31668
rect 32956 31612 33012 31668
rect 36428 31612 36484 31668
rect 36876 31612 36932 31668
rect 51100 31612 51156 31668
rect 52780 31612 52836 31668
rect 7980 31500 8036 31556
rect 50764 31500 50820 31556
rect 51548 31500 51604 31556
rect 51772 31500 51828 31556
rect 3612 31388 3668 31444
rect 6300 31388 6356 31444
rect 14252 31388 14308 31444
rect 24892 31388 24948 31444
rect 29484 31388 29540 31444
rect 32172 31388 32228 31444
rect 32844 31388 32900 31444
rect 49196 31388 49252 31444
rect 51884 31388 51940 31444
rect 54348 31388 54404 31444
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 6076 31276 6132 31332
rect 6972 31276 7028 31332
rect 9100 31276 9156 31332
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 43804 31332 43860 31388
rect 43908 31332 43964 31388
rect 44012 31332 44068 31388
rect 29820 31276 29876 31332
rect 44156 31276 44212 31332
rect 45500 31276 45556 31332
rect 52780 31276 52836 31332
rect 53228 31276 53284 31332
rect 25564 31164 25620 31220
rect 26124 31164 26180 31220
rect 27916 31164 27972 31220
rect 30716 31164 30772 31220
rect 33068 31164 33124 31220
rect 37100 31164 37156 31220
rect 47292 31164 47348 31220
rect 7308 31052 7364 31108
rect 20188 31052 20244 31108
rect 26460 31052 26516 31108
rect 44156 31052 44212 31108
rect 49084 31052 49140 31108
rect 50764 31052 50820 31108
rect 53676 31052 53732 31108
rect 5964 30940 6020 30996
rect 10444 30940 10500 30996
rect 14364 30940 14420 30996
rect 16940 30940 16996 30996
rect 17500 30940 17556 30996
rect 23100 30940 23156 30996
rect 23660 30940 23716 30996
rect 25452 30940 25508 30996
rect 30044 30940 30100 30996
rect 32732 30940 32788 30996
rect 47068 30940 47124 30996
rect 3612 30828 3668 30884
rect 10668 30828 10724 30884
rect 13132 30828 13188 30884
rect 24892 30828 24948 30884
rect 7308 30716 7364 30772
rect 8204 30716 8260 30772
rect 8876 30716 8932 30772
rect 9660 30716 9716 30772
rect 9884 30716 9940 30772
rect 14364 30716 14420 30772
rect 36204 30828 36260 30884
rect 36988 30828 37044 30884
rect 41580 30828 41636 30884
rect 52780 30828 52836 30884
rect 53116 30828 53172 30884
rect 34636 30716 34692 30772
rect 35084 30716 35140 30772
rect 36876 30716 36932 30772
rect 51548 30716 51604 30772
rect 23548 30604 23604 30660
rect 25452 30604 25508 30660
rect 44156 30604 44212 30660
rect 46732 30604 46788 30660
rect 48860 30604 48916 30660
rect 50764 30604 50820 30660
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 44464 30548 44520 30604
rect 44568 30548 44624 30604
rect 44672 30548 44728 30604
rect 2716 30492 2772 30548
rect 8988 30492 9044 30548
rect 9436 30492 9492 30548
rect 21308 30492 21364 30548
rect 47404 30492 47460 30548
rect 48300 30492 48356 30548
rect 6860 30380 6916 30436
rect 21532 30380 21588 30436
rect 22988 30380 23044 30436
rect 28364 30380 28420 30436
rect 32844 30380 32900 30436
rect 33068 30380 33124 30436
rect 36988 30380 37044 30436
rect 37548 30380 37604 30436
rect 42588 30380 42644 30436
rect 48524 30380 48580 30436
rect 50316 30380 50372 30436
rect 2492 30268 2548 30324
rect 7084 30268 7140 30324
rect 8764 30268 8820 30324
rect 12460 30268 12516 30324
rect 12684 30268 12740 30324
rect 24892 30268 24948 30324
rect 26124 30268 26180 30324
rect 31948 30268 32004 30324
rect 39676 30268 39732 30324
rect 47068 30268 47124 30324
rect 4284 30156 4340 30212
rect 4844 30156 4900 30212
rect 5628 30156 5684 30212
rect 10444 30156 10500 30212
rect 12796 30156 12852 30212
rect 13244 30156 13300 30212
rect 13804 30156 13860 30212
rect 14252 30156 14308 30212
rect 27468 30156 27524 30212
rect 27916 30156 27972 30212
rect 36092 30156 36148 30212
rect 37660 30156 37716 30212
rect 39564 30156 39620 30212
rect 40236 30156 40292 30212
rect 3500 30044 3556 30100
rect 5292 30044 5348 30100
rect 10892 30044 10948 30100
rect 18060 30044 18116 30100
rect 20188 30044 20244 30100
rect 6972 29932 7028 29988
rect 15820 29932 15876 29988
rect 20076 29932 20132 29988
rect 3052 29820 3108 29876
rect 5292 29820 5348 29876
rect 6076 29820 6132 29876
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 2604 29708 2660 29764
rect 5068 29708 5124 29764
rect 5516 29708 5572 29764
rect 8204 29708 8260 29764
rect 20076 29708 20132 29764
rect 9324 29596 9380 29652
rect 12236 29596 12292 29652
rect 2492 29484 2548 29540
rect 5964 29484 6020 29540
rect 15820 29484 15876 29540
rect 19068 29484 19124 29540
rect 1372 29260 1428 29316
rect 2604 29260 2660 29316
rect 5180 29260 5236 29316
rect 6524 29260 6580 29316
rect 17836 29372 17892 29428
rect 18508 29372 18564 29428
rect 18844 29372 18900 29428
rect 22876 30044 22932 30100
rect 26124 30044 26180 30100
rect 27356 30044 27412 30100
rect 29820 30044 29876 30100
rect 41020 30156 41076 30212
rect 45164 30044 45220 30100
rect 46172 30044 46228 30100
rect 47964 30044 48020 30100
rect 53900 30044 53956 30100
rect 27916 29932 27972 29988
rect 33628 29932 33684 29988
rect 34300 29932 34356 29988
rect 34972 29932 35028 29988
rect 44940 29932 44996 29988
rect 49756 29932 49812 29988
rect 50764 29932 50820 29988
rect 31052 29820 31108 29876
rect 34860 29820 34916 29876
rect 35420 29820 35476 29876
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 43804 29764 43860 29820
rect 43908 29764 43964 29820
rect 44012 29764 44068 29820
rect 33740 29708 33796 29764
rect 34412 29708 34468 29764
rect 34636 29708 34692 29764
rect 48524 29708 48580 29764
rect 48860 29708 48916 29764
rect 38892 29596 38948 29652
rect 48748 29596 48804 29652
rect 54908 29596 54964 29652
rect 36204 29484 36260 29540
rect 36988 29484 37044 29540
rect 45948 29484 46004 29540
rect 53452 29484 53508 29540
rect 28252 29372 28308 29428
rect 30828 29372 30884 29428
rect 22092 29260 22148 29316
rect 25228 29260 25284 29316
rect 32172 29260 32228 29316
rect 35196 29260 35252 29316
rect 2156 29148 2212 29204
rect 5964 29148 6020 29204
rect 8988 29148 9044 29204
rect 12572 29148 12628 29204
rect 34972 29148 35028 29204
rect 35420 29148 35476 29204
rect 2716 29036 2772 29092
rect 4956 29036 5012 29092
rect 12908 29036 12964 29092
rect 13692 29036 13748 29092
rect 28252 29036 28308 29092
rect 49980 29036 50036 29092
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 44464 28980 44520 29036
rect 44568 28980 44624 29036
rect 44672 28980 44728 29036
rect 3500 28924 3556 28980
rect 7196 28924 7252 28980
rect 23660 28924 23716 28980
rect 26460 28924 26516 28980
rect 32284 28924 32340 28980
rect 36204 28924 36260 28980
rect 40236 28924 40292 28980
rect 44156 28924 44212 28980
rect 49420 28924 49476 28980
rect 53788 28924 53844 28980
rect 3612 28812 3668 28868
rect 4956 28812 5012 28868
rect 23548 28812 23604 28868
rect 27916 28812 27972 28868
rect 29036 28812 29092 28868
rect 29820 28812 29876 28868
rect 35868 28812 35924 28868
rect 42252 28812 42308 28868
rect 44268 28812 44324 28868
rect 53004 28812 53060 28868
rect 55916 28812 55972 28868
rect 5964 28700 6020 28756
rect 12460 28700 12516 28756
rect 29708 28700 29764 28756
rect 37212 28700 37268 28756
rect 39004 28700 39060 28756
rect 7980 28588 8036 28644
rect 12572 28588 12628 28644
rect 22316 28588 22372 28644
rect 22540 28588 22596 28644
rect 35644 28588 35700 28644
rect 36764 28588 36820 28644
rect 39564 28588 39620 28644
rect 52892 28700 52948 28756
rect 47516 28588 47572 28644
rect 49756 28588 49812 28644
rect 8092 28476 8148 28532
rect 10556 28476 10612 28532
rect 10780 28476 10836 28532
rect 18956 28476 19012 28532
rect 21196 28476 21252 28532
rect 21532 28476 21588 28532
rect 33516 28476 33572 28532
rect 43372 28476 43428 28532
rect 44268 28476 44324 28532
rect 48636 28476 48692 28532
rect 51996 28476 52052 28532
rect 4844 28364 4900 28420
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 14364 28364 14420 28420
rect 27132 28364 27188 28420
rect 31612 28364 31668 28420
rect 34412 28364 34468 28420
rect 38444 28364 38500 28420
rect 38892 28364 38948 28420
rect 39788 28364 39844 28420
rect 52556 28364 52612 28420
rect 5852 28252 5908 28308
rect 31276 28252 31332 28308
rect 34188 28252 34244 28308
rect 35308 28252 35364 28308
rect 38108 28252 38164 28308
rect 42476 28252 42532 28308
rect 45164 28252 45220 28308
rect 47852 28252 47908 28308
rect 53340 28252 53396 28308
rect 4956 28140 5012 28196
rect 6300 28140 6356 28196
rect 7532 28140 7588 28196
rect 8540 28140 8596 28196
rect 11340 28140 11396 28196
rect 17052 28140 17108 28196
rect 5068 28028 5124 28084
rect 13356 28028 13412 28084
rect 20524 28028 20580 28084
rect 21756 28028 21812 28084
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 43804 28196 43860 28252
rect 43908 28196 43964 28252
rect 44012 28196 44068 28252
rect 32956 28140 33012 28196
rect 33628 28140 33684 28196
rect 39564 28140 39620 28196
rect 45388 28140 45444 28196
rect 31724 28028 31780 28084
rect 39228 28028 39284 28084
rect 40124 28028 40180 28084
rect 42140 28028 42196 28084
rect 51324 28028 51380 28084
rect 6300 27916 6356 27972
rect 17500 27916 17556 27972
rect 20412 27916 20468 27972
rect 21532 27916 21588 27972
rect 21868 27916 21924 27972
rect 42476 27916 42532 27972
rect 43148 27916 43204 27972
rect 45164 27916 45220 27972
rect 1260 27804 1316 27860
rect 9996 27804 10052 27860
rect 12796 27804 12852 27860
rect 14588 27804 14644 27860
rect 23100 27804 23156 27860
rect 29484 27804 29540 27860
rect 29932 27804 29988 27860
rect 39564 27804 39620 27860
rect 53340 27804 53396 27860
rect 6972 27692 7028 27748
rect 22204 27692 22260 27748
rect 41580 27692 41636 27748
rect 43372 27692 43428 27748
rect 43596 27692 43652 27748
rect 48860 27692 48916 27748
rect 55132 27692 55188 27748
rect 11228 27580 11284 27636
rect 14140 27580 14196 27636
rect 14364 27580 14420 27636
rect 17388 27580 17444 27636
rect 40572 27580 40628 27636
rect 1596 27468 1652 27524
rect 7084 27468 7140 27524
rect 20076 27468 20132 27524
rect 23100 27468 23156 27524
rect 41132 27468 41188 27524
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 4956 27356 5012 27412
rect 5292 27356 5348 27412
rect 7196 27356 7252 27412
rect 10892 27356 10948 27412
rect 22092 27356 22148 27412
rect 23212 27356 23268 27412
rect 24892 27356 24948 27412
rect 25228 27356 25284 27412
rect 28924 27356 28980 27412
rect 30268 27356 30324 27412
rect 44464 27412 44520 27468
rect 44568 27412 44624 27468
rect 44672 27412 44728 27468
rect 42140 27356 42196 27412
rect 50988 27356 51044 27412
rect 53228 27356 53284 27412
rect 54348 27356 54404 27412
rect 17052 27244 17108 27300
rect 41132 27244 41188 27300
rect 45164 27244 45220 27300
rect 12796 27132 12852 27188
rect 22316 27132 22372 27188
rect 27580 27132 27636 27188
rect 34748 27132 34804 27188
rect 38444 27132 38500 27188
rect 39564 27132 39620 27188
rect 43596 27132 43652 27188
rect 51772 27132 51828 27188
rect 4844 27020 4900 27076
rect 33516 27020 33572 27076
rect 45612 27020 45668 27076
rect 5180 26908 5236 26964
rect 5404 26908 5460 26964
rect 10444 26908 10500 26964
rect 14364 26908 14420 26964
rect 16156 26908 16212 26964
rect 22316 26908 22372 26964
rect 38892 26908 38948 26964
rect 40124 26908 40180 26964
rect 41356 26908 41412 26964
rect 12460 26796 12516 26852
rect 14924 26796 14980 26852
rect 30268 26796 30324 26852
rect 33852 26796 33908 26852
rect 34972 26796 35028 26852
rect 39004 26796 39060 26852
rect 39340 26796 39396 26852
rect 50652 26796 50708 26852
rect 5180 26684 5236 26740
rect 13132 26684 13188 26740
rect 17612 26684 17668 26740
rect 24892 26684 24948 26740
rect 32844 26684 32900 26740
rect 38108 26684 38164 26740
rect 38892 26684 38948 26740
rect 39228 26684 39284 26740
rect 45388 26684 45444 26740
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 43804 26628 43860 26684
rect 43908 26628 43964 26684
rect 44012 26628 44068 26684
rect 3500 26572 3556 26628
rect 8540 26572 8596 26628
rect 14140 26572 14196 26628
rect 15820 26572 15876 26628
rect 25900 26572 25956 26628
rect 39004 26572 39060 26628
rect 41468 26572 41524 26628
rect 44268 26572 44324 26628
rect 52556 26572 52612 26628
rect 4956 26460 5012 26516
rect 7196 26460 7252 26516
rect 16268 26460 16324 26516
rect 18956 26460 19012 26516
rect 3052 26348 3108 26404
rect 5628 26348 5684 26404
rect 6860 26348 6916 26404
rect 20076 26348 20132 26404
rect 25564 26348 25620 26404
rect 34188 26348 34244 26404
rect 39676 26348 39732 26404
rect 2716 26236 2772 26292
rect 21868 26236 21924 26292
rect 32956 26236 33012 26292
rect 44156 26348 44212 26404
rect 42700 26236 42756 26292
rect 12236 26124 12292 26180
rect 17948 26124 18004 26180
rect 26236 26124 26292 26180
rect 31164 26124 31220 26180
rect 35644 26124 35700 26180
rect 36988 26124 37044 26180
rect 39004 26124 39060 26180
rect 50092 26124 50148 26180
rect 2716 26012 2772 26068
rect 9548 26012 9604 26068
rect 38892 26012 38948 26068
rect 40460 26012 40516 26068
rect 48188 26012 48244 26068
rect 4956 25900 5012 25956
rect 5516 25900 5572 25956
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 15596 25900 15652 25956
rect 20748 25900 20804 25956
rect 23436 25900 23492 25956
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 44464 25844 44520 25900
rect 44568 25844 44624 25900
rect 44672 25844 44728 25900
rect 7532 25788 7588 25844
rect 13244 25788 13300 25844
rect 21868 25788 21924 25844
rect 22428 25788 22484 25844
rect 23100 25788 23156 25844
rect 32284 25788 32340 25844
rect 33740 25788 33796 25844
rect 34748 25788 34804 25844
rect 45388 25788 45444 25844
rect 50316 25788 50372 25844
rect 54796 25788 54852 25844
rect 1708 25676 1764 25732
rect 29372 25676 29428 25732
rect 33628 25676 33684 25732
rect 33852 25676 33908 25732
rect 43372 25676 43428 25732
rect 45500 25676 45556 25732
rect 49644 25676 49700 25732
rect 8876 25564 8932 25620
rect 9884 25564 9940 25620
rect 11564 25564 11620 25620
rect 13916 25564 13972 25620
rect 22876 25564 22932 25620
rect 23660 25564 23716 25620
rect 28252 25564 28308 25620
rect 28700 25564 28756 25620
rect 29036 25564 29092 25620
rect 33180 25564 33236 25620
rect 33516 25564 33572 25620
rect 34860 25564 34916 25620
rect 37212 25564 37268 25620
rect 53004 25564 53060 25620
rect 53900 25564 53956 25620
rect 4956 25452 5012 25508
rect 11788 25452 11844 25508
rect 12012 25452 12068 25508
rect 19404 25452 19460 25508
rect 19740 25452 19796 25508
rect 2716 25340 2772 25396
rect 7980 25340 8036 25396
rect 9548 25340 9604 25396
rect 9772 25340 9828 25396
rect 11004 25340 11060 25396
rect 1596 25228 1652 25284
rect 8540 25228 8596 25284
rect 41244 25452 41300 25508
rect 42588 25452 42644 25508
rect 51100 25452 51156 25508
rect 13692 25340 13748 25396
rect 35196 25340 35252 25396
rect 38108 25340 38164 25396
rect 50540 25340 50596 25396
rect 28812 25228 28868 25284
rect 30828 25228 30884 25284
rect 34748 25228 34804 25284
rect 39340 25228 39396 25284
rect 55804 25228 55860 25284
rect 38220 25116 38276 25172
rect 44156 25116 44212 25172
rect 44940 25116 44996 25172
rect 49420 25116 49476 25172
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 4956 25004 5012 25060
rect 5516 25004 5572 25060
rect 11676 25004 11732 25060
rect 28700 25004 28756 25060
rect 29260 25004 29316 25060
rect 19852 24892 19908 24948
rect 22092 24892 22148 24948
rect 22316 24892 22372 24948
rect 43804 25060 43860 25116
rect 43908 25060 43964 25116
rect 44012 25060 44068 25116
rect 32284 25004 32340 25060
rect 39676 25004 39732 25060
rect 41692 25004 41748 25060
rect 30492 24892 30548 24948
rect 44268 24892 44324 24948
rect 50316 24892 50372 24948
rect 1708 24780 1764 24836
rect 24892 24780 24948 24836
rect 26124 24780 26180 24836
rect 29260 24780 29316 24836
rect 33740 24780 33796 24836
rect 38220 24780 38276 24836
rect 41580 24780 41636 24836
rect 53228 24780 53284 24836
rect 2156 24668 2212 24724
rect 3388 24668 3444 24724
rect 4956 24668 5012 24724
rect 5516 24668 5572 24724
rect 5964 24668 6020 24724
rect 12908 24668 12964 24724
rect 19516 24668 19572 24724
rect 29036 24668 29092 24724
rect 31276 24668 31332 24724
rect 31500 24668 31556 24724
rect 32172 24668 32228 24724
rect 34748 24668 34804 24724
rect 50204 24668 50260 24724
rect 51660 24668 51716 24724
rect 5292 24556 5348 24612
rect 21532 24556 21588 24612
rect 21868 24556 21924 24612
rect 24892 24556 24948 24612
rect 32284 24556 32340 24612
rect 33068 24556 33124 24612
rect 34636 24556 34692 24612
rect 34972 24556 35028 24612
rect 41580 24556 41636 24612
rect 42252 24556 42308 24612
rect 51212 24556 51268 24612
rect 17836 24444 17892 24500
rect 26684 24444 26740 24500
rect 28140 24444 28196 24500
rect 38220 24444 38276 24500
rect 41132 24444 41188 24500
rect 45836 24444 45892 24500
rect 46956 24444 47012 24500
rect 49644 24444 49700 24500
rect 56476 24444 56532 24500
rect 1932 24332 1988 24388
rect 5068 24332 5124 24388
rect 5292 24332 5348 24388
rect 7980 24332 8036 24388
rect 8204 24332 8260 24388
rect 13132 24332 13188 24388
rect 14588 24332 14644 24388
rect 17612 24332 17668 24388
rect 21868 24332 21924 24388
rect 22092 24332 22148 24388
rect 27468 24332 27524 24388
rect 27916 24332 27972 24388
rect 28476 24332 28532 24388
rect 34636 24332 34692 24388
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 44464 24276 44520 24332
rect 44568 24276 44624 24332
rect 44672 24276 44728 24332
rect 49308 24332 49364 24388
rect 53452 24332 53508 24388
rect 57148 24332 57204 24388
rect 3388 24220 3444 24276
rect 4956 24220 5012 24276
rect 20076 24220 20132 24276
rect 22428 24220 22484 24276
rect 29820 24220 29876 24276
rect 39228 24220 39284 24276
rect 39676 24220 39732 24276
rect 40236 24220 40292 24276
rect 44156 24220 44212 24276
rect 56140 24220 56196 24276
rect 2604 24108 2660 24164
rect 5180 24108 5236 24164
rect 28476 24108 28532 24164
rect 33628 24108 33684 24164
rect 38220 24108 38276 24164
rect 39004 24108 39060 24164
rect 44268 24108 44324 24164
rect 9996 23996 10052 24052
rect 18508 23996 18564 24052
rect 30044 23996 30100 24052
rect 31164 23996 31220 24052
rect 53228 23996 53284 24052
rect 56812 23996 56868 24052
rect 3388 23884 3444 23940
rect 5628 23884 5684 23940
rect 6972 23884 7028 23940
rect 12684 23884 12740 23940
rect 17276 23884 17332 23940
rect 17612 23884 17668 23940
rect 22316 23884 22372 23940
rect 26348 23884 26404 23940
rect 29036 23884 29092 23940
rect 33852 23884 33908 23940
rect 41692 23884 41748 23940
rect 12236 23772 12292 23828
rect 18732 23772 18788 23828
rect 20636 23772 20692 23828
rect 20972 23772 21028 23828
rect 25228 23772 25284 23828
rect 36988 23772 37044 23828
rect 2380 23660 2436 23716
rect 9100 23660 9156 23716
rect 20412 23660 20468 23716
rect 21532 23660 21588 23716
rect 21868 23660 21924 23716
rect 27692 23660 27748 23716
rect 31612 23660 31668 23716
rect 34860 23660 34916 23716
rect 39564 23660 39620 23716
rect 56252 23660 56308 23716
rect 56812 23660 56868 23716
rect 17948 23548 18004 23604
rect 23100 23548 23156 23604
rect 25564 23548 25620 23604
rect 29260 23548 29316 23604
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 33852 23548 33908 23604
rect 41020 23548 41076 23604
rect 56364 23548 56420 23604
rect 43804 23492 43860 23548
rect 43908 23492 43964 23548
rect 44012 23492 44068 23548
rect 4284 23436 4340 23492
rect 9772 23436 9828 23492
rect 15372 23436 15428 23492
rect 17276 23436 17332 23492
rect 18732 23436 18788 23492
rect 23436 23436 23492 23492
rect 25452 23436 25508 23492
rect 32172 23436 32228 23492
rect 35420 23436 35476 23492
rect 36988 23436 37044 23492
rect 37212 23436 37268 23492
rect 41580 23436 41636 23492
rect 44156 23436 44212 23492
rect 19740 23324 19796 23380
rect 22428 23324 22484 23380
rect 23100 23324 23156 23380
rect 39676 23324 39732 23380
rect 54796 23324 54852 23380
rect 9996 23212 10052 23268
rect 11004 23212 11060 23268
rect 12012 23212 12068 23268
rect 20972 23212 21028 23268
rect 21868 23212 21924 23268
rect 4956 23100 5012 23156
rect 7196 23100 7252 23156
rect 8876 23100 8932 23156
rect 34188 23212 34244 23268
rect 38444 23212 38500 23268
rect 42476 23212 42532 23268
rect 44156 23212 44212 23268
rect 16940 23100 16996 23156
rect 18956 23100 19012 23156
rect 20300 23100 20356 23156
rect 20748 23100 20804 23156
rect 22876 23100 22932 23156
rect 39676 23100 39732 23156
rect 40572 23100 40628 23156
rect 41580 23100 41636 23156
rect 46508 23100 46564 23156
rect 47852 23100 47908 23156
rect 6524 22988 6580 23044
rect 11564 22988 11620 23044
rect 16492 22988 16548 23044
rect 30268 22988 30324 23044
rect 31164 22988 31220 23044
rect 33292 22988 33348 23044
rect 44156 22988 44212 23044
rect 45948 22988 46004 23044
rect 48748 22988 48804 23044
rect 52332 22988 52388 23044
rect 52668 22988 52724 23044
rect 8092 22876 8148 22932
rect 8540 22876 8596 22932
rect 19292 22876 19348 22932
rect 21532 22876 21588 22932
rect 22540 22876 22596 22932
rect 36540 22876 36596 22932
rect 36988 22876 37044 22932
rect 38892 22876 38948 22932
rect 49980 22876 50036 22932
rect 19740 22764 19796 22820
rect 22316 22764 22372 22820
rect 30828 22764 30884 22820
rect 34188 22764 34244 22820
rect 34860 22764 34916 22820
rect 35084 22764 35140 22820
rect 47628 22764 47684 22820
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 44464 22708 44520 22764
rect 44568 22708 44624 22764
rect 44672 22708 44728 22764
rect 5068 22652 5124 22708
rect 9772 22652 9828 22708
rect 14140 22652 14196 22708
rect 16156 22652 16212 22708
rect 16492 22652 16548 22708
rect 21308 22652 21364 22708
rect 39228 22652 39284 22708
rect 40572 22652 40628 22708
rect 44156 22652 44212 22708
rect 51100 22652 51156 22708
rect 2380 22540 2436 22596
rect 4956 22540 5012 22596
rect 7756 22540 7812 22596
rect 30268 22540 30324 22596
rect 32284 22540 32340 22596
rect 33292 22540 33348 22596
rect 36540 22540 36596 22596
rect 37212 22540 37268 22596
rect 40348 22540 40404 22596
rect 48524 22540 48580 22596
rect 2492 22428 2548 22484
rect 15260 22428 15316 22484
rect 19292 22428 19348 22484
rect 28140 22428 28196 22484
rect 30828 22428 30884 22484
rect 9660 22316 9716 22372
rect 10444 22316 10500 22372
rect 17276 22316 17332 22372
rect 22988 22316 23044 22372
rect 26124 22316 26180 22372
rect 30940 22316 30996 22372
rect 34188 22316 34244 22372
rect 34524 22316 34580 22372
rect 42588 22316 42644 22372
rect 48412 22316 48468 22372
rect 2380 22204 2436 22260
rect 5404 22092 5460 22148
rect 7644 22092 7700 22148
rect 9548 22092 9604 22148
rect 21532 22092 21588 22148
rect 22540 22092 22596 22148
rect 33292 22092 33348 22148
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 46732 21980 46788 22036
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 43804 21924 43860 21980
rect 43908 21924 43964 21980
rect 44012 21924 44068 21980
rect 12236 21868 12292 21924
rect 12460 21868 12516 21924
rect 27020 21868 27076 21924
rect 34300 21868 34356 21924
rect 34748 21868 34804 21924
rect 39564 21868 39620 21924
rect 40012 21868 40068 21924
rect 40460 21868 40516 21924
rect 40796 21868 40852 21924
rect 55692 21868 55748 21924
rect 8652 21756 8708 21812
rect 13916 21756 13972 21812
rect 14252 21756 14308 21812
rect 18732 21756 18788 21812
rect 21532 21756 21588 21812
rect 22428 21756 22484 21812
rect 40572 21756 40628 21812
rect 42140 21756 42196 21812
rect 42700 21756 42756 21812
rect 43372 21756 43428 21812
rect 45948 21756 46004 21812
rect 47068 21756 47124 21812
rect 51884 21756 51940 21812
rect 52668 21756 52724 21812
rect 54236 21756 54292 21812
rect 54684 21756 54740 21812
rect 13804 21644 13860 21700
rect 26460 21644 26516 21700
rect 35532 21644 35588 21700
rect 38892 21644 38948 21700
rect 40908 21644 40964 21700
rect 41580 21644 41636 21700
rect 3500 21532 3556 21588
rect 8876 21532 8932 21588
rect 23100 21532 23156 21588
rect 46508 21532 46564 21588
rect 49308 21532 49364 21588
rect 49868 21532 49924 21588
rect 7644 21420 7700 21476
rect 10332 21420 10388 21476
rect 14924 21420 14980 21476
rect 19628 21420 19684 21476
rect 20412 21420 20468 21476
rect 23548 21420 23604 21476
rect 26908 21420 26964 21476
rect 41580 21420 41636 21476
rect 47964 21420 48020 21476
rect 48636 21420 48692 21476
rect 18620 21308 18676 21364
rect 26348 21308 26404 21364
rect 48188 21308 48244 21364
rect 52332 21308 52388 21364
rect 10332 21196 10388 21252
rect 12796 21196 12852 21252
rect 16940 21196 16996 21252
rect 20076 21196 20132 21252
rect 20300 21196 20356 21252
rect 20748 21196 20804 21252
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 3052 21084 3108 21140
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 27468 21196 27524 21252
rect 55692 21196 55748 21252
rect 44464 21140 44520 21196
rect 44568 21140 44624 21196
rect 44672 21140 44728 21196
rect 18172 21084 18228 21140
rect 22988 21084 23044 21140
rect 26460 21084 26516 21140
rect 31276 21084 31332 21140
rect 39228 21084 39284 21140
rect 41580 21084 41636 21140
rect 41804 21084 41860 21140
rect 48636 21084 48692 21140
rect 51884 21084 51940 21140
rect 1596 20972 1652 21028
rect 3500 20972 3556 21028
rect 36764 20972 36820 21028
rect 50204 20972 50260 21028
rect 13804 20860 13860 20916
rect 17948 20860 18004 20916
rect 18620 20860 18676 20916
rect 23548 20860 23604 20916
rect 24220 20860 24276 20916
rect 25340 20860 25396 20916
rect 43596 20860 43652 20916
rect 3052 20748 3108 20804
rect 5516 20748 5572 20804
rect 6076 20748 6132 20804
rect 6300 20748 6356 20804
rect 34300 20748 34356 20804
rect 40796 20748 40852 20804
rect 42588 20748 42644 20804
rect 46620 20748 46676 20804
rect 51660 20748 51716 20804
rect 5404 20636 5460 20692
rect 23436 20636 23492 20692
rect 35980 20636 36036 20692
rect 45388 20636 45444 20692
rect 14252 20524 14308 20580
rect 18284 20524 18340 20580
rect 25116 20524 25172 20580
rect 26236 20524 26292 20580
rect 28700 20524 28756 20580
rect 29372 20524 29428 20580
rect 31724 20524 31780 20580
rect 49868 20524 49924 20580
rect 51548 20524 51604 20580
rect 6412 20412 6468 20468
rect 20972 20412 21028 20468
rect 22876 20412 22932 20468
rect 27132 20412 27188 20468
rect 28028 20412 28084 20468
rect 30044 20412 30100 20468
rect 32284 20412 32340 20468
rect 41020 20412 41076 20468
rect 41580 20412 41636 20468
rect 42028 20412 42084 20468
rect 43596 20412 43652 20468
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 43804 20356 43860 20412
rect 43908 20356 43964 20412
rect 44012 20356 44068 20412
rect 3052 20300 3108 20356
rect 23660 20300 23716 20356
rect 25228 20300 25284 20356
rect 28476 20300 28532 20356
rect 33068 20300 33124 20356
rect 37436 20300 37492 20356
rect 38892 20300 38948 20356
rect 47628 20300 47684 20356
rect 52444 20300 52500 20356
rect 8540 20188 8596 20244
rect 14140 20188 14196 20244
rect 18284 20188 18340 20244
rect 1596 20076 1652 20132
rect 7644 20076 7700 20132
rect 9884 20076 9940 20132
rect 11004 20076 11060 20132
rect 44268 20076 44324 20132
rect 48636 20076 48692 20132
rect 48860 20076 48916 20132
rect 54460 20076 54516 20132
rect 5740 19964 5796 20020
rect 10108 19964 10164 20020
rect 13580 19964 13636 20020
rect 23660 19964 23716 20020
rect 25004 19964 25060 20020
rect 26460 19964 26516 20020
rect 30044 19964 30100 20020
rect 30940 19964 30996 20020
rect 40572 19964 40628 20020
rect 3388 19852 3444 19908
rect 4844 19852 4900 19908
rect 10668 19852 10724 19908
rect 15596 19852 15652 19908
rect 23436 19852 23492 19908
rect 33852 19852 33908 19908
rect 36876 19852 36932 19908
rect 43148 19852 43204 19908
rect 47404 19852 47460 19908
rect 52668 19852 52724 19908
rect 5740 19740 5796 19796
rect 6300 19740 6356 19796
rect 13580 19740 13636 19796
rect 33516 19740 33572 19796
rect 45164 19740 45220 19796
rect 18284 19628 18340 19684
rect 27916 19628 27972 19684
rect 41132 19628 41188 19684
rect 42140 19628 42196 19684
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 44464 19572 44520 19628
rect 44568 19572 44624 19628
rect 44672 19572 44728 19628
rect 5068 19516 5124 19572
rect 6300 19516 6356 19572
rect 20076 19516 20132 19572
rect 25004 19516 25060 19572
rect 2380 19404 2436 19460
rect 35084 19404 35140 19460
rect 41020 19404 41076 19460
rect 45164 19404 45220 19460
rect 23660 19292 23716 19348
rect 31836 19292 31892 19348
rect 46620 19292 46676 19348
rect 49644 19292 49700 19348
rect 54572 19292 54628 19348
rect 7196 19180 7252 19236
rect 9324 19180 9380 19236
rect 11564 19180 11620 19236
rect 14252 19180 14308 19236
rect 19068 19180 19124 19236
rect 21420 19180 21476 19236
rect 28924 19180 28980 19236
rect 29932 19180 29988 19236
rect 34636 19180 34692 19236
rect 34972 19180 35028 19236
rect 38444 19180 38500 19236
rect 11004 19068 11060 19124
rect 47964 19180 48020 19236
rect 31836 19068 31892 19124
rect 33740 19068 33796 19124
rect 40572 19068 40628 19124
rect 44268 19068 44324 19124
rect 50316 19068 50372 19124
rect 6300 18956 6356 19012
rect 6524 18956 6580 19012
rect 13580 18956 13636 19012
rect 14252 18956 14308 19012
rect 34972 18956 35028 19012
rect 41132 18956 41188 19012
rect 51996 18956 52052 19012
rect 1484 18844 1540 18900
rect 30940 18844 30996 18900
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 7644 18732 7700 18788
rect 14252 18732 14308 18788
rect 18284 18732 18340 18788
rect 35084 18732 35140 18788
rect 41020 18732 41076 18788
rect 3164 18620 3220 18676
rect 6524 18620 6580 18676
rect 46396 18844 46452 18900
rect 51212 18844 51268 18900
rect 53452 18844 53508 18900
rect 43804 18788 43860 18844
rect 43908 18788 43964 18844
rect 44012 18788 44068 18844
rect 47964 18732 48020 18788
rect 53676 18620 53732 18676
rect 27356 18508 27412 18564
rect 34524 18508 34580 18564
rect 1260 18396 1316 18452
rect 2604 18396 2660 18452
rect 7420 18396 7476 18452
rect 7980 18396 8036 18452
rect 9100 18396 9156 18452
rect 12236 18396 12292 18452
rect 14812 18396 14868 18452
rect 15036 18396 15092 18452
rect 17164 18396 17220 18452
rect 18060 18396 18116 18452
rect 40460 18396 40516 18452
rect 40908 18396 40964 18452
rect 44268 18396 44324 18452
rect 52444 18396 52500 18452
rect 3164 18284 3220 18340
rect 4284 18284 4340 18340
rect 7084 18284 7140 18340
rect 9436 18284 9492 18340
rect 10668 18284 10724 18340
rect 12012 18284 12068 18340
rect 14252 18284 14308 18340
rect 17052 18284 17108 18340
rect 21308 18284 21364 18340
rect 28364 18284 28420 18340
rect 37100 18284 37156 18340
rect 51772 18284 51828 18340
rect 252 18060 308 18116
rect 5516 18060 5572 18116
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 12908 18172 12964 18228
rect 27244 18172 27300 18228
rect 31388 18172 31444 18228
rect 36988 18172 37044 18228
rect 37772 18172 37828 18228
rect 41020 18172 41076 18228
rect 7756 18060 7812 18116
rect 16044 18060 16100 18116
rect 25452 18060 25508 18116
rect 33740 18060 33796 18116
rect 34412 18060 34468 18116
rect 36204 18060 36260 18116
rect 42140 18060 42196 18116
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 1484 17948 1540 18004
rect 12460 17948 12516 18004
rect 14700 17948 14756 18004
rect 31500 17948 31556 18004
rect 44464 18004 44520 18060
rect 44568 18004 44624 18060
rect 44672 18004 44728 18060
rect 51548 18172 51604 18228
rect 38444 17948 38500 18004
rect 47852 17948 47908 18004
rect 53452 17948 53508 18004
rect 6188 17836 6244 17892
rect 8540 17836 8596 17892
rect 16156 17836 16212 17892
rect 31052 17836 31108 17892
rect 35308 17836 35364 17892
rect 37884 17836 37940 17892
rect 6300 17724 6356 17780
rect 12796 17724 12852 17780
rect 17164 17724 17220 17780
rect 38444 17724 38500 17780
rect 41692 17724 41748 17780
rect 47068 17724 47124 17780
rect 50204 17724 50260 17780
rect 51772 17724 51828 17780
rect 2156 17612 2212 17668
rect 3388 17612 3444 17668
rect 13916 17612 13972 17668
rect 22428 17612 22484 17668
rect 25116 17612 25172 17668
rect 30380 17612 30436 17668
rect 31052 17612 31108 17668
rect 32284 17612 32340 17668
rect 47628 17612 47684 17668
rect 1708 17500 1764 17556
rect 2716 17500 2772 17556
rect 27916 17500 27972 17556
rect 33404 17500 33460 17556
rect 33964 17500 34020 17556
rect 47292 17500 47348 17556
rect 49980 17500 50036 17556
rect 50204 17500 50260 17556
rect 3500 17388 3556 17444
rect 5068 17388 5124 17444
rect 5292 17388 5348 17444
rect 5740 17388 5796 17444
rect 6188 17388 6244 17444
rect 27468 17388 27524 17444
rect 31500 17388 31556 17444
rect 37772 17388 37828 17444
rect 38108 17388 38164 17444
rect 51436 17388 51492 17444
rect 4956 17276 5012 17332
rect 16604 17276 16660 17332
rect 45948 17276 46004 17332
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 43804 17220 43860 17276
rect 43908 17220 43964 17276
rect 44012 17220 44068 17276
rect 5964 17164 6020 17220
rect 24220 17164 24276 17220
rect 47404 17164 47460 17220
rect 1036 17052 1092 17108
rect 28140 17052 28196 17108
rect 34412 17052 34468 17108
rect 34860 17052 34916 17108
rect 37212 17052 37268 17108
rect 49084 17052 49140 17108
rect 52444 17052 52500 17108
rect 252 16940 308 16996
rect 1372 16940 1428 16996
rect 5180 16940 5236 16996
rect 3164 16828 3220 16884
rect 7756 16828 7812 16884
rect 21308 16940 21364 16996
rect 24220 16940 24276 16996
rect 25116 16940 25172 16996
rect 28812 16940 28868 16996
rect 34972 16940 35028 16996
rect 44940 16940 44996 16996
rect 45164 16940 45220 16996
rect 45836 16940 45892 16996
rect 51772 16940 51828 16996
rect 54908 16940 54964 16996
rect 25788 16828 25844 16884
rect 35420 16828 35476 16884
rect 588 16716 644 16772
rect 2940 16716 2996 16772
rect 4172 16716 4228 16772
rect 5180 16716 5236 16772
rect 6748 16716 6804 16772
rect 11116 16716 11172 16772
rect 13244 16716 13300 16772
rect 14140 16716 14196 16772
rect 16604 16716 16660 16772
rect 32844 16716 32900 16772
rect 33068 16716 33124 16772
rect 1036 16604 1092 16660
rect 7084 16604 7140 16660
rect 7644 16604 7700 16660
rect 11788 16604 11844 16660
rect 13916 16604 13972 16660
rect 35084 16604 35140 16660
rect 35420 16604 35476 16660
rect 4172 16492 4228 16548
rect 9772 16492 9828 16548
rect 11340 16492 11396 16548
rect 13692 16492 13748 16548
rect 20188 16492 20244 16548
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 40908 16828 40964 16884
rect 45948 16828 46004 16884
rect 42364 16716 42420 16772
rect 42588 16716 42644 16772
rect 43036 16716 43092 16772
rect 48524 16716 48580 16772
rect 49532 16716 49588 16772
rect 50204 16716 50260 16772
rect 53004 16604 53060 16660
rect 29708 16492 29764 16548
rect 31388 16492 31444 16548
rect 34860 16492 34916 16548
rect 35308 16492 35364 16548
rect 44268 16492 44324 16548
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 44464 16436 44520 16492
rect 44568 16436 44624 16492
rect 44672 16436 44728 16492
rect 2940 16380 2996 16436
rect 14476 16380 14532 16436
rect 20972 16380 21028 16436
rect 27020 16380 27076 16436
rect 30380 16380 30436 16436
rect 41468 16380 41524 16436
rect 44940 16380 44996 16436
rect 45612 16380 45668 16436
rect 55132 16380 55188 16436
rect 6524 16268 6580 16324
rect 22876 16268 22932 16324
rect 28700 16268 28756 16324
rect 29820 16268 29876 16324
rect 30604 16268 30660 16324
rect 32844 16268 32900 16324
rect 51996 16268 52052 16324
rect 52332 16268 52388 16324
rect 1932 16156 1988 16212
rect 7196 16156 7252 16212
rect 13132 16156 13188 16212
rect 18508 16156 18564 16212
rect 32396 16156 32452 16212
rect 33180 16156 33236 16212
rect 35084 16156 35140 16212
rect 41356 16156 41412 16212
rect 48972 16156 49028 16212
rect 3612 16044 3668 16100
rect 6972 16044 7028 16100
rect 20972 16044 21028 16100
rect 24220 16044 24276 16100
rect 31052 16044 31108 16100
rect 32284 16044 32340 16100
rect 35980 16044 36036 16100
rect 36876 16044 36932 16100
rect 45164 16044 45220 16100
rect 46508 16044 46564 16100
rect 49196 16044 49252 16100
rect 21308 15932 21364 15988
rect 23660 15932 23716 15988
rect 44940 15932 44996 15988
rect 47068 15932 47124 15988
rect 3164 15820 3220 15876
rect 3612 15820 3668 15876
rect 12012 15820 12068 15876
rect 15260 15820 15316 15876
rect 27804 15820 27860 15876
rect 31052 15820 31108 15876
rect 34412 15820 34468 15876
rect 37100 15708 37156 15764
rect 51548 15708 51604 15764
rect 51996 15708 52052 15764
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 43804 15652 43860 15708
rect 43908 15652 43964 15708
rect 44012 15652 44068 15708
rect 3052 15596 3108 15652
rect 7084 15596 7140 15652
rect 7644 15596 7700 15652
rect 9548 15596 9604 15652
rect 11452 15596 11508 15652
rect 19292 15596 19348 15652
rect 23660 15596 23716 15652
rect 29820 15596 29876 15652
rect 32284 15596 32340 15652
rect 34188 15596 34244 15652
rect 43372 15596 43428 15652
rect 44940 15596 44996 15652
rect 48188 15596 48244 15652
rect 4172 15484 4228 15540
rect 8652 15484 8708 15540
rect 21308 15484 21364 15540
rect 33180 15484 33236 15540
rect 38108 15484 38164 15540
rect 5180 15260 5236 15316
rect 38444 15372 38500 15428
rect 46508 15372 46564 15428
rect 46732 15372 46788 15428
rect 48860 15372 48916 15428
rect 53676 15372 53732 15428
rect 55356 15372 55412 15428
rect 19292 15260 19348 15316
rect 32844 15260 32900 15316
rect 33516 15260 33572 15316
rect 37548 15260 37604 15316
rect 41916 15260 41972 15316
rect 45164 15260 45220 15316
rect 45388 15260 45444 15316
rect 49420 15260 49476 15316
rect 4284 15148 4340 15204
rect 4956 15148 5012 15204
rect 9996 15148 10052 15204
rect 15372 15148 15428 15204
rect 24220 15148 24276 15204
rect 38444 15148 38500 15204
rect 5628 15036 5684 15092
rect 6972 15036 7028 15092
rect 41356 15036 41412 15092
rect 44268 15036 44324 15092
rect 44940 15036 44996 15092
rect 48860 15036 48916 15092
rect 2940 14924 2996 14980
rect 4956 14924 5012 14980
rect 6860 14924 6916 14980
rect 17164 14924 17220 14980
rect 22428 14924 22484 14980
rect 32844 14924 32900 14980
rect 37548 14924 37604 14980
rect 47628 14924 47684 14980
rect 53676 14924 53732 14980
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 5068 14812 5124 14868
rect 12124 14812 12180 14868
rect 14140 14812 14196 14868
rect 15372 14812 15428 14868
rect 30940 14812 30996 14868
rect 31164 14812 31220 14868
rect 41020 14812 41076 14868
rect 42700 14812 42756 14868
rect 44464 14868 44520 14924
rect 44568 14868 44624 14924
rect 44672 14868 44728 14924
rect 45948 14812 46004 14868
rect 49532 14812 49588 14868
rect 51436 14812 51492 14868
rect 5740 14700 5796 14756
rect 6748 14700 6804 14756
rect 8652 14700 8708 14756
rect 15036 14700 15092 14756
rect 29372 14700 29428 14756
rect 41356 14700 41412 14756
rect 41916 14700 41972 14756
rect 48188 14700 48244 14756
rect 48524 14700 48580 14756
rect 48972 14700 49028 14756
rect 51660 14700 51716 14756
rect 56588 14700 56644 14756
rect 12572 14588 12628 14644
rect 54124 14588 54180 14644
rect 5404 14476 5460 14532
rect 6300 14476 6356 14532
rect 6748 14476 6804 14532
rect 11004 14476 11060 14532
rect 12236 14476 12292 14532
rect 17836 14476 17892 14532
rect 18956 14476 19012 14532
rect 24220 14476 24276 14532
rect 31164 14476 31220 14532
rect 43148 14476 43204 14532
rect 44940 14476 44996 14532
rect 46172 14476 46228 14532
rect 17724 14364 17780 14420
rect 27244 14364 27300 14420
rect 30268 14364 30324 14420
rect 42028 14364 42084 14420
rect 43596 14364 43652 14420
rect 18956 14252 19012 14308
rect 39788 14252 39844 14308
rect 51436 14252 51492 14308
rect 21532 14140 21588 14196
rect 24220 14140 24276 14196
rect 43484 14140 43540 14196
rect 47964 14140 48020 14196
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 43804 14084 43860 14140
rect 43908 14084 43964 14140
rect 44012 14084 44068 14140
rect 52108 14140 52164 14196
rect 29260 14028 29316 14084
rect 43596 14028 43652 14084
rect 44940 14028 44996 14084
rect 46396 14028 46452 14084
rect 140 13916 196 13972
rect 3164 13916 3220 13972
rect 4956 13916 5012 13972
rect 9660 13916 9716 13972
rect 9996 13916 10052 13972
rect 10220 13916 10276 13972
rect 11228 13916 11284 13972
rect 13580 13916 13636 13972
rect 39788 13916 39844 13972
rect 32172 13804 32228 13860
rect 43372 13804 43428 13860
rect 48860 13804 48916 13860
rect 3500 13692 3556 13748
rect 6188 13692 6244 13748
rect 10444 13692 10500 13748
rect 11004 13692 11060 13748
rect 11228 13692 11284 13748
rect 14700 13692 14756 13748
rect 17612 13692 17668 13748
rect 20860 13692 20916 13748
rect 39564 13692 39620 13748
rect 47180 13692 47236 13748
rect 15372 13580 15428 13636
rect 17948 13580 18004 13636
rect 23660 13580 23716 13636
rect 29484 13580 29540 13636
rect 32060 13580 32116 13636
rect 33292 13580 33348 13636
rect 34412 13580 34468 13636
rect 37996 13580 38052 13636
rect 47852 13580 47908 13636
rect 48524 13580 48580 13636
rect 52556 13580 52612 13636
rect 1372 13468 1428 13524
rect 3052 13468 3108 13524
rect 5516 13468 5572 13524
rect 6188 13468 6244 13524
rect 6412 13468 6468 13524
rect 9548 13468 9604 13524
rect 16156 13468 16212 13524
rect 22428 13468 22484 13524
rect 32172 13468 32228 13524
rect 48412 13468 48468 13524
rect 49644 13468 49700 13524
rect 5628 13356 5684 13412
rect 7196 13356 7252 13412
rect 34860 13356 34916 13412
rect 43372 13356 43428 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 6412 13244 6468 13300
rect 11564 13244 11620 13300
rect 14924 13244 14980 13300
rect 16604 13244 16660 13300
rect 18060 13244 18116 13300
rect 23548 13244 23604 13300
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 50204 13356 50260 13412
rect 52108 13356 52164 13412
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 48300 13244 48356 13300
rect 48524 13244 48580 13300
rect 49196 13244 49252 13300
rect 3052 13132 3108 13188
rect 3276 13132 3332 13188
rect 7756 13132 7812 13188
rect 12908 13132 12964 13188
rect 23660 13132 23716 13188
rect 25676 13132 25732 13188
rect 47516 13132 47572 13188
rect 52668 13132 52724 13188
rect 54684 13132 54740 13188
rect 1708 13020 1764 13076
rect 4956 13020 5012 13076
rect 5516 13020 5572 13076
rect 5740 13020 5796 13076
rect 6300 13020 6356 13076
rect 9660 13020 9716 13076
rect 13804 13020 13860 13076
rect 14476 13020 14532 13076
rect 27020 13020 27076 13076
rect 28700 13020 28756 13076
rect 38892 13020 38948 13076
rect 45164 13020 45220 13076
rect 47404 13020 47460 13076
rect 5292 12908 5348 12964
rect 10556 12908 10612 12964
rect 12124 12908 12180 12964
rect 21532 12908 21588 12964
rect 29148 12908 29204 12964
rect 36876 12908 36932 12964
rect 41244 12908 41300 12964
rect 41804 12908 41860 12964
rect 43260 12908 43316 12964
rect 48972 12908 49028 12964
rect 52556 12908 52612 12964
rect 2156 12796 2212 12852
rect 6412 12796 6468 12852
rect 7196 12796 7252 12852
rect 16828 12796 16884 12852
rect 17276 12796 17332 12852
rect 2828 12684 2884 12740
rect 5292 12684 5348 12740
rect 8204 12684 8260 12740
rect 30044 12684 30100 12740
rect 33404 12684 33460 12740
rect 40572 12684 40628 12740
rect 43484 12684 43540 12740
rect 44940 12684 44996 12740
rect 49756 12684 49812 12740
rect 3612 12572 3668 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 11116 12572 11172 12628
rect 23660 12572 23716 12628
rect 26124 12572 26180 12628
rect 43148 12572 43204 12628
rect 46508 12572 46564 12628
rect 47292 12572 47348 12628
rect 49196 12572 49252 12628
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 364 12460 420 12516
rect 2940 12460 2996 12516
rect 3388 12460 3444 12516
rect 14924 12460 14980 12516
rect 28924 12460 28980 12516
rect 29148 12460 29204 12516
rect 40796 12460 40852 12516
rect 42140 12460 42196 12516
rect 45612 12460 45668 12516
rect 140 12348 196 12404
rect 6748 12348 6804 12404
rect 8204 12348 8260 12404
rect 11564 12348 11620 12404
rect 15372 12348 15428 12404
rect 17836 12348 17892 12404
rect 2380 12236 2436 12292
rect 4956 12236 5012 12292
rect 11788 12236 11844 12292
rect 17948 12236 18004 12292
rect 28700 12236 28756 12292
rect 28924 12236 28980 12292
rect 31836 12236 31892 12292
rect 34636 12236 34692 12292
rect 37100 12236 37156 12292
rect 140 12124 196 12180
rect 1932 12124 1988 12180
rect 3276 12124 3332 12180
rect 3500 12124 3556 12180
rect 7420 12124 7476 12180
rect 14140 12124 14196 12180
rect 33852 12124 33908 12180
rect 46620 12124 46676 12180
rect 49196 12124 49252 12180
rect 52668 12124 52724 12180
rect 6300 12012 6356 12068
rect 7868 12012 7924 12068
rect 11116 12012 11172 12068
rect 11340 12012 11396 12068
rect 17612 12012 17668 12068
rect 21980 12012 22036 12068
rect 28476 12012 28532 12068
rect 31612 12012 31668 12068
rect 31948 12012 32004 12068
rect 34524 12012 34580 12068
rect 47852 12012 47908 12068
rect 48524 12012 48580 12068
rect 6748 11900 6804 11956
rect 7308 11900 7364 11956
rect 9660 11900 9716 11956
rect 14476 11900 14532 11956
rect 23660 11900 23716 11956
rect 29148 11900 29204 11956
rect 1260 11788 1316 11844
rect 2044 11788 2100 11844
rect 9996 11788 10052 11844
rect 15372 11788 15428 11844
rect 15596 11788 15652 11844
rect 23548 11788 23604 11844
rect 26684 11788 26740 11844
rect 34188 11788 34244 11844
rect 35532 11788 35588 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 54460 12012 54516 12068
rect 45836 11900 45892 11956
rect 47292 11900 47348 11956
rect 50428 11900 50484 11956
rect 52668 11900 52724 11956
rect 53788 11900 53844 11956
rect 54124 11900 54180 11956
rect 42924 11788 42980 11844
rect 46732 11788 46788 11844
rect 49084 11788 49140 11844
rect 52108 11788 52164 11844
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 16604 11676 16660 11732
rect 24220 11676 24276 11732
rect 29036 11676 29092 11732
rect 38892 11676 38948 11732
rect 5628 11564 5684 11620
rect 9660 11564 9716 11620
rect 9996 11564 10052 11620
rect 13580 11564 13636 11620
rect 14700 11564 14756 11620
rect 15372 11564 15428 11620
rect 15596 11564 15652 11620
rect 16156 11564 16212 11620
rect 17836 11564 17892 11620
rect 25452 11564 25508 11620
rect 49532 11564 49588 11620
rect 50092 11564 50148 11620
rect 50764 11564 50820 11620
rect 56476 11564 56532 11620
rect 812 11452 868 11508
rect 4956 11452 5012 11508
rect 5404 11452 5460 11508
rect 6748 11452 6804 11508
rect 7084 11452 7140 11508
rect 16492 11452 16548 11508
rect 29932 11452 29988 11508
rect 42588 11452 42644 11508
rect 48972 11452 49028 11508
rect 52892 11452 52948 11508
rect 6972 11340 7028 11396
rect 9436 11340 9492 11396
rect 9996 11340 10052 11396
rect 33180 11340 33236 11396
rect 44156 11340 44212 11396
rect 48636 11340 48692 11396
rect 3276 11228 3332 11284
rect 5628 11228 5684 11284
rect 7868 11228 7924 11284
rect 8988 11228 9044 11284
rect 37100 11228 37156 11284
rect 39340 11228 39396 11284
rect 39564 11228 39620 11284
rect 44940 11228 44996 11284
rect 51772 11228 51828 11284
rect 18508 11116 18564 11172
rect 32172 11116 32228 11172
rect 40908 11116 40964 11172
rect 46956 11116 47012 11172
rect 812 11004 868 11060
rect 5964 11004 6020 11060
rect 9436 11004 9492 11060
rect 9660 11004 9716 11060
rect 10220 11004 10276 11060
rect 15036 11004 15092 11060
rect 22428 11004 22484 11060
rect 24220 11004 24276 11060
rect 26348 11004 26404 11060
rect 29932 11004 29988 11060
rect 40348 11004 40404 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 47628 11004 47684 11060
rect 48412 11004 48468 11060
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 53788 10892 53844 10948
rect 5180 10780 5236 10836
rect 5404 10780 5460 10836
rect 5964 10780 6020 10836
rect 6188 10780 6244 10836
rect 15260 10780 15316 10836
rect 16268 10780 16324 10836
rect 16604 10780 16660 10836
rect 12908 10668 12964 10724
rect 22428 10668 22484 10724
rect 29260 10668 29316 10724
rect 37212 10668 37268 10724
rect 48188 10668 48244 10724
rect 49420 10668 49476 10724
rect 49644 10668 49700 10724
rect 4844 10556 4900 10612
rect 15708 10556 15764 10612
rect 25004 10556 25060 10612
rect 25452 10556 25508 10612
rect 31276 10556 31332 10612
rect 49756 10556 49812 10612
rect 52780 10556 52836 10612
rect 5964 10444 6020 10500
rect 3500 10332 3556 10388
rect 4172 10332 4228 10388
rect 4844 10332 4900 10388
rect 9436 10332 9492 10388
rect 15596 10332 15652 10388
rect 15820 10332 15876 10388
rect 56252 10444 56308 10500
rect 44156 10332 44212 10388
rect 49532 10332 49588 10388
rect 49756 10332 49812 10388
rect 56140 10332 56196 10388
rect 6300 10220 6356 10276
rect 7196 10220 7252 10276
rect 7980 10220 8036 10276
rect 23660 10220 23716 10276
rect 26348 10220 26404 10276
rect 28476 10220 28532 10276
rect 32060 10220 32116 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 6860 10108 6916 10164
rect 8876 10108 8932 10164
rect 23212 10108 23268 10164
rect 9436 9996 9492 10052
rect 9660 9996 9716 10052
rect 10108 9996 10164 10052
rect 14700 9996 14756 10052
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 35980 10108 36036 10164
rect 42140 10108 42196 10164
rect 50764 10220 50820 10276
rect 53900 10108 53956 10164
rect 54796 10108 54852 10164
rect 22764 9996 22820 10052
rect 26124 9996 26180 10052
rect 33964 9996 34020 10052
rect 41468 9996 41524 10052
rect 45724 9996 45780 10052
rect 56364 9996 56420 10052
rect 19404 9884 19460 9940
rect 22092 9884 22148 9940
rect 28252 9884 28308 9940
rect 37212 9884 37268 9940
rect 49420 9884 49476 9940
rect 2492 9772 2548 9828
rect 4284 9772 4340 9828
rect 7868 9772 7924 9828
rect 21196 9772 21252 9828
rect 26684 9772 26740 9828
rect 31388 9772 31444 9828
rect 33404 9772 33460 9828
rect 34748 9772 34804 9828
rect 43036 9772 43092 9828
rect 44156 9772 44212 9828
rect 47068 9772 47124 9828
rect 9324 9660 9380 9716
rect 9660 9660 9716 9716
rect 47180 9660 47236 9716
rect 8652 9548 8708 9604
rect 13020 9548 13076 9604
rect 16268 9548 16324 9604
rect 17500 9548 17556 9604
rect 27692 9548 27748 9604
rect 31388 9548 31444 9604
rect 36428 9548 36484 9604
rect 45388 9548 45444 9604
rect 47964 9548 48020 9604
rect 2492 9436 2548 9492
rect 3388 9436 3444 9492
rect 4284 9436 4340 9492
rect 9324 9436 9380 9492
rect 13804 9436 13860 9492
rect 15260 9436 15316 9492
rect 15820 9436 15876 9492
rect 16492 9436 16548 9492
rect 17836 9436 17892 9492
rect 22876 9436 22932 9492
rect 32844 9436 32900 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 16940 9324 16996 9380
rect 20972 9324 21028 9380
rect 26572 9324 26628 9380
rect 26796 9324 26852 9380
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 35980 9324 36036 9380
rect 39004 9324 39060 9380
rect 2156 9212 2212 9268
rect 5068 9212 5124 9268
rect 5516 9212 5572 9268
rect 6188 9212 6244 9268
rect 9436 9212 9492 9268
rect 9884 9212 9940 9268
rect 14364 9212 14420 9268
rect 20748 9212 20804 9268
rect 21756 9212 21812 9268
rect 24220 9212 24276 9268
rect 26908 9212 26964 9268
rect 33404 9212 33460 9268
rect 36764 9212 36820 9268
rect 36988 9212 37044 9268
rect 43372 9212 43428 9268
rect 50764 9212 50820 9268
rect 52332 9212 52388 9268
rect 53564 9212 53620 9268
rect 1260 8988 1316 9044
rect 6748 8988 6804 9044
rect 7980 8988 8036 9044
rect 15596 8988 15652 9044
rect 27692 8988 27748 9044
rect 29036 8988 29092 9044
rect 32844 8988 32900 9044
rect 5180 8876 5236 8932
rect 53340 8876 53396 8932
rect 11564 8764 11620 8820
rect 43372 8764 43428 8820
rect 45164 8764 45220 8820
rect 5068 8652 5124 8708
rect 19852 8652 19908 8708
rect 23660 8652 23716 8708
rect 26684 8652 26740 8708
rect 38668 8652 38724 8708
rect 50540 8652 50596 8708
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 4956 8540 5012 8596
rect 13356 8540 13412 8596
rect 18060 8540 18116 8596
rect 18620 8540 18676 8596
rect 26572 8540 26628 8596
rect 32172 8540 32228 8596
rect 14476 8428 14532 8484
rect 21308 8428 21364 8484
rect 23100 8428 23156 8484
rect 3164 8204 3220 8260
rect 4284 8204 4340 8260
rect 13468 8316 13524 8372
rect 21196 8316 21252 8372
rect 23324 8316 23380 8372
rect 23548 8316 23604 8372
rect 9548 8204 9604 8260
rect 10332 8204 10388 8260
rect 16828 8204 16884 8260
rect 17388 8204 17444 8260
rect 18060 8204 18116 8260
rect 26684 8204 26740 8260
rect 29820 8204 29876 8260
rect 30380 8204 30436 8260
rect 31388 8204 31444 8260
rect 32508 8204 32564 8260
rect 33740 8204 33796 8260
rect 14700 8092 14756 8148
rect 19852 8092 19908 8148
rect 27356 8092 27412 8148
rect 34412 8092 34468 8148
rect 1484 7980 1540 8036
rect 3612 7980 3668 8036
rect 6300 7980 6356 8036
rect 6748 7980 6804 8036
rect 4172 7868 4228 7924
rect 7532 7868 7588 7924
rect 42476 8316 42532 8372
rect 36316 8204 36372 8260
rect 47964 8204 48020 8260
rect 50988 8204 51044 8260
rect 51884 7980 51940 8036
rect 32060 7868 32116 7924
rect 50764 7868 50820 7924
rect 2604 7756 2660 7812
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 6412 7756 6468 7812
rect 14364 7756 14420 7812
rect 15372 7756 15428 7812
rect 16044 7756 16100 7812
rect 16828 7756 16884 7812
rect 33740 7756 33796 7812
rect 40460 7756 40516 7812
rect 44156 7756 44212 7812
rect 48860 7756 48916 7812
rect 13468 7644 13524 7700
rect 30044 7644 30100 7700
rect 37100 7644 37156 7700
rect 40236 7644 40292 7700
rect 48300 7644 48356 7700
rect 6412 7532 6468 7588
rect 8204 7532 8260 7588
rect 15036 7532 15092 7588
rect 16492 7532 16548 7588
rect 22204 7532 22260 7588
rect 25116 7532 25172 7588
rect 26684 7532 26740 7588
rect 4956 7420 5012 7476
rect 6524 7420 6580 7476
rect 8540 7420 8596 7476
rect 9660 7420 9716 7476
rect 10108 7420 10164 7476
rect 13580 7420 13636 7476
rect 21196 7420 21252 7476
rect 25900 7420 25956 7476
rect 30940 7420 30996 7476
rect 31388 7420 31444 7476
rect 39900 7420 39956 7476
rect 40236 7420 40292 7476
rect 14924 7308 14980 7364
rect 42028 7308 42084 7364
rect 42364 7308 42420 7364
rect 51100 7308 51156 7364
rect 8652 7196 8708 7252
rect 14364 7196 14420 7252
rect 1484 7084 1540 7140
rect 9324 7084 9380 7140
rect 32732 7084 32788 7140
rect 38220 7084 38276 7140
rect 41580 7084 41636 7140
rect 44156 7084 44212 7140
rect 3388 6972 3444 7028
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 5404 6972 5460 7028
rect 31836 6860 31892 6916
rect 33068 6860 33124 6916
rect 33628 6860 33684 6916
rect 42924 6860 42980 6916
rect 45724 6860 45780 6916
rect 54124 6860 54180 6916
rect 1372 6748 1428 6804
rect 20076 6748 20132 6804
rect 22204 6748 22260 6804
rect 26908 6748 26964 6804
rect 38220 6748 38276 6804
rect 41356 6748 41412 6804
rect 9100 6636 9156 6692
rect 9996 6636 10052 6692
rect 15372 6636 15428 6692
rect 18284 6636 18340 6692
rect 24892 6636 24948 6692
rect 28364 6636 28420 6692
rect 33404 6636 33460 6692
rect 33628 6636 33684 6692
rect 41580 6636 41636 6692
rect 43036 6636 43092 6692
rect 2828 6524 2884 6580
rect 15596 6524 15652 6580
rect 16940 6524 16996 6580
rect 19740 6524 19796 6580
rect 33180 6524 33236 6580
rect 34636 6524 34692 6580
rect 39788 6524 39844 6580
rect 40124 6524 40180 6580
rect 40460 6524 40516 6580
rect 44268 6524 44324 6580
rect 45724 6636 45780 6692
rect 50652 6636 50708 6692
rect 5180 6412 5236 6468
rect 8652 6412 8708 6468
rect 18732 6412 18788 6468
rect 35084 6412 35140 6468
rect 36540 6412 36596 6468
rect 44940 6412 44996 6468
rect 52780 6412 52836 6468
rect 7084 6300 7140 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 18956 6300 19012 6356
rect 33068 6300 33124 6356
rect 34972 6300 35028 6356
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 4284 6188 4340 6244
rect 6860 6188 6916 6244
rect 9100 6188 9156 6244
rect 13356 6188 13412 6244
rect 16492 6188 16548 6244
rect 44156 6188 44212 6244
rect 45164 6188 45220 6244
rect 52780 6188 52836 6244
rect 55132 6188 55188 6244
rect 700 6076 756 6132
rect 17724 6076 17780 6132
rect 23100 6076 23156 6132
rect 11564 5964 11620 6020
rect 11788 5964 11844 6020
rect 12012 5964 12068 6020
rect 3052 5852 3108 5908
rect 6300 5852 6356 5908
rect 7980 5852 8036 5908
rect 9324 5852 9380 5908
rect 10108 5852 10164 5908
rect 15596 5852 15652 5908
rect 15820 5852 15876 5908
rect 21084 5852 21140 5908
rect 33180 5852 33236 5908
rect 33404 5852 33460 5908
rect 34860 5852 34916 5908
rect 35084 5852 35140 5908
rect 19068 5740 19124 5796
rect 27580 5740 27636 5796
rect 29372 5740 29428 5796
rect 39900 5740 39956 5796
rect 40348 5740 40404 5796
rect 44940 5740 44996 5796
rect 50876 5740 50932 5796
rect 3164 5516 3220 5572
rect 6748 5516 6804 5572
rect 11340 5516 11396 5572
rect 14700 5516 14756 5572
rect 14924 5516 14980 5572
rect 18396 5516 18452 5572
rect 27580 5516 27636 5572
rect 44268 5516 44324 5572
rect 47068 5516 47124 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 700 5404 756 5460
rect 3500 5404 3556 5460
rect 44828 5404 44884 5460
rect 19068 5292 19124 5348
rect 3500 5180 3556 5236
rect 14476 5180 14532 5236
rect 15260 5180 15316 5236
rect 34636 5292 34692 5348
rect 28252 5180 28308 5236
rect 41020 5180 41076 5236
rect 56140 5180 56196 5236
rect 2716 5068 2772 5124
rect 12684 5068 12740 5124
rect 15820 5068 15876 5124
rect 18956 5068 19012 5124
rect 20524 5068 20580 5124
rect 27020 5068 27076 5124
rect 43596 5068 43652 5124
rect 44268 5068 44324 5124
rect 44940 5068 44996 5124
rect 18732 4956 18788 5012
rect 42812 4956 42868 5012
rect 46844 4956 46900 5012
rect 49308 4956 49364 5012
rect 5628 4844 5684 4900
rect 9100 4844 9156 4900
rect 12124 4844 12180 4900
rect 13468 4844 13524 4900
rect 14588 4844 14644 4900
rect 44828 4844 44884 4900
rect 47964 4844 48020 4900
rect 50316 4844 50372 4900
rect 3612 4732 3668 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 5292 4732 5348 4788
rect 27020 4732 27076 4788
rect 31948 4732 32004 4788
rect 35980 4732 36036 4788
rect 43596 4732 43652 4788
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 18060 4620 18116 4676
rect 20300 4620 20356 4676
rect 31836 4620 31892 4676
rect 7420 4508 7476 4564
rect 7980 4508 8036 4564
rect 8652 4508 8708 4564
rect 9436 4508 9492 4564
rect 20972 4508 21028 4564
rect 45500 4508 45556 4564
rect 12124 4396 12180 4452
rect 14028 4396 14084 4452
rect 18508 4396 18564 4452
rect 21084 4396 21140 4452
rect 28252 4396 28308 4452
rect 28588 4396 28644 4452
rect 39900 4396 39956 4452
rect 10108 4284 10164 4340
rect 27916 4284 27972 4340
rect 32620 4284 32676 4340
rect 34076 4284 34132 4340
rect 35756 4284 35812 4340
rect 38556 4284 38612 4340
rect 1820 4172 1876 4228
rect 9436 4172 9492 4228
rect 3612 4060 3668 4116
rect 476 3948 532 4004
rect 4172 3948 4228 4004
rect 5964 3948 6020 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24220 4060 24276 4116
rect 35980 4060 36036 4116
rect 43596 4060 43652 4116
rect 52892 4060 52948 4116
rect 31500 3948 31556 4004
rect 44268 3948 44324 4004
rect 45388 3948 45444 4004
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 3500 3836 3556 3892
rect 9660 3836 9716 3892
rect 20188 3836 20244 3892
rect 44156 3836 44212 3892
rect 46060 3836 46116 3892
rect 812 3724 868 3780
rect 9772 3724 9828 3780
rect 11116 3724 11172 3780
rect 13020 3724 13076 3780
rect 26796 3724 26852 3780
rect 32172 3724 32228 3780
rect 53788 3724 53844 3780
rect 55356 3724 55412 3780
rect 3500 3612 3556 3668
rect 14140 3612 14196 3668
rect 19628 3612 19684 3668
rect 28140 3612 28196 3668
rect 36316 3612 36372 3668
rect 40908 3612 40964 3668
rect 45052 3612 45108 3668
rect 1484 3500 1540 3556
rect 26124 3500 26180 3556
rect 31164 3500 31220 3556
rect 3332 3388 3388 3444
rect 14028 3388 14084 3444
rect 21084 3388 21140 3444
rect 44268 3388 44324 3444
rect 2940 3276 2996 3332
rect 6860 3276 6916 3332
rect 14140 3276 14196 3332
rect 33964 3276 34020 3332
rect 43484 3276 43540 3332
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 13804 3052 13860 3108
rect 23324 3164 23380 3220
rect 25452 3164 25508 3220
rect 28364 3164 28420 3220
rect 34412 3164 34468 3220
rect 42364 3164 42420 3220
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 24220 3052 24276 3108
rect 26460 3052 26516 3108
rect 27132 3052 27188 3108
rect 35980 3052 36036 3108
rect 36204 3052 36260 3108
rect 52220 3052 52276 3108
rect 40908 2940 40964 2996
rect 7756 2828 7812 2884
rect 13020 2828 13076 2884
rect 26460 2828 26516 2884
rect 31724 2828 31780 2884
rect 48412 2828 48468 2884
rect 924 2716 980 2772
rect 8092 2716 8148 2772
rect 18508 2716 18564 2772
rect 24220 2716 24276 2772
rect 25340 2716 25396 2772
rect 33292 2716 33348 2772
rect 33740 2716 33796 2772
rect 34188 2716 34244 2772
rect 35196 2716 35252 2772
rect 36316 2716 36372 2772
rect 36652 2716 36708 2772
rect 37324 2716 37380 2772
rect 39116 2716 39172 2772
rect 39564 2716 39620 2772
rect 42140 2716 42196 2772
rect 6860 2604 6916 2660
rect 8652 2604 8708 2660
rect 19180 2604 19236 2660
rect 23436 2604 23492 2660
rect 29036 2604 29092 2660
rect 32060 2604 32116 2660
rect 38892 2604 38948 2660
rect 40348 2604 40404 2660
rect 48748 2604 48804 2660
rect 13020 2492 13076 2548
rect 18284 2492 18340 2548
rect 45276 2492 45332 2548
rect 48412 2492 48468 2548
rect 32060 2380 32116 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 2828 2268 2884 2324
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 24220 2268 24276 2324
rect 25340 2268 25396 2324
rect 6188 2156 6244 2212
rect 9660 2156 9716 2212
rect 19516 2156 19572 2212
rect 20076 2156 20132 2212
rect 22876 2156 22932 2212
rect 25228 2156 25284 2212
rect 26236 2156 26292 2212
rect 36092 2156 36148 2212
rect 38332 2156 38388 2212
rect 40684 2156 40740 2212
rect 43260 2156 43316 2212
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 46284 2156 46340 2212
rect 48076 2156 48132 2212
rect 18284 2044 18340 2100
rect 10220 1932 10276 1988
rect 12908 1932 12964 1988
rect 15036 1932 15092 1988
rect 25340 1932 25396 1988
rect 2940 1820 2996 1876
rect 48188 1820 48244 1876
rect 18620 1708 18676 1764
rect 19180 1708 19236 1764
rect 35980 1708 36036 1764
rect 40908 1708 40964 1764
rect 6076 1596 6132 1652
rect 8316 1596 8372 1652
rect 9212 1596 9268 1652
rect 11452 1596 11508 1652
rect 12348 1596 12404 1652
rect 13244 1596 13300 1652
rect 14252 1596 14308 1652
rect 14812 1596 14868 1652
rect 15932 1596 15988 1652
rect 16380 1596 16436 1652
rect 16828 1596 16884 1652
rect 17276 1596 17332 1652
rect 18172 1596 18228 1652
rect 20412 1596 20468 1652
rect 20748 1596 20804 1652
rect 23548 1596 23604 1652
rect 24220 1596 24276 1652
rect 38780 1596 38836 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 1148 1484 1204 1540
rect 1596 1484 1652 1540
rect 8204 1484 8260 1540
rect 8988 1484 9044 1540
rect 11676 1484 11732 1540
rect 15036 1484 15092 1540
rect 19964 1484 20020 1540
rect 588 1372 644 1428
rect 16380 1372 16436 1428
rect 16604 1372 16660 1428
rect 4284 1260 4340 1316
rect 8428 1260 8484 1316
rect 13020 1260 13076 1316
rect 30156 1260 30212 1316
rect 1036 1148 1092 1204
rect 2268 1148 2324 1204
rect 4172 1148 4228 1204
rect 4844 1148 4900 1204
rect 5852 1148 5908 1204
rect 7868 1148 7924 1204
rect 8764 1148 8820 1204
rect 9884 1148 9940 1204
rect 31052 1148 31108 1204
rect 37660 1148 37716 1204
rect 39452 1148 39508 1204
rect 11564 1036 11620 1092
rect 16380 1036 16436 1092
rect 52332 1036 52388 1092
rect 13916 924 13972 980
rect 21644 924 21700 980
rect 4284 812 4340 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 13692 812 13748 868
rect 23324 812 23380 868
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 6636 700 6692 756
rect 11900 700 11956 756
rect 15484 700 15540 756
rect 20636 700 20692 756
rect 22652 700 22708 756
rect 22876 700 22932 756
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 47740 700 47796 756
rect 2156 588 2212 644
rect 2492 588 2548 644
rect 54012 588 54068 644
rect 13020 364 13076 420
rect 15148 364 15204 420
rect 7756 252 7812 308
rect 12908 140 12964 196
rect 39788 140 39844 196
rect 10780 28 10836 84
rect 22876 28 22932 84
rect 32732 28 32788 84
rect 36764 28 36820 84
<< metal4 >>
rect 476 56756 532 56766
rect 252 56308 308 56318
rect 140 54964 196 54974
rect 140 13972 196 54908
rect 252 18116 308 56252
rect 252 16996 308 18060
rect 252 16930 308 16940
rect 364 46452 420 46462
rect 140 13906 196 13916
rect 364 12516 420 46396
rect 364 12450 420 12460
rect 140 12404 196 12414
rect 140 12180 196 12348
rect 140 12114 196 12124
rect 476 4004 532 56700
rect 3776 56476 4096 57456
rect 3388 56420 3444 56430
rect 2940 56084 2996 56094
rect 812 55860 868 55870
rect 700 50036 756 50046
rect 700 42980 756 49980
rect 812 48804 868 55804
rect 1708 55412 1764 55422
rect 1372 54516 1428 54526
rect 1260 54068 1316 54078
rect 812 48738 868 48748
rect 1148 50372 1204 50382
rect 924 46564 980 46574
rect 700 41698 756 42924
rect 588 41642 756 41698
rect 812 43988 868 43998
rect 588 36820 644 41642
rect 812 41636 868 43932
rect 700 41412 756 41422
rect 700 38836 756 41356
rect 700 38770 756 38780
rect 588 36754 644 36764
rect 476 3938 532 3948
rect 588 16772 644 16782
rect 588 1428 644 16716
rect 812 11508 868 41580
rect 812 11442 868 11452
rect 812 11060 868 11070
rect 700 6132 756 6142
rect 700 5460 756 6076
rect 700 5394 756 5404
rect 812 3780 868 11004
rect 812 3714 868 3724
rect 924 2772 980 46508
rect 1148 46004 1204 50316
rect 1148 45938 1204 45948
rect 1036 44996 1092 45006
rect 1036 39358 1092 44940
rect 1148 43204 1204 43214
rect 1148 40292 1204 43148
rect 1148 39620 1204 40236
rect 1148 39554 1204 39564
rect 1036 39302 1204 39358
rect 1036 39172 1092 39182
rect 1036 17108 1092 39116
rect 1036 17042 1092 17052
rect 924 2706 980 2716
rect 1036 16660 1092 16670
rect 588 1362 644 1372
rect 1036 1204 1092 16604
rect 1148 1540 1204 39302
rect 1260 32452 1316 54012
rect 1260 32386 1316 32396
rect 1372 29316 1428 54460
rect 1596 51604 1652 51614
rect 1596 49700 1652 51548
rect 1596 49140 1652 49644
rect 1596 49074 1652 49084
rect 1708 48898 1764 55356
rect 2492 54404 2548 54414
rect 1932 52948 1988 52958
rect 1932 51828 1988 52892
rect 1932 51762 1988 51772
rect 2380 51156 2436 51166
rect 1484 48842 1764 48898
rect 1820 50484 1876 50494
rect 1484 37268 1540 48842
rect 1708 48468 1764 48478
rect 1708 47796 1764 48412
rect 1596 43988 1652 43998
rect 1596 43428 1652 43932
rect 1596 43362 1652 43372
rect 1596 41860 1652 41870
rect 1596 38164 1652 41804
rect 1708 41188 1764 47740
rect 1820 44578 1876 50428
rect 2044 49924 2100 49934
rect 1932 49140 1988 49150
rect 1932 47012 1988 49084
rect 2044 48468 2100 49868
rect 2268 49812 2324 49822
rect 2268 49028 2324 49756
rect 2268 48962 2324 48972
rect 2380 49476 2436 51100
rect 2044 48402 2100 48412
rect 2380 48244 2436 49420
rect 2380 48178 2436 48188
rect 1932 46946 1988 46956
rect 2492 46378 2548 54348
rect 2828 52948 2884 52958
rect 2268 46322 2548 46378
rect 2604 52836 2660 52846
rect 2604 52164 2660 52780
rect 2044 46004 2100 46014
rect 2044 44772 2100 45948
rect 2044 44706 2100 44716
rect 1820 44522 1988 44578
rect 1708 41122 1764 41132
rect 1932 44436 1988 44522
rect 1596 38098 1652 38108
rect 1820 39060 1876 39070
rect 1484 37202 1540 37212
rect 1372 29250 1428 29260
rect 1708 32452 1764 32462
rect 1260 27860 1316 27870
rect 1260 18452 1316 27804
rect 1596 27524 1652 27534
rect 1596 25284 1652 27468
rect 1596 21028 1652 25228
rect 1708 25732 1764 32396
rect 1708 24836 1764 25676
rect 1708 24770 1764 24780
rect 1596 20962 1652 20972
rect 1596 20132 1652 20142
rect 1260 18386 1316 18396
rect 1484 18900 1540 18910
rect 1484 18004 1540 18844
rect 1372 16996 1428 17006
rect 1372 13524 1428 16940
rect 1260 11844 1316 11854
rect 1260 9044 1316 11788
rect 1260 8978 1316 8988
rect 1372 6804 1428 13468
rect 1484 8036 1540 17948
rect 1484 7970 1540 7980
rect 1372 6738 1428 6748
rect 1484 7140 1540 7150
rect 1484 3556 1540 7084
rect 1484 3490 1540 3500
rect 1148 1474 1204 1484
rect 1596 1540 1652 20076
rect 1708 17556 1764 17566
rect 1708 13076 1764 17500
rect 1708 13010 1764 13020
rect 1820 4228 1876 39004
rect 1932 33908 1988 44380
rect 2268 42532 2324 46322
rect 2604 44578 2660 52108
rect 2716 50932 2772 50942
rect 2716 49364 2772 50876
rect 2716 49298 2772 49308
rect 2268 42466 2324 42476
rect 2380 44522 2660 44578
rect 2716 49140 2772 49150
rect 2380 41524 2436 44522
rect 2604 44436 2660 44446
rect 2044 41188 2100 41198
rect 2044 39060 2100 41132
rect 2044 38994 2100 39004
rect 2268 39956 2324 39966
rect 2268 38276 2324 39900
rect 2268 38210 2324 38220
rect 2044 37940 2100 37950
rect 2044 36708 2100 37884
rect 2044 36642 2100 36652
rect 2156 37380 2212 37390
rect 1932 33842 1988 33852
rect 2044 33460 2100 33470
rect 1932 24388 1988 24398
rect 1932 16212 1988 24332
rect 1932 12180 1988 16156
rect 1932 12114 1988 12124
rect 2044 11844 2100 33404
rect 2156 31892 2212 37324
rect 2156 31826 2212 31836
rect 2268 33796 2324 33806
rect 2156 29204 2212 29214
rect 2156 24724 2212 29148
rect 2156 24658 2212 24668
rect 2156 17668 2212 17678
rect 2156 12852 2212 17612
rect 2156 12786 2212 12796
rect 2044 11778 2100 11788
rect 1820 4162 1876 4172
rect 2156 9268 2212 9278
rect 1596 1474 1652 1484
rect 1036 1138 1092 1148
rect 2156 644 2212 9212
rect 2268 1204 2324 33740
rect 2380 23716 2436 41468
rect 2492 41748 2548 41758
rect 2492 38948 2548 41692
rect 2492 38882 2548 38892
rect 2492 34020 2548 34030
rect 2492 30324 2548 33964
rect 2492 30258 2548 30268
rect 2604 29764 2660 44380
rect 2716 33572 2772 49084
rect 2716 33506 2772 33516
rect 2716 32228 2772 32238
rect 2716 30548 2772 32172
rect 2716 30482 2772 30492
rect 2604 29698 2660 29708
rect 2380 23650 2436 23660
rect 2492 29540 2548 29550
rect 2380 22596 2436 22606
rect 2380 22260 2436 22540
rect 2380 19460 2436 22204
rect 2380 12292 2436 19404
rect 2380 12226 2436 12236
rect 2492 22484 2548 29484
rect 2604 29316 2660 29326
rect 2604 24164 2660 29260
rect 2716 29092 2772 29102
rect 2716 26292 2772 29036
rect 2716 26226 2772 26236
rect 2716 26068 2772 26078
rect 2716 25396 2772 26012
rect 2716 25330 2772 25340
rect 2604 24098 2660 24108
rect 2492 9828 2548 22428
rect 2492 9762 2548 9772
rect 2604 18452 2660 18462
rect 2268 1138 2324 1148
rect 2492 9492 2548 9502
rect 2156 578 2212 588
rect 2492 644 2548 9436
rect 2604 7812 2660 18396
rect 2604 7746 2660 7756
rect 2716 17556 2772 17566
rect 2716 5124 2772 17500
rect 2828 12740 2884 52892
rect 2940 42196 2996 56028
rect 3052 55300 3108 55310
rect 3052 44578 3108 55244
rect 3276 55300 3332 55310
rect 3164 53060 3220 53070
rect 3164 48804 3220 53004
rect 3276 52836 3332 55244
rect 3388 54852 3444 56364
rect 3388 54786 3444 54796
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 3776 54908 4096 56420
rect 4436 55692 4756 57456
rect 6188 57204 6244 57214
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 5068 56308 5124 56318
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 3612 54068 3668 54078
rect 3276 52770 3332 52780
rect 3388 53844 3444 53854
rect 3388 53508 3444 53788
rect 3388 51940 3444 53452
rect 3500 53396 3556 53406
rect 3500 52388 3556 53340
rect 3500 52322 3556 52332
rect 3388 51492 3444 51884
rect 3388 51426 3444 51436
rect 3612 51380 3668 54012
rect 3612 51314 3668 51324
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 4284 55076 4340 55086
rect 3776 51772 4096 53284
rect 4172 53284 4228 53294
rect 4172 52948 4228 53228
rect 4172 52882 4228 52892
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3388 51156 3444 51166
rect 3164 48738 3220 48748
rect 3276 50484 3332 50494
rect 3164 48468 3220 48478
rect 3164 44758 3220 48412
rect 3276 45668 3332 50428
rect 3388 49252 3444 51100
rect 3388 49186 3444 49196
rect 3500 50932 3556 50942
rect 3500 49028 3556 50876
rect 3776 50204 4096 51716
rect 4172 52052 4228 52062
rect 4172 51716 4228 51996
rect 4172 51650 4228 51660
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3500 48962 3556 48972
rect 3612 49364 3668 49374
rect 3612 47796 3668 49308
rect 3612 47730 3668 47740
rect 3776 48636 4096 50148
rect 4284 49078 4340 55020
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3388 47348 3444 47358
rect 3388 46788 3444 47292
rect 3776 47068 4096 48580
rect 4172 49022 4340 49078
rect 4436 54124 4756 55636
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 4956 55636 5012 55646
rect 4956 49978 5012 55580
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4172 47684 4228 49022
rect 4172 47618 4228 47628
rect 4284 48916 4340 48926
rect 3388 46722 3444 46732
rect 3612 47012 3668 47022
rect 3612 46788 3668 46956
rect 3612 46722 3668 46732
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3388 46452 3444 46462
rect 3388 45892 3444 46396
rect 3388 45826 3444 45836
rect 3500 46004 3556 46014
rect 3276 45108 3332 45612
rect 3276 45042 3332 45052
rect 3388 45108 3444 45118
rect 3164 44702 3332 44758
rect 3052 44522 3220 44578
rect 2940 42130 2996 42140
rect 3052 41524 3108 41534
rect 3052 40404 3108 41468
rect 3052 40338 3108 40348
rect 3052 39620 3108 39630
rect 2940 38724 2996 38734
rect 2940 37940 2996 38668
rect 2940 16772 2996 37884
rect 3052 36372 3108 39564
rect 3052 36306 3108 36316
rect 3052 35252 3108 35262
rect 3052 29876 3108 35196
rect 3052 29810 3108 29820
rect 3052 26404 3108 26414
rect 3052 21140 3108 26348
rect 3052 21074 3108 21084
rect 3052 20804 3108 20814
rect 3052 20356 3108 20748
rect 3052 20290 3108 20300
rect 3164 18676 3220 44522
rect 3276 44324 3332 44702
rect 3276 44258 3332 44268
rect 3164 18340 3220 18620
rect 3164 18274 3220 18284
rect 3276 43540 3332 43550
rect 2940 16706 2996 16716
rect 3164 16884 3220 16894
rect 2940 16436 2996 16446
rect 2940 14980 2996 16380
rect 3164 15876 3220 16828
rect 3164 15810 3220 15820
rect 2940 14914 2996 14924
rect 3052 15652 3108 15662
rect 3052 13524 3108 15596
rect 3052 13458 3108 13468
rect 3164 13972 3220 13982
rect 2828 12674 2884 12684
rect 3052 13188 3108 13198
rect 2940 12516 2996 12526
rect 2716 5058 2772 5068
rect 2828 6580 2884 6590
rect 2828 2324 2884 6524
rect 2828 2258 2884 2268
rect 2940 3332 2996 12460
rect 3052 5908 3108 13132
rect 3164 8260 3220 13916
rect 3276 13188 3332 43484
rect 3388 43092 3444 45052
rect 3388 43026 3444 43036
rect 3500 42756 3556 45948
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3612 45220 3668 45230
rect 3612 43540 3668 45164
rect 3612 43474 3668 43484
rect 3776 43932 4096 45444
rect 4284 45332 4340 48860
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3500 42690 3556 42700
rect 3612 42868 3668 42878
rect 3388 42532 3444 42542
rect 3388 40852 3444 42476
rect 3388 35812 3444 40796
rect 3500 42420 3556 42430
rect 3500 39060 3556 42364
rect 3612 41524 3668 42812
rect 3612 41458 3668 41468
rect 3776 42364 4096 43876
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3500 38994 3556 39004
rect 3612 40964 3668 40974
rect 3388 35746 3444 35756
rect 3500 37604 3556 37614
rect 3388 31892 3444 31902
rect 3388 26398 3444 31836
rect 3500 30100 3556 37548
rect 3612 32788 3668 40908
rect 3612 32722 3668 32732
rect 3776 40796 4096 42308
rect 4172 45220 4228 45230
rect 4172 41860 4228 45164
rect 4284 44436 4340 45276
rect 4284 44370 4340 44380
rect 4436 47852 4756 49364
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 4844 49922 5012 49978
rect 4844 45220 4900 49922
rect 4844 45154 4900 45164
rect 4956 49700 5012 49710
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4284 44212 4340 44222
rect 4284 43204 4340 44156
rect 4284 43138 4340 43148
rect 4436 43148 4756 44660
rect 4844 44884 4900 44894
rect 4844 43540 4900 44828
rect 4844 43474 4900 43484
rect 4172 41794 4228 41804
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 4436 41580 4756 43092
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 4172 41524 4228 41534
rect 4172 40740 4228 41468
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 4172 40674 4228 40684
rect 4284 41076 4340 41086
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 4172 40068 4228 40078
rect 4172 39284 4228 40012
rect 4172 39218 4228 39228
rect 3776 37660 4096 39172
rect 4284 38458 4340 41020
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 4172 38402 4340 38458
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4436 38444 4756 39956
rect 4844 42420 4900 42430
rect 4844 39172 4900 42364
rect 4844 39106 4900 39116
rect 4956 38836 5012 49644
rect 5068 49140 5124 56252
rect 5964 54404 6020 54414
rect 5852 52724 5908 52734
rect 5404 50820 5460 50830
rect 5068 49074 5124 49084
rect 5292 50708 5348 50718
rect 5180 48916 5236 48926
rect 5068 48468 5124 48478
rect 5068 47098 5124 48412
rect 5180 47348 5236 48860
rect 5180 47282 5236 47292
rect 5068 47042 5236 47098
rect 5180 46340 5236 47042
rect 5068 45556 5124 45566
rect 5068 44212 5124 45500
rect 5180 44660 5236 46284
rect 5180 44594 5236 44604
rect 5068 44146 5124 44156
rect 4956 38770 5012 38780
rect 5068 41860 5124 41870
rect 4172 37604 4228 38402
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4172 37538 4228 37548
rect 4284 37716 4340 37726
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3776 34524 4096 36036
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 3776 32956 4096 34468
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3612 32452 3668 32462
rect 3612 31892 3668 32396
rect 3612 31826 3668 31836
rect 3612 31444 3668 31454
rect 3612 30884 3668 31388
rect 3612 30818 3668 30828
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3500 30034 3556 30044
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 3500 28980 3556 28990
rect 3500 26628 3556 28924
rect 3500 26562 3556 26572
rect 3612 28868 3668 28878
rect 3388 26342 3556 26398
rect 3388 24724 3444 24734
rect 3388 24276 3444 24668
rect 3388 24210 3444 24220
rect 3388 23940 3444 23950
rect 3388 19908 3444 23884
rect 3500 21588 3556 26342
rect 3500 21028 3556 21532
rect 3500 20962 3556 20972
rect 3388 19842 3444 19852
rect 3276 13122 3332 13132
rect 3388 17668 3444 17678
rect 3388 12516 3444 17612
rect 3500 17444 3556 17454
rect 3500 15958 3556 17388
rect 3612 16100 3668 28812
rect 3612 16034 3668 16044
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3776 25116 4096 26628
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 3776 23548 4096 25060
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3776 20412 4096 21924
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 3776 18844 4096 20356
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3500 15902 3668 15958
rect 3612 15876 3668 15902
rect 3388 12450 3444 12460
rect 3500 13748 3556 13758
rect 3276 12180 3332 12190
rect 3276 11458 3332 12124
rect 3500 12180 3556 13692
rect 3612 12628 3668 15820
rect 3612 12562 3668 12572
rect 3776 15708 4096 17220
rect 4172 37156 4228 37166
rect 4172 16772 4228 37100
rect 4284 36932 4340 37660
rect 4284 36866 4340 36876
rect 4436 36876 4756 38388
rect 5068 38388 5124 41804
rect 5180 40740 5236 40750
rect 5180 38724 5236 40684
rect 5292 38836 5348 50652
rect 5292 38770 5348 38780
rect 5180 38658 5236 38668
rect 4956 37604 5012 37614
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4844 37156 4900 37166
rect 4844 36932 4900 37100
rect 4844 36866 4900 36876
rect 4436 35308 4756 36820
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4284 34132 4340 34142
rect 4284 33796 4340 34076
rect 4284 33730 4340 33740
rect 4436 33740 4756 35252
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 4284 32900 4340 32910
rect 4284 31780 4340 32844
rect 4284 30212 4340 31724
rect 4284 30146 4340 30156
rect 4436 32172 4756 33684
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4844 33796 4900 33806
rect 4844 30212 4900 33740
rect 4844 30146 4900 30156
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4956 29092 5012 37548
rect 5068 37558 5124 38332
rect 5292 37716 5348 37726
rect 5068 37502 5236 37558
rect 5068 37268 5124 37278
rect 5068 36820 5124 37212
rect 5068 36754 5124 36764
rect 5180 31780 5236 37502
rect 5292 35364 5348 37660
rect 5292 35298 5348 35308
rect 5180 31714 5236 31724
rect 5292 34020 5348 34030
rect 5292 30100 5348 33964
rect 5292 30034 5348 30044
rect 5292 29876 5348 29886
rect 4956 28868 5012 29036
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4844 28420 4900 28430
rect 4844 27076 4900 28364
rect 4956 28196 5012 28812
rect 4956 28130 5012 28140
rect 5068 29764 5124 29774
rect 5068 28084 5124 29708
rect 4844 27010 4900 27020
rect 4956 27412 5012 27422
rect 4956 26938 5012 27356
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4172 16706 4228 16716
rect 4284 23492 4340 23502
rect 4284 18340 4340 23436
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 3776 14140 4096 15652
rect 4172 16548 4228 16558
rect 4172 15540 4228 16492
rect 4172 15474 4228 15484
rect 4284 15418 4340 18284
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3776 12572 4096 14084
rect 3500 12114 3556 12124
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3276 11402 3444 11458
rect 3276 11284 3332 11294
rect 3276 9298 3332 11228
rect 3388 9492 3444 11402
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3388 9426 3444 9436
rect 3500 10388 3556 10398
rect 3276 9242 3444 9298
rect 3164 8194 3220 8204
rect 3388 7028 3444 9242
rect 3500 8038 3556 10332
rect 3776 9436 4096 10948
rect 4172 15362 4340 15418
rect 4436 22764 4756 24276
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4844 26882 5012 26938
rect 4844 20098 4900 26882
rect 4956 26516 5012 26526
rect 4956 25956 5012 26460
rect 4956 25890 5012 25900
rect 4956 25508 5012 25518
rect 4956 25060 5012 25452
rect 4956 24994 5012 25004
rect 4956 24724 5012 24734
rect 4956 24276 5012 24668
rect 5068 24388 5124 28028
rect 5180 29316 5236 29326
rect 5180 26964 5236 29260
rect 5292 27412 5348 29820
rect 5292 27346 5348 27356
rect 5180 26898 5236 26908
rect 5404 26964 5460 50764
rect 5516 48804 5572 48814
rect 5516 41860 5572 48748
rect 5740 46788 5796 46798
rect 5740 46452 5796 46732
rect 5628 46004 5684 46014
rect 5628 45332 5684 45948
rect 5628 45266 5684 45276
rect 5516 41794 5572 41804
rect 5628 44996 5684 45006
rect 5628 41698 5684 44940
rect 5740 43540 5796 46396
rect 5740 43474 5796 43484
rect 5516 41642 5684 41698
rect 5516 37940 5572 41642
rect 5628 41188 5684 41198
rect 5628 39358 5684 41132
rect 5740 40516 5796 40526
rect 5740 39620 5796 40460
rect 5740 39554 5796 39564
rect 5628 39302 5796 39358
rect 5516 37156 5572 37884
rect 5516 37090 5572 37100
rect 5628 38052 5684 38062
rect 5516 34244 5572 34254
rect 5516 29764 5572 34188
rect 5628 33572 5684 37996
rect 5740 36148 5796 39302
rect 5740 36082 5796 36092
rect 5628 30212 5684 33516
rect 5628 30146 5684 30156
rect 5740 35812 5796 35822
rect 5516 29698 5572 29708
rect 5068 24322 5124 24332
rect 5180 26740 5236 26750
rect 4956 24210 5012 24220
rect 5180 24164 5236 26684
rect 5292 24612 5348 24622
rect 5292 24388 5348 24556
rect 5292 24322 5348 24332
rect 5180 24098 5236 24108
rect 4956 23156 5012 23166
rect 4956 22596 5012 23100
rect 4956 22530 5012 22540
rect 5068 22708 5124 22718
rect 4844 20042 5012 20098
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 4436 16492 4756 18004
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4172 10388 4228 15362
rect 4172 10322 4228 10332
rect 4284 15204 4340 15214
rect 4284 9828 4340 15148
rect 4284 9762 4340 9772
rect 4436 14924 4756 16436
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 4436 13356 4756 14868
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 4844 19908 4900 19918
rect 4844 10612 4900 19852
rect 4956 17332 5012 20042
rect 5068 19572 5124 22652
rect 5068 17444 5124 19516
rect 5404 22148 5460 26908
rect 5628 26404 5684 26414
rect 5516 25956 5572 25966
rect 5516 25060 5572 25900
rect 5516 24994 5572 25004
rect 5404 20692 5460 22092
rect 5516 24724 5572 24734
rect 5516 20804 5572 24668
rect 5628 23940 5684 26348
rect 5628 23874 5684 23884
rect 5516 20738 5572 20748
rect 5068 17378 5124 17388
rect 5292 17444 5348 17454
rect 4956 15204 5012 17276
rect 5180 16996 5236 17006
rect 5180 16772 5236 16940
rect 5180 16706 5236 16716
rect 4956 15138 5012 15148
rect 5180 15316 5236 15326
rect 4956 14980 5012 14990
rect 4956 13972 5012 14924
rect 4956 13906 5012 13916
rect 5068 14868 5124 14878
rect 4956 13076 5012 13086
rect 4956 12292 5012 13020
rect 4956 12226 5012 12236
rect 4844 10546 4900 10556
rect 4956 11508 5012 11518
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3612 8038 3668 8046
rect 3500 8036 3668 8038
rect 3500 7982 3612 8036
rect 3612 7970 3668 7980
rect 3388 6962 3444 6972
rect 3776 7868 4096 9380
rect 4284 9492 4340 9502
rect 4284 8260 4340 9436
rect 4284 8194 4340 8204
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3052 5842 3108 5852
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3164 5572 3220 5582
rect 3220 5516 3556 5518
rect 3164 5462 3556 5516
rect 3500 5460 3556 5462
rect 3500 5394 3556 5404
rect 3500 5236 3556 5246
rect 3500 3892 3556 5180
rect 3612 4788 3668 4798
rect 3612 4116 3668 4732
rect 3612 4050 3668 4060
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3500 3826 3556 3836
rect 3500 3668 3556 3678
rect 3500 3538 3556 3612
rect 3332 3482 3556 3538
rect 3332 3444 3388 3482
rect 3332 3378 3388 3388
rect 2940 1876 2996 3276
rect 2940 1810 2996 1820
rect 3776 3164 4096 4676
rect 4172 7924 4228 7934
rect 4172 4004 4228 7868
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4172 3938 4228 3948
rect 4284 6244 4340 6254
rect 4284 3718 4340 6188
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 2492 578 2548 588
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4172 3662 4340 3718
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4172 1204 4228 3662
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4172 1138 4228 1148
rect 4284 1316 4340 1326
rect 4284 868 4340 1260
rect 4284 802 4340 812
rect 4436 812 4756 2324
rect 4844 10388 4900 10398
rect 4844 1204 4900 10332
rect 4956 8758 5012 11452
rect 5068 9268 5124 14812
rect 5180 10836 5236 15260
rect 5292 12964 5348 17388
rect 5404 14532 5460 20636
rect 5740 20020 5796 35756
rect 5740 19954 5796 19964
rect 5852 28308 5908 52668
rect 5964 52052 6020 54348
rect 6076 53284 6132 53294
rect 6076 52724 6132 53228
rect 6076 52658 6132 52668
rect 5964 36372 6020 51996
rect 6076 50372 6132 50382
rect 6076 49252 6132 50316
rect 6188 49364 6244 57148
rect 22764 57204 22820 57214
rect 21308 57092 21364 57102
rect 16492 56980 16548 56990
rect 13356 55748 13412 55758
rect 9436 55524 9492 55534
rect 6860 55412 6916 55422
rect 6188 49298 6244 49308
rect 6412 53956 6468 53966
rect 6076 49186 6132 49196
rect 5964 36306 6020 36316
rect 6076 47684 6132 47694
rect 6076 35924 6132 47628
rect 6300 45332 6356 45342
rect 6188 45220 6244 45230
rect 6188 44436 6244 45164
rect 6300 44772 6356 45276
rect 6300 44706 6356 44716
rect 6188 44370 6244 44380
rect 6076 35858 6132 35868
rect 6188 39060 6244 39070
rect 5964 35252 6020 35262
rect 5964 33124 6020 35196
rect 5964 30996 6020 33068
rect 6076 35140 6132 35150
rect 6076 31332 6132 35084
rect 6076 31266 6132 31276
rect 5964 30930 6020 30940
rect 6076 29876 6132 29886
rect 5964 29540 6020 29550
rect 5964 29204 6020 29484
rect 5964 29138 6020 29148
rect 5740 19796 5796 19806
rect 5404 14466 5460 14476
rect 5516 18116 5572 18126
rect 5516 14338 5572 18060
rect 5740 17444 5796 19740
rect 5740 17378 5796 17388
rect 5292 12898 5348 12908
rect 5404 14282 5572 14338
rect 5628 15092 5684 15102
rect 5180 10770 5236 10780
rect 5292 12740 5348 12750
rect 5068 9202 5124 9212
rect 5180 8932 5236 8942
rect 4956 8708 5124 8758
rect 4956 8702 5068 8708
rect 5068 8642 5124 8652
rect 4956 8596 5012 8606
rect 4956 7476 5012 8540
rect 4956 7410 5012 7420
rect 5180 6468 5236 8876
rect 5180 6402 5236 6412
rect 5292 4788 5348 12684
rect 5404 11508 5460 14282
rect 5628 13618 5684 15036
rect 5516 13562 5684 13618
rect 5740 14756 5796 14766
rect 5516 13524 5572 13562
rect 5516 13458 5572 13468
rect 5628 13412 5684 13422
rect 5404 11442 5460 11452
rect 5516 13076 5572 13086
rect 5404 10836 5460 10846
rect 5404 7028 5460 10780
rect 5516 9268 5572 13020
rect 5628 11620 5684 13356
rect 5740 13076 5796 14700
rect 5740 13010 5796 13020
rect 5628 11554 5684 11564
rect 5852 11458 5908 28252
rect 5964 28756 6020 28766
rect 5964 24724 6020 28700
rect 5964 24658 6020 24668
rect 6076 20998 6132 29820
rect 5964 20942 6132 20998
rect 5964 17220 6020 20942
rect 5964 17154 6020 17164
rect 6076 20804 6132 20814
rect 5740 11402 5908 11458
rect 5516 9202 5572 9212
rect 5628 11284 5684 11294
rect 5404 6962 5460 6972
rect 5628 4900 5684 11228
rect 5740 11098 5796 11402
rect 5740 11042 5908 11098
rect 5628 4834 5684 4844
rect 5292 4722 5348 4732
rect 4844 1138 4900 1148
rect 5852 1204 5908 11042
rect 5964 11060 6020 11070
rect 5964 10836 6020 11004
rect 5964 10770 6020 10780
rect 5964 10500 6020 10510
rect 5964 4004 6020 10444
rect 5964 3938 6020 3948
rect 6076 1652 6132 20748
rect 6188 17892 6244 39004
rect 6300 36820 6356 36830
rect 6300 35476 6356 36764
rect 6300 35410 6356 35420
rect 6412 34580 6468 53900
rect 6636 53620 6692 53630
rect 6636 52276 6692 53564
rect 6636 52210 6692 52220
rect 6748 52836 6804 52846
rect 6412 34514 6468 34524
rect 6524 51156 6580 51166
rect 6412 32116 6468 32126
rect 6300 31444 6356 31454
rect 6300 28196 6356 31388
rect 6300 28130 6356 28140
rect 6300 27972 6356 27982
rect 6300 20804 6356 27916
rect 6300 20738 6356 20748
rect 6412 20638 6468 32060
rect 6524 29316 6580 51100
rect 6748 49140 6804 52780
rect 6748 49074 6804 49084
rect 6748 47124 6804 47134
rect 6636 45444 6692 45454
rect 6636 44212 6692 45388
rect 6636 44146 6692 44156
rect 6636 43316 6692 43326
rect 6636 41878 6692 43260
rect 6748 43204 6804 47068
rect 6748 43138 6804 43148
rect 6636 41822 6804 41878
rect 6524 29250 6580 29260
rect 6636 35476 6692 35486
rect 6300 20582 6468 20638
rect 6524 23044 6580 23054
rect 6300 19796 6356 20582
rect 6300 19572 6356 19740
rect 6300 19506 6356 19516
rect 6412 20468 6468 20478
rect 6188 17826 6244 17836
rect 6300 19012 6356 19022
rect 6300 17780 6356 18956
rect 6188 17444 6244 17454
rect 6188 13748 6244 17388
rect 6188 13682 6244 13692
rect 6300 14532 6356 17724
rect 6412 16138 6468 20412
rect 6524 19012 6580 22988
rect 6524 18946 6580 18956
rect 6524 18676 6580 18686
rect 6524 16324 6580 18620
rect 6524 16258 6580 16268
rect 6412 16082 6580 16138
rect 6188 13524 6244 13534
rect 6188 10836 6244 13468
rect 6300 13076 6356 14476
rect 6412 13524 6468 13534
rect 6412 13300 6468 13468
rect 6412 13234 6468 13244
rect 6300 13010 6356 13020
rect 6412 12852 6468 12862
rect 6188 10770 6244 10780
rect 6300 12068 6356 12078
rect 6300 10276 6356 12012
rect 6300 10210 6356 10220
rect 6188 9268 6244 9278
rect 6188 2212 6244 9212
rect 6300 8036 6356 8046
rect 6300 5908 6356 7980
rect 6412 7812 6468 12796
rect 6412 7588 6468 7756
rect 6412 7522 6468 7532
rect 6524 7476 6580 16082
rect 6524 7410 6580 7420
rect 6300 5842 6356 5852
rect 6188 2146 6244 2156
rect 6076 1586 6132 1596
rect 5852 1138 5908 1148
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 6636 756 6692 35420
rect 6748 18838 6804 41822
rect 6860 36708 6916 55356
rect 8204 55300 8260 55310
rect 7644 54180 7700 54190
rect 7308 53844 7364 53854
rect 6972 53508 7028 53518
rect 6972 52948 7028 53452
rect 7308 53060 7364 53788
rect 7308 52994 7364 53004
rect 7420 53396 7476 53406
rect 6972 52882 7028 52892
rect 7308 52052 7364 52062
rect 7084 51044 7140 51054
rect 6972 45556 7028 45566
rect 6972 43988 7028 45500
rect 7084 44578 7140 50988
rect 7084 44522 7252 44578
rect 6972 43922 7028 43932
rect 7084 43540 7140 43550
rect 6972 43316 7028 43326
rect 6972 41412 7028 43260
rect 6972 41346 7028 41356
rect 6860 36642 6916 36652
rect 6972 40852 7028 40862
rect 6972 35364 7028 40796
rect 6972 35298 7028 35308
rect 7084 33012 7140 43484
rect 7196 35140 7252 44522
rect 7308 42756 7364 51996
rect 7420 51492 7476 53340
rect 7420 51426 7476 51436
rect 7308 39956 7364 42700
rect 7308 39890 7364 39900
rect 7420 47124 7476 47134
rect 7420 46004 7476 47068
rect 7196 33908 7252 35084
rect 7196 33842 7252 33852
rect 7084 32946 7140 32956
rect 7196 32564 7252 32574
rect 7084 32340 7140 32350
rect 6972 31332 7028 31342
rect 6860 30436 6916 30446
rect 6860 26404 6916 30380
rect 6972 29988 7028 31276
rect 6972 29922 7028 29932
rect 7084 30324 7140 32284
rect 6860 26338 6916 26348
rect 6972 27748 7028 27758
rect 6972 23940 7028 27692
rect 7084 27524 7140 30268
rect 7196 28980 7252 32508
rect 7308 31108 7364 31118
rect 7308 30772 7364 31052
rect 7308 30706 7364 30716
rect 7196 28914 7252 28924
rect 7084 27458 7140 27468
rect 7196 27412 7252 27422
rect 7196 26516 7252 27356
rect 7196 26450 7252 26460
rect 6972 23874 7028 23884
rect 7196 23156 7252 23166
rect 7196 19236 7252 23100
rect 7196 19170 7252 19180
rect 6748 18782 7364 18838
rect 7084 18340 7140 18350
rect 6748 16772 6804 16782
rect 6748 14756 6804 16716
rect 7084 16660 7140 18284
rect 7084 16594 7140 16604
rect 7196 16212 7252 16222
rect 6972 16100 7028 16110
rect 6972 15092 7028 16044
rect 6748 14532 6804 14700
rect 6748 14466 6804 14476
rect 6860 14980 6916 14990
rect 6748 12404 6804 12414
rect 6748 11956 6804 12348
rect 6748 11890 6804 11900
rect 6748 11508 6804 11518
rect 6748 9044 6804 11452
rect 6860 10558 6916 14924
rect 6972 11396 7028 15036
rect 7084 15652 7140 15662
rect 7084 11508 7140 15596
rect 7196 13412 7252 16156
rect 7196 13346 7252 13356
rect 7084 11442 7140 11452
rect 7196 12852 7252 12862
rect 6972 11330 7028 11340
rect 6860 10502 7140 10558
rect 6748 8978 6804 8988
rect 6860 10164 6916 10174
rect 6748 8036 6804 8046
rect 6748 5572 6804 7980
rect 6860 6244 6916 10108
rect 7084 6356 7140 10502
rect 7196 10276 7252 12796
rect 7196 10210 7252 10220
rect 7308 11956 7364 18782
rect 7420 18452 7476 45948
rect 7532 45668 7588 45678
rect 7532 44212 7588 45612
rect 7532 44146 7588 44156
rect 7532 32452 7588 32462
rect 7532 28196 7588 32396
rect 7532 28130 7588 28140
rect 7420 18386 7476 18396
rect 7532 25844 7588 25854
rect 7084 6290 7140 6300
rect 6860 6178 6916 6188
rect 7308 6058 7364 11900
rect 6748 5506 6804 5516
rect 6860 6002 7364 6058
rect 7420 12180 7476 12190
rect 6860 3332 6916 6002
rect 7420 4564 7476 12124
rect 7532 7924 7588 25788
rect 7644 22148 7700 54124
rect 7868 54180 7924 54190
rect 7868 52724 7924 54124
rect 7868 52658 7924 52668
rect 8092 52388 8148 52398
rect 7868 50596 7924 50606
rect 7756 48020 7812 48030
rect 7756 47236 7812 47964
rect 7756 47170 7812 47180
rect 7868 47124 7924 50540
rect 7868 47058 7924 47068
rect 7980 49476 8036 49486
rect 7980 48356 8036 49420
rect 7756 46676 7812 46686
rect 7756 38612 7812 46620
rect 7980 44100 8036 48300
rect 7980 44034 8036 44044
rect 7756 38546 7812 38556
rect 7868 43988 7924 43998
rect 7868 38276 7924 43932
rect 7868 37604 7924 38220
rect 7868 37538 7924 37548
rect 7980 38836 8036 38846
rect 7980 37044 8036 38780
rect 7868 35924 7924 35934
rect 7756 34580 7812 34590
rect 7756 22596 7812 34524
rect 7756 22530 7812 22540
rect 7644 22082 7700 22092
rect 7644 21476 7700 21486
rect 7644 20458 7700 21420
rect 7644 20402 7812 20458
rect 7644 20132 7700 20142
rect 7644 18788 7700 20076
rect 7644 16660 7700 18732
rect 7756 18116 7812 20402
rect 7756 18050 7812 18060
rect 7644 15652 7700 16604
rect 7644 15586 7700 15596
rect 7756 16884 7812 16894
rect 7756 13188 7812 16828
rect 7756 13122 7812 13132
rect 7868 12068 7924 35868
rect 7980 35476 8036 36988
rect 7980 35410 8036 35420
rect 7980 33348 8036 33358
rect 7980 32452 8036 33292
rect 7980 32386 8036 32396
rect 7980 32116 8036 32126
rect 7980 31556 8036 32060
rect 7980 31490 8036 31500
rect 7980 28644 8036 28654
rect 7980 25396 8036 28588
rect 8092 28532 8148 52332
rect 8204 30772 8260 55244
rect 8540 55300 8596 55310
rect 8428 53956 8484 53966
rect 8428 53172 8484 53900
rect 8428 53106 8484 53116
rect 8428 51380 8484 51390
rect 8428 49812 8484 51324
rect 8428 49746 8484 49756
rect 8204 30706 8260 30716
rect 8316 45220 8372 45230
rect 8092 28466 8148 28476
rect 8204 29764 8260 29774
rect 7980 25330 8036 25340
rect 7980 24388 8036 24398
rect 7980 18452 8036 24332
rect 8204 24388 8260 29708
rect 8204 24322 8260 24332
rect 7980 18386 8036 18396
rect 8092 22932 8148 22942
rect 7868 11284 7924 12012
rect 7868 11218 7924 11228
rect 7980 10276 8036 10286
rect 7532 7858 7588 7868
rect 7868 9828 7924 9838
rect 7420 4498 7476 4508
rect 6860 2660 6916 3276
rect 6860 2594 6916 2604
rect 7756 2884 7812 2894
rect 6636 690 6692 700
rect 7756 308 7812 2828
rect 7868 1204 7924 9772
rect 7980 9044 8036 10220
rect 7980 8978 8036 8988
rect 7980 5908 8036 5918
rect 7980 4564 8036 5852
rect 7980 4498 8036 4508
rect 8092 2772 8148 22876
rect 8204 12740 8260 12750
rect 8204 12404 8260 12684
rect 8204 12338 8260 12348
rect 8092 2706 8148 2716
rect 8204 7588 8260 7598
rect 8204 1540 8260 7532
rect 8316 1652 8372 45164
rect 8428 41188 8484 41198
rect 8428 38836 8484 41132
rect 8428 38770 8484 38780
rect 8428 37716 8484 37726
rect 8428 35812 8484 37660
rect 8428 35746 8484 35756
rect 8428 35588 8484 35598
rect 8428 34916 8484 35532
rect 8428 34850 8484 34860
rect 8316 1586 8372 1596
rect 8428 33012 8484 33022
rect 8428 32340 8484 32956
rect 8204 1474 8260 1484
rect 8428 1316 8484 32284
rect 8540 28196 8596 55244
rect 8988 54404 9044 54414
rect 8652 53284 8708 53294
rect 8652 36372 8708 53228
rect 8988 52388 9044 54348
rect 8988 52322 9044 52332
rect 8764 50372 8820 50382
rect 8764 44324 8820 50316
rect 9100 49812 9156 49822
rect 8764 44258 8820 44268
rect 8988 45668 9044 45678
rect 8652 36306 8708 36316
rect 8764 43876 8820 43886
rect 8764 41860 8820 43820
rect 8988 42868 9044 45612
rect 8988 42802 9044 42812
rect 8764 34804 8820 41804
rect 8876 41636 8932 41646
rect 8876 40964 8932 41580
rect 8876 40898 8932 40908
rect 8876 39844 8932 39854
rect 8876 35924 8932 39788
rect 8876 35858 8932 35868
rect 8764 34738 8820 34748
rect 8988 34468 9044 34478
rect 8876 30772 8932 30782
rect 8540 28130 8596 28140
rect 8764 30324 8820 30334
rect 8540 26628 8596 26638
rect 8540 25284 8596 26572
rect 8540 25218 8596 25228
rect 8540 22932 8596 22942
rect 8540 20244 8596 22876
rect 8540 20178 8596 20188
rect 8652 21812 8708 21822
rect 8652 20098 8708 21756
rect 8540 20042 8708 20098
rect 8540 17892 8596 20042
rect 8540 7476 8596 17836
rect 8652 15540 8708 15550
rect 8652 14756 8708 15484
rect 8652 14690 8708 14700
rect 8540 7410 8596 7420
rect 8652 9604 8708 9614
rect 8652 7252 8708 9548
rect 8652 6468 8708 7196
rect 8652 6402 8708 6412
rect 8652 4564 8708 4574
rect 8652 2660 8708 4508
rect 8652 2594 8708 2604
rect 8428 1250 8484 1260
rect 7868 1138 7924 1148
rect 8764 1204 8820 30268
rect 8876 25620 8932 30716
rect 8988 30548 9044 34412
rect 9100 34020 9156 49756
rect 9212 47684 9268 47694
rect 9212 39844 9268 47628
rect 9212 39778 9268 39788
rect 9324 42308 9380 42318
rect 9324 36838 9380 42252
rect 9436 37044 9492 55468
rect 9660 55524 9716 55534
rect 9548 43092 9604 43102
rect 9548 41524 9604 43036
rect 9548 41458 9604 41468
rect 9548 40964 9604 40974
rect 9548 39844 9604 40908
rect 9548 39778 9604 39788
rect 9548 39508 9604 39518
rect 9548 38724 9604 39452
rect 9548 38658 9604 38668
rect 9436 36978 9492 36988
rect 9324 36782 9492 36838
rect 9436 35812 9492 36782
rect 9660 36596 9716 55468
rect 10444 55300 10500 55310
rect 9660 36530 9716 36540
rect 9772 54292 9828 54302
rect 9436 35746 9492 35756
rect 9100 33238 9156 33964
rect 9436 35588 9492 35598
rect 9100 33182 9268 33238
rect 8988 30482 9044 30492
rect 9100 31332 9156 31342
rect 8876 25554 8932 25564
rect 8988 29204 9044 29214
rect 8876 23156 8932 23166
rect 8876 21588 8932 23100
rect 8876 21522 8932 21532
rect 8988 20998 9044 29148
rect 9100 23716 9156 31276
rect 9100 23650 9156 23660
rect 8876 20942 9044 20998
rect 8876 10164 8932 20942
rect 9100 18452 9156 18462
rect 8876 10098 8932 10108
rect 8988 11284 9044 11294
rect 8988 1540 9044 11228
rect 9100 6692 9156 18396
rect 9100 6626 9156 6636
rect 9100 6244 9156 6254
rect 9100 4900 9156 6188
rect 9100 4834 9156 4844
rect 9212 1652 9268 33182
rect 9436 30548 9492 35532
rect 9436 30482 9492 30492
rect 9548 32228 9604 32238
rect 9324 29652 9380 29662
rect 9548 29638 9604 32172
rect 9324 19236 9380 29596
rect 9324 19170 9380 19180
rect 9436 29582 9604 29638
rect 9660 30772 9716 30782
rect 9436 18340 9492 29582
rect 9548 26068 9604 26078
rect 9548 25396 9604 26012
rect 9548 25330 9604 25340
rect 9660 22372 9716 30716
rect 9772 25396 9828 54236
rect 9996 53396 10052 53406
rect 9996 46116 10052 53340
rect 9996 46050 10052 46060
rect 10108 51940 10164 51950
rect 9884 45892 9940 45902
rect 9884 39732 9940 45836
rect 9884 38164 9940 39676
rect 9884 38098 9940 38108
rect 9996 41188 10052 41198
rect 9996 34804 10052 41132
rect 9996 34738 10052 34748
rect 9996 34244 10052 34254
rect 9884 31780 9940 31790
rect 9884 30772 9940 31724
rect 9884 30706 9940 30716
rect 9996 27860 10052 34188
rect 9996 27794 10052 27804
rect 9772 25330 9828 25340
rect 9884 25620 9940 25630
rect 9772 23492 9828 23502
rect 9772 22708 9828 23436
rect 9772 22642 9828 22652
rect 9660 22306 9716 22316
rect 9436 18274 9492 18284
rect 9548 22148 9604 22158
rect 9548 15652 9604 22092
rect 9884 22078 9940 25564
rect 9996 24052 10052 24062
rect 9996 23268 10052 23996
rect 9996 23202 10052 23212
rect 9548 15586 9604 15596
rect 9660 22022 9940 22078
rect 9660 14338 9716 22022
rect 10108 20998 10164 51884
rect 10220 49812 10276 49822
rect 10220 46676 10276 49756
rect 10332 48020 10388 48030
rect 10332 47124 10388 47964
rect 10332 47058 10388 47068
rect 10220 46610 10276 46620
rect 10332 38836 10388 38846
rect 10332 37156 10388 38780
rect 10332 37018 10388 37100
rect 10220 36962 10388 37018
rect 10220 35218 10276 36962
rect 10220 35162 10388 35218
rect 10332 31668 10388 35162
rect 10332 31602 10388 31612
rect 10444 30996 10500 55244
rect 13132 55076 13188 55086
rect 12796 54740 12852 54750
rect 12460 53732 12516 53742
rect 11564 53620 11620 53630
rect 10668 53284 10724 53294
rect 10668 52276 10724 53228
rect 10668 52210 10724 52220
rect 10668 51268 10724 51278
rect 10668 49140 10724 51212
rect 10668 49074 10724 49084
rect 10892 49924 10948 49934
rect 10892 48244 10948 49868
rect 11340 49252 11396 49262
rect 10892 48178 10948 48188
rect 11004 48692 11060 48702
rect 10892 46452 10948 46462
rect 10780 44884 10836 44894
rect 10556 43876 10612 43886
rect 10556 42196 10612 43820
rect 10556 42130 10612 42140
rect 10444 30930 10500 30940
rect 10556 40404 10612 40414
rect 10444 30212 10500 30222
rect 10444 26964 10500 30156
rect 10556 28532 10612 40348
rect 10668 40180 10724 40190
rect 10668 39844 10724 40124
rect 10668 39778 10724 39788
rect 10780 38836 10836 44828
rect 10892 41636 10948 46396
rect 11004 46018 11060 48636
rect 11228 48580 11284 48590
rect 11228 47684 11284 48524
rect 11228 47618 11284 47628
rect 11340 46340 11396 49196
rect 11004 45962 11172 46018
rect 11116 45556 11172 45962
rect 11116 45298 11172 45500
rect 11004 45242 11172 45298
rect 11004 44772 11060 45242
rect 11004 44706 11060 44716
rect 10892 41570 10948 41580
rect 11116 44660 11172 44670
rect 10780 38770 10836 38780
rect 10892 39284 10948 39294
rect 10892 38612 10948 39228
rect 10892 38546 10948 38556
rect 11004 33908 11060 33918
rect 10556 28466 10612 28476
rect 10668 30884 10724 30894
rect 10668 28378 10724 30828
rect 10892 30100 10948 30110
rect 10444 26898 10500 26908
rect 10556 28322 10724 28378
rect 10780 28532 10836 28542
rect 10444 22372 10500 22382
rect 10332 21476 10388 21486
rect 10332 21252 10388 21420
rect 10108 20942 10276 20998
rect 9884 20132 9940 20142
rect 9436 14282 9716 14338
rect 9772 16548 9828 16558
rect 9436 11396 9492 14282
rect 9660 13972 9716 13982
rect 9436 11330 9492 11340
rect 9548 13524 9604 13534
rect 9436 11060 9492 11070
rect 9436 10388 9492 11004
rect 9436 10322 9492 10332
rect 9436 10052 9492 10062
rect 9324 9716 9380 9726
rect 9324 9492 9380 9660
rect 9324 9426 9380 9436
rect 9436 9268 9492 9996
rect 9324 7140 9380 7150
rect 9324 5908 9380 7084
rect 9324 5842 9380 5852
rect 9436 4564 9492 9212
rect 9548 8260 9604 13468
rect 9660 13076 9716 13916
rect 9660 11956 9716 13020
rect 9660 11890 9716 11900
rect 9660 11620 9716 11630
rect 9660 11060 9716 11564
rect 9660 10994 9716 11004
rect 9660 10052 9716 10062
rect 9660 9716 9716 9996
rect 9660 9650 9716 9660
rect 9548 8194 9604 8204
rect 9436 4228 9492 4508
rect 9436 4162 9492 4172
rect 9660 7476 9716 7486
rect 9660 3892 9716 7420
rect 9660 2212 9716 3836
rect 9772 3780 9828 16492
rect 9884 9268 9940 20076
rect 10108 20020 10164 20030
rect 9996 15204 10052 15214
rect 9996 13972 10052 15148
rect 9996 13906 10052 13916
rect 9996 11844 10052 11854
rect 9996 11620 10052 11788
rect 9996 11554 10052 11564
rect 9884 9202 9940 9212
rect 9996 11396 10052 11406
rect 9996 9118 10052 11340
rect 10108 10052 10164 19964
rect 10220 13972 10276 20942
rect 10220 13906 10276 13916
rect 10108 9986 10164 9996
rect 10220 11060 10276 11070
rect 9772 3714 9828 3724
rect 9884 9062 10052 9118
rect 9660 2146 9716 2156
rect 9212 1586 9268 1596
rect 8988 1474 9044 1484
rect 8764 1138 8820 1148
rect 9884 1204 9940 9062
rect 10108 7476 10164 7486
rect 9996 6692 10052 6702
rect 9996 4618 10052 6636
rect 10108 5908 10164 7420
rect 10108 5842 10164 5852
rect 9996 4562 10164 4618
rect 10108 4340 10164 4562
rect 10108 4274 10164 4284
rect 10220 1988 10276 11004
rect 10332 8260 10388 21196
rect 10444 13748 10500 22316
rect 10444 13682 10500 13692
rect 10556 12964 10612 28322
rect 10668 19908 10724 19918
rect 10668 18340 10724 19852
rect 10668 18274 10724 18284
rect 10556 12898 10612 12908
rect 10332 8194 10388 8204
rect 10220 1922 10276 1932
rect 9884 1138 9940 1148
rect 7756 242 7812 252
rect 10780 84 10836 28476
rect 10892 27412 10948 30044
rect 10892 27346 10948 27356
rect 11004 25678 11060 33852
rect 10892 25622 11060 25678
rect 10892 21178 10948 25622
rect 11004 25396 11060 25406
rect 11004 23268 11060 25340
rect 11004 23202 11060 23212
rect 10892 21122 11060 21178
rect 11004 20132 11060 21122
rect 11004 19124 11060 20076
rect 11004 19058 11060 19068
rect 11116 16772 11172 44604
rect 11228 44324 11284 44334
rect 11228 27636 11284 44268
rect 11340 38388 11396 46284
rect 11452 48244 11508 48254
rect 11452 45668 11508 48188
rect 11452 40180 11508 45612
rect 11452 40114 11508 40124
rect 11340 38322 11396 38332
rect 11340 35364 11396 35374
rect 11340 32900 11396 35308
rect 11340 32834 11396 32844
rect 11452 33348 11508 33358
rect 11452 32564 11508 33292
rect 11452 32498 11508 32508
rect 11228 27570 11284 27580
rect 11340 28196 11396 28206
rect 11116 16706 11172 16716
rect 11340 16548 11396 28140
rect 11564 25620 11620 53564
rect 11564 25554 11620 25564
rect 11676 53508 11732 53518
rect 11676 25318 11732 53452
rect 12124 52388 12180 52398
rect 12124 51604 12180 52332
rect 12012 50036 12068 50046
rect 12012 49812 12068 49980
rect 12012 49746 12068 49756
rect 11788 45892 11844 45902
rect 11788 39732 11844 45836
rect 11900 42868 11956 42878
rect 11900 40978 11956 42812
rect 12012 42084 12068 42094
rect 12012 41188 12068 42028
rect 12012 41122 12068 41132
rect 11900 40922 12068 40978
rect 11788 35812 11844 39676
rect 11788 35746 11844 35756
rect 11900 40404 11956 40414
rect 11788 33908 11844 33918
rect 11788 25508 11844 33852
rect 11788 25442 11844 25452
rect 11676 25262 11844 25318
rect 11676 25060 11732 25070
rect 11340 16482 11396 16492
rect 11564 23044 11620 23054
rect 11564 19236 11620 22988
rect 11452 15652 11508 15662
rect 11004 14532 11060 14542
rect 11004 13748 11060 14476
rect 11004 8578 11060 13692
rect 11228 13972 11284 13982
rect 11228 13748 11284 13916
rect 11228 13682 11284 13692
rect 11116 12628 11172 12638
rect 11116 12068 11172 12572
rect 11116 12002 11172 12012
rect 11340 12068 11396 12078
rect 11004 8522 11172 8578
rect 11116 3780 11172 8522
rect 11340 5572 11396 12012
rect 11340 5506 11396 5516
rect 11116 3714 11172 3724
rect 11452 1652 11508 15596
rect 11564 13300 11620 19180
rect 11564 13234 11620 13244
rect 11564 12404 11620 12414
rect 11564 8820 11620 12348
rect 11564 8754 11620 8764
rect 11452 1586 11508 1596
rect 11564 6020 11620 6030
rect 11564 1092 11620 5964
rect 11676 1540 11732 25004
rect 11788 16660 11844 25262
rect 11788 16594 11844 16604
rect 11788 12292 11844 12302
rect 11788 6020 11844 12236
rect 11788 5954 11844 5964
rect 11676 1474 11732 1484
rect 11564 1026 11620 1036
rect 11900 756 11956 40348
rect 12012 37716 12068 40922
rect 12012 25508 12068 37660
rect 12012 25442 12068 25452
rect 12012 23268 12068 23278
rect 12012 18340 12068 23212
rect 12012 18274 12068 18284
rect 12012 15876 12068 15886
rect 12012 6020 12068 15820
rect 12124 14868 12180 51548
rect 12348 50708 12404 50718
rect 12348 50484 12404 50652
rect 12348 50418 12404 50428
rect 12460 50372 12516 53676
rect 12460 49028 12516 50316
rect 12460 48962 12516 48972
rect 12684 51268 12740 51278
rect 12684 50484 12740 51212
rect 12348 48356 12404 48366
rect 12236 46116 12292 46126
rect 12236 40404 12292 46060
rect 12236 40338 12292 40348
rect 12236 32564 12292 32574
rect 12236 32004 12292 32508
rect 12236 31938 12292 31948
rect 12236 29652 12292 29662
rect 12236 26180 12292 29596
rect 12236 26114 12292 26124
rect 12236 23828 12292 23838
rect 12236 21924 12292 23772
rect 12236 21858 12292 21868
rect 12124 12964 12180 14812
rect 12236 18452 12292 18462
rect 12236 14532 12292 18396
rect 12236 14466 12292 14476
rect 12124 12898 12180 12908
rect 12012 5954 12068 5964
rect 12124 4900 12180 4910
rect 12124 4452 12180 4844
rect 12124 4386 12180 4396
rect 12348 1652 12404 48300
rect 12684 44578 12740 50428
rect 12796 48692 12852 54684
rect 12796 48626 12852 48636
rect 13020 47124 13076 47134
rect 12908 46676 12964 46686
rect 12908 46116 12964 46620
rect 12908 46050 12964 46060
rect 12684 44522 12852 44578
rect 12684 43764 12740 43774
rect 12460 42644 12516 42654
rect 12460 40740 12516 42588
rect 12460 40674 12516 40684
rect 12572 42420 12628 42430
rect 12460 40292 12516 40302
rect 12460 39060 12516 40236
rect 12572 39508 12628 42364
rect 12572 39442 12628 39452
rect 12460 38994 12516 39004
rect 12684 38388 12740 43708
rect 12684 37716 12740 38332
rect 12684 37650 12740 37660
rect 12460 34244 12516 34254
rect 12460 30324 12516 34188
rect 12460 29278 12516 30268
rect 12684 30324 12740 30334
rect 12460 29222 12628 29278
rect 12460 28756 12516 29222
rect 12572 29204 12628 29222
rect 12572 29138 12628 29148
rect 12460 26852 12516 28700
rect 12460 26786 12516 26796
rect 12572 28644 12628 28654
rect 12460 21924 12516 21934
rect 12460 18004 12516 21868
rect 12460 17938 12516 17948
rect 12572 14644 12628 28588
rect 12684 23940 12740 30268
rect 12796 30212 12852 44522
rect 12908 43764 12964 43774
rect 12908 31780 12964 43708
rect 13020 42196 13076 47068
rect 13020 42130 13076 42140
rect 13020 40292 13076 40302
rect 13020 39844 13076 40236
rect 13020 39778 13076 39788
rect 12908 31714 12964 31724
rect 13020 39508 13076 39518
rect 12796 30146 12852 30156
rect 12908 29092 12964 29102
rect 12796 27860 12852 27870
rect 12796 27188 12852 27804
rect 12796 27122 12852 27132
rect 12684 23874 12740 23884
rect 12908 24724 12964 29036
rect 12908 22438 12964 24668
rect 12572 14578 12628 14588
rect 12684 22382 12964 22438
rect 12684 5124 12740 22382
rect 12796 21252 12852 21262
rect 12796 17780 12852 21196
rect 12796 17714 12852 17724
rect 12908 18228 12964 18238
rect 12908 13188 12964 18172
rect 12908 13122 12964 13132
rect 12684 5058 12740 5068
rect 12908 10724 12964 10734
rect 12348 1586 12404 1596
rect 12908 1988 12964 10668
rect 13020 9604 13076 39452
rect 13132 39284 13188 55020
rect 13356 54628 13412 55692
rect 14812 55636 14868 55646
rect 14812 55300 14868 55580
rect 14812 55234 14868 55244
rect 15596 55300 15652 55310
rect 15596 55198 15652 55244
rect 15372 55142 15652 55198
rect 13356 54562 13412 54572
rect 13468 55076 13524 55086
rect 13132 39218 13188 39228
rect 13244 53172 13300 53182
rect 13132 38836 13188 38846
rect 13132 38052 13188 38780
rect 13132 36820 13188 37996
rect 13132 36754 13188 36764
rect 13132 30884 13188 30894
rect 13132 26740 13188 30828
rect 13244 30212 13300 53116
rect 13468 48020 13524 55020
rect 15372 55076 15428 55142
rect 15372 55010 15428 55020
rect 14476 54292 14532 54302
rect 14028 54180 14084 54190
rect 13804 53732 13860 53742
rect 13580 53060 13636 53070
rect 13580 51716 13636 53004
rect 13580 51650 13636 51660
rect 13468 47954 13524 47964
rect 13580 49588 13636 49598
rect 13468 47796 13524 47806
rect 13356 44436 13412 44446
rect 13356 42868 13412 44380
rect 13468 44324 13524 47740
rect 13580 44660 13636 49532
rect 13580 44594 13636 44604
rect 13692 48020 13748 48030
rect 13468 44258 13524 44268
rect 13356 42802 13412 42812
rect 13468 43652 13524 43662
rect 13468 41188 13524 43596
rect 13580 42084 13636 42094
rect 13580 41300 13636 42028
rect 13580 41234 13636 41244
rect 13468 41122 13524 41132
rect 13356 39508 13412 39518
rect 13356 33908 13412 39452
rect 13580 36708 13636 36718
rect 13580 36148 13636 36652
rect 13580 36082 13636 36092
rect 13356 33842 13412 33852
rect 13580 35028 13636 35038
rect 13244 30146 13300 30156
rect 13468 33348 13524 33358
rect 13132 26674 13188 26684
rect 13356 28084 13412 28094
rect 13356 25858 13412 28028
rect 13244 25844 13412 25858
rect 13300 25802 13412 25844
rect 13244 25778 13300 25788
rect 13132 24388 13188 24398
rect 13132 16212 13188 24332
rect 13132 16146 13188 16156
rect 13244 16772 13300 16782
rect 13020 3780 13076 9548
rect 13020 3714 13076 3724
rect 13020 2884 13076 2894
rect 13020 2548 13076 2828
rect 13020 2482 13076 2492
rect 11900 690 11956 700
rect 12908 196 12964 1932
rect 13244 1652 13300 16716
rect 13356 8596 13412 8606
rect 13356 6244 13412 8540
rect 13356 6178 13412 6188
rect 13468 8372 13524 33292
rect 13580 20020 13636 34972
rect 13692 34132 13748 47964
rect 13804 46564 13860 53676
rect 13804 41300 13860 46508
rect 13804 41234 13860 41244
rect 13916 45220 13972 45230
rect 13692 32340 13748 34076
rect 13916 33572 13972 45164
rect 13916 33506 13972 33516
rect 13692 32274 13748 32284
rect 13916 32564 13972 32574
rect 13804 30212 13860 30222
rect 13692 29092 13748 29102
rect 13692 25396 13748 29036
rect 13692 25330 13748 25340
rect 13804 21700 13860 30156
rect 13916 25620 13972 32508
rect 13916 25554 13972 25564
rect 13804 21634 13860 21644
rect 13916 21812 13972 21822
rect 13580 19796 13636 19964
rect 13580 19730 13636 19740
rect 13804 20916 13860 20926
rect 13580 19012 13636 19022
rect 13580 13972 13636 18956
rect 13580 13906 13636 13916
rect 13692 16548 13748 16558
rect 13468 7700 13524 8316
rect 13468 4900 13524 7644
rect 13580 11620 13636 11630
rect 13580 7476 13636 11564
rect 13580 7410 13636 7420
rect 13468 4834 13524 4844
rect 13244 1586 13300 1596
rect 13020 1316 13076 1326
rect 13020 420 13076 1260
rect 13692 868 13748 16492
rect 13804 13076 13860 20860
rect 13916 17668 13972 21756
rect 13916 17602 13972 17612
rect 13804 13010 13860 13020
rect 13916 16660 13972 16670
rect 13804 9492 13860 9502
rect 13804 3108 13860 9436
rect 13804 3042 13860 3052
rect 13916 980 13972 16604
rect 14028 4452 14084 54124
rect 14252 53732 14308 53742
rect 14252 53284 14308 53676
rect 14252 53218 14308 53228
rect 14252 52164 14308 52174
rect 14252 51828 14308 52108
rect 14252 51762 14308 51772
rect 14252 47012 14308 47022
rect 14252 46676 14308 46956
rect 14252 46610 14308 46620
rect 14252 46116 14308 46126
rect 14140 40964 14196 40974
rect 14140 39508 14196 40908
rect 14140 39442 14196 39452
rect 14252 39358 14308 46060
rect 14140 39302 14308 39358
rect 14364 41300 14420 41310
rect 14140 32340 14196 39302
rect 14252 38164 14308 38174
rect 14252 34468 14308 38108
rect 14364 35588 14420 41244
rect 14364 35522 14420 35532
rect 14252 34402 14308 34412
rect 14252 34132 14308 34142
rect 14252 33796 14308 34076
rect 14252 33730 14308 33740
rect 14140 32274 14196 32284
rect 14252 31444 14308 31454
rect 14252 30212 14308 31388
rect 14364 30996 14420 31006
rect 14364 30772 14420 30940
rect 14364 30706 14420 30716
rect 14252 30146 14308 30156
rect 14364 28420 14420 28430
rect 14140 27636 14196 27646
rect 14140 26628 14196 27580
rect 14364 27636 14420 28364
rect 14364 27570 14420 27580
rect 14140 26562 14196 26572
rect 14364 26964 14420 26974
rect 14140 22708 14196 22718
rect 14140 20244 14196 22652
rect 14140 20178 14196 20188
rect 14252 21812 14308 21822
rect 14252 20580 14308 21756
rect 14252 19236 14308 20524
rect 14252 19170 14308 19180
rect 14252 19012 14308 19022
rect 14252 18788 14308 18956
rect 14252 18722 14308 18732
rect 14252 18340 14308 18350
rect 14140 16772 14196 16782
rect 14140 14868 14196 16716
rect 14140 14802 14196 14812
rect 14028 4386 14084 4396
rect 14140 12180 14196 12190
rect 14140 3668 14196 12124
rect 14140 3602 14196 3612
rect 14028 3482 14196 3538
rect 14028 3444 14084 3482
rect 14028 3378 14084 3388
rect 14140 3332 14196 3482
rect 14140 3266 14196 3276
rect 14252 1652 14308 18284
rect 14364 9268 14420 26908
rect 14476 16436 14532 54236
rect 15148 54292 15204 54302
rect 14924 52164 14980 52174
rect 14924 51828 14980 52108
rect 14924 51762 14980 51772
rect 15036 51268 15092 51278
rect 15036 50708 15092 51212
rect 15036 50642 15092 50652
rect 14588 49252 14644 49262
rect 14588 46788 14644 49196
rect 15036 49028 15092 49038
rect 15036 47796 15092 48972
rect 14588 46722 14644 46732
rect 14812 47012 14868 47022
rect 14588 46452 14644 46462
rect 14588 42238 14644 46396
rect 14812 46116 14868 46956
rect 15036 46788 15092 47740
rect 14812 46050 14868 46060
rect 14924 46564 14980 46574
rect 14924 46004 14980 46508
rect 14924 45938 14980 45948
rect 14700 45108 14756 45118
rect 14700 42420 14756 45052
rect 14700 42354 14756 42364
rect 14588 42182 14756 42238
rect 14588 39732 14644 39742
rect 14588 38724 14644 39676
rect 14588 38658 14644 38668
rect 14588 38500 14644 38510
rect 14588 37828 14644 38444
rect 14700 38052 14756 42182
rect 14700 37986 14756 37996
rect 14812 42196 14868 42206
rect 14588 37762 14644 37772
rect 14812 34804 14868 42140
rect 14812 34738 14868 34748
rect 14924 36596 14980 36606
rect 14588 34132 14644 34142
rect 14588 27860 14644 34076
rect 14588 27794 14644 27804
rect 14700 32340 14756 32350
rect 14476 16370 14532 16380
rect 14588 24388 14644 24398
rect 14476 13076 14532 13086
rect 14476 11956 14532 13020
rect 14476 11890 14532 11900
rect 14364 9202 14420 9212
rect 14476 8484 14532 8494
rect 14364 7812 14420 7822
rect 14364 7252 14420 7756
rect 14364 7186 14420 7196
rect 14476 5236 14532 8428
rect 14476 5170 14532 5180
rect 14588 4900 14644 24332
rect 14700 18004 14756 32284
rect 14924 26852 14980 36540
rect 14924 26786 14980 26796
rect 14924 21476 14980 21486
rect 14700 13748 14756 17948
rect 14700 13682 14756 13692
rect 14812 18452 14868 18462
rect 14700 11620 14756 11630
rect 14700 10052 14756 11564
rect 14700 9986 14756 9996
rect 14700 8148 14756 8158
rect 14700 5572 14756 8092
rect 14700 5506 14756 5516
rect 14588 4834 14644 4844
rect 14252 1586 14308 1596
rect 14812 1652 14868 18396
rect 14924 13300 14980 21420
rect 15036 18452 15092 46732
rect 15036 18386 15092 18396
rect 14924 13234 14980 13244
rect 15036 14756 15092 14766
rect 14924 12516 14980 12526
rect 14924 8938 14980 12460
rect 15036 11060 15092 14700
rect 15036 10994 15092 11004
rect 14924 8882 15092 8938
rect 15036 7588 15092 8882
rect 15036 7522 15092 7532
rect 14924 7364 14980 7374
rect 14924 5572 14980 7308
rect 14924 5506 14980 5516
rect 14812 1586 14868 1596
rect 15036 1988 15092 1998
rect 15036 1540 15092 1932
rect 15036 1474 15092 1484
rect 13916 914 13972 924
rect 13692 802 13748 812
rect 13020 354 13076 364
rect 15148 420 15204 54236
rect 15372 54292 15428 54302
rect 15260 50596 15316 50606
rect 15260 22484 15316 50540
rect 15372 38612 15428 54236
rect 15596 53172 15652 53182
rect 15596 52678 15652 53116
rect 16268 52948 16324 52958
rect 16268 52858 16324 52892
rect 15708 52836 16324 52858
rect 15764 52802 16324 52836
rect 15708 52770 15764 52780
rect 15596 52622 15988 52678
rect 15484 51380 15540 51390
rect 15484 49140 15540 51324
rect 15484 49074 15540 49084
rect 15372 38546 15428 38556
rect 15484 48692 15540 48702
rect 15372 38388 15428 38398
rect 15372 36148 15428 38332
rect 15372 36082 15428 36092
rect 15372 34244 15428 34254
rect 15372 33796 15428 34188
rect 15372 33730 15428 33740
rect 15260 15876 15316 22428
rect 15260 15810 15316 15820
rect 15372 23492 15428 23502
rect 15372 15204 15428 23436
rect 15372 15138 15428 15148
rect 15372 14868 15428 14878
rect 15372 13636 15428 14812
rect 15372 13570 15428 13580
rect 15372 12404 15428 12414
rect 15372 11844 15428 12348
rect 15372 11778 15428 11788
rect 15372 11620 15428 11630
rect 15260 10836 15316 10846
rect 15260 9492 15316 10780
rect 15260 9426 15316 9436
rect 15372 8038 15428 11564
rect 15260 7982 15428 8038
rect 15260 5236 15316 7982
rect 15372 7812 15428 7822
rect 15372 6692 15428 7756
rect 15372 6626 15428 6636
rect 15260 5170 15316 5180
rect 15484 756 15540 48636
rect 15932 46452 15988 52622
rect 16380 52612 16436 52622
rect 15932 46386 15988 46396
rect 16044 49028 16100 49038
rect 16044 45108 16100 48972
rect 16044 45042 16100 45052
rect 16268 44996 16324 45006
rect 15820 43540 15876 43550
rect 15820 42420 15876 43484
rect 15820 42354 15876 42364
rect 16268 40740 16324 44940
rect 16268 40674 16324 40684
rect 15932 39284 15988 39294
rect 15596 38612 15652 38622
rect 15596 34692 15652 38556
rect 15596 34626 15652 34636
rect 15708 37044 15764 37054
rect 15596 33796 15652 33806
rect 15596 25956 15652 33740
rect 15708 32788 15764 36988
rect 15708 32722 15764 32732
rect 15820 29988 15876 29998
rect 15820 29540 15876 29932
rect 15820 29474 15876 29484
rect 15596 25890 15652 25900
rect 15820 26628 15876 26638
rect 15596 19908 15652 19918
rect 15596 11844 15652 19852
rect 15596 11778 15652 11788
rect 15596 11620 15652 11630
rect 15596 10388 15652 11564
rect 15596 10322 15652 10332
rect 15708 10612 15764 10622
rect 15708 10198 15764 10556
rect 15596 10142 15764 10198
rect 15820 10388 15876 26572
rect 15596 9044 15652 10142
rect 15820 9492 15876 10332
rect 15820 9426 15876 9436
rect 15596 8978 15652 8988
rect 15596 6580 15652 6590
rect 15596 5908 15652 6524
rect 15596 5842 15652 5852
rect 15820 5908 15876 5918
rect 15820 5124 15876 5852
rect 15820 5058 15876 5068
rect 15932 1652 15988 39228
rect 16156 34468 16212 34478
rect 16156 26964 16212 34412
rect 16156 26898 16212 26908
rect 16268 32564 16324 32574
rect 16268 26516 16324 32508
rect 16156 22708 16212 22718
rect 16044 18116 16100 18126
rect 16044 7812 16100 18060
rect 16156 17892 16212 22652
rect 16156 13524 16212 17836
rect 16156 13458 16212 13468
rect 16268 11998 16324 26460
rect 16156 11942 16324 11998
rect 16156 11620 16212 11942
rect 16156 11554 16212 11564
rect 16268 10836 16324 10846
rect 16268 9604 16324 10780
rect 16268 9538 16324 9548
rect 16044 7746 16100 7756
rect 15932 1586 15988 1596
rect 16380 1652 16436 52556
rect 16492 49700 16548 56924
rect 19740 55300 19796 55310
rect 18284 55076 18340 55086
rect 18284 55018 18340 55020
rect 18284 54962 18452 55018
rect 17724 53172 17780 53182
rect 17724 52948 17780 53116
rect 17724 52882 17780 52892
rect 16716 52622 17108 52678
rect 16716 52388 16772 52622
rect 16716 52322 16772 52332
rect 16940 52388 16996 52398
rect 16940 51058 16996 52332
rect 17052 52276 17108 52622
rect 17052 52210 17108 52220
rect 18172 52612 18228 52622
rect 16828 51002 16996 51058
rect 16828 50260 16884 51002
rect 16828 50194 16884 50204
rect 16492 49634 16548 49644
rect 16940 49812 16996 49822
rect 16492 48692 16548 48702
rect 16492 47348 16548 48636
rect 16492 33460 16548 47292
rect 16828 48132 16884 48142
rect 16828 46340 16884 48076
rect 16828 46274 16884 46284
rect 16940 44436 16996 49756
rect 16940 43540 16996 44380
rect 16940 43474 16996 43484
rect 17052 49700 17108 49710
rect 17052 49140 17108 49644
rect 16716 42980 16772 42990
rect 16492 33394 16548 33404
rect 16604 40292 16660 40302
rect 16492 23044 16548 23054
rect 16492 22708 16548 22988
rect 16492 22642 16548 22652
rect 16604 17332 16660 40236
rect 16716 39732 16772 42924
rect 16716 39666 16772 39676
rect 16828 40964 16884 40974
rect 16828 33796 16884 40908
rect 16828 33730 16884 33740
rect 16940 40404 16996 40414
rect 16940 32788 16996 40348
rect 17052 34132 17108 49084
rect 18172 49588 18228 52556
rect 17500 48580 17556 48590
rect 17164 47572 17220 47582
rect 17164 42980 17220 47516
rect 17164 42914 17220 42924
rect 17276 46452 17332 46462
rect 17276 42778 17332 46396
rect 17500 46378 17556 48524
rect 18060 47684 18116 47694
rect 17500 46322 17668 46378
rect 17052 34066 17108 34076
rect 17164 42722 17332 42778
rect 17500 46228 17556 46238
rect 16940 32722 16996 32732
rect 16828 32564 16884 32574
rect 16604 17266 16660 17276
rect 16716 31892 16772 31902
rect 16604 16772 16660 16782
rect 16604 13300 16660 16716
rect 16604 13234 16660 13244
rect 16604 11732 16660 11742
rect 16492 11508 16548 11518
rect 16492 9492 16548 11452
rect 16604 10836 16660 11676
rect 16604 10770 16660 10780
rect 16492 9426 16548 9436
rect 16716 9298 16772 31836
rect 16828 12852 16884 32508
rect 16940 30996 16996 31006
rect 16940 23338 16996 30940
rect 17052 28196 17108 28206
rect 17052 27300 17108 28140
rect 17052 27234 17108 27244
rect 16940 23282 17108 23338
rect 16940 23156 16996 23166
rect 16940 21252 16996 23100
rect 16940 21186 16996 21196
rect 17052 18340 17108 23282
rect 17164 18452 17220 42722
rect 17500 40078 17556 46172
rect 17612 45220 17668 46322
rect 17612 45154 17668 45164
rect 17276 40022 17556 40078
rect 17612 42868 17668 42878
rect 17276 23940 17332 40022
rect 17388 36932 17444 36942
rect 17388 35700 17444 36876
rect 17388 35634 17444 35644
rect 17612 35588 17668 42812
rect 17612 35522 17668 35532
rect 17724 37268 17780 37278
rect 17724 35028 17780 37212
rect 17388 34020 17444 34030
rect 17388 33348 17444 33964
rect 17388 33282 17444 33292
rect 17388 32452 17444 32462
rect 17388 27636 17444 32396
rect 17500 32116 17556 32126
rect 17500 30996 17556 32060
rect 17500 30930 17556 30940
rect 17388 27570 17444 27580
rect 17500 27972 17556 27982
rect 17276 23874 17332 23884
rect 17276 23492 17332 23502
rect 17276 22372 17332 23436
rect 17276 22306 17332 22316
rect 17500 20998 17556 27916
rect 17612 26740 17668 26750
rect 17612 24388 17668 26684
rect 17612 24322 17668 24332
rect 17164 18386 17220 18396
rect 17388 20942 17556 20998
rect 17612 23940 17668 23950
rect 17052 18274 17108 18284
rect 17164 17780 17220 17790
rect 17164 14980 17220 17724
rect 17164 14914 17220 14924
rect 16828 12786 16884 12796
rect 17276 12852 17332 12862
rect 16604 9242 16772 9298
rect 16940 9380 16996 9390
rect 16492 7588 16548 7598
rect 16492 6244 16548 7532
rect 16492 6178 16548 6188
rect 16380 1586 16436 1596
rect 16380 1428 16436 1438
rect 16380 1092 16436 1372
rect 16604 1428 16660 9242
rect 16828 8260 16884 8270
rect 16828 7812 16884 8204
rect 16828 1652 16884 7756
rect 16940 6580 16996 9324
rect 16940 6514 16996 6524
rect 16828 1586 16884 1596
rect 17276 1652 17332 12796
rect 17388 8260 17444 20942
rect 17612 20818 17668 23884
rect 17500 20762 17668 20818
rect 17500 9604 17556 20762
rect 17724 14420 17780 34972
rect 17836 31780 17892 31790
rect 17836 29428 17892 31724
rect 17836 24500 17892 29372
rect 18060 30100 18116 47628
rect 18172 46452 18228 49532
rect 18172 46386 18228 46396
rect 18172 44548 18228 44558
rect 18172 40292 18228 44492
rect 18172 38724 18228 40236
rect 18172 38658 18228 38668
rect 18284 34244 18340 34254
rect 18284 32676 18340 34188
rect 18284 32610 18340 32620
rect 17836 24434 17892 24444
rect 17948 26180 18004 26190
rect 17948 23604 18004 26124
rect 17948 23538 18004 23548
rect 17948 20916 18004 20926
rect 17612 13748 17668 13758
rect 17612 12068 17668 13692
rect 17612 12002 17668 12012
rect 17500 9538 17556 9548
rect 17388 8194 17444 8204
rect 17724 6132 17780 14364
rect 17836 14532 17892 14542
rect 17836 12404 17892 14476
rect 17836 12338 17892 12348
rect 17948 13636 18004 20860
rect 18060 18452 18116 30044
rect 18284 31780 18340 31790
rect 18284 22798 18340 31724
rect 18060 18386 18116 18396
rect 18172 22742 18340 22798
rect 18172 21140 18228 22742
rect 17948 12292 18004 13580
rect 17948 12226 18004 12236
rect 18060 13300 18116 13310
rect 17836 11620 17892 11630
rect 17836 9492 17892 11564
rect 17836 9426 17892 9436
rect 17724 6066 17780 6076
rect 18060 8596 18116 13244
rect 18060 8260 18116 8540
rect 18060 4676 18116 8204
rect 18060 4610 18116 4620
rect 17276 1586 17332 1596
rect 18172 1652 18228 21084
rect 18284 20580 18340 20590
rect 18284 20244 18340 20524
rect 18284 20178 18340 20188
rect 18284 19684 18340 19694
rect 18284 18788 18340 19628
rect 18284 18722 18340 18732
rect 18284 6692 18340 6702
rect 18284 2548 18340 6636
rect 18396 5572 18452 54962
rect 18620 54404 18676 54414
rect 18508 49476 18564 49486
rect 18508 47236 18564 49420
rect 18508 47170 18564 47180
rect 18620 44996 18676 54348
rect 18620 44930 18676 44940
rect 18732 54068 18788 54078
rect 18508 43988 18564 43998
rect 18508 41748 18564 43932
rect 18508 41682 18564 41692
rect 18508 33124 18564 33134
rect 18508 29428 18564 33068
rect 18508 29362 18564 29372
rect 18508 24052 18564 24062
rect 18508 16212 18564 23996
rect 18732 23828 18788 54012
rect 19628 52724 19684 52734
rect 19180 52164 19236 52174
rect 18844 49812 18900 49822
rect 18844 31618 18900 49756
rect 18956 49588 19012 49598
rect 18956 44660 19012 49532
rect 19180 48916 19236 52108
rect 19180 48850 19236 48860
rect 18956 44594 19012 44604
rect 19180 48020 19236 48030
rect 18956 42532 19012 42542
rect 18956 38164 19012 42476
rect 18956 38098 19012 38108
rect 18956 33796 19012 33806
rect 18956 32788 19012 33740
rect 18956 32722 19012 32732
rect 18844 31562 19124 31618
rect 19068 29540 19124 31562
rect 18732 23762 18788 23772
rect 18844 29428 18900 29438
rect 18732 23492 18788 23502
rect 18732 21812 18788 23436
rect 18732 21746 18788 21756
rect 18620 21364 18676 21374
rect 18620 20916 18676 21308
rect 18620 20850 18676 20860
rect 18508 16138 18564 16156
rect 18508 16082 18676 16138
rect 18396 5506 18452 5516
rect 18508 11172 18564 11182
rect 18508 4452 18564 11116
rect 18508 2772 18564 4396
rect 18508 2706 18564 2716
rect 18620 8596 18676 16082
rect 18284 2100 18340 2492
rect 18284 2034 18340 2044
rect 18620 1764 18676 8540
rect 18844 8398 18900 29372
rect 18956 28532 19012 28542
rect 18956 26516 19012 28476
rect 18956 26450 19012 26460
rect 18956 23156 19012 23166
rect 18956 14532 19012 23100
rect 19068 19236 19124 29484
rect 19068 19170 19124 19180
rect 18956 14308 19012 14476
rect 18956 14242 19012 14252
rect 18844 8342 19012 8398
rect 18732 6468 18788 6478
rect 18732 5012 18788 6412
rect 18956 6356 19012 8342
rect 18956 5124 19012 6300
rect 19068 5796 19124 5806
rect 19068 5348 19124 5740
rect 19068 5282 19124 5292
rect 18956 5058 19012 5068
rect 18732 4946 18788 4956
rect 18620 1698 18676 1708
rect 19180 2660 19236 47964
rect 19292 43316 19348 43326
rect 19292 41412 19348 43260
rect 19292 41346 19348 41356
rect 19516 41972 19572 41982
rect 19404 25508 19460 25518
rect 19292 22932 19348 22942
rect 19292 22484 19348 22876
rect 19292 22418 19348 22428
rect 19292 15652 19348 15662
rect 19292 15316 19348 15596
rect 19292 15250 19348 15260
rect 19404 9940 19460 25452
rect 19404 9874 19460 9884
rect 19516 24724 19572 41916
rect 19180 1764 19236 2604
rect 19516 2212 19572 24668
rect 19628 21476 19684 52668
rect 19740 50148 19796 55244
rect 20636 54852 20692 54862
rect 19964 54068 20020 54078
rect 19740 50082 19796 50092
rect 19852 53172 19908 53182
rect 19852 52724 19908 53116
rect 19852 49252 19908 52668
rect 19852 49186 19908 49196
rect 19964 52612 20020 54012
rect 20188 54068 20244 54078
rect 20188 53620 20244 54012
rect 20188 53554 20244 53564
rect 19852 48468 19908 48478
rect 19852 43540 19908 48412
rect 19852 43474 19908 43484
rect 19852 40292 19908 40302
rect 19740 35588 19796 35598
rect 19740 34468 19796 35532
rect 19740 25508 19796 34412
rect 19740 25442 19796 25452
rect 19852 24948 19908 40236
rect 19852 24882 19908 24892
rect 19740 23380 19796 23390
rect 19740 22820 19796 23324
rect 19740 22754 19796 22764
rect 19628 21410 19684 21420
rect 19852 8708 19908 8718
rect 19852 8148 19908 8652
rect 19852 8082 19908 8092
rect 19740 6580 19796 6590
rect 19740 6418 19796 6524
rect 19628 6362 19796 6418
rect 19628 3668 19684 6362
rect 19964 3898 20020 52556
rect 20300 53396 20356 53406
rect 20076 48020 20132 48030
rect 20076 43764 20132 47964
rect 20076 42868 20132 43708
rect 20076 42802 20132 42812
rect 20300 42420 20356 53340
rect 20300 42354 20356 42364
rect 20636 47460 20692 54796
rect 20860 54180 20916 54190
rect 20860 50260 20916 54124
rect 21084 53620 21140 53630
rect 20860 50194 20916 50204
rect 20972 52052 21028 52062
rect 20636 37198 20692 47404
rect 20524 37142 20692 37198
rect 20748 48916 20804 48926
rect 20188 31108 20244 31118
rect 20188 30100 20244 31052
rect 20076 29988 20132 29998
rect 20076 29764 20132 29932
rect 20076 27524 20132 29708
rect 20076 27458 20132 27468
rect 20076 26404 20132 26414
rect 20076 24276 20132 26348
rect 20076 24210 20132 24220
rect 20076 21252 20132 21262
rect 20076 19572 20132 21196
rect 20076 19506 20132 19516
rect 20188 16548 20244 30044
rect 20524 28084 20580 37142
rect 20636 35140 20692 35150
rect 20636 32900 20692 35084
rect 20636 32834 20692 32844
rect 20524 28018 20580 28028
rect 20412 27972 20468 27982
rect 20412 23716 20468 27916
rect 20748 25956 20804 48860
rect 20972 48580 21028 51996
rect 20972 48244 21028 48524
rect 20972 48178 21028 48188
rect 20860 44324 20916 44334
rect 20860 40438 20916 44268
rect 20972 44100 21028 44110
rect 20972 43204 21028 44044
rect 20972 43138 21028 43148
rect 20972 42644 21028 42654
rect 20972 40628 21028 42588
rect 20972 40562 21028 40572
rect 20860 40382 21028 40438
rect 20972 38388 21028 40382
rect 20748 25858 20804 25900
rect 20412 23650 20468 23660
rect 20524 25802 20804 25858
rect 20860 36484 20916 36494
rect 20300 23156 20356 23166
rect 20300 21252 20356 23100
rect 20300 21186 20356 21196
rect 20412 21476 20468 21486
rect 20188 16482 20244 16492
rect 19628 3602 19684 3612
rect 19852 3842 20020 3898
rect 20076 6804 20132 6814
rect 20076 3898 20132 6748
rect 20300 4676 20356 4686
rect 20188 3898 20244 3902
rect 20076 3892 20244 3898
rect 20076 3842 20188 3892
rect 19852 3538 19908 3842
rect 20188 3826 20244 3836
rect 20300 3538 20356 4620
rect 19852 3482 20020 3538
rect 19516 2146 19572 2156
rect 19180 1698 19236 1708
rect 18172 1586 18228 1596
rect 19964 1540 20020 3482
rect 20076 3482 20356 3538
rect 20076 2212 20132 3482
rect 20076 2146 20132 2156
rect 20412 1652 20468 21420
rect 20524 5124 20580 25802
rect 20524 5058 20580 5068
rect 20636 23828 20692 23838
rect 20412 1586 20468 1596
rect 19964 1474 20020 1484
rect 16604 1362 16660 1372
rect 16380 1026 16436 1036
rect 15484 690 15540 700
rect 20636 756 20692 23772
rect 20748 23156 20804 23166
rect 20748 21252 20804 23100
rect 20748 21186 20804 21196
rect 20860 13748 20916 36428
rect 20972 23828 21028 38332
rect 20972 23762 21028 23772
rect 20972 23268 21028 23278
rect 20972 20468 21028 23212
rect 20972 20402 21028 20412
rect 20972 16436 21028 16446
rect 20972 16100 21028 16380
rect 20972 16034 21028 16044
rect 20860 13682 20916 13692
rect 20972 9380 21028 9390
rect 20748 9268 20804 9278
rect 20748 1652 20804 9212
rect 20972 4564 21028 9324
rect 21084 5908 21140 53564
rect 21196 46004 21252 46014
rect 21196 45668 21252 45948
rect 21196 45602 21252 45612
rect 21196 45108 21252 45118
rect 21196 44660 21252 45052
rect 21196 44594 21252 44604
rect 21308 43988 21364 57036
rect 21980 55972 22036 55982
rect 21644 55300 21700 55310
rect 21532 52164 21588 52174
rect 21308 43922 21364 43932
rect 21420 48020 21476 48030
rect 21420 43858 21476 47964
rect 21196 43802 21476 43858
rect 21532 46004 21588 52108
rect 21196 32004 21252 43802
rect 21308 42420 21364 42430
rect 21308 32452 21364 42364
rect 21532 35038 21588 45948
rect 21420 34982 21588 35038
rect 21420 34580 21476 34982
rect 21420 34514 21476 34524
rect 21532 34804 21588 34814
rect 21308 32386 21364 32396
rect 21420 33460 21476 33470
rect 21196 31938 21252 31948
rect 21308 30548 21364 30558
rect 21196 28532 21252 28542
rect 21196 9828 21252 28476
rect 21308 22708 21364 30492
rect 21308 22642 21364 22652
rect 21420 19236 21476 33404
rect 21532 30436 21588 34748
rect 21532 30370 21588 30380
rect 21532 28532 21588 28542
rect 21532 27972 21588 28476
rect 21532 27906 21588 27916
rect 21532 24612 21588 24622
rect 21532 23716 21588 24556
rect 21532 23650 21588 23660
rect 21532 22932 21588 22942
rect 21532 22148 21588 22876
rect 21532 22082 21588 22092
rect 21420 19170 21476 19180
rect 21532 21812 21588 21822
rect 21308 18340 21364 18350
rect 21308 16996 21364 18284
rect 21308 16930 21364 16940
rect 21196 9762 21252 9772
rect 21308 15988 21364 15998
rect 21308 15540 21364 15932
rect 21308 8484 21364 15484
rect 21532 14196 21588 21756
rect 21532 12964 21588 14140
rect 21532 12898 21588 12908
rect 21308 8418 21364 8428
rect 21196 8372 21252 8382
rect 21196 7476 21252 8316
rect 21196 7410 21252 7420
rect 21084 5842 21140 5852
rect 20972 4498 21028 4508
rect 21084 4452 21140 4462
rect 21084 3444 21140 4396
rect 21084 3378 21140 3388
rect 20748 1586 20804 1596
rect 21644 980 21700 55244
rect 21980 48356 22036 55916
rect 22540 55300 22596 55310
rect 21980 48290 22036 48300
rect 22092 53732 22148 53742
rect 21980 46564 22036 46574
rect 21980 45220 22036 46508
rect 22092 45892 22148 53676
rect 22316 52724 22372 52734
rect 22204 49140 22260 49150
rect 22204 48916 22260 49084
rect 22204 48850 22260 48860
rect 22092 45826 22148 45836
rect 21868 32788 21924 32798
rect 21756 28084 21812 28094
rect 21756 9268 21812 28028
rect 21868 27972 21924 32732
rect 21868 27906 21924 27916
rect 21868 26292 21924 26302
rect 21868 25844 21924 26236
rect 21868 25778 21924 25788
rect 21868 24612 21924 24622
rect 21868 24388 21924 24556
rect 21868 24322 21924 24332
rect 21868 23716 21924 23726
rect 21868 23268 21924 23660
rect 21868 23202 21924 23212
rect 21980 12068 22036 45164
rect 22204 44884 22260 44894
rect 22204 36820 22260 44828
rect 22316 40964 22372 52668
rect 22316 40898 22372 40908
rect 22428 49588 22484 49598
rect 22316 40740 22372 40750
rect 22316 39956 22372 40684
rect 22316 39890 22372 39900
rect 22204 36754 22260 36764
rect 22428 36478 22484 49532
rect 22540 45220 22596 55244
rect 22540 45154 22596 45164
rect 22652 50260 22708 50270
rect 22092 36422 22484 36478
rect 22540 44996 22596 45006
rect 22092 29316 22148 36422
rect 22540 36298 22596 44940
rect 22092 29250 22148 29260
rect 22316 36242 22596 36298
rect 22316 28644 22372 36242
rect 22428 36036 22484 36046
rect 22428 35028 22484 35980
rect 22428 34962 22484 34972
rect 22316 28578 22372 28588
rect 22540 28644 22596 28654
rect 22204 27748 22260 27758
rect 22092 27412 22148 27422
rect 22092 24948 22148 27356
rect 22092 24882 22148 24892
rect 21980 12002 22036 12012
rect 22092 24388 22148 24398
rect 22092 9940 22148 24332
rect 22092 9874 22148 9884
rect 21756 9202 21812 9212
rect 22204 7588 22260 27692
rect 22316 27188 22372 27198
rect 22316 26964 22372 27132
rect 22316 26898 22372 26908
rect 22428 25844 22484 25854
rect 22316 24948 22372 24958
rect 22316 23940 22372 24892
rect 22428 24276 22484 25788
rect 22428 24210 22484 24220
rect 22316 23874 22372 23884
rect 22540 23518 22596 28588
rect 22316 23462 22596 23518
rect 22316 22820 22372 23462
rect 22316 22754 22372 22764
rect 22428 23380 22484 23390
rect 22428 21812 22484 23324
rect 22540 22932 22596 22942
rect 22540 22148 22596 22876
rect 22540 22082 22596 22092
rect 22428 21746 22484 21756
rect 22428 17668 22484 17678
rect 22428 14980 22484 17612
rect 22428 13524 22484 14924
rect 22428 13458 22484 13468
rect 22428 11060 22484 11070
rect 22428 10724 22484 11004
rect 22428 10658 22484 10668
rect 22204 6804 22260 7532
rect 22204 6738 22260 6748
rect 21644 914 21700 924
rect 20636 690 20692 700
rect 22652 756 22708 50204
rect 22764 47124 22820 57148
rect 23776 56476 24096 57456
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23436 54292 23492 54302
rect 22764 47058 22820 47068
rect 22988 53732 23044 53742
rect 22764 46900 22820 46910
rect 22764 45668 22820 46844
rect 22764 45602 22820 45612
rect 22764 42308 22820 42318
rect 22764 40068 22820 42252
rect 22764 40002 22820 40012
rect 22876 41748 22932 41758
rect 22876 35476 22932 41692
rect 22876 35410 22932 35420
rect 22764 35252 22820 35262
rect 22764 10052 22820 35196
rect 22876 34132 22932 34142
rect 22876 33908 22932 34076
rect 22876 33842 22932 33852
rect 22988 33124 23044 53676
rect 23324 53508 23380 53518
rect 23100 51716 23156 51726
rect 23100 50372 23156 51660
rect 23100 50306 23156 50316
rect 23212 51156 23268 51166
rect 23212 49588 23268 51100
rect 23212 49522 23268 49532
rect 23212 46116 23268 46126
rect 22988 33058 23044 33068
rect 23100 45892 23156 45902
rect 23100 42756 23156 45836
rect 22876 32900 22932 32910
rect 22876 32116 22932 32844
rect 22876 32050 22932 32060
rect 23100 31780 23156 42700
rect 23212 41524 23268 46060
rect 23212 40516 23268 41468
rect 23212 40450 23268 40460
rect 23212 39732 23268 39742
rect 23212 33460 23268 39676
rect 23212 33394 23268 33404
rect 23100 31714 23156 31724
rect 23100 30996 23156 31006
rect 22988 30436 23044 30446
rect 22876 30100 22932 30110
rect 22876 25620 22932 30044
rect 22876 25554 22932 25564
rect 22876 23156 22932 23166
rect 22876 20468 22932 23100
rect 22988 22372 23044 30380
rect 23100 27860 23156 30940
rect 23100 27524 23156 27804
rect 23100 27458 23156 27468
rect 23212 27412 23268 27422
rect 23100 25844 23156 25854
rect 23100 23604 23156 25788
rect 23100 23538 23156 23548
rect 22988 21140 23044 22316
rect 23100 23380 23156 23390
rect 23100 21588 23156 23324
rect 23100 21522 23156 21532
rect 22988 21074 23044 21084
rect 22876 16324 22932 20412
rect 22876 16258 22932 16268
rect 23212 10164 23268 27356
rect 23212 10098 23268 10108
rect 22764 9986 22820 9996
rect 22876 9492 22932 9502
rect 22876 2212 22932 9436
rect 23100 8484 23156 8494
rect 23100 6132 23156 8428
rect 23324 8372 23380 53452
rect 23436 41076 23492 54236
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 24436 55692 24756 57456
rect 38444 57092 38500 57102
rect 27804 56868 27860 56878
rect 27132 56084 27188 56094
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 25900 55972 25956 55982
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 23776 51772 24096 53284
rect 24220 53284 24276 53294
rect 24220 52612 24276 53228
rect 24220 52546 24276 52556
rect 24436 52556 24756 54068
rect 25788 55524 25844 55534
rect 25564 53844 25620 53854
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 23660 51044 23716 51054
rect 23548 50932 23604 50942
rect 23548 48468 23604 50876
rect 23660 50260 23716 50988
rect 23660 50194 23716 50204
rect 23776 50204 24096 51716
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 25228 53620 25284 53630
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23548 48402 23604 48412
rect 23660 49812 23716 49822
rect 23436 41010 23492 41020
rect 23548 45220 23604 45230
rect 23436 37156 23492 37166
rect 23436 34468 23492 37100
rect 23436 34402 23492 34412
rect 23548 31668 23604 45164
rect 23660 35476 23716 49756
rect 23660 35410 23716 35420
rect 23776 48636 24096 50148
rect 24220 50596 24276 50606
rect 24220 50036 24276 50540
rect 24220 49970 24276 49980
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 24220 49588 24276 49598
rect 24220 48580 24276 49532
rect 24220 41972 24276 48524
rect 24220 41906 24276 41916
rect 24436 49420 24756 50932
rect 25004 52388 25060 52398
rect 25004 50596 25060 52332
rect 25004 50530 25060 50540
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 25228 49700 25284 53564
rect 25228 47638 25284 49644
rect 25340 50708 25396 50718
rect 25340 48468 25396 50652
rect 25340 48402 25396 48412
rect 25228 47582 25396 47638
rect 25116 46676 25172 46686
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 25004 46564 25060 46574
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 24220 41076 24276 41086
rect 24220 38388 24276 41020
rect 24220 38322 24276 38332
rect 24436 40012 24756 41524
rect 24892 45892 24948 45902
rect 24892 40292 24948 45836
rect 25004 43876 25060 46508
rect 25004 43810 25060 43820
rect 24892 40226 24948 40236
rect 25004 43540 25060 43550
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 24436 36876 24756 38388
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 23776 34524 24096 36036
rect 24220 36820 24276 36830
rect 24220 36036 24276 36764
rect 24220 35970 24276 35980
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 23660 34468 23716 34478
rect 23660 33124 23716 34412
rect 23660 33058 23716 33068
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23548 31602 23604 31612
rect 23660 32228 23716 32238
rect 23660 30996 23716 32172
rect 23660 30930 23716 30940
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23548 30660 23604 30670
rect 23548 28868 23604 30604
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 23436 25956 23492 25966
rect 23436 23492 23492 25900
rect 23436 23426 23492 23436
rect 23548 21476 23604 28812
rect 23660 28980 23716 28990
rect 23660 25620 23716 28924
rect 23660 25554 23716 25564
rect 23776 28252 24096 29764
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23548 21410 23604 21420
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 23548 20916 23604 20926
rect 23324 8306 23380 8316
rect 23436 20692 23492 20702
rect 23436 19908 23492 20636
rect 23100 6066 23156 6076
rect 22876 2146 22932 2156
rect 23324 3220 23380 3230
rect 23324 868 23380 3164
rect 23436 2660 23492 19852
rect 23548 13300 23604 20860
rect 23776 20412 24096 21924
rect 24220 35476 24276 35486
rect 24220 20916 24276 35420
rect 24220 20850 24276 20860
rect 24436 35308 24756 36820
rect 24892 37268 24948 37278
rect 24892 36820 24948 37212
rect 24892 36754 24948 36764
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24892 34468 24948 34478
rect 24892 34244 24948 34412
rect 24892 34178 24948 34188
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24892 34020 24948 34030
rect 24892 33796 24948 33964
rect 24892 33730 24948 33740
rect 24436 32172 24756 33684
rect 24892 32900 24948 32910
rect 24892 32564 24948 32844
rect 24892 32498 24948 32508
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24892 31444 24948 31454
rect 24892 30884 24948 31388
rect 24892 30818 24948 30828
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 24892 30324 24948 30334
rect 24892 27412 24948 30268
rect 24892 27346 24948 27356
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24892 26740 24948 26750
rect 24892 24836 24948 26684
rect 24892 24770 24948 24780
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 23660 20356 23716 20366
rect 23660 20020 23716 20300
rect 23660 19954 23716 19964
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23660 19348 23716 19358
rect 23660 15988 23716 19292
rect 23660 15922 23716 15932
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 24436 19628 24756 21140
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 23776 15708 24096 17220
rect 24220 17220 24276 17230
rect 24220 16996 24276 17164
rect 24220 16930 24276 16940
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 23660 15652 23716 15662
rect 23660 13636 23716 15596
rect 23660 13570 23716 13580
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 23776 14140 24096 15652
rect 24220 16100 24276 16110
rect 24220 15204 24276 16044
rect 24220 15138 24276 15148
rect 24436 14924 24756 16436
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 24220 14532 24276 14542
rect 24220 14196 24276 14476
rect 24220 14130 24276 14140
rect 23548 13234 23604 13244
rect 23660 13188 23716 13198
rect 23660 12898 23716 13132
rect 23548 12842 23716 12898
rect 23548 11844 23604 12842
rect 23660 12628 23716 12638
rect 23660 11956 23716 12572
rect 23660 11890 23716 11900
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23548 11778 23604 11788
rect 23776 11004 24096 12516
rect 24436 13356 24756 14868
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 24220 11732 24276 11742
rect 24220 11060 24276 11676
rect 24220 10994 24276 11004
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23660 10276 23716 10286
rect 23660 8708 23716 10220
rect 23660 8642 23716 8652
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23436 2594 23492 2604
rect 23548 8372 23604 8382
rect 23548 1652 23604 8316
rect 23548 1586 23604 1596
rect 23776 7868 24096 9380
rect 24436 10220 24756 11732
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 24220 9268 24276 9278
rect 24220 4116 24276 9212
rect 24220 4050 24276 4060
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24892 24612 24948 24622
rect 24892 6692 24948 24556
rect 25004 20278 25060 43484
rect 25116 38836 25172 46620
rect 25228 45556 25284 45566
rect 25228 42532 25284 45500
rect 25228 42466 25284 42476
rect 25228 39396 25284 39406
rect 25228 39060 25284 39340
rect 25228 38994 25284 39004
rect 25116 38388 25172 38780
rect 25116 38322 25172 38332
rect 25116 37604 25172 37614
rect 25116 35476 25172 37548
rect 25116 35410 25172 35420
rect 25228 36036 25284 36046
rect 25116 33796 25172 33806
rect 25116 20580 25172 33740
rect 25228 29316 25284 35980
rect 25228 29250 25284 29260
rect 25228 27412 25284 27422
rect 25228 23828 25284 27356
rect 25228 23762 25284 23772
rect 25116 20514 25172 20524
rect 25340 20916 25396 47582
rect 25564 45780 25620 53788
rect 25564 45714 25620 45724
rect 25676 48132 25732 48142
rect 25452 45444 25508 45454
rect 25452 42084 25508 45388
rect 25452 42018 25508 42028
rect 25452 38948 25508 38958
rect 25452 38612 25508 38892
rect 25452 38546 25508 38556
rect 25564 35140 25620 35150
rect 25452 34804 25508 34814
rect 25452 30996 25508 34748
rect 25564 31220 25620 35084
rect 25676 34916 25732 48076
rect 25676 34850 25732 34860
rect 25564 31154 25620 31164
rect 25676 32452 25732 32462
rect 25452 30660 25508 30940
rect 25452 30594 25508 30604
rect 25564 26404 25620 26414
rect 25564 23604 25620 26348
rect 25564 23538 25620 23548
rect 25228 20356 25284 20366
rect 25004 20222 25172 20278
rect 25004 20020 25060 20030
rect 25004 19572 25060 19964
rect 25004 10612 25060 19516
rect 25116 17668 25172 20222
rect 25116 17602 25172 17612
rect 25004 10546 25060 10556
rect 25116 16996 25172 17006
rect 25116 7588 25172 16940
rect 25116 7522 25172 7532
rect 24892 6626 24948 6636
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 23776 1596 24096 3108
rect 24220 3108 24276 3118
rect 24220 2772 24276 3052
rect 24220 2706 24276 2716
rect 24436 2380 24756 3892
rect 23324 802 23380 812
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 24220 2324 24276 2334
rect 24220 1652 24276 2268
rect 24220 1586 24276 1596
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 22652 690 22708 700
rect 22876 756 22932 766
rect 15148 354 15204 364
rect 12908 130 12964 140
rect 10780 18 10836 28
rect 22876 84 22932 700
rect 22876 18 22932 28
rect 23776 0 24096 1540
rect 24436 812 24756 2324
rect 25228 2212 25284 20300
rect 25340 2772 25396 20860
rect 25452 23492 25508 23502
rect 25452 18116 25508 23436
rect 25452 18050 25508 18060
rect 25676 13188 25732 32396
rect 25788 16884 25844 55468
rect 25900 52388 25956 55916
rect 26460 55860 26516 55870
rect 25900 52322 25956 52332
rect 26124 52612 26180 52622
rect 25900 52164 25956 52174
rect 25900 44772 25956 52108
rect 26124 48132 26180 52556
rect 26460 50484 26516 55804
rect 26908 55300 26964 55310
rect 26684 54404 26740 54414
rect 26460 50418 26516 50428
rect 26572 52388 26628 52398
rect 26124 48066 26180 48076
rect 26572 48692 26628 52332
rect 26460 47460 26516 47470
rect 26460 47124 26516 47404
rect 26460 47058 26516 47068
rect 25900 33124 25956 44716
rect 26572 41188 26628 48636
rect 26684 44660 26740 54348
rect 26796 53844 26852 53854
rect 26796 53396 26852 53788
rect 26796 53330 26852 53340
rect 26684 44594 26740 44604
rect 26796 50372 26852 50382
rect 26796 48916 26852 50316
rect 26572 41122 26628 41132
rect 26684 44100 26740 44110
rect 26124 39620 26180 39630
rect 26124 33238 26180 39564
rect 26684 39620 26740 44044
rect 26796 39732 26852 48860
rect 26908 44100 26964 55244
rect 27020 46788 27076 46798
rect 27020 44212 27076 46732
rect 27020 44146 27076 44156
rect 26908 44034 26964 44044
rect 27020 40404 27076 40414
rect 26796 39666 26852 39676
rect 26908 40180 26964 40190
rect 26684 39554 26740 39564
rect 25900 33058 25956 33068
rect 26012 33182 26180 33238
rect 26348 39508 26404 39518
rect 25900 32788 25956 32798
rect 25900 32004 25956 32732
rect 25900 31938 25956 31948
rect 25788 16818 25844 16828
rect 25900 26628 25956 26638
rect 25676 13122 25732 13132
rect 25452 11620 25508 11630
rect 25452 10612 25508 11564
rect 25452 10546 25508 10556
rect 25900 7476 25956 26572
rect 25900 7410 25956 7420
rect 26012 3358 26068 33182
rect 26236 31892 26292 31902
rect 26124 31220 26180 31230
rect 26124 30324 26180 31164
rect 26124 30258 26180 30268
rect 26124 30100 26180 30110
rect 26124 24836 26180 30044
rect 26236 26180 26292 31836
rect 26236 26114 26292 26124
rect 26124 24770 26180 24780
rect 26348 23940 26404 39452
rect 26908 38998 26964 40124
rect 26684 38942 26964 38998
rect 27020 39172 27076 40348
rect 26572 33124 26628 33134
rect 26572 31892 26628 33068
rect 26572 31826 26628 31836
rect 26460 31108 26516 31118
rect 26460 28980 26516 31052
rect 26460 28914 26516 28924
rect 26124 22372 26180 22382
rect 26124 12628 26180 22316
rect 26348 21364 26404 23884
rect 26684 24500 26740 38942
rect 26908 38724 26964 38734
rect 26908 37604 26964 38668
rect 26908 37538 26964 37548
rect 26348 21298 26404 21308
rect 26460 21700 26516 21710
rect 26460 21140 26516 21644
rect 26460 21074 26516 21084
rect 26124 12562 26180 12572
rect 26236 20580 26292 20590
rect 26124 10052 26180 10062
rect 26124 3556 26180 9996
rect 26124 3490 26180 3500
rect 25452 3302 26068 3358
rect 25452 3220 25508 3302
rect 25452 3154 25508 3164
rect 25340 2706 25396 2716
rect 25228 2146 25284 2156
rect 25340 2324 25396 2334
rect 25340 1988 25396 2268
rect 26236 2212 26292 20524
rect 26460 20020 26516 20030
rect 26348 11060 26404 11070
rect 26348 10276 26404 11004
rect 26348 10210 26404 10220
rect 26460 3108 26516 19964
rect 26684 14338 26740 24444
rect 26572 14282 26740 14338
rect 26796 36932 26852 36942
rect 26572 9380 26628 14282
rect 26796 14158 26852 36876
rect 27020 28918 27076 39116
rect 27132 36372 27188 56028
rect 27580 55524 27636 55534
rect 27244 54292 27300 54302
rect 27244 43204 27300 54236
rect 27468 46116 27524 46126
rect 27244 43138 27300 43148
rect 27356 44996 27412 45006
rect 27132 36306 27188 36316
rect 27244 37268 27300 37278
rect 26684 14102 26852 14158
rect 26908 28862 27076 28918
rect 27132 34692 27188 34702
rect 26908 21476 26964 28862
rect 27132 28420 27188 34636
rect 27132 28354 27188 28364
rect 26684 11844 26740 14102
rect 26684 11778 26740 11788
rect 26908 13078 26964 21420
rect 27020 21924 27076 21934
rect 27020 16436 27076 21868
rect 27020 16370 27076 16380
rect 27132 20468 27188 20478
rect 27020 13078 27076 13086
rect 26908 13076 27076 13078
rect 26908 13022 27020 13076
rect 26684 9828 26740 9838
rect 26684 9658 26740 9772
rect 26684 9602 26852 9658
rect 26572 8596 26628 9324
rect 26796 9380 26852 9602
rect 26572 8530 26628 8540
rect 26684 8708 26740 8718
rect 26684 8260 26740 8652
rect 26684 7588 26740 8204
rect 26684 7522 26740 7532
rect 26796 3780 26852 9324
rect 26908 9268 26964 13022
rect 27020 13010 27076 13020
rect 26908 6804 26964 9212
rect 26908 6738 26964 6748
rect 27020 5124 27076 5134
rect 27020 4788 27076 5068
rect 27020 4722 27076 4732
rect 26796 3714 26852 3724
rect 26460 2884 26516 3052
rect 27132 3108 27188 20412
rect 27244 18228 27300 37212
rect 27356 36036 27412 44940
rect 27468 42308 27524 46060
rect 27468 42242 27524 42252
rect 27356 35970 27412 35980
rect 27356 33908 27412 33918
rect 27356 30100 27412 33852
rect 27356 30034 27412 30044
rect 27468 30212 27524 30222
rect 27468 24388 27524 30156
rect 27580 27188 27636 55468
rect 27692 48692 27748 48702
rect 27692 38276 27748 48636
rect 27692 38210 27748 38220
rect 27580 27122 27636 27132
rect 27692 34916 27748 34926
rect 27468 24322 27524 24332
rect 27692 23716 27748 34860
rect 27692 23650 27748 23660
rect 27468 21252 27524 21262
rect 27244 14420 27300 18172
rect 27244 14354 27300 14364
rect 27356 18564 27412 18574
rect 27356 8148 27412 18508
rect 27468 17444 27524 21196
rect 27468 17378 27524 17388
rect 27804 15876 27860 56812
rect 34972 56420 35028 56430
rect 31724 56084 31780 56094
rect 29596 55860 29652 55870
rect 28812 55748 28868 55758
rect 28028 55524 28084 55534
rect 27916 54292 27972 54302
rect 27916 45444 27972 54236
rect 27916 45378 27972 45388
rect 27916 33124 27972 33134
rect 27916 31668 27972 33068
rect 27916 31602 27972 31612
rect 27916 31220 27972 31230
rect 27916 30212 27972 31164
rect 27916 30146 27972 30156
rect 27916 29988 27972 29998
rect 27916 28868 27972 29932
rect 27916 28802 27972 28812
rect 27916 24388 27972 24398
rect 27916 19684 27972 24332
rect 28028 20468 28084 55468
rect 28588 51044 28644 51054
rect 28140 50148 28196 50158
rect 28140 49364 28196 50092
rect 28140 49298 28196 49308
rect 28364 48580 28420 48590
rect 28364 47684 28420 48524
rect 28364 47618 28420 47628
rect 28476 47460 28532 47470
rect 28252 47012 28308 47022
rect 28140 46564 28196 46574
rect 28140 44660 28196 46508
rect 28140 44594 28196 44604
rect 28140 41188 28196 41198
rect 28140 24500 28196 41132
rect 28252 37156 28308 46956
rect 28364 46004 28420 46014
rect 28364 43092 28420 45948
rect 28364 43026 28420 43036
rect 28364 42868 28420 42878
rect 28364 42308 28420 42812
rect 28364 42242 28420 42252
rect 28252 37090 28308 37100
rect 28364 30436 28420 30446
rect 28252 29428 28308 29438
rect 28252 29092 28308 29372
rect 28252 29026 28308 29036
rect 28140 22484 28196 24444
rect 28140 22418 28196 22428
rect 28252 25620 28308 25630
rect 28028 20402 28084 20412
rect 27916 19618 27972 19628
rect 27804 15810 27860 15820
rect 27916 17556 27972 17566
rect 27692 9604 27748 9614
rect 27692 9044 27748 9548
rect 27692 8978 27748 8988
rect 27356 8082 27412 8092
rect 27580 5796 27636 5806
rect 27580 5572 27636 5740
rect 27580 5506 27636 5516
rect 27916 4340 27972 17500
rect 27916 4274 27972 4284
rect 28140 17108 28196 17118
rect 28140 3668 28196 17052
rect 28252 9940 28308 25564
rect 28364 18340 28420 30380
rect 28476 24388 28532 47404
rect 28588 46918 28644 50988
rect 28588 46862 28756 46918
rect 28700 46738 28756 46862
rect 28476 24322 28532 24332
rect 28588 46682 28756 46738
rect 28588 39396 28644 46682
rect 28476 24164 28532 24174
rect 28476 20356 28532 24108
rect 28476 20290 28532 20300
rect 28364 18274 28420 18284
rect 28476 12068 28532 12078
rect 28476 10276 28532 12012
rect 28476 10210 28532 10220
rect 28252 9874 28308 9884
rect 28364 6692 28420 6702
rect 28252 5236 28308 5246
rect 28252 4452 28308 5180
rect 28252 4386 28308 4396
rect 28140 3602 28196 3612
rect 28364 3220 28420 6636
rect 28588 4452 28644 39340
rect 28700 35252 28756 35262
rect 28700 31668 28756 35196
rect 28700 31602 28756 31612
rect 28812 28918 28868 55692
rect 29372 55524 29428 55534
rect 29036 52724 29092 52734
rect 29036 49812 29092 52668
rect 29036 49746 29092 49756
rect 29260 50596 29316 50606
rect 29260 47460 29316 50540
rect 29260 47394 29316 47404
rect 29036 46788 29092 46798
rect 28924 46452 28980 46462
rect 28924 46116 28980 46396
rect 29036 46340 29092 46732
rect 29036 46274 29092 46284
rect 28924 46050 28980 46060
rect 28700 28862 28868 28918
rect 28924 44324 28980 44334
rect 28700 25620 28756 28862
rect 28700 25554 28756 25564
rect 28924 27412 28980 44268
rect 29372 44212 29428 55468
rect 29484 52052 29540 52062
rect 29484 50372 29540 51996
rect 29484 50306 29540 50316
rect 29484 48244 29540 48254
rect 29484 47638 29540 48188
rect 29596 47796 29652 55804
rect 30044 55860 30100 55870
rect 29708 52388 29764 52398
rect 29708 52164 29764 52332
rect 29708 52098 29764 52108
rect 30044 51380 30100 55804
rect 30716 55524 30772 55534
rect 29820 51268 29876 51278
rect 29596 47730 29652 47740
rect 29708 49588 29764 49598
rect 29484 47582 29652 47638
rect 29372 44146 29428 44156
rect 29484 47460 29540 47470
rect 29148 42532 29204 42542
rect 29148 41860 29204 42476
rect 29148 41794 29204 41804
rect 29036 41188 29092 41198
rect 29036 40516 29092 41132
rect 29484 41188 29540 47404
rect 29484 41122 29540 41132
rect 29596 47236 29652 47582
rect 29596 40798 29652 47180
rect 29708 43764 29764 49532
rect 29708 43698 29764 43708
rect 29820 45668 29876 51212
rect 30044 51156 30100 51324
rect 30044 51090 30100 51100
rect 30156 55412 30212 55422
rect 29820 40964 29876 45612
rect 29820 40898 29876 40908
rect 29932 50484 29988 50494
rect 29596 40742 29876 40798
rect 29036 40450 29092 40460
rect 29260 38724 29316 38734
rect 29036 38052 29092 38062
rect 29036 28868 29092 37996
rect 29036 28802 29092 28812
rect 29148 35476 29204 35486
rect 28812 25284 28868 25294
rect 28700 25060 28756 25070
rect 28700 20580 28756 25004
rect 28700 20514 28756 20524
rect 28812 16996 28868 25228
rect 28924 19236 28980 27356
rect 29036 25620 29092 25630
rect 29036 24724 29092 25564
rect 29036 24658 29092 24668
rect 28924 19170 28980 19180
rect 29036 23940 29092 23950
rect 28812 16930 28868 16940
rect 28700 16324 28756 16334
rect 28700 13076 28756 16268
rect 28700 12292 28756 13020
rect 28700 12226 28756 12236
rect 28924 12516 28980 12526
rect 28924 12292 28980 12460
rect 28924 12226 28980 12236
rect 29036 11732 29092 23884
rect 29148 12964 29204 35420
rect 29260 25060 29316 38668
rect 29372 38388 29428 38398
rect 29372 32452 29428 38332
rect 29820 35476 29876 40742
rect 29932 37156 29988 50428
rect 30044 50148 30100 50158
rect 30044 48718 30100 50092
rect 30156 48898 30212 55356
rect 30492 55412 30548 55422
rect 30380 54852 30436 54862
rect 30268 51380 30324 51390
rect 30268 50820 30324 51324
rect 30268 50754 30324 50764
rect 30380 49140 30436 54796
rect 30380 49074 30436 49084
rect 30156 48842 30324 48898
rect 30044 48662 30212 48718
rect 29932 37090 29988 37100
rect 30044 48468 30100 48478
rect 29820 35410 29876 35420
rect 29932 36932 29988 36942
rect 29932 36372 29988 36876
rect 29932 32878 29988 36316
rect 30044 35700 30100 48412
rect 30156 46788 30212 48662
rect 30268 47348 30324 48842
rect 30268 47282 30324 47292
rect 30380 48020 30436 48030
rect 30156 44996 30212 46732
rect 30156 44930 30212 44940
rect 30380 36372 30436 47964
rect 30380 36306 30436 36316
rect 30044 35634 30100 35644
rect 30380 33572 30436 33582
rect 29932 32822 30212 32878
rect 29372 25732 29428 32396
rect 29708 32340 29764 32350
rect 29484 31444 29540 31454
rect 29484 27860 29540 31388
rect 29484 27794 29540 27804
rect 29708 28756 29764 32284
rect 29820 31332 29876 31342
rect 29820 30100 29876 31276
rect 30044 30996 30100 31006
rect 30044 30898 30100 30940
rect 29820 30034 29876 30044
rect 29932 30842 30100 30898
rect 29372 25666 29428 25676
rect 29260 24994 29316 25004
rect 29260 24836 29316 24846
rect 29260 23604 29316 24780
rect 29260 23538 29316 23548
rect 29372 20580 29428 20590
rect 29372 14878 29428 20524
rect 29708 16548 29764 28700
rect 29820 28868 29876 28878
rect 29820 24276 29876 28812
rect 29820 24210 29876 24220
rect 29932 27860 29988 30842
rect 29932 20098 29988 27804
rect 30044 24052 30100 24062
rect 30044 20468 30100 23996
rect 30044 20402 30100 20412
rect 29932 20042 30100 20098
rect 30044 20020 30100 20042
rect 30044 19954 30100 19964
rect 29708 16482 29764 16492
rect 29932 19236 29988 19246
rect 29820 16324 29876 16334
rect 29820 15652 29876 16268
rect 29372 14822 29540 14878
rect 29372 14756 29428 14766
rect 29148 12898 29204 12908
rect 29260 14084 29316 14094
rect 29148 12516 29204 12526
rect 29148 11956 29204 12460
rect 29148 11890 29204 11900
rect 29036 11666 29092 11676
rect 29260 10724 29316 14028
rect 29260 10658 29316 10668
rect 28588 4386 28644 4396
rect 29036 9044 29092 9054
rect 28364 3154 28420 3164
rect 27132 3042 27188 3052
rect 26460 2818 26516 2828
rect 29036 2660 29092 8988
rect 29372 5796 29428 14700
rect 29484 13636 29540 14822
rect 29484 13570 29540 13580
rect 29820 8260 29876 15596
rect 29932 11508 29988 19180
rect 29932 11060 29988 11452
rect 29932 10994 29988 11004
rect 30044 12740 30100 12750
rect 29820 8194 29876 8204
rect 30044 7700 30100 12684
rect 30044 7634 30100 7644
rect 29372 5730 29428 5740
rect 29036 2594 29092 2604
rect 26236 2146 26292 2156
rect 25340 1922 25396 1932
rect 30156 1316 30212 32822
rect 30268 27412 30324 27422
rect 30268 26852 30324 27356
rect 30268 26786 30324 26796
rect 30268 23044 30324 23054
rect 30268 22596 30324 22988
rect 30268 22530 30324 22540
rect 30380 17668 30436 33516
rect 30492 24948 30548 55356
rect 30604 53508 30660 53518
rect 30604 49588 30660 53452
rect 30604 49522 30660 49532
rect 30604 49252 30660 49262
rect 30604 48580 30660 49196
rect 30604 48514 30660 48524
rect 30492 24882 30548 24892
rect 30604 44548 30660 44558
rect 30604 41748 30660 44492
rect 30716 44324 30772 55468
rect 30828 55412 30884 55422
rect 30828 52164 30884 55356
rect 31500 53732 31556 53742
rect 31164 53508 31220 53518
rect 31164 52836 31220 53452
rect 31164 52770 31220 52780
rect 30828 52098 30884 52108
rect 31164 51380 31220 51390
rect 30940 50708 30996 50718
rect 30940 50158 30996 50652
rect 30828 50102 30996 50158
rect 30828 46676 30884 50102
rect 31164 49438 31220 51324
rect 31500 50158 31556 53676
rect 30940 49382 31220 49438
rect 30940 49364 30996 49382
rect 30940 49298 30996 49308
rect 30828 46116 30884 46620
rect 30828 46050 30884 46060
rect 30716 44258 30772 44268
rect 30828 45892 30884 45902
rect 30380 17578 30436 17612
rect 30268 17522 30436 17578
rect 30268 14420 30324 17522
rect 30268 14354 30324 14364
rect 30380 16436 30436 16446
rect 30380 8260 30436 16380
rect 30604 16324 30660 41692
rect 30716 39284 30772 39294
rect 30716 33460 30772 39228
rect 30828 38612 30884 45836
rect 31052 45332 31108 45342
rect 30828 38546 30884 38556
rect 30940 41188 30996 41198
rect 30716 33394 30772 33404
rect 30828 38164 30884 38174
rect 30716 31220 30772 31230
rect 30716 29098 30772 31164
rect 30828 29428 30884 38108
rect 30940 34916 30996 41132
rect 31052 38052 31108 45276
rect 31164 41972 31220 49382
rect 31164 41906 31220 41916
rect 31276 50102 31556 50158
rect 31612 50148 31668 50158
rect 31276 48020 31332 50102
rect 31612 49798 31668 50092
rect 31500 49742 31668 49798
rect 31388 49364 31444 49374
rect 31388 48244 31444 49308
rect 31388 48178 31444 48188
rect 31500 48580 31556 49742
rect 31276 43652 31332 47964
rect 31276 41338 31332 43596
rect 31388 46340 31444 46350
rect 31388 42084 31444 46284
rect 31500 44100 31556 48524
rect 31500 44034 31556 44044
rect 31612 46900 31668 46910
rect 31388 42018 31444 42028
rect 31276 41282 31556 41338
rect 31388 41076 31444 41086
rect 31388 40516 31444 41020
rect 31388 40450 31444 40460
rect 31500 38612 31556 41282
rect 31500 38546 31556 38556
rect 31052 37986 31108 37996
rect 31612 36148 31668 46844
rect 30940 34850 30996 34860
rect 31500 34916 31556 34926
rect 31164 33572 31220 33582
rect 30828 29278 30884 29372
rect 31052 29876 31108 29886
rect 30828 29222 30996 29278
rect 30716 29042 30884 29098
rect 30828 25284 30884 29042
rect 30828 25218 30884 25228
rect 30828 22820 30884 22830
rect 30828 22484 30884 22764
rect 30828 22418 30884 22428
rect 30940 22372 30996 29222
rect 30940 22306 30996 22316
rect 30940 20020 30996 20030
rect 30940 18900 30996 19964
rect 30940 18834 30996 18844
rect 31052 17892 31108 29820
rect 31164 26180 31220 33516
rect 31276 28308 31332 28318
rect 31276 28198 31332 28252
rect 31276 28142 31444 28198
rect 31164 24052 31220 26124
rect 31164 23986 31220 23996
rect 31276 24724 31332 24734
rect 31052 17668 31108 17836
rect 31052 17602 31108 17612
rect 31164 23044 31220 23054
rect 30604 16258 30660 16268
rect 31052 16100 31108 16110
rect 31052 15876 31108 16044
rect 30380 8194 30436 8204
rect 30940 14868 30996 14878
rect 30940 7476 30996 14812
rect 30940 7410 30996 7420
rect 30156 1250 30212 1260
rect 31052 1204 31108 15820
rect 31164 14868 31220 22988
rect 31164 14802 31220 14812
rect 31276 21140 31332 24668
rect 31164 14532 31220 14542
rect 31164 3556 31220 14476
rect 31276 10612 31332 21084
rect 31388 18228 31444 28142
rect 31500 24724 31556 34860
rect 31612 28420 31668 36092
rect 31724 32878 31780 56028
rect 32508 56084 32564 56094
rect 32284 55860 32340 55870
rect 32172 55300 32228 55310
rect 31836 53172 31892 53182
rect 31836 37604 31892 53116
rect 32172 49364 32228 55244
rect 32172 49298 32228 49308
rect 32284 48468 32340 55804
rect 32396 54852 32452 54862
rect 32396 54292 32452 54796
rect 32396 54226 32452 54236
rect 32284 48402 32340 48412
rect 32396 50596 32452 50606
rect 32396 47796 32452 50540
rect 31948 46788 32004 46798
rect 31948 45444 32004 46732
rect 31948 45378 32004 45388
rect 32060 41972 32116 41982
rect 32060 40516 32116 41916
rect 32396 41972 32452 47740
rect 32396 41906 32452 41916
rect 31836 37538 31892 37548
rect 31948 38612 32004 38622
rect 31948 37268 32004 38556
rect 31948 37202 32004 37212
rect 31836 35028 31892 35038
rect 31836 33236 31892 34972
rect 31836 33170 31892 33180
rect 31948 34692 32004 34702
rect 31724 32822 31892 32878
rect 31612 28354 31668 28364
rect 31724 32564 31780 32574
rect 31724 28084 31780 32508
rect 31724 28018 31780 28028
rect 31500 24658 31556 24668
rect 31388 18162 31444 18172
rect 31612 23716 31668 23726
rect 31500 18004 31556 18014
rect 31500 17444 31556 17948
rect 31500 17378 31556 17388
rect 31276 10546 31332 10556
rect 31388 16548 31444 16558
rect 31388 10018 31444 16492
rect 31612 12068 31668 23660
rect 31612 12002 31668 12012
rect 31724 20580 31780 20590
rect 31388 9962 31556 10018
rect 31388 9828 31444 9838
rect 31388 9604 31444 9772
rect 31388 9538 31444 9548
rect 31388 8260 31444 8270
rect 31388 7476 31444 8204
rect 31388 7410 31444 7420
rect 31500 4004 31556 9962
rect 31500 3938 31556 3948
rect 31164 3490 31220 3500
rect 31724 2884 31780 20524
rect 31836 19348 31892 32822
rect 31948 30324 32004 34636
rect 31948 30258 32004 30268
rect 31836 19282 31892 19292
rect 31836 19124 31892 19134
rect 31836 12292 31892 19068
rect 32060 13636 32116 40460
rect 32508 34020 32564 56028
rect 33404 56084 33460 56094
rect 32732 55300 32788 55310
rect 32620 52276 32676 52286
rect 32620 51268 32676 52220
rect 32620 51202 32676 51212
rect 32732 51380 32788 55244
rect 33180 55188 33236 55198
rect 32732 50820 32788 51324
rect 32732 50754 32788 50764
rect 32844 54628 32900 54638
rect 32844 47796 32900 54572
rect 33068 54292 33124 54302
rect 32844 47730 32900 47740
rect 32956 52164 33012 52174
rect 32844 46676 32900 46686
rect 32844 46116 32900 46620
rect 32844 46050 32900 46060
rect 32956 43428 33012 52108
rect 32956 42532 33012 43372
rect 32956 42466 33012 42476
rect 32508 33954 32564 33964
rect 32620 41972 32676 41982
rect 32396 32788 32452 32798
rect 32172 31444 32228 31454
rect 32172 29316 32228 31388
rect 32172 24724 32228 29260
rect 32284 28980 32340 28990
rect 32284 25844 32340 28924
rect 32284 25060 32340 25788
rect 32284 24994 32340 25004
rect 32172 24658 32228 24668
rect 32284 24612 32340 24622
rect 32060 13570 32116 13580
rect 32172 23492 32228 23502
rect 32172 13860 32228 23436
rect 32284 22596 32340 24556
rect 32284 22530 32340 22540
rect 32284 20468 32340 20478
rect 32284 17668 32340 20412
rect 32284 17602 32340 17612
rect 32396 16212 32452 32732
rect 32396 16146 32452 16156
rect 32508 32564 32564 32574
rect 32284 16100 32340 16110
rect 32284 15652 32340 16044
rect 32284 15586 32340 15596
rect 32172 13524 32228 13804
rect 32172 13458 32228 13468
rect 31836 12226 31892 12236
rect 31948 12068 32004 12078
rect 31836 6916 31892 6926
rect 31836 4676 31892 6860
rect 31948 4788 32004 12012
rect 32172 11172 32228 11182
rect 32060 10276 32116 10286
rect 32060 7924 32116 10220
rect 32060 7858 32116 7868
rect 32172 8596 32228 11116
rect 31948 4722 32004 4732
rect 31836 4610 31892 4620
rect 32172 3780 32228 8540
rect 32508 8260 32564 32508
rect 32508 8194 32564 8204
rect 32620 4340 32676 41916
rect 33068 33124 33124 54236
rect 33180 47348 33236 55132
rect 33292 54964 33348 54974
rect 33292 52500 33348 54908
rect 33292 52434 33348 52444
rect 33180 47282 33236 47292
rect 33292 50932 33348 50942
rect 33068 33058 33124 33068
rect 33180 43428 33236 43438
rect 32956 31892 33012 31902
rect 32956 31668 33012 31836
rect 32844 31444 32900 31454
rect 32732 30996 32788 31006
rect 32732 12718 32788 30940
rect 32844 30436 32900 31388
rect 32844 26740 32900 30380
rect 32956 28378 33012 31612
rect 33068 31220 33124 31230
rect 33068 30436 33124 31164
rect 33068 30370 33124 30380
rect 32956 28322 33124 28378
rect 32844 26674 32900 26684
rect 32956 28196 33012 28206
rect 32956 26292 33012 28140
rect 32956 26226 33012 26236
rect 33068 24612 33124 28322
rect 33180 25620 33236 43372
rect 33292 39172 33348 50876
rect 33292 39106 33348 39116
rect 33180 25554 33236 25564
rect 33292 35700 33348 35710
rect 33068 24546 33124 24556
rect 33292 23044 33348 35644
rect 33292 22978 33348 22988
rect 33292 22596 33348 22606
rect 33292 22148 33348 22540
rect 33292 22082 33348 22092
rect 33068 20356 33124 20366
rect 32844 16772 32900 16782
rect 32844 16324 32900 16716
rect 33068 16772 33124 20300
rect 33068 16706 33124 16716
rect 33404 17556 33460 56028
rect 34748 56084 34804 56094
rect 34300 55860 34356 55870
rect 33852 55412 33908 55422
rect 33516 51156 33572 51166
rect 33516 38724 33572 51100
rect 33740 45444 33796 45454
rect 33628 45108 33684 45118
rect 33628 41076 33684 45052
rect 33628 41010 33684 41020
rect 33516 38500 33572 38668
rect 33516 38434 33572 38444
rect 33740 38388 33796 45388
rect 33740 38322 33796 38332
rect 33628 37492 33684 37502
rect 33628 35700 33684 37436
rect 33628 35634 33684 35644
rect 33852 34020 33908 55356
rect 34188 55412 34244 55422
rect 33964 51380 34020 51390
rect 33964 48580 34020 51324
rect 33964 48514 34020 48524
rect 34076 49364 34132 49374
rect 34076 47684 34132 49308
rect 34188 49252 34244 55356
rect 34300 49364 34356 55804
rect 34524 55524 34580 55534
rect 34300 49298 34356 49308
rect 34412 52164 34468 52174
rect 34188 49186 34244 49196
rect 34076 47618 34132 47628
rect 34412 44758 34468 52108
rect 34300 44702 34468 44758
rect 34076 44100 34132 44110
rect 34076 41972 34132 44044
rect 33852 33954 33908 33964
rect 33964 41076 34020 41086
rect 33964 40740 34020 41020
rect 33516 33124 33572 33134
rect 33516 28532 33572 33068
rect 33516 27076 33572 28476
rect 33628 29988 33684 29998
rect 33628 28196 33684 29932
rect 33628 28130 33684 28140
rect 33740 29764 33796 29774
rect 33516 27010 33572 27020
rect 33740 25844 33796 29708
rect 33740 25778 33796 25788
rect 33852 26852 33908 26862
rect 33628 25732 33684 25742
rect 32844 16258 32900 16268
rect 33180 16212 33236 16222
rect 33180 15540 33236 16156
rect 33180 15474 33236 15484
rect 32844 15316 32900 15326
rect 32844 14980 32900 15260
rect 32844 14914 32900 14924
rect 33292 13636 33348 13646
rect 32732 12662 32900 12718
rect 32844 9492 32900 12662
rect 32844 9044 32900 9436
rect 32844 8978 32900 8988
rect 33180 11396 33236 11406
rect 32620 4274 32676 4284
rect 32732 7140 32788 7150
rect 32172 3714 32228 3724
rect 31724 2818 31780 2828
rect 32060 2660 32116 2670
rect 32060 2436 32116 2604
rect 32060 2370 32116 2380
rect 31052 1138 31108 1148
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 32732 84 32788 7084
rect 33068 6916 33124 6926
rect 33068 6356 33124 6860
rect 33068 6290 33124 6300
rect 33180 6580 33236 11340
rect 33180 5908 33236 6524
rect 33180 5842 33236 5852
rect 33292 2772 33348 13580
rect 33404 12740 33460 17500
rect 33516 25620 33572 25630
rect 33516 19796 33572 25564
rect 33628 24164 33684 25676
rect 33852 25732 33908 26796
rect 33852 25666 33908 25676
rect 33628 24098 33684 24108
rect 33740 24836 33796 24846
rect 33516 15316 33572 19740
rect 33740 19124 33796 24780
rect 33852 23940 33908 23950
rect 33852 23604 33908 23884
rect 33852 23538 33908 23548
rect 33740 19058 33796 19068
rect 33852 19908 33908 19918
rect 33516 15250 33572 15260
rect 33740 18116 33796 18126
rect 33404 12674 33460 12684
rect 33404 9828 33460 9838
rect 33404 9268 33460 9772
rect 33404 9202 33460 9212
rect 33740 8260 33796 18060
rect 33852 12180 33908 19852
rect 33964 17556 34020 40684
rect 33964 17490 34020 17500
rect 33852 12114 33908 12124
rect 33740 8194 33796 8204
rect 33964 10052 34020 10062
rect 33740 7812 33796 7822
rect 33628 6916 33684 6926
rect 33404 6692 33460 6702
rect 33404 5908 33460 6636
rect 33628 6692 33684 6860
rect 33628 6626 33684 6636
rect 33404 5842 33460 5852
rect 33292 2706 33348 2716
rect 33740 2772 33796 7756
rect 33964 3332 34020 9996
rect 34076 4340 34132 41916
rect 34300 40740 34356 44702
rect 34300 40674 34356 40684
rect 34412 42868 34468 42878
rect 34188 35476 34244 35486
rect 34188 29818 34244 35420
rect 34300 34468 34356 34478
rect 34300 29988 34356 34412
rect 34300 29922 34356 29932
rect 34188 29762 34356 29818
rect 34188 28308 34244 28318
rect 34188 26404 34244 28252
rect 34188 26338 34244 26348
rect 34188 23268 34244 23278
rect 34188 22820 34244 23212
rect 34188 22754 34244 22764
rect 34188 22372 34244 22382
rect 34188 15652 34244 22316
rect 34300 21924 34356 29762
rect 34412 29764 34468 42812
rect 34412 29698 34468 29708
rect 34300 21858 34356 21868
rect 34412 28420 34468 28430
rect 34188 15586 34244 15596
rect 34300 20804 34356 20814
rect 34300 13798 34356 20748
rect 34412 18116 34468 28364
rect 34524 22372 34580 55468
rect 34636 52276 34692 52286
rect 34636 49700 34692 52220
rect 34636 49634 34692 49644
rect 34636 49140 34692 49150
rect 34636 46900 34692 49084
rect 34636 46834 34692 46844
rect 34636 46116 34692 46126
rect 34636 30772 34692 46060
rect 34748 41524 34804 56028
rect 34860 51156 34916 51166
rect 34860 48356 34916 51100
rect 34972 50036 35028 56364
rect 35756 55860 35812 55870
rect 35196 55748 35252 55758
rect 34972 49970 35028 49980
rect 35084 53956 35140 53966
rect 35084 52500 35140 53900
rect 35084 48804 35140 52444
rect 35084 48738 35140 48748
rect 34860 48290 34916 48300
rect 34860 47348 34916 47358
rect 34860 45444 34916 47292
rect 34860 45378 34916 45388
rect 34972 47012 35028 47022
rect 34748 41458 34804 41468
rect 34860 42980 34916 42990
rect 34636 30706 34692 30716
rect 34748 40068 34804 40078
rect 34636 29764 34692 29774
rect 34636 25138 34692 29708
rect 34748 27188 34804 40012
rect 34860 39284 34916 42924
rect 34972 40292 35028 46956
rect 35084 42532 35140 42542
rect 35084 40852 35140 42476
rect 35196 41076 35252 55692
rect 35420 55524 35476 55534
rect 35308 48356 35364 48366
rect 35308 48132 35364 48300
rect 35308 48066 35364 48076
rect 35420 44578 35476 55468
rect 35532 53844 35588 53854
rect 35532 46116 35588 53788
rect 35532 46050 35588 46060
rect 35644 46452 35700 46462
rect 35196 41010 35252 41020
rect 35308 44522 35476 44578
rect 35532 45444 35588 45454
rect 35084 40786 35140 40796
rect 34972 40226 35028 40236
rect 34860 36820 34916 39228
rect 35196 39844 35252 39854
rect 35196 38500 35252 39788
rect 35196 38434 35252 38444
rect 34860 36754 34916 36764
rect 35196 36148 35252 36158
rect 35084 30772 35140 30782
rect 34972 29988 35028 29998
rect 34748 27122 34804 27132
rect 34860 29876 34916 29886
rect 34748 25844 34804 25854
rect 34748 25284 34804 25788
rect 34748 25218 34804 25228
rect 34860 25620 34916 29820
rect 34972 29204 35028 29932
rect 34972 29138 35028 29148
rect 34636 25082 34804 25138
rect 34748 24724 34804 25082
rect 34748 24658 34804 24668
rect 34636 24612 34692 24622
rect 34636 24388 34692 24556
rect 34636 24322 34692 24332
rect 34860 23716 34916 25564
rect 34972 26852 35028 26862
rect 34972 24612 35028 26796
rect 34972 24546 35028 24556
rect 34860 23650 34916 23660
rect 34524 22306 34580 22316
rect 34860 22820 34916 22830
rect 34748 21924 34804 21934
rect 34636 19236 34692 19246
rect 34412 18050 34468 18060
rect 34524 18564 34580 18574
rect 34412 17108 34468 17118
rect 34412 15876 34468 17052
rect 34412 15810 34468 15820
rect 34300 13742 34468 13798
rect 34412 13636 34468 13742
rect 34076 4274 34132 4284
rect 34188 11844 34244 11854
rect 33964 3266 34020 3276
rect 33740 2706 33796 2716
rect 34188 2772 34244 11788
rect 34412 8148 34468 13580
rect 34524 12068 34580 18508
rect 34636 12292 34692 19180
rect 34636 12226 34692 12236
rect 34524 12002 34580 12012
rect 34748 9828 34804 21868
rect 34860 17108 34916 22764
rect 35084 22820 35140 30716
rect 35084 22754 35140 22764
rect 35196 29316 35252 36092
rect 35308 33908 35364 44522
rect 35420 42644 35476 42654
rect 35420 39732 35476 42588
rect 35420 39666 35476 39676
rect 35532 38948 35588 45388
rect 35644 40740 35700 46396
rect 35644 40674 35700 40684
rect 35308 33842 35364 33852
rect 35420 35364 35476 35374
rect 35196 25396 35252 29260
rect 35308 32452 35364 32462
rect 35308 32228 35364 32396
rect 35308 28308 35364 32172
rect 35420 29876 35476 35308
rect 35420 29810 35476 29820
rect 35308 28242 35364 28252
rect 35420 29204 35476 29214
rect 35084 19460 35140 19470
rect 34860 17042 34916 17052
rect 34972 19236 35028 19246
rect 34972 19012 35028 19180
rect 34972 16996 35028 18956
rect 35084 18788 35140 19404
rect 35084 18722 35140 18732
rect 35196 17758 35252 25340
rect 35420 23492 35476 29148
rect 35420 23426 35476 23436
rect 35532 21700 35588 38892
rect 35644 28644 35700 28654
rect 35644 26180 35700 28588
rect 35644 26114 35700 26124
rect 34972 16930 35028 16940
rect 35084 17702 35252 17758
rect 35308 17892 35364 17902
rect 35084 16858 35140 17702
rect 34972 16802 35140 16858
rect 34860 16548 34916 16558
rect 34860 13412 34916 16492
rect 34972 15958 35028 16802
rect 35084 16660 35140 16670
rect 35084 16212 35140 16604
rect 35308 16548 35364 17836
rect 35420 16884 35476 16894
rect 35420 16660 35476 16828
rect 35420 16594 35476 16604
rect 35308 16482 35364 16492
rect 35084 16146 35140 16156
rect 34972 15902 35252 15958
rect 34860 13346 34916 13356
rect 34748 9762 34804 9772
rect 34412 3220 34468 8092
rect 34636 6580 34692 6590
rect 34636 5348 34692 6524
rect 35084 6468 35140 6478
rect 34972 6356 35028 6366
rect 34972 6238 35028 6300
rect 34860 6182 35028 6238
rect 34860 5908 34916 6182
rect 34860 5842 34916 5852
rect 35084 5908 35140 6412
rect 35084 5842 35140 5852
rect 34636 5282 34692 5292
rect 34412 3154 34468 3164
rect 34188 2706 34244 2716
rect 35196 2772 35252 15902
rect 35532 11844 35588 21644
rect 35532 11778 35588 11788
rect 35756 4340 35812 55804
rect 37324 55860 37380 55870
rect 36316 55412 36372 55422
rect 35868 52948 35924 52958
rect 35868 52276 35924 52892
rect 35868 38388 35924 52220
rect 36092 46452 36148 46462
rect 35980 46116 36036 46126
rect 35980 42532 36036 46060
rect 35980 42466 36036 42476
rect 36092 40516 36148 46396
rect 35868 38322 35924 38332
rect 35980 40180 36036 40190
rect 35980 35476 36036 40124
rect 36092 37380 36148 40460
rect 36092 37314 36148 37324
rect 35980 35410 36036 35420
rect 36204 32788 36260 32798
rect 35868 32676 35924 32686
rect 35868 28868 35924 32620
rect 36204 30884 36260 32732
rect 36204 30818 36260 30828
rect 35868 28802 35924 28812
rect 36092 30212 36148 30222
rect 35980 20692 36036 20702
rect 35980 16100 36036 20636
rect 35980 16034 36036 16044
rect 35980 10164 36036 10174
rect 35980 9380 36036 10108
rect 35980 9314 36036 9324
rect 35756 4274 35812 4284
rect 35980 4788 36036 4798
rect 35980 4116 36036 4732
rect 35980 4050 36036 4060
rect 35196 2706 35252 2716
rect 35980 3108 36036 3118
rect 35980 1764 36036 3052
rect 36092 2212 36148 30156
rect 36204 29540 36260 29550
rect 36204 28980 36260 29484
rect 36204 28914 36260 28924
rect 36204 18116 36260 18126
rect 36204 3108 36260 18060
rect 36316 8260 36372 55356
rect 36540 54628 36596 54638
rect 36540 50148 36596 54572
rect 36876 54292 36932 54302
rect 36540 50082 36596 50092
rect 36652 54068 36708 54078
rect 36540 41188 36596 41198
rect 36540 31892 36596 41132
rect 36540 31826 36596 31836
rect 36428 31668 36484 31678
rect 36428 9604 36484 31612
rect 36428 9538 36484 9548
rect 36540 22932 36596 22942
rect 36540 22596 36596 22876
rect 36316 8194 36372 8204
rect 36540 6468 36596 22540
rect 36540 6402 36596 6412
rect 36204 3042 36260 3052
rect 36316 3668 36372 3678
rect 36316 2772 36372 3612
rect 36316 2706 36372 2716
rect 36652 2772 36708 54012
rect 36876 54068 36932 54236
rect 36876 54002 36932 54012
rect 36764 53844 36820 53854
rect 36764 46676 36820 53788
rect 37100 49588 37156 49598
rect 37100 47012 37156 49532
rect 37100 46946 37156 46956
rect 36764 46340 36820 46620
rect 36764 46274 36820 46284
rect 37212 43764 37268 43774
rect 36764 41524 36820 41534
rect 36764 38948 36820 41468
rect 36764 38882 36820 38892
rect 37212 37198 37268 43708
rect 37100 37142 37268 37198
rect 37100 35364 37156 37142
rect 37100 35298 37156 35308
rect 37212 35476 37268 35486
rect 36988 35028 37044 35038
rect 36876 31892 36932 31902
rect 36876 31668 36932 31836
rect 36876 31602 36932 31612
rect 36988 30884 37044 34972
rect 37100 33348 37156 33358
rect 37100 32340 37156 33292
rect 37100 32274 37156 32284
rect 36988 30818 37044 30828
rect 37100 31220 37156 31230
rect 36876 30772 36932 30782
rect 36764 28644 36820 28654
rect 36764 21028 36820 28588
rect 36764 20962 36820 20972
rect 36876 19908 36932 30716
rect 36988 30436 37044 30446
rect 36988 29540 37044 30380
rect 36988 29474 37044 29484
rect 36988 26180 37044 26190
rect 36988 23828 37044 26124
rect 36988 23762 37044 23772
rect 36988 23492 37044 23502
rect 36988 22932 37044 23436
rect 36988 22866 37044 22876
rect 36876 19842 36932 19852
rect 37100 18340 37156 31164
rect 37212 28756 37268 35420
rect 37212 25620 37268 28700
rect 37212 25554 37268 25564
rect 37100 18274 37156 18284
rect 37212 23492 37268 23502
rect 37212 22596 37268 23436
rect 36988 18228 37044 18238
rect 36876 16100 36932 16110
rect 36876 12964 36932 16044
rect 36876 12898 36932 12908
rect 36652 2706 36708 2716
rect 36764 9268 36820 9278
rect 36092 2146 36148 2156
rect 35980 1698 36036 1708
rect 32732 18 32788 28
rect 36764 84 36820 9212
rect 36988 9268 37044 18172
rect 37212 17108 37268 22540
rect 37212 17042 37268 17052
rect 37100 15764 37156 15774
rect 37100 12292 37156 15708
rect 37100 12226 37156 12236
rect 36988 9202 37044 9212
rect 37100 11284 37156 11294
rect 37100 7700 37156 11228
rect 37212 10724 37268 10734
rect 37212 9940 37268 10668
rect 37212 9874 37268 9884
rect 37100 7634 37156 7644
rect 37324 2772 37380 55804
rect 38332 55524 38388 55534
rect 37884 55412 37940 55422
rect 37772 54852 37828 54862
rect 37436 52724 37492 52734
rect 37436 52276 37492 52668
rect 37436 52210 37492 52220
rect 37548 50372 37604 50382
rect 37436 41860 37492 41870
rect 37436 36708 37492 41804
rect 37548 40516 37604 50316
rect 37772 50372 37828 54796
rect 37772 50306 37828 50316
rect 37772 46004 37828 46014
rect 37660 45892 37716 45902
rect 37660 42980 37716 45836
rect 37660 42914 37716 42924
rect 37772 43316 37828 45948
rect 37548 40450 37604 40460
rect 37436 36642 37492 36652
rect 37548 36484 37604 36494
rect 37436 32340 37492 32350
rect 37436 20356 37492 32284
rect 37548 30436 37604 36428
rect 37660 35028 37716 35038
rect 37660 31780 37716 34972
rect 37660 31714 37716 31724
rect 37548 30370 37604 30380
rect 37436 20290 37492 20300
rect 37660 30212 37716 30222
rect 37548 15316 37604 15326
rect 37548 14980 37604 15260
rect 37548 14914 37604 14924
rect 37324 2706 37380 2716
rect 37660 1204 37716 30156
rect 37772 18228 37828 43260
rect 37772 17444 37828 18172
rect 37884 17892 37940 55356
rect 38220 51268 38276 51278
rect 38220 49476 38276 51212
rect 38220 49410 38276 49420
rect 38220 47908 38276 47918
rect 38220 43876 38276 47852
rect 38220 43810 38276 43820
rect 38220 42308 38276 42318
rect 38220 36596 38276 42252
rect 38220 36530 38276 36540
rect 38108 33908 38164 33918
rect 38108 33778 38164 33852
rect 37996 33722 38164 33778
rect 37996 33058 38052 33722
rect 38108 33348 38164 33358
rect 38108 33238 38164 33292
rect 38108 33182 38276 33238
rect 37996 33002 38164 33058
rect 37884 17826 37940 17836
rect 37996 32340 38052 32350
rect 37772 17378 37828 17388
rect 37996 13636 38052 32284
rect 38108 28308 38164 33002
rect 38220 32676 38276 33182
rect 38220 32610 38276 32620
rect 38108 28242 38164 28252
rect 38108 26740 38164 26750
rect 38108 25396 38164 26684
rect 38108 25330 38164 25340
rect 38220 25172 38276 25182
rect 38220 24836 38276 25116
rect 38220 24770 38276 24780
rect 38220 24500 38276 24510
rect 38220 24164 38276 24444
rect 38220 24098 38276 24108
rect 38108 17444 38164 17454
rect 38108 15540 38164 17388
rect 38108 15474 38164 15484
rect 37996 13570 38052 13580
rect 38220 7140 38276 7150
rect 38220 6804 38276 7084
rect 38220 6738 38276 6748
rect 38332 2212 38388 55468
rect 38444 49812 38500 57036
rect 43776 56476 44096 57456
rect 42812 56420 42868 56430
rect 42364 56084 42420 56094
rect 38444 49746 38500 49756
rect 38556 55860 38612 55870
rect 38444 49476 38500 49486
rect 38444 43764 38500 49420
rect 38444 43698 38500 43708
rect 38444 35252 38500 35262
rect 38444 33460 38500 35196
rect 38444 33394 38500 33404
rect 38444 28420 38500 28430
rect 38444 27188 38500 28364
rect 38444 27122 38500 27132
rect 38444 23268 38500 23278
rect 38444 19236 38500 23212
rect 38444 19170 38500 19180
rect 38444 18004 38500 18014
rect 38444 17780 38500 17948
rect 38444 17714 38500 17724
rect 38444 15428 38500 15438
rect 38444 15204 38500 15372
rect 38444 15138 38500 15148
rect 38556 4340 38612 55804
rect 39116 55860 39172 55870
rect 38780 54628 38836 54638
rect 38668 45220 38724 45230
rect 38668 44100 38724 45164
rect 38668 44034 38724 44044
rect 38668 42532 38724 42542
rect 38668 35140 38724 42476
rect 38668 35074 38724 35084
rect 38668 31780 38724 31790
rect 38668 8708 38724 31724
rect 38668 8642 38724 8652
rect 38556 4274 38612 4284
rect 38332 2146 38388 2156
rect 38780 1652 38836 54572
rect 38892 50484 38948 50494
rect 38892 49798 38948 50428
rect 38892 49742 39060 49798
rect 38892 49588 38948 49598
rect 38892 39284 38948 49532
rect 39004 41300 39060 49742
rect 39004 41234 39060 41244
rect 38892 39218 38948 39228
rect 39004 35252 39060 35262
rect 38892 33124 38948 33134
rect 38892 29652 38948 33068
rect 39004 32228 39060 35196
rect 39004 32162 39060 32172
rect 38892 29586 38948 29596
rect 39004 28756 39060 28766
rect 38892 28420 38948 28430
rect 38892 26964 38948 28364
rect 38892 26898 38948 26908
rect 39004 26852 39060 28700
rect 39004 26786 39060 26796
rect 38892 26740 38948 26750
rect 38892 26068 38948 26684
rect 39004 26628 39060 26638
rect 39004 26180 39060 26572
rect 39004 26114 39060 26124
rect 38892 26002 38948 26012
rect 39004 24164 39060 24174
rect 38892 22932 38948 22942
rect 38892 21700 38948 22876
rect 38892 21634 38948 21644
rect 38892 20356 38948 20366
rect 38892 13076 38948 20300
rect 38892 13010 38948 13020
rect 38892 11732 38948 11742
rect 38892 2660 38948 11676
rect 39004 9380 39060 24108
rect 39004 9314 39060 9324
rect 39116 2772 39172 55804
rect 41468 55636 41524 55646
rect 40236 55524 40292 55534
rect 39452 55412 39508 55422
rect 39228 46116 39284 46126
rect 39228 44884 39284 46060
rect 39228 44818 39284 44828
rect 39340 43876 39396 43886
rect 39340 42756 39396 43820
rect 39340 42690 39396 42700
rect 39228 32452 39284 32462
rect 39228 32116 39284 32396
rect 39228 32050 39284 32060
rect 39340 31892 39396 31902
rect 39228 28084 39284 28094
rect 39228 26740 39284 28028
rect 39228 26674 39284 26684
rect 39340 26852 39396 31836
rect 39340 26038 39396 26796
rect 39228 25982 39396 26038
rect 39228 24276 39284 25982
rect 39228 24210 39284 24220
rect 39340 25284 39396 25294
rect 39228 22708 39284 22718
rect 39228 21140 39284 22652
rect 39228 21074 39284 21084
rect 39340 11284 39396 25228
rect 39340 11218 39396 11228
rect 39116 2706 39172 2716
rect 38892 2594 38948 2604
rect 38780 1586 38836 1596
rect 37660 1138 37716 1148
rect 39452 1204 39508 55356
rect 39900 54628 39956 54638
rect 39564 45892 39620 45902
rect 39564 45220 39620 45836
rect 39564 45154 39620 45164
rect 39788 45556 39844 45566
rect 39788 43876 39844 45500
rect 39788 43810 39844 43820
rect 39676 39284 39732 39294
rect 39676 38612 39732 39228
rect 39676 38546 39732 38556
rect 39564 38276 39620 38286
rect 39564 37268 39620 38220
rect 39564 37202 39620 37212
rect 39788 37268 39844 37278
rect 39676 35588 39732 35598
rect 39676 34804 39732 35532
rect 39676 34738 39732 34748
rect 39564 34580 39620 34590
rect 39564 30212 39620 34524
rect 39676 33684 39732 33694
rect 39676 33348 39732 33628
rect 39676 33282 39732 33292
rect 39564 28644 39620 30156
rect 39564 28578 39620 28588
rect 39676 32004 39732 32014
rect 39676 30324 39732 31948
rect 39564 28196 39620 28206
rect 39676 28198 39732 30268
rect 39788 28420 39844 37212
rect 39788 28354 39844 28364
rect 39900 34916 39956 54572
rect 40124 51156 40180 51166
rect 40012 47012 40068 47022
rect 40012 44996 40068 46956
rect 40124 46564 40180 51100
rect 40124 46498 40180 46508
rect 40012 44930 40068 44940
rect 39676 28142 39844 28198
rect 39564 27860 39620 28140
rect 39564 27794 39620 27804
rect 39564 27188 39620 27198
rect 39564 23716 39620 27132
rect 39676 26404 39732 26414
rect 39676 25060 39732 26348
rect 39676 24276 39732 25004
rect 39676 24210 39732 24220
rect 39564 23650 39620 23660
rect 39676 23380 39732 23390
rect 39676 23156 39732 23324
rect 39676 23090 39732 23100
rect 39564 21924 39620 21934
rect 39564 13748 39620 21868
rect 39788 20998 39844 28142
rect 39900 21178 39956 34860
rect 40012 40068 40068 40078
rect 40012 21924 40068 40012
rect 40124 39508 40180 39518
rect 40124 39284 40180 39452
rect 40124 39218 40180 39228
rect 40124 36036 40180 36046
rect 40124 33460 40180 35980
rect 40124 33394 40180 33404
rect 40236 30212 40292 55468
rect 40684 55412 40740 55422
rect 40460 54292 40516 54302
rect 40348 52276 40404 52286
rect 40348 51268 40404 52220
rect 40348 51202 40404 51212
rect 40348 44660 40404 44670
rect 40348 42868 40404 44604
rect 40460 43092 40516 54236
rect 40460 43026 40516 43036
rect 40572 52276 40628 52286
rect 40572 46564 40628 52220
rect 40348 42802 40404 42812
rect 40348 39060 40404 39070
rect 40348 34692 40404 39004
rect 40572 36932 40628 46508
rect 40572 36866 40628 36876
rect 40348 34626 40404 34636
rect 40236 30146 40292 30156
rect 40348 34132 40404 34142
rect 40236 28980 40292 28990
rect 40124 28084 40180 28094
rect 40124 26964 40180 28028
rect 40124 26898 40180 26908
rect 40236 24276 40292 28924
rect 40236 24210 40292 24220
rect 40012 21858 40068 21868
rect 40348 22596 40404 34076
rect 40460 33908 40516 33918
rect 40460 26068 40516 33852
rect 40460 26002 40516 26012
rect 40572 27636 40628 27646
rect 40572 23156 40628 27580
rect 40572 23090 40628 23100
rect 39900 21122 40180 21178
rect 39788 20942 39956 20998
rect 39788 14308 39844 14318
rect 39788 13972 39844 14252
rect 39788 13906 39844 13916
rect 39564 13682 39620 13692
rect 39564 11284 39620 11294
rect 39564 2772 39620 11228
rect 39900 7476 39956 20942
rect 39900 7410 39956 7420
rect 39564 2706 39620 2716
rect 39788 6580 39844 6590
rect 39452 1138 39508 1148
rect 39788 196 39844 6524
rect 40124 6580 40180 21122
rect 40348 11060 40404 22540
rect 40572 22708 40628 22718
rect 40460 21924 40516 21934
rect 40460 18452 40516 21868
rect 40572 21812 40628 22652
rect 40572 21746 40628 21756
rect 40460 18386 40516 18396
rect 40572 20020 40628 20030
rect 40572 19124 40628 19964
rect 40572 12740 40628 19068
rect 40572 12674 40628 12684
rect 40348 10994 40404 11004
rect 40460 7812 40516 7822
rect 40236 7700 40292 7710
rect 40236 7476 40292 7644
rect 40236 7410 40292 7420
rect 40124 6514 40180 6524
rect 40460 6580 40516 7756
rect 40460 6514 40516 6524
rect 39900 5796 39956 5806
rect 39900 4452 39956 5740
rect 39900 4386 39956 4396
rect 40348 5796 40404 5806
rect 40348 2660 40404 5740
rect 40348 2594 40404 2604
rect 40684 2212 40740 55356
rect 41356 55076 41412 55086
rect 40908 54516 40964 54526
rect 40796 52052 40852 52062
rect 40796 48692 40852 51996
rect 40796 48626 40852 48636
rect 40908 44578 40964 54460
rect 41356 52500 41412 55020
rect 41356 52434 41412 52444
rect 41356 49812 41412 49822
rect 40796 44522 40964 44578
rect 41020 47012 41076 47022
rect 41020 45332 41076 46956
rect 40796 22078 40852 44522
rect 41020 44398 41076 45276
rect 40908 44342 41076 44398
rect 41244 44436 41300 44446
rect 40908 41412 40964 44342
rect 41020 43204 41076 43214
rect 41020 41972 41076 43148
rect 41244 42868 41300 44380
rect 41020 41906 41076 41916
rect 41132 42644 41188 42654
rect 40908 41346 40964 41356
rect 41132 36372 41188 42588
rect 41244 41636 41300 42812
rect 41356 42532 41412 49756
rect 41356 42466 41412 42476
rect 41244 37380 41300 41580
rect 41356 38500 41412 38510
rect 41356 38164 41412 38444
rect 41356 38098 41412 38108
rect 41244 37314 41300 37324
rect 41356 36932 41412 36942
rect 41132 36306 41188 36316
rect 41244 36820 41300 36830
rect 40908 35700 40964 35710
rect 40908 31892 40964 35644
rect 40908 31826 40964 31836
rect 41020 30212 41076 30222
rect 41020 23604 41076 30156
rect 41132 27524 41188 27534
rect 41132 27300 41188 27468
rect 41132 27234 41188 27244
rect 41244 25678 41300 36764
rect 41356 26964 41412 36876
rect 41468 32564 41524 55580
rect 41804 52724 41860 52734
rect 41580 51044 41636 51054
rect 41580 48916 41636 50988
rect 41804 50260 41860 52668
rect 41804 50194 41860 50204
rect 41916 51268 41972 51278
rect 41580 48850 41636 48860
rect 41804 49700 41860 49710
rect 41804 47998 41860 49644
rect 41916 48244 41972 51212
rect 42140 49700 42196 49710
rect 41916 48178 41972 48188
rect 42028 49476 42084 49486
rect 41804 47942 41972 47998
rect 41804 46676 41860 46686
rect 41692 46452 41748 46462
rect 41580 46340 41636 46350
rect 41580 42868 41636 46284
rect 41580 42802 41636 42812
rect 41580 40180 41636 40190
rect 41580 39844 41636 40124
rect 41580 33012 41636 39788
rect 41692 36932 41748 46396
rect 41804 45108 41860 46620
rect 41916 45892 41972 47942
rect 41916 45826 41972 45836
rect 41804 45042 41860 45052
rect 42028 44884 42084 49420
rect 41804 44436 41860 44446
rect 41804 38276 41860 44380
rect 41916 41300 41972 41310
rect 41916 38500 41972 41244
rect 41916 38434 41972 38444
rect 41804 37918 41860 38220
rect 41804 37862 41972 37918
rect 41692 36866 41748 36876
rect 41804 37716 41860 37726
rect 41580 32946 41636 32956
rect 41468 32498 41524 32508
rect 41692 31780 41748 31790
rect 41580 30884 41636 30894
rect 41580 27748 41636 30828
rect 41580 27682 41636 27692
rect 41412 26908 41524 26938
rect 41356 26882 41524 26908
rect 41468 26628 41524 26882
rect 41244 25622 41412 25678
rect 41244 25508 41300 25518
rect 41020 23538 41076 23548
rect 41132 24500 41188 24510
rect 40796 22022 40964 22078
rect 40796 21924 40852 21934
rect 40796 20804 40852 21868
rect 40908 21700 40964 22022
rect 40908 21634 40964 21644
rect 40796 12516 40852 20748
rect 41020 20468 41076 20478
rect 41020 19460 41076 20412
rect 41020 19394 41076 19404
rect 41132 19684 41188 24444
rect 41132 19012 41188 19628
rect 41132 18946 41188 18956
rect 41020 18788 41076 18798
rect 40908 18452 40964 18462
rect 40908 16884 40964 18396
rect 41020 18228 41076 18732
rect 41020 18162 41076 18172
rect 40908 16818 40964 16828
rect 40796 12450 40852 12460
rect 41020 14868 41076 14878
rect 40908 11172 40964 11182
rect 40908 3668 40964 11116
rect 41020 5236 41076 14812
rect 41244 12964 41300 25452
rect 41356 16212 41412 25622
rect 41356 16146 41412 16156
rect 41468 16436 41524 26572
rect 41692 25060 41748 31724
rect 41692 24994 41748 25004
rect 41580 24836 41636 24846
rect 41580 24612 41636 24780
rect 41580 24546 41636 24556
rect 41692 23940 41748 23950
rect 41580 23492 41636 23502
rect 41580 23156 41636 23436
rect 41580 23090 41636 23100
rect 41580 21700 41636 21710
rect 41580 21476 41636 21644
rect 41580 21410 41636 21420
rect 41580 21140 41636 21150
rect 41580 20468 41636 21084
rect 41580 20402 41636 20412
rect 41692 17780 41748 23884
rect 41804 21140 41860 37660
rect 41916 37268 41972 37862
rect 41916 37202 41972 37212
rect 41804 21074 41860 21084
rect 41916 33012 41972 33022
rect 41692 17714 41748 17724
rect 41356 15092 41412 15102
rect 41356 14756 41412 15036
rect 41356 14690 41412 14700
rect 41244 12898 41300 12908
rect 41468 10052 41524 16380
rect 41916 15598 41972 32956
rect 41468 9986 41524 9996
rect 41804 15542 41972 15598
rect 42028 20468 42084 44828
rect 42140 38388 42196 49644
rect 42252 45444 42308 45454
rect 42252 45108 42308 45388
rect 42252 45042 42308 45052
rect 42140 37716 42196 38332
rect 42140 37650 42196 37660
rect 42252 43092 42308 43102
rect 42252 35476 42308 43036
rect 42252 35410 42308 35420
rect 42252 28868 42308 28878
rect 42140 28084 42196 28094
rect 42140 27412 42196 28028
rect 42140 27346 42196 27356
rect 42252 24612 42308 28812
rect 41804 12964 41860 15542
rect 41916 15316 41972 15326
rect 41916 14756 41972 15260
rect 41916 14690 41972 14700
rect 41804 9838 41860 12908
rect 41356 9782 41860 9838
rect 42028 14420 42084 20412
rect 42140 21812 42196 21822
rect 42140 19684 42196 21756
rect 42140 19618 42196 19628
rect 41356 6804 41412 9782
rect 42028 7364 42084 14364
rect 42140 18116 42196 18126
rect 42140 12516 42196 18060
rect 42252 16498 42308 24556
rect 42364 16772 42420 56028
rect 42700 53060 42756 53070
rect 42476 46452 42532 46462
rect 42476 46198 42532 46396
rect 42476 46142 42644 46198
rect 42476 46004 42532 46014
rect 42476 36708 42532 45948
rect 42588 45332 42644 46142
rect 42588 45266 42644 45276
rect 42700 44660 42756 53004
rect 42700 44594 42756 44604
rect 42588 40516 42644 40526
rect 42588 39732 42644 40460
rect 42588 39666 42644 39676
rect 42476 36642 42532 36652
rect 42700 37380 42756 37390
rect 42700 36596 42756 37324
rect 42700 33236 42756 36540
rect 42700 33170 42756 33180
rect 42700 33012 42756 33022
rect 42588 30436 42644 30446
rect 42476 28308 42532 28318
rect 42476 27972 42532 28252
rect 42476 23268 42532 27916
rect 42588 25508 42644 30380
rect 42700 26292 42756 32956
rect 42700 26226 42756 26236
rect 42588 25442 42644 25452
rect 42476 23202 42532 23212
rect 42588 22372 42644 22382
rect 42588 20804 42644 22316
rect 42588 20738 42644 20748
rect 42700 21812 42756 21822
rect 42364 16706 42420 16716
rect 42588 16772 42644 16782
rect 42252 16442 42532 16498
rect 42140 12450 42196 12460
rect 42028 7298 42084 7308
rect 42140 10164 42196 10174
rect 41356 6738 41412 6748
rect 41580 7140 41636 7150
rect 41580 6692 41636 7084
rect 41580 6626 41636 6636
rect 41020 5170 41076 5180
rect 40908 3602 40964 3612
rect 40684 2146 40740 2156
rect 40908 2996 40964 3006
rect 40908 1764 40964 2940
rect 42140 2772 42196 10108
rect 42476 8372 42532 16442
rect 42588 11508 42644 16716
rect 42700 14868 42756 21756
rect 42700 14802 42756 14812
rect 42588 11442 42644 11452
rect 42476 8306 42532 8316
rect 42364 7364 42420 7374
rect 42364 3220 42420 7308
rect 42812 5012 42868 56364
rect 43776 56420 43804 56476
rect 43860 56420 43908 56476
rect 43964 56420 44012 56476
rect 44068 56420 44096 56476
rect 43036 55972 43092 55982
rect 43036 52388 43092 55916
rect 43036 52322 43092 52332
rect 43260 55636 43316 55646
rect 43148 50372 43204 50382
rect 43148 49700 43204 50316
rect 43148 49634 43204 49644
rect 43148 47908 43204 47918
rect 42924 44660 42980 44670
rect 42924 11998 42980 44604
rect 43148 43204 43204 47852
rect 43148 43138 43204 43148
rect 43036 35588 43092 35598
rect 43036 16772 43092 35532
rect 43148 27972 43204 27982
rect 43148 19908 43204 27916
rect 43148 19842 43204 19852
rect 43036 16706 43092 16716
rect 43260 15418 43316 55580
rect 43776 54908 44096 56420
rect 44268 56868 44324 56878
rect 44156 56308 44212 56318
rect 44156 55748 44212 56252
rect 44156 55682 44212 55692
rect 43484 54852 43540 54862
rect 43372 54068 43428 54078
rect 43372 53284 43428 54012
rect 43484 53956 43540 54796
rect 43484 53890 43540 53900
rect 43776 54852 43804 54908
rect 43860 54852 43908 54908
rect 43964 54852 44012 54908
rect 44068 54852 44096 54908
rect 43372 53218 43428 53228
rect 43596 53844 43652 53854
rect 43372 52724 43428 52734
rect 43372 51156 43428 52668
rect 43372 50484 43428 51100
rect 43372 50418 43428 50428
rect 43484 51044 43540 51054
rect 43372 47012 43428 47022
rect 43372 28532 43428 46956
rect 43372 28466 43428 28476
rect 43372 27748 43428 27758
rect 43372 25732 43428 27692
rect 43372 25666 43428 25676
rect 43372 21812 43428 21822
rect 43372 15652 43428 21756
rect 43372 15586 43428 15596
rect 43036 15362 43316 15418
rect 43036 12358 43092 15362
rect 43148 14532 43204 14542
rect 43148 13258 43204 14476
rect 43484 14196 43540 50988
rect 43596 50596 43652 53788
rect 43596 50530 43652 50540
rect 43776 53340 44096 54852
rect 43776 53284 43804 53340
rect 43860 53284 43908 53340
rect 43964 53284 44012 53340
rect 44068 53284 44096 53340
rect 43776 51772 44096 53284
rect 43776 51716 43804 51772
rect 43860 51716 43908 51772
rect 43964 51716 44012 51772
rect 44068 51716 44096 51772
rect 43776 50204 44096 51716
rect 43776 50148 43804 50204
rect 43860 50148 43908 50204
rect 43964 50148 44012 50204
rect 44068 50148 44096 50204
rect 44156 55300 44212 55310
rect 44156 50260 44212 55244
rect 44268 51044 44324 56812
rect 44268 50978 44324 50988
rect 44436 55692 44756 57456
rect 46844 57428 46900 57438
rect 45276 57316 45332 57326
rect 44436 55636 44464 55692
rect 44520 55636 44568 55692
rect 44624 55636 44672 55692
rect 44728 55636 44756 55692
rect 44436 54124 44756 55636
rect 44436 54068 44464 54124
rect 44520 54068 44568 54124
rect 44624 54068 44672 54124
rect 44728 54068 44756 54124
rect 44436 52556 44756 54068
rect 44436 52500 44464 52556
rect 44520 52500 44568 52556
rect 44624 52500 44672 52556
rect 44728 52500 44756 52556
rect 44436 50988 44756 52500
rect 44436 50932 44464 50988
rect 44520 50932 44568 50988
rect 44624 50932 44672 50988
rect 44728 50932 44756 50988
rect 44156 50194 44212 50204
rect 44268 50596 44324 50606
rect 43776 48636 44096 50148
rect 43776 48580 43804 48636
rect 43860 48580 43908 48636
rect 43964 48580 44012 48636
rect 44068 48580 44096 48636
rect 43596 47908 43652 47918
rect 43596 47684 43652 47852
rect 43596 47618 43652 47628
rect 43596 47460 43652 47470
rect 43596 41188 43652 47404
rect 43596 41122 43652 41132
rect 43776 47068 44096 48580
rect 44156 48916 44212 48926
rect 44156 48580 44212 48860
rect 44156 48514 44212 48524
rect 43776 47012 43804 47068
rect 43860 47012 43908 47068
rect 43964 47012 44012 47068
rect 44068 47012 44096 47068
rect 44268 47572 44324 50540
rect 43776 45500 44096 47012
rect 44156 47012 44212 47022
rect 44156 46340 44212 46956
rect 44156 46274 44212 46284
rect 43776 45444 43804 45500
rect 43860 45444 43908 45500
rect 43964 45444 44012 45500
rect 44068 45444 44096 45500
rect 43776 43932 44096 45444
rect 43776 43876 43804 43932
rect 43860 43876 43908 43932
rect 43964 43876 44012 43932
rect 44068 43876 44096 43932
rect 43776 42364 44096 43876
rect 44156 44212 44212 44222
rect 44156 43876 44212 44156
rect 44156 43810 44212 43820
rect 43776 42308 43804 42364
rect 43860 42308 43908 42364
rect 43964 42308 44012 42364
rect 44068 42308 44096 42364
rect 43776 40796 44096 42308
rect 44156 42308 44212 42318
rect 44156 41636 44212 42252
rect 44156 41570 44212 41580
rect 43776 40740 43804 40796
rect 43860 40740 43908 40796
rect 43964 40740 44012 40796
rect 44068 40740 44096 40796
rect 43776 39228 44096 40740
rect 43776 39172 43804 39228
rect 43860 39172 43908 39228
rect 43964 39172 44012 39228
rect 44068 39172 44096 39228
rect 43776 37660 44096 39172
rect 43776 37604 43804 37660
rect 43860 37604 43908 37660
rect 43964 37604 44012 37660
rect 44068 37604 44096 37660
rect 43596 37044 43652 37054
rect 43596 36036 43652 36988
rect 43596 35970 43652 35980
rect 43776 36092 44096 37604
rect 44156 41188 44212 41198
rect 44156 36932 44212 41132
rect 44156 36866 44212 36876
rect 43776 36036 43804 36092
rect 43860 36036 43908 36092
rect 43964 36036 44012 36092
rect 44068 36036 44096 36092
rect 43776 34524 44096 36036
rect 43776 34468 43804 34524
rect 43860 34468 43908 34524
rect 43964 34468 44012 34524
rect 44068 34468 44096 34524
rect 43596 33348 43652 33358
rect 43596 32452 43652 33292
rect 43596 32386 43652 32396
rect 43776 32956 44096 34468
rect 43776 32900 43804 32956
rect 43860 32900 43908 32956
rect 43964 32900 44012 32956
rect 44068 32900 44096 32956
rect 43776 31388 44096 32900
rect 43776 31332 43804 31388
rect 43860 31332 43908 31388
rect 43964 31332 44012 31388
rect 44068 31332 44096 31388
rect 43776 29820 44096 31332
rect 44156 32228 44212 32238
rect 44156 31332 44212 32172
rect 44156 31266 44212 31276
rect 44156 31108 44212 31118
rect 44156 30660 44212 31052
rect 44156 30594 44212 30604
rect 43776 29764 43804 29820
rect 43860 29764 43908 29820
rect 43964 29764 44012 29820
rect 44068 29764 44096 29820
rect 43776 28252 44096 29764
rect 43776 28196 43804 28252
rect 43860 28196 43908 28252
rect 43964 28196 44012 28252
rect 44068 28196 44096 28252
rect 43596 27748 43652 27758
rect 43596 27188 43652 27692
rect 43596 27122 43652 27132
rect 43776 26684 44096 28196
rect 43776 26628 43804 26684
rect 43860 26628 43908 26684
rect 43964 26628 44012 26684
rect 44068 26628 44096 26684
rect 43776 25116 44096 26628
rect 44156 28980 44212 28990
rect 44156 26404 44212 28924
rect 44268 28868 44324 47516
rect 44268 28802 44324 28812
rect 44436 49420 44756 50932
rect 44436 49364 44464 49420
rect 44520 49364 44568 49420
rect 44624 49364 44672 49420
rect 44728 49364 44756 49420
rect 44436 47852 44756 49364
rect 44436 47796 44464 47852
rect 44520 47796 44568 47852
rect 44624 47796 44672 47852
rect 44728 47796 44756 47852
rect 44436 46284 44756 47796
rect 44436 46228 44464 46284
rect 44520 46228 44568 46284
rect 44624 46228 44672 46284
rect 44728 46228 44756 46284
rect 44436 44716 44756 46228
rect 44436 44660 44464 44716
rect 44520 44660 44568 44716
rect 44624 44660 44672 44716
rect 44728 44660 44756 44716
rect 44436 43148 44756 44660
rect 44436 43092 44464 43148
rect 44520 43092 44568 43148
rect 44624 43092 44672 43148
rect 44728 43092 44756 43148
rect 44436 41580 44756 43092
rect 44436 41524 44464 41580
rect 44520 41524 44568 41580
rect 44624 41524 44672 41580
rect 44728 41524 44756 41580
rect 44436 40012 44756 41524
rect 44436 39956 44464 40012
rect 44520 39956 44568 40012
rect 44624 39956 44672 40012
rect 44728 39956 44756 40012
rect 44436 38444 44756 39956
rect 44436 38388 44464 38444
rect 44520 38388 44568 38444
rect 44624 38388 44672 38444
rect 44728 38388 44756 38444
rect 44436 36876 44756 38388
rect 44436 36820 44464 36876
rect 44520 36820 44568 36876
rect 44624 36820 44672 36876
rect 44728 36820 44756 36876
rect 44436 35308 44756 36820
rect 44436 35252 44464 35308
rect 44520 35252 44568 35308
rect 44624 35252 44672 35308
rect 44728 35252 44756 35308
rect 44436 33740 44756 35252
rect 44436 33684 44464 33740
rect 44520 33684 44568 33740
rect 44624 33684 44672 33740
rect 44728 33684 44756 33740
rect 44436 32172 44756 33684
rect 44436 32116 44464 32172
rect 44520 32116 44568 32172
rect 44624 32116 44672 32172
rect 44728 32116 44756 32172
rect 44436 30604 44756 32116
rect 44436 30548 44464 30604
rect 44520 30548 44568 30604
rect 44624 30548 44672 30604
rect 44728 30548 44756 30604
rect 44436 29036 44756 30548
rect 44436 28980 44464 29036
rect 44520 28980 44568 29036
rect 44624 28980 44672 29036
rect 44728 28980 44756 29036
rect 44268 28532 44324 28542
rect 44268 26628 44324 28476
rect 44268 26562 44324 26572
rect 44436 27468 44756 28980
rect 44436 27412 44464 27468
rect 44520 27412 44568 27468
rect 44624 27412 44672 27468
rect 44728 27412 44756 27468
rect 44156 26338 44212 26348
rect 44436 25900 44756 27412
rect 44436 25844 44464 25900
rect 44520 25844 44568 25900
rect 44624 25844 44672 25900
rect 44728 25844 44756 25900
rect 43776 25060 43804 25116
rect 43860 25060 43908 25116
rect 43964 25060 44012 25116
rect 44068 25060 44096 25116
rect 43776 23548 44096 25060
rect 44156 25172 44212 25182
rect 44156 24276 44212 25116
rect 44156 23698 44212 24220
rect 44268 24948 44324 24958
rect 44268 24164 44324 24892
rect 44268 24098 44324 24108
rect 44436 24332 44756 25844
rect 44436 24276 44464 24332
rect 44520 24276 44568 24332
rect 44624 24276 44672 24332
rect 44728 24276 44756 24332
rect 44156 23642 44324 23698
rect 43776 23492 43804 23548
rect 43860 23492 43908 23548
rect 43964 23492 44012 23548
rect 44068 23492 44096 23548
rect 43776 21980 44096 23492
rect 44156 23492 44212 23502
rect 44156 23268 44212 23436
rect 44156 23202 44212 23212
rect 44156 23044 44212 23054
rect 44156 22708 44212 22988
rect 44156 22642 44212 22652
rect 43776 21924 43804 21980
rect 43860 21924 43908 21980
rect 43964 21924 44012 21980
rect 44068 21924 44096 21980
rect 43596 20916 43652 20926
rect 43596 20468 43652 20860
rect 43596 20402 43652 20412
rect 43776 20412 44096 21924
rect 44268 21358 44324 23642
rect 43776 20356 43804 20412
rect 43860 20356 43908 20412
rect 43964 20356 44012 20412
rect 44068 20356 44096 20412
rect 43776 18844 44096 20356
rect 43776 18788 43804 18844
rect 43860 18788 43908 18844
rect 43964 18788 44012 18844
rect 44068 18788 44096 18844
rect 43776 17276 44096 18788
rect 43776 17220 43804 17276
rect 43860 17220 43908 17276
rect 43964 17220 44012 17276
rect 44068 17220 44096 17276
rect 43776 15708 44096 17220
rect 43776 15652 43804 15708
rect 43860 15652 43908 15708
rect 43964 15652 44012 15708
rect 44068 15652 44096 15708
rect 43484 14130 43540 14140
rect 43596 14420 43652 14430
rect 43596 14084 43652 14364
rect 43596 14018 43652 14028
rect 43776 14140 44096 15652
rect 43776 14084 43804 14140
rect 43860 14084 43908 14140
rect 43964 14084 44012 14140
rect 44068 14084 44096 14140
rect 43372 13860 43428 13870
rect 43372 13412 43428 13804
rect 43372 13346 43428 13356
rect 43148 13202 43652 13258
rect 43260 12964 43316 12974
rect 43260 12898 43316 12908
rect 43260 12842 43540 12898
rect 43484 12740 43540 12842
rect 43484 12674 43540 12684
rect 43148 12628 43204 12638
rect 43148 12538 43204 12572
rect 43148 12482 43540 12538
rect 43036 12302 43316 12358
rect 42924 11942 43092 11998
rect 42924 11844 42980 11854
rect 42924 6916 42980 11788
rect 42924 6850 42980 6860
rect 43036 9828 43092 11942
rect 43036 6692 43092 9772
rect 43036 6626 43092 6636
rect 42812 4946 42868 4956
rect 42364 3154 42420 3164
rect 42140 2706 42196 2716
rect 43260 2212 43316 12302
rect 43372 9268 43428 9278
rect 43372 8820 43428 9212
rect 43372 8754 43428 8764
rect 43484 3332 43540 12482
rect 43596 5124 43652 13202
rect 43596 5058 43652 5068
rect 43776 12572 44096 14084
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 43776 11004 44096 12516
rect 44156 21302 44324 21358
rect 44436 22764 44756 24276
rect 44436 22708 44464 22764
rect 44520 22708 44568 22764
rect 44624 22708 44672 22764
rect 44728 22708 44756 22764
rect 44156 11396 44212 21302
rect 44436 21196 44756 22708
rect 44436 21140 44464 21196
rect 44520 21140 44568 21196
rect 44624 21140 44672 21196
rect 44728 21140 44756 21196
rect 44268 20132 44324 20142
rect 44268 19124 44324 20076
rect 44268 19058 44324 19068
rect 44436 19628 44756 21140
rect 44436 19572 44464 19628
rect 44520 19572 44568 19628
rect 44624 19572 44672 19628
rect 44728 19572 44756 19628
rect 44268 18452 44324 18462
rect 44268 16548 44324 18396
rect 44268 16482 44324 16492
rect 44436 18060 44756 19572
rect 44436 18004 44464 18060
rect 44520 18004 44568 18060
rect 44624 18004 44672 18060
rect 44728 18004 44756 18060
rect 44436 16492 44756 18004
rect 44436 16436 44464 16492
rect 44520 16436 44568 16492
rect 44624 16436 44672 16492
rect 44728 16436 44756 16492
rect 44156 11330 44212 11340
rect 44268 15092 44324 15102
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 43776 9436 44096 10948
rect 44156 10388 44212 10398
rect 44156 9828 44212 10332
rect 44156 9762 44212 9772
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 43776 6300 44096 7812
rect 44156 7812 44212 7822
rect 44156 7140 44212 7756
rect 44156 7074 44212 7084
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 44268 6580 44324 15036
rect 43596 4788 43652 4798
rect 43596 4116 43652 4732
rect 43596 4050 43652 4060
rect 43776 4732 44096 6244
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 43484 3266 43540 3276
rect 43260 2146 43316 2156
rect 43776 3164 44096 4676
rect 44156 6244 44212 6254
rect 44156 3892 44212 6188
rect 44268 5572 44324 6524
rect 44268 5124 44324 5516
rect 44268 5058 44324 5068
rect 44436 14924 44756 16436
rect 44436 14868 44464 14924
rect 44520 14868 44568 14924
rect 44624 14868 44672 14924
rect 44728 14868 44756 14924
rect 44436 13356 44756 14868
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44156 3826 44212 3836
rect 44268 4004 44324 4014
rect 44268 3444 44324 3948
rect 44268 3378 44324 3388
rect 44436 3948 44756 5460
rect 44828 56644 44884 56654
rect 44828 5460 44884 56588
rect 44940 55860 44996 55870
rect 44940 38500 44996 55804
rect 44940 38434 44996 38444
rect 45052 55636 45108 55646
rect 44940 32788 44996 32798
rect 44940 32452 44996 32732
rect 44940 32386 44996 32396
rect 44940 29988 44996 29998
rect 44940 25172 44996 29932
rect 44940 25106 44996 25116
rect 44940 16996 44996 17006
rect 44940 16436 44996 16940
rect 44940 16370 44996 16380
rect 44940 15988 44996 15998
rect 44940 15652 44996 15932
rect 44940 15586 44996 15596
rect 44940 15092 44996 15102
rect 44940 14532 44996 15036
rect 44940 14466 44996 14476
rect 44940 14084 44996 14094
rect 44940 12740 44996 14028
rect 44940 12674 44996 12684
rect 44940 11284 44996 11294
rect 44940 6468 44996 11228
rect 44940 6402 44996 6412
rect 44828 4900 44884 5404
rect 44940 5796 44996 5806
rect 44940 5124 44996 5740
rect 44940 5058 44996 5068
rect 44828 4834 44884 4844
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 40908 1698 40964 1708
rect 39788 130 39844 140
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 36764 18 36820 28
rect 43776 0 44096 1540
rect 44436 2380 44756 3892
rect 45052 3668 45108 55580
rect 45164 53172 45220 53182
rect 45164 51492 45220 53116
rect 45164 51426 45220 51436
rect 45164 50260 45220 50270
rect 45164 46564 45220 50204
rect 45164 46498 45220 46508
rect 45164 42980 45220 42990
rect 45164 41188 45220 42924
rect 45164 41122 45220 41132
rect 45164 40068 45220 40078
rect 45164 39732 45220 40012
rect 45164 39666 45220 39676
rect 45164 38724 45220 38734
rect 45164 30100 45220 38668
rect 45164 30034 45220 30044
rect 45164 28308 45220 28318
rect 45164 27972 45220 28252
rect 45164 27300 45220 27916
rect 45164 27234 45220 27244
rect 45164 19796 45220 19806
rect 45164 19460 45220 19740
rect 45164 19394 45220 19404
rect 45164 16996 45220 17006
rect 45164 16100 45220 16940
rect 45164 16034 45220 16044
rect 45164 15316 45220 15326
rect 45164 13076 45220 15260
rect 45164 13010 45220 13020
rect 45164 8820 45220 8830
rect 45164 6244 45220 8764
rect 45164 6178 45220 6188
rect 45052 3602 45108 3612
rect 45276 2548 45332 57260
rect 46844 57092 46900 57372
rect 46844 57026 46900 57036
rect 48524 57428 48580 57438
rect 46284 56196 46340 56206
rect 45948 55972 46004 55982
rect 45500 55636 45556 55646
rect 45388 54852 45444 54862
rect 45388 49028 45444 54796
rect 45388 48962 45444 48972
rect 45388 42308 45444 42318
rect 45388 39956 45444 42252
rect 45388 39890 45444 39900
rect 45500 38458 45556 55580
rect 45724 53060 45780 53070
rect 45612 52164 45668 52174
rect 45612 45444 45668 52108
rect 45724 49438 45780 53004
rect 45948 53060 46004 55916
rect 45948 52994 46004 53004
rect 46060 55524 46116 55534
rect 45948 51380 46004 51390
rect 45948 50484 46004 51324
rect 45948 50418 46004 50428
rect 45724 49382 45892 49438
rect 45724 49252 45780 49262
rect 45724 48804 45780 49196
rect 45836 48916 45892 49382
rect 45836 48850 45892 48860
rect 45724 48738 45780 48748
rect 45612 45378 45668 45388
rect 45836 44436 45892 44446
rect 45836 42644 45892 44380
rect 45836 42578 45892 42588
rect 45948 39508 46004 39518
rect 45948 38836 46004 39452
rect 45948 38770 46004 38780
rect 45500 38402 45780 38458
rect 45612 32564 45668 32574
rect 45500 31332 45556 31342
rect 45388 28196 45444 28206
rect 45388 26740 45444 28140
rect 45388 25844 45444 26684
rect 45388 25778 45444 25788
rect 45500 25732 45556 31276
rect 45612 27076 45668 32508
rect 45612 27010 45668 27020
rect 45500 25666 45556 25676
rect 45724 20998 45780 38402
rect 45836 37940 45892 37950
rect 45836 31780 45892 37884
rect 45836 31714 45892 31724
rect 45948 33572 46004 33582
rect 45948 29540 46004 33516
rect 45500 20942 45780 20998
rect 45836 24500 45892 24510
rect 45388 20692 45444 20702
rect 45388 15316 45444 20636
rect 45388 15250 45444 15260
rect 45388 9604 45444 9614
rect 45388 4004 45444 9548
rect 45500 4564 45556 20942
rect 45836 17578 45892 24444
rect 45948 23044 46004 29484
rect 45948 22978 46004 22988
rect 45724 17522 45892 17578
rect 45948 21812 46004 21822
rect 45612 16436 45668 16446
rect 45612 12516 45668 16380
rect 45612 12450 45668 12460
rect 45724 10052 45780 17522
rect 45948 17332 46004 21756
rect 45948 17266 46004 17276
rect 45836 16996 45892 17006
rect 45836 11956 45892 16940
rect 45948 16884 46004 16894
rect 45948 14868 46004 16828
rect 45948 14802 46004 14812
rect 45836 11890 45892 11900
rect 45724 9986 45780 9996
rect 45724 6916 45780 6926
rect 45724 6692 45780 6860
rect 45724 6626 45780 6636
rect 45500 4498 45556 4508
rect 45388 3938 45444 3948
rect 46060 3892 46116 55468
rect 46172 54516 46228 54526
rect 46172 35252 46228 54460
rect 46172 35186 46228 35196
rect 46172 30100 46228 30110
rect 46172 14532 46228 30044
rect 46172 14466 46228 14476
rect 46060 3826 46116 3836
rect 45276 2482 45332 2492
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 46284 2212 46340 56140
rect 47404 55860 47460 55870
rect 46844 55524 46900 55534
rect 46396 55300 46452 55310
rect 46396 35476 46452 55244
rect 46620 48916 46676 48926
rect 46620 42868 46676 48860
rect 46508 41972 46564 41982
rect 46508 36820 46564 41916
rect 46508 36754 46564 36764
rect 46396 34132 46452 35420
rect 46396 34066 46452 34076
rect 46508 36260 46564 36270
rect 46508 23156 46564 36204
rect 46508 23090 46564 23100
rect 46508 21588 46564 21598
rect 46396 18900 46452 18910
rect 46396 14084 46452 18844
rect 46508 16100 46564 21532
rect 46620 20804 46676 42812
rect 46732 36820 46788 36830
rect 46732 36036 46788 36764
rect 46732 35970 46788 35980
rect 46732 34804 46788 34814
rect 46732 33572 46788 34748
rect 46732 33506 46788 33516
rect 46732 30660 46788 30670
rect 46732 22036 46788 30604
rect 46732 21970 46788 21980
rect 46620 20738 46676 20748
rect 46508 16034 46564 16044
rect 46620 19348 46676 19358
rect 46396 14018 46452 14028
rect 46508 15428 46564 15438
rect 46508 12628 46564 15372
rect 46508 12562 46564 12572
rect 46620 12180 46676 19292
rect 46620 12114 46676 12124
rect 46732 15428 46788 15438
rect 46732 11844 46788 15372
rect 46732 11778 46788 11788
rect 46844 5012 46900 55468
rect 47292 55524 47348 55534
rect 46956 46452 47012 46462
rect 46956 41972 47012 46396
rect 46956 41906 47012 41916
rect 47180 46340 47236 46350
rect 46956 41188 47012 41198
rect 46956 36260 47012 41132
rect 46956 36194 47012 36204
rect 47068 39956 47124 39966
rect 47068 39396 47124 39900
rect 47180 39844 47236 46284
rect 47180 39778 47236 39788
rect 46956 34692 47012 34702
rect 46956 34244 47012 34636
rect 46956 34178 47012 34188
rect 47068 31892 47124 39340
rect 47292 38724 47348 55468
rect 47292 38658 47348 38668
rect 47404 36820 47460 55804
rect 48188 54964 48244 54974
rect 47404 36754 47460 36764
rect 47516 53732 47572 53742
rect 47516 36148 47572 53676
rect 48188 47638 48244 54908
rect 48524 54740 48580 57372
rect 55804 56756 55860 56766
rect 48524 54674 48580 54684
rect 48636 56532 48692 56542
rect 48524 54068 48580 54078
rect 48524 53620 48580 54012
rect 48524 53554 48580 53564
rect 48300 52724 48356 52734
rect 48300 48244 48356 52668
rect 48636 52612 48692 56476
rect 52444 56532 52500 56542
rect 52108 55860 52164 55870
rect 48972 55524 49028 55534
rect 48636 52546 48692 52556
rect 48860 54068 48916 54078
rect 48300 48178 48356 48188
rect 48412 52500 48468 52510
rect 47964 47582 48244 47638
rect 47964 47348 48020 47582
rect 47964 47282 48020 47292
rect 48188 47348 48244 47358
rect 47628 45332 47684 45342
rect 47628 42196 47684 45276
rect 47628 42130 47684 42140
rect 47852 43428 47908 43438
rect 47292 35476 47348 35486
rect 47292 34804 47348 35420
rect 47292 34738 47348 34748
rect 47180 34356 47236 34366
rect 47180 33908 47236 34300
rect 47180 33842 47236 33852
rect 47292 34244 47348 34254
rect 47292 33684 47348 34188
rect 47292 33618 47348 33628
rect 47516 33598 47572 36092
rect 47852 38500 47908 43372
rect 48076 42308 48132 42318
rect 47740 35252 47796 35262
rect 47404 33542 47572 33598
rect 47628 33628 47684 33638
rect 47068 31826 47124 31836
rect 47292 32564 47348 32574
rect 47292 31220 47348 32508
rect 47292 31154 47348 31164
rect 47068 30996 47124 31006
rect 47068 30324 47124 30940
rect 47068 30258 47124 30268
rect 47404 30548 47460 33542
rect 46956 24500 47012 24510
rect 46956 11172 47012 24444
rect 47068 21812 47124 21822
rect 47068 17780 47124 21756
rect 47404 19908 47460 30492
rect 47628 32004 47684 33572
rect 47404 19842 47460 19852
rect 47516 28644 47572 28654
rect 47068 17714 47124 17724
rect 47292 17556 47348 17566
rect 46956 11106 47012 11116
rect 47068 15988 47124 15998
rect 47068 10198 47124 15932
rect 47292 15598 47348 17500
rect 47180 15542 47348 15598
rect 47404 17220 47460 17230
rect 47180 13748 47236 15542
rect 47180 13682 47236 13692
rect 47404 13076 47460 17164
rect 47516 13188 47572 28588
rect 47628 22820 47684 31948
rect 47628 22754 47684 22764
rect 47628 20356 47684 20366
rect 47628 17668 47684 20300
rect 47628 17602 47684 17612
rect 47516 13122 47572 13132
rect 47628 14980 47684 14990
rect 47404 13010 47460 13020
rect 47292 12628 47348 12638
rect 47292 11956 47348 12572
rect 47292 11890 47348 11900
rect 47628 11060 47684 14924
rect 47628 10994 47684 11004
rect 47068 10142 47236 10198
rect 47068 9828 47124 9838
rect 47068 5572 47124 9772
rect 47180 9716 47236 10142
rect 47180 9650 47236 9660
rect 47068 5506 47124 5516
rect 46844 4946 46900 4956
rect 46284 2146 46340 2156
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
rect 47740 756 47796 35196
rect 47852 28308 47908 38444
rect 47964 41748 48020 41758
rect 47964 40964 48020 41692
rect 47964 33684 48020 40908
rect 48076 40404 48132 42252
rect 48076 40338 48132 40348
rect 47964 33618 48020 33628
rect 48076 38724 48132 38734
rect 47964 32228 48020 32238
rect 47964 30100 48020 32172
rect 47964 30034 48020 30044
rect 47852 28242 47908 28252
rect 47852 23156 47908 23166
rect 47852 18004 47908 23100
rect 47964 21476 48020 21486
rect 47964 19236 48020 21420
rect 47964 19170 48020 19180
rect 47852 17938 47908 17948
rect 47964 18788 48020 18798
rect 47964 14196 48020 18732
rect 47964 14130 48020 14140
rect 47852 13636 47908 13646
rect 47852 12068 47908 13580
rect 47852 12002 47908 12012
rect 47964 9604 48020 9614
rect 47964 8260 48020 9548
rect 47964 4900 48020 8204
rect 47964 4834 48020 4844
rect 48076 2212 48132 38668
rect 48188 26068 48244 47292
rect 48188 26002 48244 26012
rect 48300 47012 48356 47022
rect 48300 46452 48356 46956
rect 48300 30548 48356 46396
rect 48412 38164 48468 52444
rect 48860 52500 48916 54012
rect 48860 52434 48916 52444
rect 48524 50596 48580 50606
rect 48524 44996 48580 50540
rect 48748 50260 48804 50270
rect 48524 44930 48580 44940
rect 48636 48916 48692 48926
rect 48524 43988 48580 43998
rect 48524 42980 48580 43932
rect 48524 42914 48580 42924
rect 48524 40516 48580 40526
rect 48524 39396 48580 40460
rect 48524 39330 48580 39340
rect 48412 38098 48468 38108
rect 48524 35364 48580 35374
rect 48188 21364 48244 21374
rect 48188 15652 48244 21308
rect 48188 15586 48244 15596
rect 48076 2146 48132 2156
rect 48188 14756 48244 14766
rect 48188 10724 48244 14700
rect 48188 1876 48244 10668
rect 48300 13300 48356 30492
rect 48412 33572 48468 33582
rect 48412 22372 48468 33516
rect 48524 30436 48580 35308
rect 48636 34020 48692 48860
rect 48748 48356 48804 50204
rect 48748 48290 48804 48300
rect 48748 46340 48804 46350
rect 48748 45556 48804 46284
rect 48748 45490 48804 45500
rect 48860 45668 48916 45678
rect 48748 44436 48804 44446
rect 48748 43988 48804 44380
rect 48748 43922 48804 43932
rect 48860 41524 48916 45612
rect 48860 41458 48916 41468
rect 48636 33954 48692 33964
rect 48748 36484 48804 36494
rect 48524 30370 48580 30380
rect 48412 22306 48468 22316
rect 48524 29764 48580 29774
rect 48524 22596 48580 29708
rect 48748 29652 48804 36428
rect 48860 30660 48916 30670
rect 48860 29764 48916 30604
rect 48860 29698 48916 29708
rect 48748 29586 48804 29596
rect 48524 16772 48580 22540
rect 48636 28532 48692 28542
rect 48636 21476 48692 28476
rect 48860 27748 48916 27758
rect 48636 21140 48692 21420
rect 48636 21074 48692 21084
rect 48748 23044 48804 23054
rect 48524 16706 48580 16716
rect 48636 20132 48692 20142
rect 48524 14756 48580 14766
rect 48524 13636 48580 14700
rect 48524 13570 48580 13580
rect 48300 7700 48356 13244
rect 48412 13524 48468 13534
rect 48412 11060 48468 13468
rect 48524 13300 48580 13310
rect 48524 12068 48580 13244
rect 48524 12002 48580 12012
rect 48636 11396 48692 20076
rect 48636 11330 48692 11340
rect 48412 10994 48468 11004
rect 48300 7634 48356 7644
rect 48412 2884 48468 2894
rect 48412 2548 48468 2828
rect 48748 2660 48804 22988
rect 48860 20132 48916 27692
rect 48860 20066 48916 20076
rect 48972 20098 49028 55468
rect 49420 55524 49476 55534
rect 49196 52724 49252 52734
rect 49196 48468 49252 52668
rect 49196 48402 49252 48412
rect 49308 48244 49364 48254
rect 49084 47124 49140 47134
rect 49084 46228 49140 47068
rect 49084 46162 49140 46172
rect 49196 46900 49252 46910
rect 49084 46004 49140 46014
rect 49084 36372 49140 45948
rect 49196 45892 49252 46844
rect 49196 45826 49252 45836
rect 49196 44996 49252 45006
rect 49196 42644 49252 44940
rect 49196 42578 49252 42588
rect 49196 41748 49252 41758
rect 49196 37044 49252 41692
rect 49308 40292 49364 48188
rect 49420 46788 49476 55468
rect 49980 55524 50036 55534
rect 49644 52052 49700 52062
rect 49420 46722 49476 46732
rect 49532 50484 49588 50494
rect 49532 46004 49588 50428
rect 49644 50372 49700 51996
rect 49644 50306 49700 50316
rect 49868 51604 49924 51614
rect 49644 46900 49700 46910
rect 49644 46738 49700 46844
rect 49644 46682 49812 46738
rect 49532 45938 49588 45948
rect 49644 46452 49700 46462
rect 49308 39172 49364 40236
rect 49308 39106 49364 39116
rect 49308 38276 49364 38286
rect 49308 37828 49364 38220
rect 49308 37762 49364 37772
rect 49196 36978 49252 36988
rect 49084 36306 49140 36316
rect 49308 33572 49364 33582
rect 49084 33348 49140 33358
rect 49084 31108 49140 33292
rect 49196 32340 49252 32350
rect 49196 31444 49252 32284
rect 49196 31378 49252 31388
rect 49084 31042 49140 31052
rect 49308 24388 49364 33516
rect 49420 32788 49476 32798
rect 49420 28980 49476 32732
rect 49420 28914 49476 28924
rect 49644 25732 49700 46396
rect 49756 45556 49812 46682
rect 49868 46340 49924 51548
rect 49980 49252 50036 55468
rect 50876 55524 50932 55534
rect 50092 54516 50148 54526
rect 50092 53060 50148 54460
rect 50092 52994 50148 53004
rect 50764 53732 50820 53742
rect 50092 51604 50148 51614
rect 50092 50932 50148 51548
rect 50204 51492 50260 51502
rect 50204 51156 50260 51436
rect 50204 51090 50260 51100
rect 50316 51380 50372 51390
rect 50316 50878 50372 51324
rect 50092 50866 50148 50876
rect 50204 50822 50372 50878
rect 50428 50932 50484 50942
rect 50204 50820 50260 50822
rect 50204 50754 50260 50764
rect 49980 49186 50036 49196
rect 50092 47796 50148 47806
rect 49868 46274 49924 46284
rect 49980 47572 50036 47582
rect 49756 45490 49812 45500
rect 49868 46004 49924 46014
rect 49756 44884 49812 44894
rect 49756 29988 49812 44828
rect 49868 41636 49924 45948
rect 49868 41570 49924 41580
rect 49868 41300 49924 41310
rect 49868 40628 49924 41244
rect 49868 40562 49924 40572
rect 49756 29922 49812 29932
rect 49868 39172 49924 39182
rect 49644 25666 49700 25676
rect 49756 28644 49812 28654
rect 49308 24322 49364 24332
rect 49420 25172 49476 25182
rect 49308 21588 49364 21598
rect 48972 20042 49140 20098
rect 49084 17108 49140 20042
rect 48972 16212 49028 16222
rect 48860 15428 48916 15438
rect 48860 15092 48916 15372
rect 48860 15026 48916 15036
rect 48972 14756 49028 16156
rect 48972 14690 49028 14700
rect 48860 13860 48916 13870
rect 48860 7812 48916 13804
rect 48972 12964 49028 12974
rect 48972 11508 49028 12908
rect 49084 11844 49140 17052
rect 49196 16100 49252 16110
rect 49196 13300 49252 16044
rect 49196 13234 49252 13244
rect 49196 12628 49252 12638
rect 49196 12180 49252 12572
rect 49196 12114 49252 12124
rect 49084 11778 49140 11788
rect 48972 11442 49028 11452
rect 48860 7746 48916 7756
rect 49308 5012 49364 21532
rect 49420 15316 49476 25116
rect 49644 24500 49700 24510
rect 49644 19348 49700 24444
rect 49420 15250 49476 15260
rect 49532 16772 49588 16782
rect 49532 14868 49588 16716
rect 49532 14802 49588 14812
rect 49644 13524 49700 19292
rect 49644 13458 49700 13468
rect 49756 12740 49812 28588
rect 49868 21588 49924 39116
rect 49980 33236 50036 47516
rect 50092 43764 50148 47740
rect 50092 43698 50148 43708
rect 50204 47124 50260 47134
rect 50204 42868 50260 47068
rect 50316 46788 50372 46798
rect 50316 44996 50372 46732
rect 50428 45332 50484 50876
rect 50540 50820 50596 50830
rect 50540 46004 50596 50764
rect 50764 50708 50820 53676
rect 50652 50372 50708 50382
rect 50652 47012 50708 50316
rect 50652 46946 50708 46956
rect 50540 45938 50596 45948
rect 50428 45266 50484 45276
rect 50316 44930 50372 44940
rect 50372 43204 50428 43214
rect 50372 43138 50428 43148
rect 50372 43082 50484 43138
rect 50428 42958 50484 43082
rect 50428 42902 50596 42958
rect 50204 42802 50260 42812
rect 50540 42756 50596 42902
rect 50540 42690 50596 42700
rect 50428 42532 50484 42542
rect 50428 42418 50484 42476
rect 50204 42362 50484 42418
rect 50204 42196 50260 42362
rect 50204 42130 50260 42140
rect 50428 42196 50484 42206
rect 50204 41076 50260 41086
rect 50204 40516 50260 41020
rect 50204 40450 50260 40460
rect 50316 40964 50372 40974
rect 50092 39060 50148 39070
rect 50092 37380 50148 39004
rect 50316 38998 50372 40908
rect 50428 40964 50484 42140
rect 50428 40898 50484 40908
rect 50540 40628 50596 40638
rect 50428 40068 50484 40078
rect 50428 39284 50484 40012
rect 50428 39218 50484 39228
rect 50204 38942 50372 38998
rect 50428 39060 50484 39070
rect 50204 38836 50260 38942
rect 50204 38770 50260 38780
rect 50092 37314 50148 37324
rect 50428 35700 50484 39004
rect 50540 37268 50596 40572
rect 50652 39284 50708 39294
rect 50652 38724 50708 39228
rect 50652 38658 50708 38668
rect 50540 37202 50596 37212
rect 50652 37156 50708 37166
rect 50204 34804 50260 34814
rect 49980 33170 50036 33180
rect 50092 33348 50148 33358
rect 49980 32676 50036 32686
rect 49980 29092 50036 32620
rect 49980 29026 50036 29036
rect 50092 26180 50148 33292
rect 50204 33236 50260 34748
rect 50204 33170 50260 33180
rect 50316 34580 50372 34590
rect 50316 30436 50372 34524
rect 50316 30370 50372 30380
rect 50092 26114 50148 26124
rect 50316 25844 50372 25854
rect 50316 24948 50372 25788
rect 50316 24882 50372 24892
rect 50204 24724 50260 24734
rect 49868 20580 49924 21532
rect 49868 20514 49924 20524
rect 49980 22932 50036 22942
rect 49980 20458 50036 22876
rect 50204 21028 50260 24668
rect 50204 20962 50260 20972
rect 49868 20402 50036 20458
rect 49868 17218 49924 20402
rect 50428 19378 50484 35644
rect 50540 37044 50596 37054
rect 50540 25396 50596 36988
rect 50652 34468 50708 37100
rect 50764 37044 50820 50652
rect 50764 36978 50820 36988
rect 50652 34402 50708 34412
rect 50764 36372 50820 36382
rect 50652 34244 50708 34254
rect 50652 33236 50708 34188
rect 50652 33170 50708 33180
rect 50540 25330 50596 25340
rect 50652 33012 50708 33022
rect 50652 26852 50708 32956
rect 50764 31556 50820 36316
rect 50764 31490 50820 31500
rect 50764 31108 50820 31118
rect 50764 30660 50820 31052
rect 50764 30594 50820 30604
rect 50204 19322 50484 19378
rect 50204 18838 50260 19322
rect 50316 19124 50372 19134
rect 50316 19018 50372 19068
rect 50316 18962 50596 19018
rect 50204 18782 50484 18838
rect 50092 17882 50372 17938
rect 50092 17758 50148 17882
rect 49980 17702 50148 17758
rect 50204 17780 50260 17790
rect 49980 17556 50036 17702
rect 49980 17490 50036 17500
rect 50204 17556 50260 17724
rect 50204 17490 50260 17500
rect 49868 17162 50148 17218
rect 49756 12674 49812 12684
rect 49532 11620 49588 11630
rect 49532 10738 49588 11564
rect 50092 11620 50148 17162
rect 50204 16772 50260 16782
rect 50204 13412 50260 16716
rect 50204 13346 50260 13356
rect 50092 11554 50148 11564
rect 49420 10724 49476 10734
rect 49420 9940 49476 10668
rect 49532 10724 49700 10738
rect 49532 10682 49644 10724
rect 49532 10388 49588 10682
rect 49644 10658 49700 10668
rect 49532 10322 49588 10332
rect 49756 10612 49812 10622
rect 49756 10388 49812 10556
rect 49756 10322 49812 10332
rect 49420 9874 49476 9884
rect 49308 4946 49364 4956
rect 50316 4900 50372 17882
rect 50428 11956 50484 18782
rect 50428 11890 50484 11900
rect 50540 8708 50596 18962
rect 50540 8642 50596 8652
rect 50652 6692 50708 26796
rect 50764 29988 50820 29998
rect 50764 11620 50820 29932
rect 50764 10276 50820 11564
rect 50764 10210 50820 10220
rect 50764 9268 50820 9278
rect 50764 7924 50820 9212
rect 50764 7858 50820 7868
rect 50652 6626 50708 6636
rect 50876 5796 50932 55468
rect 51436 55188 51492 55198
rect 51100 53508 51156 53518
rect 50988 52836 51044 52846
rect 50988 52276 51044 52780
rect 50988 52210 51044 52220
rect 51100 51598 51156 53452
rect 50988 51542 51156 51598
rect 51324 53060 51380 53070
rect 50988 44324 51044 51542
rect 51212 50932 51268 50942
rect 51212 50596 51268 50876
rect 51212 50530 51268 50540
rect 51212 49700 51268 49710
rect 50988 44258 51044 44268
rect 51100 48916 51156 48926
rect 50988 43428 51044 43438
rect 50988 42980 51044 43372
rect 50988 42914 51044 42924
rect 51100 40438 51156 48860
rect 51212 48244 51268 49644
rect 51212 48178 51268 48188
rect 51324 47796 51380 53004
rect 51436 50372 51492 55132
rect 51996 54740 52052 54750
rect 51436 50306 51492 50316
rect 51548 53732 51604 53742
rect 51324 47730 51380 47740
rect 51436 47348 51492 47358
rect 50988 40404 51156 40438
rect 51044 40382 51156 40404
rect 51212 46340 51268 46350
rect 50988 40338 51044 40348
rect 51100 35252 51156 35262
rect 50988 35140 51044 35150
rect 50988 32228 51044 35084
rect 51100 33796 51156 35196
rect 51100 33730 51156 33740
rect 50988 32162 51044 32172
rect 51100 33572 51156 33582
rect 51100 33012 51156 33516
rect 51100 31668 51156 32956
rect 51100 31602 51156 31612
rect 50988 27412 51044 27422
rect 50988 8260 51044 27356
rect 50988 8194 51044 8204
rect 51100 25508 51156 25518
rect 51100 22708 51156 25452
rect 51100 7364 51156 22652
rect 51212 24612 51268 46284
rect 51436 44996 51492 47292
rect 51436 44930 51492 44940
rect 51436 44324 51492 44334
rect 51324 43428 51380 43438
rect 51324 28084 51380 43372
rect 51324 28018 51380 28028
rect 51212 18900 51268 24556
rect 51212 18834 51268 18844
rect 51436 17444 51492 44268
rect 51548 41524 51604 53676
rect 51884 52276 51940 52286
rect 51548 41458 51604 41468
rect 51660 51380 51716 51390
rect 51660 40068 51716 51324
rect 51772 49476 51828 49486
rect 51772 42308 51828 49420
rect 51772 42242 51828 42252
rect 51884 46228 51940 52220
rect 51996 50484 52052 54684
rect 51996 50418 52052 50428
rect 51660 40002 51716 40012
rect 51548 37156 51604 37166
rect 51548 35364 51604 37100
rect 51548 35298 51604 35308
rect 51660 36932 51716 36942
rect 51548 31556 51604 31566
rect 51548 30772 51604 31500
rect 51548 30706 51604 30716
rect 51660 24724 51716 36876
rect 51772 36596 51828 36606
rect 51772 35252 51828 36540
rect 51884 35364 51940 46172
rect 51884 35298 51940 35308
rect 51996 45444 52052 45454
rect 51772 35186 51828 35196
rect 51884 34132 51940 34142
rect 51772 32564 51828 32574
rect 51772 32004 51828 32508
rect 51772 31938 51828 31948
rect 51884 32116 51940 34076
rect 51772 31556 51828 31566
rect 51772 27188 51828 31500
rect 51884 31444 51940 32060
rect 51884 31378 51940 31388
rect 51996 28532 52052 45388
rect 52108 42756 52164 55804
rect 52444 55558 52500 56476
rect 52332 55502 52500 55558
rect 54348 55860 54404 55870
rect 52332 50596 52388 55502
rect 52444 55412 52500 55422
rect 52444 50932 52500 55356
rect 54012 55300 54068 55310
rect 53788 53956 53844 53966
rect 53564 53900 53788 53938
rect 53564 53882 53844 53900
rect 52444 50866 52500 50876
rect 52556 53732 52612 53742
rect 52332 50530 52388 50540
rect 52108 42690 52164 42700
rect 52220 50372 52276 50382
rect 52108 42196 52164 42206
rect 52108 36260 52164 42140
rect 52108 36194 52164 36204
rect 51996 28466 52052 28476
rect 52108 34580 52164 34590
rect 51772 27122 51828 27132
rect 51660 24658 51716 24668
rect 51884 21812 51940 21822
rect 51884 21140 51940 21756
rect 51660 20804 51716 20814
rect 51436 17378 51492 17388
rect 51548 20580 51604 20590
rect 51548 18228 51604 20524
rect 51548 15764 51604 18172
rect 51548 15698 51604 15708
rect 51436 14868 51492 14878
rect 51436 14308 51492 14812
rect 51660 14756 51716 20748
rect 51772 18340 51828 18350
rect 51772 17780 51828 18284
rect 51772 17714 51828 17724
rect 51660 14690 51716 14700
rect 51772 16996 51828 17006
rect 51436 14242 51492 14252
rect 51772 11284 51828 16940
rect 51772 11218 51828 11228
rect 51884 8036 51940 21084
rect 51996 19018 52052 19022
rect 52108 19018 52164 34524
rect 51996 19012 52164 19018
rect 52052 18962 52164 19012
rect 51996 18946 52052 18956
rect 51996 16324 52052 16334
rect 51996 15764 52052 16268
rect 51996 15698 52052 15708
rect 52108 14196 52164 18962
rect 52108 14130 52164 14140
rect 52108 13412 52164 13422
rect 52108 11844 52164 13356
rect 52108 11778 52164 11788
rect 51884 7970 51940 7980
rect 51100 7298 51156 7308
rect 50876 5730 50932 5740
rect 50316 4834 50372 4844
rect 52220 3108 52276 50316
rect 52556 50260 52612 53676
rect 53452 53284 53508 53294
rect 53116 52500 53172 52510
rect 52668 52052 52724 52062
rect 52668 50932 52724 51996
rect 52668 50866 52724 50876
rect 52780 51492 52836 51502
rect 52780 50698 52836 51436
rect 52556 50194 52612 50204
rect 52668 50642 52836 50698
rect 52332 49588 52388 49598
rect 52332 23044 52388 49532
rect 52556 49588 52612 49598
rect 52444 47460 52500 47470
rect 52444 43092 52500 47404
rect 52444 43026 52500 43036
rect 52444 42756 52500 42766
rect 52444 40964 52500 42700
rect 52444 40898 52500 40908
rect 52444 39396 52500 39406
rect 52444 35924 52500 39340
rect 52444 35858 52500 35868
rect 52332 22978 52388 22988
rect 52444 32900 52500 32910
rect 52332 21364 52388 21374
rect 52332 16324 52388 21308
rect 52444 20356 52500 32844
rect 52556 32116 52612 49532
rect 52668 47124 52724 50642
rect 52668 47058 52724 47068
rect 52780 50484 52836 50494
rect 52668 43540 52724 43550
rect 52668 42308 52724 43484
rect 52668 42242 52724 42252
rect 52556 32050 52612 32060
rect 52668 41300 52724 41310
rect 52556 28420 52612 28430
rect 52556 26628 52612 28364
rect 52556 26562 52612 26572
rect 52668 23044 52724 41244
rect 52780 36596 52836 50428
rect 53004 50484 53060 50494
rect 52892 50260 52948 50270
rect 52892 42644 52948 50204
rect 53004 47684 53060 50428
rect 53116 48356 53172 52444
rect 53116 48290 53172 48300
rect 53340 48580 53396 48590
rect 53004 47618 53060 47628
rect 53004 46788 53060 46798
rect 53004 43876 53060 46732
rect 53116 46676 53172 46686
rect 53116 45668 53172 46620
rect 53116 45602 53172 45612
rect 53004 43810 53060 43820
rect 53116 45332 53172 45342
rect 53116 43678 53172 45276
rect 52892 42578 52948 42588
rect 53004 43622 53172 43678
rect 53228 43876 53284 43886
rect 52892 42308 52948 42318
rect 52892 39844 52948 42252
rect 52892 39778 52948 39788
rect 52780 36530 52836 36540
rect 52892 37044 52948 37054
rect 52780 34804 52836 34814
rect 52780 33684 52836 34748
rect 52892 34580 52948 36988
rect 52892 34514 52948 34524
rect 52780 33618 52836 33628
rect 52892 33460 52948 33470
rect 52892 32878 52948 33404
rect 53004 33124 53060 43622
rect 53004 33058 53060 33068
rect 53116 41636 53172 41646
rect 52892 32822 53060 32878
rect 52892 32676 52948 32686
rect 52780 31668 52836 31678
rect 52780 31332 52836 31612
rect 52780 31266 52836 31276
rect 52668 21812 52724 22988
rect 52668 21746 52724 21756
rect 52780 30884 52836 30894
rect 52444 20290 52500 20300
rect 52668 19908 52724 19918
rect 52444 18452 52500 18462
rect 52444 17108 52500 18396
rect 52444 17042 52500 17052
rect 52332 16258 52388 16268
rect 52556 13636 52612 13646
rect 52556 12964 52612 13580
rect 52668 13188 52724 19852
rect 52668 13122 52724 13132
rect 52556 12898 52612 12908
rect 52668 12180 52724 12190
rect 52668 11956 52724 12124
rect 52668 11890 52724 11900
rect 52780 10612 52836 30828
rect 52892 28756 52948 32620
rect 53004 28868 53060 32822
rect 53116 30884 53172 41580
rect 53228 37380 53284 43820
rect 53340 40852 53396 48524
rect 53340 40786 53396 40796
rect 53340 40516 53396 40526
rect 53340 39620 53396 40460
rect 53452 40180 53508 53228
rect 53564 50820 53620 53882
rect 53900 53732 53956 53742
rect 53564 50754 53620 50764
rect 53676 51156 53732 51166
rect 53676 48916 53732 51100
rect 53676 48850 53732 48860
rect 53788 48244 53844 48254
rect 53676 47684 53732 47694
rect 53564 44772 53620 44782
rect 53564 43540 53620 44716
rect 53564 43474 53620 43484
rect 53452 40114 53508 40124
rect 53564 43316 53620 43326
rect 53340 38052 53396 39564
rect 53340 37986 53396 37996
rect 53228 37314 53284 37324
rect 53340 36484 53396 36494
rect 53340 33684 53396 36428
rect 53340 33618 53396 33628
rect 53452 35252 53508 35262
rect 53340 33124 53396 33134
rect 53116 30818 53172 30828
rect 53228 31332 53284 31342
rect 53004 28802 53060 28812
rect 52892 28690 52948 28700
rect 53228 27412 53284 31276
rect 53340 28558 53396 33068
rect 53452 31780 53508 35196
rect 53452 29540 53508 31724
rect 53452 29474 53508 29484
rect 53340 28502 53508 28558
rect 53004 25620 53060 25630
rect 53004 16660 53060 25564
rect 53228 24836 53284 27356
rect 53228 24052 53284 24780
rect 53228 23986 53284 23996
rect 53340 28308 53396 28318
rect 53340 27860 53396 28252
rect 53004 16594 53060 16604
rect 52780 10546 52836 10556
rect 52892 11508 52948 11518
rect 52220 3042 52276 3052
rect 52332 9268 52388 9278
rect 48748 2594 48804 2604
rect 48412 2482 48468 2492
rect 48188 1810 48244 1820
rect 52332 1092 52388 9212
rect 52780 6468 52836 6478
rect 52780 6244 52836 6412
rect 52780 6178 52836 6188
rect 52892 4116 52948 11452
rect 53340 8932 53396 27804
rect 53452 24388 53508 28502
rect 53452 24322 53508 24332
rect 53452 18900 53508 18910
rect 53452 18004 53508 18844
rect 53452 17938 53508 17948
rect 53564 9268 53620 43260
rect 53676 42868 53732 47628
rect 53788 45556 53844 48188
rect 53788 45490 53844 45500
rect 53676 42802 53732 42812
rect 53788 44884 53844 44894
rect 53788 42308 53844 44828
rect 53900 44436 53956 53676
rect 53900 44370 53956 44380
rect 53788 42242 53844 42252
rect 53900 44212 53956 44222
rect 53788 42084 53844 42094
rect 53676 41748 53732 41758
rect 53676 31108 53732 41692
rect 53788 39396 53844 42028
rect 53788 39330 53844 39340
rect 53900 38276 53956 44156
rect 53900 38210 53956 38220
rect 53676 31042 53732 31052
rect 53788 37044 53844 37054
rect 53788 28980 53844 36988
rect 53900 33348 53956 33358
rect 53900 30100 53956 33292
rect 53900 30034 53956 30044
rect 53676 18676 53732 18686
rect 53676 15428 53732 18620
rect 53676 14980 53732 15372
rect 53676 14914 53732 14924
rect 53788 11956 53844 28924
rect 53788 11890 53844 11900
rect 53900 25620 53956 25630
rect 53564 9202 53620 9212
rect 53788 10948 53844 10958
rect 53340 8866 53396 8876
rect 52892 4050 52948 4060
rect 53788 3780 53844 10892
rect 53900 10164 53956 25564
rect 53900 10098 53956 10108
rect 53788 3714 53844 3724
rect 52332 1026 52388 1036
rect 47740 690 47796 700
rect 54012 644 54068 55244
rect 54124 52164 54180 52174
rect 54124 44884 54180 52108
rect 54236 51716 54292 51726
rect 54236 51156 54292 51660
rect 54236 51090 54292 51100
rect 54124 44818 54180 44828
rect 54236 50708 54292 50718
rect 54124 44324 54180 44334
rect 54124 37492 54180 44268
rect 54124 37426 54180 37436
rect 54124 34132 54180 34142
rect 54124 33238 54180 34076
rect 54236 33460 54292 50652
rect 54348 44398 54404 55804
rect 55580 55860 55636 55870
rect 54684 54516 54740 54526
rect 54460 51380 54516 51390
rect 54460 50878 54516 51324
rect 54460 50822 54628 50878
rect 54460 50148 54516 50158
rect 54460 44772 54516 50092
rect 54460 44706 54516 44716
rect 54348 44342 54516 44398
rect 54348 44100 54404 44110
rect 54348 41300 54404 44044
rect 54348 41234 54404 41244
rect 54348 40964 54404 40974
rect 54348 39284 54404 40908
rect 54348 39218 54404 39228
rect 54460 38998 54516 44342
rect 54572 42980 54628 50822
rect 54684 43652 54740 54460
rect 55468 54292 55524 54302
rect 55244 52948 55300 52958
rect 55132 51716 55188 51726
rect 54796 50822 54964 50878
rect 54796 50820 54852 50822
rect 54796 50754 54852 50764
rect 54796 50596 54852 50606
rect 54796 44212 54852 50540
rect 54908 48356 54964 50822
rect 54908 48290 54964 48300
rect 55020 50820 55076 50830
rect 55020 47796 55076 50764
rect 55020 47730 55076 47740
rect 55020 47012 55076 47022
rect 54908 46004 54964 46014
rect 54908 45780 54964 45948
rect 54908 45714 54964 45724
rect 54796 44146 54852 44156
rect 54908 44884 54964 44894
rect 54684 43586 54740 43596
rect 54796 43764 54852 43774
rect 54796 43092 54852 43708
rect 54796 43026 54852 43036
rect 54572 42914 54628 42924
rect 54348 38942 54516 38998
rect 54796 42644 54852 42654
rect 54348 37604 54404 38942
rect 54684 38612 54740 38622
rect 54348 37538 54404 37548
rect 54572 38388 54628 38398
rect 54236 33394 54292 33404
rect 54460 37044 54516 37054
rect 54124 33182 54292 33238
rect 54124 31892 54180 31902
rect 54124 14644 54180 31836
rect 54236 21812 54292 33182
rect 54348 31444 54404 31454
rect 54348 27412 54404 31388
rect 54348 27346 54404 27356
rect 54236 21746 54292 21756
rect 54124 14578 54180 14588
rect 54460 20132 54516 36988
rect 54460 12068 54516 20076
rect 54572 19348 54628 38332
rect 54684 32788 54740 38556
rect 54796 36372 54852 42588
rect 54796 36306 54852 36316
rect 54684 32722 54740 32732
rect 54796 35812 54852 35822
rect 54796 25844 54852 35756
rect 54796 25778 54852 25788
rect 54908 29652 54964 44828
rect 55020 44100 55076 46956
rect 55020 44034 55076 44044
rect 55020 43652 55076 43662
rect 55020 43204 55076 43596
rect 55020 34020 55076 43148
rect 55132 37380 55188 51660
rect 55244 37492 55300 52892
rect 55356 51604 55412 51614
rect 55356 50932 55412 51548
rect 55356 50866 55412 50876
rect 55356 45444 55412 45454
rect 55356 42084 55412 45388
rect 55356 42018 55412 42028
rect 55468 41748 55524 54236
rect 55580 42420 55636 55804
rect 55580 42354 55636 42364
rect 55692 54292 55748 54302
rect 55468 41682 55524 41692
rect 55580 42084 55636 42094
rect 55356 41412 55412 41422
rect 55356 37828 55412 41356
rect 55356 37762 55412 37772
rect 55244 37426 55300 37436
rect 55356 37604 55412 37614
rect 55132 37314 55188 37324
rect 55020 33954 55076 33964
rect 55132 37156 55188 37166
rect 54796 23380 54852 23390
rect 54572 19282 54628 19292
rect 54684 21812 54740 21822
rect 54684 13188 54740 21756
rect 54684 13122 54740 13132
rect 54460 12002 54516 12012
rect 54124 11956 54180 11966
rect 54124 6916 54180 11900
rect 54796 10164 54852 23324
rect 54908 16996 54964 29596
rect 55132 27748 55188 37100
rect 55356 35700 55412 37548
rect 55356 35634 55412 35644
rect 55580 35700 55636 42028
rect 55692 39956 55748 54236
rect 55804 49700 55860 56700
rect 55804 49634 55860 49644
rect 56924 52724 56980 52734
rect 56588 49588 56644 49598
rect 56028 49476 56084 49486
rect 55804 46900 55860 46910
rect 55804 46116 55860 46844
rect 55804 46050 55860 46060
rect 56028 42868 56084 49420
rect 56252 46676 56308 46686
rect 56140 45332 56196 45342
rect 56140 43876 56196 45276
rect 56140 43810 56196 43820
rect 56028 42802 56084 42812
rect 56140 43540 56196 43550
rect 56140 42084 56196 43484
rect 56140 42018 56196 42028
rect 55692 39890 55748 39900
rect 55804 41188 55860 41198
rect 55580 35634 55636 35644
rect 55132 27682 55188 27692
rect 55804 25284 55860 41132
rect 56140 39620 56196 39630
rect 55916 33236 55972 33246
rect 55916 28868 55972 33180
rect 55916 28802 55972 28812
rect 55804 25218 55860 25228
rect 56140 24276 56196 39564
rect 56252 36820 56308 46620
rect 56476 45220 56532 45230
rect 56364 41412 56420 41422
rect 56364 38388 56420 41356
rect 56364 38322 56420 38332
rect 56252 36754 56308 36764
rect 56476 35812 56532 45164
rect 56476 35746 56532 35756
rect 56140 24210 56196 24220
rect 56476 24500 56532 24510
rect 56252 23716 56308 23726
rect 55692 21924 55748 21934
rect 55692 21252 55748 21868
rect 55692 21186 55748 21196
rect 54908 16930 54964 16940
rect 54796 10098 54852 10108
rect 55132 16436 55188 16446
rect 54124 6850 54180 6860
rect 55132 6244 55188 16380
rect 55132 6178 55188 6188
rect 55356 15428 55412 15438
rect 55356 3780 55412 15372
rect 56252 10500 56308 23660
rect 56252 10434 56308 10444
rect 56364 23604 56420 23614
rect 56140 10388 56196 10398
rect 56140 5236 56196 10332
rect 56364 10052 56420 23548
rect 56476 11620 56532 24444
rect 56588 14756 56644 49532
rect 56812 42084 56868 42094
rect 56700 38724 56756 38734
rect 56700 38276 56756 38668
rect 56812 38388 56868 42028
rect 56812 38322 56868 38332
rect 56700 38210 56756 38220
rect 56924 36596 56980 52668
rect 57260 51604 57316 51614
rect 57148 51156 57204 51166
rect 57036 41188 57092 41198
rect 57036 36820 57092 41132
rect 57036 36754 57092 36764
rect 56924 36530 56980 36540
rect 57148 34804 57204 51100
rect 57260 35252 57316 51548
rect 57260 35186 57316 35196
rect 57372 43540 57428 43550
rect 57148 34738 57204 34748
rect 57372 24418 57428 43484
rect 57148 24388 57428 24418
rect 57204 24362 57428 24388
rect 57148 24322 57204 24332
rect 56812 24052 56868 24062
rect 56812 23716 56868 23996
rect 56812 23650 56868 23660
rect 56588 14690 56644 14700
rect 56476 11554 56532 11564
rect 56364 9986 56420 9996
rect 56140 5170 56196 5180
rect 55356 3714 55412 3724
rect 54012 578 54068 588
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0859_
timestamp 1486834041
transform -1 0 35952 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0860_
timestamp 1486834041
transform 1 0 42784 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0861_
timestamp 1486834041
transform 1 0 13664 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0862_
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0863_
timestamp 1486834041
transform 1 0 35504 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0864_
timestamp 1486834041
transform 1 0 36288 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0865_
timestamp 1486834041
transform -1 0 12432 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0866_
timestamp 1486834041
transform -1 0 13776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0867_
timestamp 1486834041
transform -1 0 19376 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0868_
timestamp 1486834041
transform 1 0 31136 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0869_
timestamp 1486834041
transform -1 0 28224 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0870_
timestamp 1486834041
transform 1 0 18480 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0871_
timestamp 1486834041
transform 1 0 18928 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0872_
timestamp 1486834041
transform -1 0 21952 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0873_
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0874_
timestamp 1486834041
transform 1 0 35504 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0875_
timestamp 1486834041
transform 1 0 32368 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0876_
timestamp 1486834041
transform -1 0 34720 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0877_
timestamp 1486834041
transform 1 0 35504 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0878_
timestamp 1486834041
transform -1 0 16352 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0879_
timestamp 1486834041
transform 1 0 16464 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0880_
timestamp 1486834041
transform 1 0 4144 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0881_
timestamp 1486834041
transform -1 0 9184 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0882_
timestamp 1486834041
transform -1 0 52976 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0883_
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0884_
timestamp 1486834041
transform 1 0 11984 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0885_
timestamp 1486834041
transform -1 0 42448 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0886_
timestamp 1486834041
transform -1 0 50400 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0887_
timestamp 1486834041
transform 1 0 47824 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0888_
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0889_
timestamp 1486834041
transform -1 0 13104 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0890_
timestamp 1486834041
transform -1 0 8176 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0891_
timestamp 1486834041
transform 1 0 28672 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0892_
timestamp 1486834041
transform 1 0 18368 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0893_
timestamp 1486834041
transform 1 0 18816 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0894_
timestamp 1486834041
transform -1 0 9184 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0895_
timestamp 1486834041
transform -1 0 8848 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0896_
timestamp 1486834041
transform 1 0 20608 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0897_
timestamp 1486834041
transform -1 0 25200 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0898_
timestamp 1486834041
transform -1 0 16688 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0899_
timestamp 1486834041
transform -1 0 16688 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0900_
timestamp 1486834041
transform 1 0 16240 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0901_
timestamp 1486834041
transform 1 0 20496 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0902_
timestamp 1486834041
transform 1 0 4704 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0903_
timestamp 1486834041
transform 1 0 3248 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0904_
timestamp 1486834041
transform 1 0 31584 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0905_
timestamp 1486834041
transform 1 0 3136 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0906_
timestamp 1486834041
transform -1 0 6160 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0907_
timestamp 1486834041
transform 1 0 51184 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0908_
timestamp 1486834041
transform -1 0 52192 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0909_
timestamp 1486834041
transform -1 0 56560 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0910_
timestamp 1486834041
transform -1 0 12096 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0911_
timestamp 1486834041
transform -1 0 9184 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0912_
timestamp 1486834041
transform 1 0 7616 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0913_
timestamp 1486834041
transform 1 0 8064 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0914_
timestamp 1486834041
transform -1 0 6832 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0915_
timestamp 1486834041
transform -1 0 6608 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0916_
timestamp 1486834041
transform 1 0 12768 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0917_
timestamp 1486834041
transform 1 0 54096 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0918_
timestamp 1486834041
transform 1 0 42672 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0919_
timestamp 1486834041
transform 1 0 42672 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0920_
timestamp 1486834041
transform 1 0 38416 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0921_
timestamp 1486834041
transform 1 0 15008 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0922_
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0923_
timestamp 1486834041
transform 1 0 19824 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0924_
timestamp 1486834041
transform 1 0 25088 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0925_
timestamp 1486834041
transform -1 0 8512 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0926_
timestamp 1486834041
transform 1 0 30912 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0927_
timestamp 1486834041
transform -1 0 43120 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0928_
timestamp 1486834041
transform -1 0 45024 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0929_
timestamp 1486834041
transform 1 0 3136 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0930_
timestamp 1486834041
transform -1 0 6160 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0931_
timestamp 1486834041
transform 1 0 11760 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0932_
timestamp 1486834041
transform 1 0 11088 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0933_
timestamp 1486834041
transform 1 0 3136 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0934_
timestamp 1486834041
transform 1 0 3136 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0935_
timestamp 1486834041
transform -1 0 12432 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0936_
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0937_
timestamp 1486834041
transform -1 0 12992 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0938_
timestamp 1486834041
transform 1 0 17024 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0939_
timestamp 1486834041
transform 1 0 19264 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0940_
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0941_
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0942_
timestamp 1486834041
transform -1 0 20272 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0943_
timestamp 1486834041
transform 1 0 18928 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0944_
timestamp 1486834041
transform 1 0 22848 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0945_
timestamp 1486834041
transform 1 0 19040 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0946_
timestamp 1486834041
transform -1 0 18928 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0947_
timestamp 1486834041
transform 1 0 18928 0 1 13328
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0948_
timestamp 1486834041
transform -1 0 48944 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0949_
timestamp 1486834041
transform 1 0 32368 0 -1 25872
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0950_
timestamp 1486834041
transform 1 0 31472 0 -1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0951_
timestamp 1486834041
transform -1 0 35504 0 1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0952_
timestamp 1486834041
transform 1 0 32592 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0953_
timestamp 1486834041
transform 1 0 32256 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0954_
timestamp 1486834041
transform 1 0 26096 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0955_
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0956_
timestamp 1486834041
transform 1 0 24528 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0957_
timestamp 1486834041
transform 1 0 26656 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0958_
timestamp 1486834041
transform 1 0 24528 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0959_
timestamp 1486834041
transform 1 0 25424 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0960_
timestamp 1486834041
transform 1 0 25536 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0961_
timestamp 1486834041
transform -1 0 26432 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _0962_
timestamp 1486834041
transform 1 0 26432 0 -1 5488
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0963_
timestamp 1486834041
transform 1 0 32256 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0964_
timestamp 1486834041
transform 1 0 26768 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0965_
timestamp 1486834041
transform 1 0 44128 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0966_
timestamp 1486834041
transform 1 0 15232 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0967_
timestamp 1486834041
transform -1 0 16352 0 -1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0968_
timestamp 1486834041
transform 1 0 15120 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0969_
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0970_
timestamp 1486834041
transform 1 0 16240 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0971_
timestamp 1486834041
transform -1 0 16240 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0972_
timestamp 1486834041
transform -1 0 17136 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0973_
timestamp 1486834041
transform 1 0 17472 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0974_
timestamp 1486834041
transform -1 0 16352 0 -1 10192
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0975_
timestamp 1486834041
transform 1 0 41888 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0976_
timestamp 1486834041
transform 1 0 43008 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0977_
timestamp 1486834041
transform -1 0 13776 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0978_
timestamp 1486834041
transform 1 0 10640 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0979_
timestamp 1486834041
transform -1 0 15120 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0980_
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0981_
timestamp 1486834041
transform -1 0 12432 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0982_
timestamp 1486834041
transform -1 0 14784 0 -1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0983_
timestamp 1486834041
transform -1 0 12768 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0984_
timestamp 1486834041
transform -1 0 10640 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0985_
timestamp 1486834041
transform 1 0 11312 0 1 5488
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0986_
timestamp 1486834041
transform 1 0 19824 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0987_
timestamp 1486834041
transform 1 0 27888 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0988_
timestamp 1486834041
transform 1 0 45920 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0989_
timestamp 1486834041
transform 1 0 46032 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0990_
timestamp 1486834041
transform -1 0 49616 0 -1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0991_
timestamp 1486834041
transform -1 0 56336 0 1 3920
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0992_
timestamp 1486834041
transform -1 0 36512 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0993_
timestamp 1486834041
transform -1 0 37296 0 1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0994_
timestamp 1486834041
transform 1 0 32368 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0995_
timestamp 1486834041
transform 1 0 31920 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0996_
timestamp 1486834041
transform -1 0 33376 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0997_
timestamp 1486834041
transform 1 0 35280 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0998_
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0999_
timestamp 1486834041
transform 1 0 34496 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1000_
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1001_
timestamp 1486834041
transform 1 0 33376 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1002_
timestamp 1486834041
transform -1 0 33936 0 -1 7056
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1003_
timestamp 1486834041
transform 1 0 33936 0 -1 7056
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1004_
timestamp 1486834041
transform 1 0 36176 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1005_
timestamp 1486834041
transform -1 0 36624 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1006_
timestamp 1486834041
transform -1 0 37744 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1007_
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1008_
timestamp 1486834041
transform 1 0 20048 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1009_
timestamp 1486834041
transform 1 0 35728 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1010_
timestamp 1486834041
transform 1 0 36400 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1011_
timestamp 1486834041
transform 1 0 37744 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1012_
timestamp 1486834041
transform 1 0 38976 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1013_
timestamp 1486834041
transform -1 0 18144 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1014_
timestamp 1486834041
transform 1 0 20608 0 1 2352
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1015_
timestamp 1486834041
transform 1 0 19600 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1016_
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1017_
timestamp 1486834041
transform -1 0 20272 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1018_
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1019_
timestamp 1486834041
transform -1 0 23072 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1020_
timestamp 1486834041
transform -1 0 22064 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1021_
timestamp 1486834041
transform 1 0 19376 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1022_
timestamp 1486834041
transform -1 0 20272 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1023_
timestamp 1486834041
transform 1 0 20384 0 -1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1024_
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1025_
timestamp 1486834041
transform -1 0 20272 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1026_
timestamp 1486834041
transform -1 0 23296 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1027_
timestamp 1486834041
transform 1 0 18144 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1028_
timestamp 1486834041
transform -1 0 22848 0 1 2352
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1029_
timestamp 1486834041
transform 1 0 28336 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1030_
timestamp 1486834041
transform -1 0 37296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1031_
timestamp 1486834041
transform 1 0 37856 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1032_
timestamp 1486834041
transform 1 0 38528 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1033_
timestamp 1486834041
transform 1 0 37856 0 -1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1034_
timestamp 1486834041
transform 1 0 53872 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1035_
timestamp 1486834041
transform 1 0 53536 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1036_
timestamp 1486834041
transform -1 0 8512 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1037_
timestamp 1486834041
transform -1 0 14560 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1038_
timestamp 1486834041
transform -1 0 8512 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1039_
timestamp 1486834041
transform 1 0 7616 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1040_
timestamp 1486834041
transform -1 0 8848 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1041_
timestamp 1486834041
transform 1 0 7616 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1042_
timestamp 1486834041
transform -1 0 7616 0 1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1043_
timestamp 1486834041
transform -1 0 4928 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1044_
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1045_
timestamp 1486834041
transform 1 0 40096 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1046_
timestamp 1486834041
transform 1 0 25424 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1047_
timestamp 1486834041
transform -1 0 16352 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1048_
timestamp 1486834041
transform 1 0 14784 0 -1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1049_
timestamp 1486834041
transform 1 0 14896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1050_
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1051_
timestamp 1486834041
transform 1 0 14784 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1052_
timestamp 1486834041
transform 1 0 15792 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1053_
timestamp 1486834041
transform -1 0 17136 0 -1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1054_
timestamp 1486834041
transform -1 0 14784 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1055_
timestamp 1486834041
transform 1 0 15344 0 -1 7056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1056_
timestamp 1486834041
transform 1 0 28448 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1057_
timestamp 1486834041
transform 1 0 41216 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1058_
timestamp 1486834041
transform -1 0 43792 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1059_
timestamp 1486834041
transform 1 0 44016 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1060_
timestamp 1486834041
transform -1 0 51632 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1061_
timestamp 1486834041
transform 1 0 53872 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1062_
timestamp 1486834041
transform -1 0 51632 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1063_
timestamp 1486834041
transform 1 0 51408 0 -1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1064_
timestamp 1486834041
transform 1 0 50736 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1065_
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1066_
timestamp 1486834041
transform 1 0 51856 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1067_
timestamp 1486834041
transform 1 0 51744 0 -1 13328
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1068_
timestamp 1486834041
transform -1 0 52528 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1069_
timestamp 1486834041
transform 1 0 49728 0 -1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1070_
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1071_
timestamp 1486834041
transform 1 0 49952 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1072_
timestamp 1486834041
transform -1 0 48272 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1073_
timestamp 1486834041
transform 1 0 48272 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1074_
timestamp 1486834041
transform 1 0 48832 0 1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1075_
timestamp 1486834041
transform 1 0 46704 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1076_
timestamp 1486834041
transform -1 0 49056 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1077_
timestamp 1486834041
transform 1 0 46144 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1078_
timestamp 1486834041
transform 1 0 45248 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1079_
timestamp 1486834041
transform 1 0 43232 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1080_
timestamp 1486834041
transform 1 0 44688 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1081_
timestamp 1486834041
transform 1 0 46256 0 1 16464
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1082_
timestamp 1486834041
transform 1 0 47152 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1083_
timestamp 1486834041
transform 1 0 50624 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1084_
timestamp 1486834041
transform 1 0 34832 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1085_
timestamp 1486834041
transform 1 0 52752 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1086_
timestamp 1486834041
transform 1 0 44912 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1087_
timestamp 1486834041
transform 1 0 53424 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1088_
timestamp 1486834041
transform 1 0 52752 0 -1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1089_
timestamp 1486834041
transform -1 0 53312 0 -1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1090_
timestamp 1486834041
transform 1 0 47040 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1091_
timestamp 1486834041
transform -1 0 55552 0 -1 19600
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1092_
timestamp 1486834041
transform 1 0 47264 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1093_
timestamp 1486834041
transform -1 0 55440 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1094_
timestamp 1486834041
transform -1 0 53200 0 1 18032
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1095_
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1096_
timestamp 1486834041
transform 1 0 46816 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1097_
timestamp 1486834041
transform -1 0 48048 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1098_
timestamp 1486834041
transform 1 0 48048 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1099_
timestamp 1486834041
transform 1 0 47040 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1100_
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1101_
timestamp 1486834041
transform 1 0 47936 0 -1 13328
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _1102_
timestamp 1486834041
transform 1 0 50400 0 -1 16464
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1103_
timestamp 1486834041
transform -1 0 55888 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1104_
timestamp 1486834041
transform -1 0 53312 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1105_
timestamp 1486834041
transform -1 0 51520 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1106_
timestamp 1486834041
transform 1 0 55328 0 1 21168
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1107_
timestamp 1486834041
transform 1 0 51744 0 -1 21168
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _1108_
timestamp 1486834041
transform 1 0 53872 0 -1 18032
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1109_
timestamp 1486834041
transform -1 0 56560 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1110_
timestamp 1486834041
transform 1 0 53872 0 -1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1111_
timestamp 1486834041
transform 1 0 52192 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1112_
timestamp 1486834041
transform -1 0 53536 0 1 19600
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1113_
timestamp 1486834041
transform 1 0 49952 0 1 25872
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1114_
timestamp 1486834041
transform 1 0 8848 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1486834041
transform 1 0 5936 0 -1 55664
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1116_
timestamp 1486834041
transform 1 0 9184 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1117_
timestamp 1486834041
transform -1 0 8512 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1118_
timestamp 1486834041
transform -1 0 12432 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1119_
timestamp 1486834041
transform -1 0 13216 0 1 38416
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1120_
timestamp 1486834041
transform 1 0 8960 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1122_
timestamp 1486834041
transform -1 0 10752 0 1 46256
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1123_
timestamp 1486834041
transform 1 0 43456 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1124_
timestamp 1486834041
transform 1 0 26432 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1125_
timestamp 1486834041
transform 1 0 20496 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1126_
timestamp 1486834041
transform -1 0 21504 0 1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1127_
timestamp 1486834041
transform 1 0 21168 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1128_
timestamp 1486834041
transform -1 0 21392 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1129_
timestamp 1486834041
transform 1 0 20496 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1130_
timestamp 1486834041
transform 1 0 20608 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1131_
timestamp 1486834041
transform -1 0 21168 0 1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1132_
timestamp 1486834041
transform -1 0 21952 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1133_
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1134_
timestamp 1486834041
transform -1 0 40656 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1135_
timestamp 1486834041
transform -1 0 34496 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1136_
timestamp 1486834041
transform 1 0 23744 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1137_
timestamp 1486834041
transform 1 0 40208 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1138_
timestamp 1486834041
transform -1 0 55552 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1139_
timestamp 1486834041
transform 1 0 16688 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1140_
timestamp 1486834041
transform -1 0 17136 0 -1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1141_
timestamp 1486834041
transform -1 0 20272 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1142_
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1143_
timestamp 1486834041
transform -1 0 21616 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1144_
timestamp 1486834041
transform -1 0 20384 0 -1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1145_
timestamp 1486834041
transform 1 0 19376 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1146_
timestamp 1486834041
transform -1 0 20272 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1147_
timestamp 1486834041
transform -1 0 19824 0 -1 29008
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1148_
timestamp 1486834041
transform 1 0 15344 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1149_
timestamp 1486834041
transform -1 0 21392 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1150_
timestamp 1486834041
transform 1 0 15008 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1151_
timestamp 1486834041
transform 1 0 15120 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1152_
timestamp 1486834041
transform -1 0 21056 0 1 46256
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1153_
timestamp 1486834041
transform -1 0 16352 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1154_
timestamp 1486834041
transform -1 0 16352 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1155_
timestamp 1486834041
transform 1 0 15008 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1156_
timestamp 1486834041
transform -1 0 17136 0 -1 44688
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1157_
timestamp 1486834041
transform 1 0 15344 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1158_
timestamp 1486834041
transform 1 0 15344 0 -1 49392
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1159_
timestamp 1486834041
transform 1 0 23296 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1160_
timestamp 1486834041
transform 1 0 27104 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1161_
timestamp 1486834041
transform 1 0 26432 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1162_
timestamp 1486834041
transform -1 0 51632 0 1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1163_
timestamp 1486834041
transform 1 0 53088 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1164_
timestamp 1486834041
transform -1 0 53536 0 1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1165_
timestamp 1486834041
transform 1 0 41104 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1166_
timestamp 1486834041
transform 1 0 43344 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1167_
timestamp 1486834041
transform 1 0 26320 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1168_
timestamp 1486834041
transform 1 0 50736 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1169_
timestamp 1486834041
transform 1 0 50288 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1170_
timestamp 1486834041
transform 1 0 48832 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1171_
timestamp 1486834041
transform -1 0 49168 0 -1 14896
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1172_
timestamp 1486834041
transform 1 0 50736 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1173_
timestamp 1486834041
transform 1 0 49616 0 -1 32144
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1174_
timestamp 1486834041
transform -1 0 41440 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1175_
timestamp 1486834041
transform -1 0 34384 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1176_
timestamp 1486834041
transform 1 0 3360 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1177_
timestamp 1486834041
transform 1 0 2240 0 -1 39984
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1178_
timestamp 1486834041
transform 1 0 1008 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1179_
timestamp 1486834041
transform 1 0 3696 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1180_
timestamp 1486834041
transform 1 0 2800 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1181_
timestamp 1486834041
transform 1 0 3472 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1182_
timestamp 1486834041
transform -1 0 3696 0 1 49392
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1183_
timestamp 1486834041
transform 1 0 3696 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1184_
timestamp 1486834041
transform 1 0 4816 0 1 39984
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1185_
timestamp 1486834041
transform 1 0 40992 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1186_
timestamp 1486834041
transform -1 0 39536 0 -1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1187_
timestamp 1486834041
transform 1 0 38416 0 1 27440
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1188_
timestamp 1486834041
transform 1 0 39536 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1189_
timestamp 1486834041
transform 1 0 38640 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1190_
timestamp 1486834041
transform 1 0 38752 0 1 24304
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1191_
timestamp 1486834041
transform 1 0 38976 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1192_
timestamp 1486834041
transform 1 0 38640 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1193_
timestamp 1486834041
transform -1 0 53648 0 1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1194_
timestamp 1486834041
transform -1 0 51520 0 1 43120
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1195_
timestamp 1486834041
transform 1 0 32144 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1196_
timestamp 1486834041
transform 1 0 29680 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1197_
timestamp 1486834041
transform 1 0 8176 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1198_
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1199_
timestamp 1486834041
transform 1 0 3136 0 1 38416
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1200_
timestamp 1486834041
transform -1 0 8512 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1201_
timestamp 1486834041
transform 1 0 8736 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1202_
timestamp 1486834041
transform -1 0 9968 0 -1 36848
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1203_
timestamp 1486834041
transform 1 0 8064 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1204_
timestamp 1486834041
transform -1 0 8512 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1205_
timestamp 1486834041
transform -1 0 10192 0 -1 38416
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1206_
timestamp 1486834041
transform -1 0 46144 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1207_
timestamp 1486834041
transform 1 0 35840 0 -1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1208_
timestamp 1486834041
transform 1 0 36176 0 1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1209_
timestamp 1486834041
transform -1 0 36288 0 -1 24304
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1486834041
transform -1 0 35952 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1211_
timestamp 1486834041
transform 1 0 36176 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1212_
timestamp 1486834041
transform 1 0 40096 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1213_
timestamp 1486834041
transform 1 0 16688 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1214_
timestamp 1486834041
transform -1 0 16688 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1215_
timestamp 1486834041
transform 1 0 8288 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1216_
timestamp 1486834041
transform -1 0 8512 0 -1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1217_
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1218_
timestamp 1486834041
transform 1 0 9968 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1219_
timestamp 1486834041
transform 1 0 8064 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1220_
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1221_
timestamp 1486834041
transform 1 0 7392 0 -1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1222_
timestamp 1486834041
transform 1 0 9296 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1223_
timestamp 1486834041
transform 1 0 8960 0 -1 30576
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1224_
timestamp 1486834041
transform 1 0 22960 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1225_
timestamp 1486834041
transform 1 0 26320 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1226_
timestamp 1486834041
transform 1 0 24080 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1227_
timestamp 1486834041
transform 1 0 50064 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1228_
timestamp 1486834041
transform 1 0 54096 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1229_
timestamp 1486834041
transform -1 0 44576 0 1 47824
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1230_
timestamp 1486834041
transform -1 0 51632 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1231_
timestamp 1486834041
transform 1 0 48496 0 1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1232_
timestamp 1486834041
transform 1 0 50624 0 -1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1233_
timestamp 1486834041
transform -1 0 50624 0 -1 41552
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1234_
timestamp 1486834041
transform 1 0 27888 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1235_
timestamp 1486834041
transform 1 0 14672 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1236_
timestamp 1486834041
transform 1 0 40320 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1237_
timestamp 1486834041
transform 1 0 3136 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1238_
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1239_
timestamp 1486834041
transform 1 0 2240 0 -1 33712
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1240_
timestamp 1486834041
transform 1 0 3696 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1241_
timestamp 1486834041
transform -1 0 4592 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1242_
timestamp 1486834041
transform 1 0 4144 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1243_
timestamp 1486834041
transform -1 0 8288 0 -1 35280
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1244_
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1245_
timestamp 1486834041
transform -1 0 4144 0 -1 35280
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1246_
timestamp 1486834041
transform 1 0 23632 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1247_
timestamp 1486834041
transform 1 0 40880 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1248_
timestamp 1486834041
transform 1 0 41216 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1249_
timestamp 1486834041
transform 1 0 40096 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1250_
timestamp 1486834041
transform -1 0 53200 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1251_
timestamp 1486834041
transform 1 0 53760 0 -1 44688
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1252_
timestamp 1486834041
transform 1 0 53536 0 -1 43120
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1253_
timestamp 1486834041
transform 1 0 52080 0 -1 44688
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1254_
timestamp 1486834041
transform 1 0 51072 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1255_
timestamp 1486834041
transform 1 0 50512 0 1 47824
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1256_
timestamp 1486834041
transform 1 0 52192 0 1 46256
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1257_
timestamp 1486834041
transform 1 0 54432 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1258_
timestamp 1486834041
transform 1 0 51856 0 1 44688
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1259_
timestamp 1486834041
transform 1 0 50400 0 -1 44688
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1260_
timestamp 1486834041
transform 1 0 48272 0 -1 50960
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1261_
timestamp 1486834041
transform 1 0 1008 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1262_
timestamp 1486834041
transform 1 0 3920 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1263_
timestamp 1486834041
transform 1 0 7056 0 -1 39984
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1264_
timestamp 1486834041
transform 1 0 3696 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1265_
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1266_
timestamp 1486834041
transform -1 0 22176 0 1 55664
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1267_
timestamp 1486834041
transform 1 0 2352 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1268_
timestamp 1486834041
transform 1 0 3360 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1269_
timestamp 1486834041
transform 1 0 3584 0 1 46256
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1270_
timestamp 1486834041
transform -1 0 45920 0 1 33712
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1271_
timestamp 1486834041
transform 1 0 42560 0 1 36848
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1272_
timestamp 1486834041
transform 1 0 45920 0 1 33712
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1273_
timestamp 1486834041
transform 1 0 46816 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1274_
timestamp 1486834041
transform -1 0 47600 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1275_
timestamp 1486834041
transform 1 0 42560 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1276_
timestamp 1486834041
transform -1 0 47600 0 -1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1277_
timestamp 1486834041
transform 1 0 18704 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1278_
timestamp 1486834041
transform -1 0 19376 0 -1 35280
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1279_
timestamp 1486834041
transform 1 0 18816 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1280_
timestamp 1486834041
transform -1 0 20272 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1281_
timestamp 1486834041
transform 1 0 19376 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1282_
timestamp 1486834041
transform 1 0 20608 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1283_
timestamp 1486834041
transform -1 0 21056 0 1 33712
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1284_
timestamp 1486834041
transform -1 0 20160 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1285_
timestamp 1486834041
transform -1 0 20384 0 -1 35280
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1286_
timestamp 1486834041
transform 1 0 40096 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1287_
timestamp 1486834041
transform 1 0 29120 0 1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1288_
timestamp 1486834041
transform 1 0 29792 0 -1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1289_
timestamp 1486834041
transform -1 0 28112 0 1 30576
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1290_
timestamp 1486834041
transform 1 0 28672 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1291_
timestamp 1486834041
transform 1 0 46144 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1292_
timestamp 1486834041
transform -1 0 47152 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1293_
timestamp 1486834041
transform 1 0 47936 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1294_
timestamp 1486834041
transform 1 0 49056 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1295_
timestamp 1486834041
transform -1 0 50064 0 1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1296_
timestamp 1486834041
transform 1 0 51072 0 1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1297_
timestamp 1486834041
transform 1 0 54432 0 1 32144
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1298_
timestamp 1486834041
transform 1 0 51856 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1299_
timestamp 1486834041
transform -1 0 56112 0 1 33712
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1300_
timestamp 1486834041
transform 1 0 55776 0 -1 30576
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1301_
timestamp 1486834041
transform 1 0 52528 0 1 32144
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1302_
timestamp 1486834041
transform 1 0 51520 0 -1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1303_
timestamp 1486834041
transform 1 0 52080 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1304_
timestamp 1486834041
transform 1 0 32256 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1305_
timestamp 1486834041
transform 1 0 31808 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1306_
timestamp 1486834041
transform -1 0 35840 0 1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1307_
timestamp 1486834041
transform 1 0 31472 0 -1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1308_
timestamp 1486834041
transform -1 0 35952 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1309_
timestamp 1486834041
transform -1 0 34160 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1310_
timestamp 1486834041
transform 1 0 32256 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1311_
timestamp 1486834041
transform 1 0 31136 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1312_
timestamp 1486834041
transform 1 0 34160 0 1 29008
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1313_
timestamp 1486834041
transform 1 0 36176 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1314_
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1315_
timestamp 1486834041
transform 1 0 29120 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1316_
timestamp 1486834041
transform 1 0 40208 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1317_
timestamp 1486834041
transform 1 0 2912 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1318_
timestamp 1486834041
transform 1 0 3136 0 1 41552
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1319_
timestamp 1486834041
transform 1 0 3248 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1320_
timestamp 1486834041
transform -1 0 4368 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1321_
timestamp 1486834041
transform -1 0 4592 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1322_
timestamp 1486834041
transform 1 0 4368 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1323_
timestamp 1486834041
transform -1 0 3696 0 -1 55664
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1324_
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1325_
timestamp 1486834041
transform -1 0 4480 0 1 43120
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1326_
timestamp 1486834041
transform 1 0 28000 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1327_
timestamp 1486834041
transform 1 0 40208 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1486834041
transform 1 0 40544 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1329_
timestamp 1486834041
transform -1 0 44464 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1330_
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1331_
timestamp 1486834041
transform -1 0 43792 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1332_
timestamp 1486834041
transform 1 0 44352 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1333_
timestamp 1486834041
transform -1 0 52976 0 1 29008
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1334_
timestamp 1486834041
transform -1 0 54768 0 -1 29008
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1335_
timestamp 1486834041
transform 1 0 54432 0 1 22736
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1336_
timestamp 1486834041
transform 1 0 55776 0 -1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1337_
timestamp 1486834041
transform -1 0 55440 0 -1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1338_
timestamp 1486834041
transform 1 0 52528 0 -1 29008
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1339_
timestamp 1486834041
transform 1 0 51856 0 1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1340_
timestamp 1486834041
transform 1 0 54656 0 -1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1341_
timestamp 1486834041
transform 1 0 50064 0 1 29008
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1342_
timestamp 1486834041
transform 1 0 51184 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1343_
timestamp 1486834041
transform 1 0 47936 0 -1 29008
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1344_
timestamp 1486834041
transform 1 0 51856 0 1 43120
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1345_
timestamp 1486834041
transform 1 0 38752 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1346_
timestamp 1486834041
transform -1 0 42896 0 1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1347_
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1348_
timestamp 1486834041
transform -1 0 43792 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1349_
timestamp 1486834041
transform 1 0 39088 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1350_
timestamp 1486834041
transform -1 0 39872 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1351_
timestamp 1486834041
transform 1 0 44016 0 1 43120
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1352_
timestamp 1486834041
transform -1 0 40544 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1353_
timestamp 1486834041
transform 1 0 42560 0 1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1354_
timestamp 1486834041
transform 1 0 42336 0 -1 41552
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1355_
timestamp 1486834041
transform 1 0 39536 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1356_
timestamp 1486834041
transform -1 0 46704 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1357_
timestamp 1486834041
transform 1 0 42448 0 1 44688
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1358_
timestamp 1486834041
transform -1 0 43008 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1359_
timestamp 1486834041
transform 1 0 42896 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1360_
timestamp 1486834041
transform -1 0 44240 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1361_
timestamp 1486834041
transform 1 0 42448 0 -1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1362_
timestamp 1486834041
transform -1 0 43344 0 1 19600
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1363_
timestamp 1486834041
transform -1 0 43792 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1364_
timestamp 1486834041
transform 1 0 46592 0 -1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1365_
timestamp 1486834041
transform -1 0 43792 0 1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1366_
timestamp 1486834041
transform 1 0 47936 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1367_
timestamp 1486834041
transform 1 0 46256 0 -1 49392
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1486834041
transform -1 0 49840 0 1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1369_
timestamp 1486834041
transform 1 0 45360 0 -1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1370_
timestamp 1486834041
transform 1 0 48608 0 1 43120
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_
timestamp 1486834041
transform -1 0 43568 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1372_
timestamp 1486834041
transform -1 0 45696 0 1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1373_
timestamp 1486834041
transform 1 0 46032 0 -1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1374_
timestamp 1486834041
transform 1 0 45472 0 -1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1375_
timestamp 1486834041
transform 1 0 46480 0 -1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1376_
timestamp 1486834041
transform -1 0 45472 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1377_
timestamp 1486834041
transform -1 0 56560 0 1 44688
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1378_
timestamp 1486834041
transform 1 0 47936 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1379_
timestamp 1486834041
transform 1 0 38976 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1380_
timestamp 1486834041
transform 1 0 11200 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1381_
timestamp 1486834041
transform -1 0 10192 0 1 52528
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1382_
timestamp 1486834041
transform 1 0 11424 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1383_
timestamp 1486834041
transform 1 0 12992 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1384_
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1385_
timestamp 1486834041
transform -1 0 14896 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1386_
timestamp 1486834041
transform -1 0 22288 0 1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1387_
timestamp 1486834041
transform -1 0 12432 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1388_
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1389_
timestamp 1486834041
transform 1 0 36176 0 1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1390_
timestamp 1486834041
transform 1 0 36176 0 1 39984
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1391_
timestamp 1486834041
transform -1 0 35952 0 1 39984
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1392_
timestamp 1486834041
transform -1 0 37072 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1393_
timestamp 1486834041
transform 1 0 36624 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1394_
timestamp 1486834041
transform 1 0 34496 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1395_
timestamp 1486834041
transform 1 0 13888 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1396_
timestamp 1486834041
transform 1 0 15904 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1397_
timestamp 1486834041
transform 1 0 39312 0 -1 39984
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1398_
timestamp 1486834041
transform 1 0 37856 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1399_
timestamp 1486834041
transform 1 0 34272 0 1 41552
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1400_
timestamp 1486834041
transform 1 0 40320 0 1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1401_
timestamp 1486834041
transform 1 0 41440 0 1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1402_
timestamp 1486834041
transform 1 0 38976 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1403_
timestamp 1486834041
transform -1 0 35504 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1404_
timestamp 1486834041
transform 1 0 24416 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1405_
timestamp 1486834041
transform -1 0 20160 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1406_
timestamp 1486834041
transform 1 0 16688 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1407_
timestamp 1486834041
transform 1 0 19824 0 -1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1408_
timestamp 1486834041
transform -1 0 21056 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1409_
timestamp 1486834041
transform 1 0 15568 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1410_
timestamp 1486834041
transform 1 0 16912 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1411_
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1412_
timestamp 1486834041
transform -1 0 16352 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1413_
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1414_
timestamp 1486834041
transform 1 0 35056 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1415_
timestamp 1486834041
transform 1 0 28560 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1416_
timestamp 1486834041
transform 1 0 32368 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1417_
timestamp 1486834041
transform -1 0 32704 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1418_
timestamp 1486834041
transform 1 0 26320 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1419_
timestamp 1486834041
transform 1 0 13440 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1420_
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1421_
timestamp 1486834041
transform -1 0 24528 0 1 50960
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1422_
timestamp 1486834041
transform 1 0 24528 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1423_
timestamp 1486834041
transform 1 0 26320 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1424_
timestamp 1486834041
transform 1 0 23296 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1425_
timestamp 1486834041
transform 1 0 24752 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1426_
timestamp 1486834041
transform -1 0 25984 0 1 55664
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1427_
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1428_
timestamp 1486834041
transform 1 0 25312 0 -1 54096
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1429_
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1430_
timestamp 1486834041
transform 1 0 27776 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1431_
timestamp 1486834041
transform 1 0 26768 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1432_
timestamp 1486834041
transform 1 0 36176 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1433_
timestamp 1486834041
transform 1 0 32256 0 -1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1434_
timestamp 1486834041
transform 1 0 30352 0 -1 49392
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1435_
timestamp 1486834041
transform 1 0 36960 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1436_
timestamp 1486834041
transform 1 0 27104 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1437_
timestamp 1486834041
transform 1 0 12992 0 1 13328
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1438_
timestamp 1486834041
transform 1 0 15232 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1439_
timestamp 1486834041
transform 1 0 16576 0 -1 18032
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1440_
timestamp 1486834041
transform 1 0 13216 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1441_
timestamp 1486834041
transform 1 0 35280 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1442_
timestamp 1486834041
transform 1 0 6048 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1443_
timestamp 1486834041
transform -1 0 4592 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1444_
timestamp 1486834041
transform 1 0 5040 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1445_
timestamp 1486834041
transform -1 0 6048 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1446_
timestamp 1486834041
transform -1 0 8512 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1447_
timestamp 1486834041
transform -1 0 7616 0 -1 38416
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1448_
timestamp 1486834041
transform 1 0 6160 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1449_
timestamp 1486834041
transform -1 0 6496 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1450_
timestamp 1486834041
transform -1 0 6160 0 1 50960
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1451_
timestamp 1486834041
transform 1 0 19152 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1452_
timestamp 1486834041
transform 1 0 37408 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1453_
timestamp 1486834041
transform 1 0 36176 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1454_
timestamp 1486834041
transform 1 0 31472 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1455_
timestamp 1486834041
transform 1 0 34048 0 -1 55664
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1456_
timestamp 1486834041
transform -1 0 35616 0 1 54096
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1457_
timestamp 1486834041
transform 1 0 38416 0 1 54096
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1458_
timestamp 1486834041
transform 1 0 36288 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1459_
timestamp 1486834041
transform 1 0 37520 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1460_
timestamp 1486834041
transform -1 0 36288 0 -1 50960
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1461_
timestamp 1486834041
transform -1 0 38416 0 -1 55664
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1462_
timestamp 1486834041
transform 1 0 40432 0 -1 54096
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1463_
timestamp 1486834041
transform 1 0 38304 0 -1 44688
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1486834041
transform -1 0 37632 0 -1 41552
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1465_
timestamp 1486834041
transform -1 0 35952 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1466_
timestamp 1486834041
transform -1 0 35952 0 1 46256
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1467_
timestamp 1486834041
transform 1 0 34832 0 1 41552
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1468_
timestamp 1486834041
transform 1 0 39200 0 1 43120
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1469_
timestamp 1486834041
transform -1 0 37408 0 1 47824
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1470_
timestamp 1486834041
transform 1 0 26768 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1471_
timestamp 1486834041
transform -1 0 38304 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1472_
timestamp 1486834041
transform 1 0 32480 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1473_
timestamp 1486834041
transform 1 0 29008 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1474_
timestamp 1486834041
transform 1 0 29456 0 1 46256
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1475_
timestamp 1486834041
transform 1 0 30352 0 -1 44688
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1476_
timestamp 1486834041
transform -1 0 32032 0 -1 47824
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1477_
timestamp 1486834041
transform 1 0 34496 0 -1 52528
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1478_
timestamp 1486834041
transform 1 0 30352 0 -1 46256
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1479_
timestamp 1486834041
transform -1 0 30464 0 1 49392
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1480_
timestamp 1486834041
transform 1 0 30240 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1481_
timestamp 1486834041
transform 1 0 36176 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1482_
timestamp 1486834041
transform -1 0 32032 0 -1 49392
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1483_
timestamp 1486834041
transform 1 0 34608 0 1 52528
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1486834041
transform 1 0 38192 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1485_
timestamp 1486834041
transform 1 0 34272 0 -1 47824
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1486_
timestamp 1486834041
transform -1 0 32032 0 -1 44688
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1487_
timestamp 1486834041
transform -1 0 32032 0 -1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1488_
timestamp 1486834041
transform 1 0 32480 0 1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1489_
timestamp 1486834041
transform 1 0 36736 0 -1 44688
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1490_
timestamp 1486834041
transform 1 0 34720 0 1 47824
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1491_
timestamp 1486834041
transform 1 0 35168 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1492_
timestamp 1486834041
transform 1 0 36176 0 1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1493_
timestamp 1486834041
transform -1 0 34272 0 -1 47824
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1494_
timestamp 1486834041
transform -1 0 43008 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1495_
timestamp 1486834041
transform 1 0 41888 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1496_
timestamp 1486834041
transform -1 0 18368 0 -1 47824
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1497_
timestamp 1486834041
transform 1 0 18592 0 1 49392
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1498_
timestamp 1486834041
transform 1 0 16688 0 -1 49392
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1499_
timestamp 1486834041
transform 1 0 13888 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1500_
timestamp 1486834041
transform 1 0 10752 0 1 44688
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1501_
timestamp 1486834041
transform -1 0 12432 0 1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1502_
timestamp 1486834041
transform 1 0 47936 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1503_
timestamp 1486834041
transform 1 0 47040 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1504_
timestamp 1486834041
transform 1 0 44240 0 1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1505_
timestamp 1486834041
transform 1 0 47040 0 1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1506_
timestamp 1486834041
transform 1 0 48272 0 1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1507_
timestamp 1486834041
transform -1 0 50736 0 1 32144
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1508_
timestamp 1486834041
transform 1 0 43232 0 1 35280
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1509_
timestamp 1486834041
transform -1 0 55552 0 1 35280
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1510_
timestamp 1486834041
transform 1 0 52976 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1511_
timestamp 1486834041
transform 1 0 52976 0 -1 39984
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1512_
timestamp 1486834041
transform -1 0 53312 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1513_
timestamp 1486834041
transform 1 0 55776 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1514_
timestamp 1486834041
transform 1 0 53536 0 -1 36848
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1515_
timestamp 1486834041
transform -1 0 55216 0 -1 39984
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1516_
timestamp 1486834041
transform 1 0 55440 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1517_
timestamp 1486834041
transform -1 0 54432 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1518_
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1519_
timestamp 1486834041
transform 1 0 45920 0 -1 7056
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1520_
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1521_
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1522_
timestamp 1486834041
transform 1 0 50176 0 1 33712
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1523_
timestamp 1486834041
transform 1 0 51856 0 1 38416
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1524_
timestamp 1486834041
transform 1 0 55552 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1525_
timestamp 1486834041
transform 1 0 53984 0 -1 35280
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1526_
timestamp 1486834041
transform 1 0 50400 0 1 38416
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1527_
timestamp 1486834041
transform 1 0 55776 0 -1 35280
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1528_
timestamp 1486834041
transform -1 0 55552 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1529_
timestamp 1486834041
transform -1 0 51520 0 1 39984
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1530_
timestamp 1486834041
transform -1 0 53088 0 1 35280
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1531_
timestamp 1486834041
transform 1 0 48496 0 1 38416
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1532_
timestamp 1486834041
transform 1 0 8848 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1533_
timestamp 1486834041
transform 1 0 10192 0 -1 43120
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1534_
timestamp 1486834041
transform 1 0 10416 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1535_
timestamp 1486834041
transform -1 0 8512 0 -1 43120
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1536_
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1537_
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1538_
timestamp 1486834041
transform 1 0 3808 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1486834041
transform -1 0 3808 0 -1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1540_
timestamp 1486834041
transform -1 0 4816 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1541_
timestamp 1486834041
transform -1 0 4592 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1542_
timestamp 1486834041
transform 1 0 3808 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1486834041
transform -1 0 3808 0 -1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1544_
timestamp 1486834041
transform 1 0 4816 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1545_
timestamp 1486834041
transform -1 0 4592 0 1 25872
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1546_
timestamp 1486834041
transform 1 0 6608 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1547_
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1548_
timestamp 1486834041
transform 1 0 4928 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1549_
timestamp 1486834041
transform 1 0 5264 0 1 24304
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1550_
timestamp 1486834041
transform 1 0 7280 0 -1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1551_
timestamp 1486834041
transform 1 0 7392 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1552_
timestamp 1486834041
transform 1 0 6720 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1553_
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1554_
timestamp 1486834041
transform -1 0 6720 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1555_
timestamp 1486834041
transform 1 0 3920 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1556_
timestamp 1486834041
transform 1 0 3808 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1557_
timestamp 1486834041
transform 1 0 2800 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1558_
timestamp 1486834041
transform 1 0 3136 0 1 33712
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1559_
timestamp 1486834041
transform 1 0 4816 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1560_
timestamp 1486834041
transform -1 0 4592 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1486834041
transform -1 0 6048 0 1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1562_
timestamp 1486834041
transform 1 0 3472 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1563_
timestamp 1486834041
transform -1 0 4480 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1564_
timestamp 1486834041
transform 1 0 3584 0 1 32144
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1565_
timestamp 1486834041
transform 1 0 12432 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1566_
timestamp 1486834041
transform 1 0 11088 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1486834041
transform 1 0 12208 0 -1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1486834041
transform -1 0 13552 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1569_
timestamp 1486834041
transform 1 0 13552 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1570_
timestamp 1486834041
transform 1 0 12768 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1486834041
transform -1 0 12432 0 1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1572_
timestamp 1486834041
transform -1 0 12432 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1573_
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1574_
timestamp 1486834041
transform 1 0 8064 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1575_
timestamp 1486834041
transform 1 0 9520 0 1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1576_
timestamp 1486834041
transform 1 0 7616 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1577_
timestamp 1486834041
transform 1 0 10080 0 1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1578_
timestamp 1486834041
transform 1 0 8400 0 1 27440
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1579_
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1580_
timestamp 1486834041
transform -1 0 10752 0 1 44688
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1581_
timestamp 1486834041
transform 1 0 10976 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1582_
timestamp 1486834041
transform 1 0 11088 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1583_
timestamp 1486834041
transform 1 0 6832 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1584_
timestamp 1486834041
transform -1 0 6496 0 1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1585_
timestamp 1486834041
transform 1 0 4928 0 1 43120
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1486834041
transform 1 0 7952 0 -1 44688
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1587_
timestamp 1486834041
transform 1 0 8848 0 1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1588_
timestamp 1486834041
transform 1 0 8400 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1589_
timestamp 1486834041
transform -1 0 9968 0 -1 43120
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1590_
timestamp 1486834041
transform -1 0 13776 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1591_
timestamp 1486834041
transform 1 0 3136 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1592_
timestamp 1486834041
transform -1 0 2016 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1593_
timestamp 1486834041
transform 1 0 3360 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1594_
timestamp 1486834041
transform -1 0 4592 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1595_
timestamp 1486834041
transform 1 0 5600 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1596_
timestamp 1486834041
transform -1 0 5488 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1597_
timestamp 1486834041
transform 1 0 4928 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1486834041
transform -1 0 2688 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1599_
timestamp 1486834041
transform 1 0 3136 0 1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1600_
timestamp 1486834041
transform -1 0 8512 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1601_
timestamp 1486834041
transform 1 0 5376 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1602_
timestamp 1486834041
transform -1 0 5264 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1603_
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1604_
timestamp 1486834041
transform 1 0 7056 0 1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1605_
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1606_
timestamp 1486834041
transform 1 0 5824 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1607_
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1608_
timestamp 1486834041
transform 1 0 5376 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1609_
timestamp 1486834041
transform -1 0 7840 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1486834041
transform -1 0 9296 0 -1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1611_
timestamp 1486834041
transform 1 0 9744 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1612_
timestamp 1486834041
transform 1 0 11312 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1613_
timestamp 1486834041
transform 1 0 10080 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1486834041
transform 1 0 11200 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1615_
timestamp 1486834041
transform 1 0 9968 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1616_
timestamp 1486834041
transform 1 0 11872 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1617_
timestamp 1486834041
transform 1 0 8848 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1618_
timestamp 1486834041
transform -1 0 9968 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1619_
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1620_
timestamp 1486834041
transform 1 0 8848 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1621_
timestamp 1486834041
transform 1 0 9632 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1622_
timestamp 1486834041
transform -1 0 13664 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1486834041
transform -1 0 12320 0 1 19600
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1624_
timestamp 1486834041
transform 1 0 10640 0 1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1625_
timestamp 1486834041
transform 1 0 8848 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1626_
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1486834041
transform 1 0 10976 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1628_
timestamp 1486834041
transform 1 0 9184 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1629_
timestamp 1486834041
transform -1 0 9632 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1630_
timestamp 1486834041
transform 1 0 10976 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1631_
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1486834041
transform -1 0 16352 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1633_
timestamp 1486834041
transform 1 0 15680 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1634_
timestamp 1486834041
transform -1 0 15680 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1635_
timestamp 1486834041
transform 1 0 16464 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1636_
timestamp 1486834041
transform 1 0 19264 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1637_
timestamp 1486834041
transform 1 0 16576 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1638_
timestamp 1486834041
transform -1 0 17584 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1639_
timestamp 1486834041
transform 1 0 16688 0 1 25872
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1640_
timestamp 1486834041
transform 1 0 4928 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1641_
timestamp 1486834041
transform 1 0 4592 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1642_
timestamp 1486834041
transform 1 0 4928 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1643_
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1644_
timestamp 1486834041
transform 1 0 1344 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1645_
timestamp 1486834041
transform -1 0 18704 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1646_
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1647_
timestamp 1486834041
transform -1 0 17920 0 1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1648_
timestamp 1486834041
transform 1 0 2576 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1649_
timestamp 1486834041
transform 1 0 3136 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1650_
timestamp 1486834041
transform -1 0 2576 0 -1 22736
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1651_
timestamp 1486834041
transform 1 0 16688 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1652_
timestamp 1486834041
transform 1 0 16688 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1653_
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1654_
timestamp 1486834041
transform 1 0 9968 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1655_
timestamp 1486834041
transform 1 0 9856 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1656_
timestamp 1486834041
transform 1 0 6832 0 -1 33712
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1657_
timestamp 1486834041
transform 1 0 28336 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1658_
timestamp 1486834041
transform 1 0 28000 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1659_
timestamp 1486834041
transform -1 0 31920 0 -1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1660_
timestamp 1486834041
transform 1 0 37744 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1661_
timestamp 1486834041
transform 1 0 37072 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1662_
timestamp 1486834041
transform -1 0 39872 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1663_
timestamp 1486834041
transform 1 0 30576 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1664_
timestamp 1486834041
transform 1 0 30464 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1665_
timestamp 1486834041
transform -1 0 33936 0 -1 2352
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1486834041
transform 1 0 31472 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1667_
timestamp 1486834041
transform -1 0 35280 0 1 18032
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1668_
timestamp 1486834041
transform 1 0 30576 0 -1 19600
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1486834041
transform -1 0 32032 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1670_
timestamp 1486834041
transform 1 0 32368 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1671_
timestamp 1486834041
transform -1 0 34160 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1672_
timestamp 1486834041
transform -1 0 35392 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1673_
timestamp 1486834041
transform 1 0 43344 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1674_
timestamp 1486834041
transform 1 0 20608 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1675_
timestamp 1486834041
transform 1 0 20608 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1676_
timestamp 1486834041
transform 1 0 18592 0 1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1677_
timestamp 1486834041
transform 1 0 20608 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1678_
timestamp 1486834041
transform 1 0 20608 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1679_
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1680_
timestamp 1486834041
transform -1 0 20608 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1681_
timestamp 1486834041
transform 1 0 21840 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1682_
timestamp 1486834041
transform 1 0 21504 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1683_
timestamp 1486834041
transform 1 0 20384 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1684_
timestamp 1486834041
transform 1 0 19600 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1685_
timestamp 1486834041
transform 1 0 20496 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1686_
timestamp 1486834041
transform 1 0 28112 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1687_
timestamp 1486834041
transform 1 0 28336 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1688_
timestamp 1486834041
transform -1 0 31584 0 -1 39984
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1689_
timestamp 1486834041
transform 1 0 34496 0 -1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1690_
timestamp 1486834041
transform 1 0 35056 0 -1 32144
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1486834041
transform 1 0 35392 0 1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1692_
timestamp 1486834041
transform -1 0 37632 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1693_
timestamp 1486834041
transform 1 0 38416 0 1 32144
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1694_
timestamp 1486834041
transform 1 0 36176 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1486834041
transform 1 0 38080 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1696_
timestamp 1486834041
transform -1 0 55552 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1697_
timestamp 1486834041
transform 1 0 30800 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1698_
timestamp 1486834041
transform 1 0 30464 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1699_
timestamp 1486834041
transform -1 0 32032 0 -1 43120
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1700_
timestamp 1486834041
transform 1 0 14224 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1701_
timestamp 1486834041
transform 1 0 14336 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1702_
timestamp 1486834041
transform -1 0 16352 0 -1 38416
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1703_
timestamp 1486834041
transform 1 0 26544 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1704_
timestamp 1486834041
transform 1 0 26544 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1705_
timestamp 1486834041
transform 1 0 24864 0 -1 49392
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1706_
timestamp 1486834041
transform -1 0 26320 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1707_
timestamp 1486834041
transform -1 0 26320 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1708_
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1709_
timestamp 1486834041
transform 1 0 29008 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1710_
timestamp 1486834041
transform 1 0 28448 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1711_
timestamp 1486834041
transform 1 0 28896 0 1 54096
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1712_
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1713_
timestamp 1486834041
transform 1 0 24080 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1714_
timestamp 1486834041
transform 1 0 22512 0 -1 38416
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1715_
timestamp 1486834041
transform -1 0 4592 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1716_
timestamp 1486834041
transform 1 0 1008 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1717_
timestamp 1486834041
transform -1 0 4928 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1718_
timestamp 1486834041
transform 1 0 1792 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1719_
timestamp 1486834041
transform -1 0 41440 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1720_
timestamp 1486834041
transform -1 0 39760 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1721_
timestamp 1486834041
transform 1 0 32704 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1722_
timestamp 1486834041
transform 1 0 31808 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1723_
timestamp 1486834041
transform 1 0 23408 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1724_
timestamp 1486834041
transform 1 0 24528 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1725_
timestamp 1486834041
transform 1 0 22848 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1726_
timestamp 1486834041
transform 1 0 23408 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1727_
timestamp 1486834041
transform 1 0 36288 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1728_
timestamp 1486834041
transform 1 0 38080 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1729_
timestamp 1486834041
transform 1 0 11648 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1730_
timestamp 1486834041
transform 1 0 42000 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1731_
timestamp 1486834041
transform 1 0 12656 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1732_
timestamp 1486834041
transform 1 0 12992 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1733_
timestamp 1486834041
transform 1 0 12768 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1734_
timestamp 1486834041
transform 1 0 12656 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1735_
timestamp 1486834041
transform -1 0 4928 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1736_
timestamp 1486834041
transform 1 0 1008 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1737_
timestamp 1486834041
transform -1 0 4592 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1738_
timestamp 1486834041
transform -1 0 4592 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1739_
timestamp 1486834041
transform -1 0 35840 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1740_
timestamp 1486834041
transform -1 0 35840 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1486834041
transform 1 0 39200 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1742_
timestamp 1486834041
transform -1 0 41328 0 1 18032
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1743_
timestamp 1486834041
transform -1 0 40992 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1744_
timestamp 1486834041
transform 1 0 42336 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1745_
timestamp 1486834041
transform 1 0 40656 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1746_
timestamp 1486834041
transform 1 0 39872 0 1 21168
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1747_
timestamp 1486834041
transform 1 0 36848 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1748_
timestamp 1486834041
transform 1 0 38752 0 -1 21168
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1749_
timestamp 1486834041
transform 1 0 41328 0 -1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1750_
timestamp 1486834041
transform -1 0 42336 0 -1 21168
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1751_
timestamp 1486834041
transform 1 0 28784 0 -1 55664
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1752_
timestamp 1486834041
transform 1 0 40096 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1753_
timestamp 1486834041
transform -1 0 42336 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1754_
timestamp 1486834041
transform -1 0 42000 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1755_
timestamp 1486834041
transform 1 0 40208 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1756_
timestamp 1486834041
transform 1 0 43008 0 1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1757_
timestamp 1486834041
transform 1 0 38976 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1758_
timestamp 1486834041
transform 1 0 40320 0 -1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1759_
timestamp 1486834041
transform 1 0 41552 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1760_
timestamp 1486834041
transform 1 0 42336 0 -1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1761_
timestamp 1486834041
transform 1 0 40544 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1762_
timestamp 1486834041
transform 1 0 40992 0 1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1763_
timestamp 1486834041
transform -1 0 43008 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1764_
timestamp 1486834041
transform -1 0 50400 0 -1 52528
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1765_
timestamp 1486834041
transform -1 0 44912 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1766_
timestamp 1486834041
transform -1 0 46032 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1767_
timestamp 1486834041
transform -1 0 45136 0 1 50960
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1768_
timestamp 1486834041
transform 1 0 45808 0 -1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1486834041
transform 1 0 46928 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1770_
timestamp 1486834041
transform 1 0 50064 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1771_
timestamp 1486834041
transform 1 0 49504 0 1 18032
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1772_
timestamp 1486834041
transform 1 0 49056 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1773_
timestamp 1486834041
transform 1 0 48496 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1774_
timestamp 1486834041
transform 1 0 51072 0 1 21168
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1775_
timestamp 1486834041
transform 1 0 53424 0 -1 24304
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1776_
timestamp 1486834041
transform 1 0 51856 0 1 24304
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1777_
timestamp 1486834041
transform 1 0 46592 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1778_
timestamp 1486834041
transform 1 0 47152 0 -1 29008
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1779_
timestamp 1486834041
transform 1 0 45136 0 1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1780_
timestamp 1486834041
transform 1 0 44800 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1781_
timestamp 1486834041
transform 1 0 47040 0 -1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1782_
timestamp 1486834041
transform 1 0 51856 0 1 27440
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1783_
timestamp 1486834041
transform 1 0 46032 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1784_
timestamp 1486834041
transform 1 0 47936 0 -1 38416
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1785_
timestamp 1486834041
transform 1 0 47936 0 -1 39984
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1486834041
transform 1 0 46816 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1787_
timestamp 1486834041
transform 1 0 48832 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1788_
timestamp 1486834041
transform -1 0 47712 0 -1 38416
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1789_
timestamp 1486834041
transform 1 0 48048 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1790_
timestamp 1486834041
transform 1 0 23632 0 1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1486834041
transform 1 0 44016 0 1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1792_
timestamp 1486834041
transform -1 0 51632 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1793_
timestamp 1486834041
transform 1 0 52528 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1794_
timestamp 1486834041
transform 1 0 49504 0 1 50960
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1795_
timestamp 1486834041
transform -1 0 49168 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1486834041
transform 1 0 46256 0 1 46256
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1797_
timestamp 1486834041
transform 1 0 43232 0 1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1798_
timestamp 1486834041
transform -1 0 48272 0 1 49392
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1799_
timestamp 1486834041
transform 1 0 49168 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1800_
timestamp 1486834041
transform 1 0 47936 0 -1 49392
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1801_
timestamp 1486834041
transform 1 0 42336 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1486834041
transform 1 0 28336 0 1 54096
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1803_
timestamp 1486834041
transform 1 0 28448 0 1 50960
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1804_
timestamp 1486834041
transform -1 0 44912 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1805_
timestamp 1486834041
transform 1 0 44912 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1806_
timestamp 1486834041
transform 1 0 42560 0 1 50960
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1807_
timestamp 1486834041
transform -1 0 55552 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1808_
timestamp 1486834041
transform -1 0 55440 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1809_
timestamp 1486834041
transform 1 0 53648 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1810_
timestamp 1486834041
transform 1 0 53088 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1811_
timestamp 1486834041
transform 1 0 53312 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1812_
timestamp 1486834041
transform 1 0 54096 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1813_
timestamp 1486834041
transform 1 0 53312 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1814_
timestamp 1486834041
transform 1 0 52864 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1815_
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1816_
timestamp 1486834041
transform 1 0 49840 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1817_
timestamp 1486834041
transform -1 0 53760 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1818_
timestamp 1486834041
transform -1 0 51520 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1819_
timestamp 1486834041
transform 1 0 49504 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1820_
timestamp 1486834041
transform 1 0 50064 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1821_
timestamp 1486834041
transform -1 0 54432 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1822_
timestamp 1486834041
transform 1 0 49952 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1823_
timestamp 1486834041
transform -1 0 50288 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1824_
timestamp 1486834041
transform -1 0 50736 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1825_
timestamp 1486834041
transform 1 0 47824 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1826_
timestamp 1486834041
transform 1 0 51184 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1827_
timestamp 1486834041
transform -1 0 55552 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1828_
timestamp 1486834041
transform -1 0 55328 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1829_
timestamp 1486834041
transform 1 0 54208 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1830_
timestamp 1486834041
transform -1 0 54320 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1831_
timestamp 1486834041
transform 1 0 53872 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1832_
timestamp 1486834041
transform -1 0 54096 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1833_
timestamp 1486834041
transform 1 0 51632 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1834_
timestamp 1486834041
transform 1 0 53088 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1835_
timestamp 1486834041
transform 1 0 50512 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1836_
timestamp 1486834041
transform 1 0 49392 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1837_
timestamp 1486834041
transform 1 0 53312 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1838_
timestamp 1486834041
transform 1 0 53536 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1839_
timestamp 1486834041
transform 1 0 53312 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1840_
timestamp 1486834041
transform 1 0 49392 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1841_
timestamp 1486834041
transform 1 0 49392 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1842_
timestamp 1486834041
transform 1 0 49280 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1843_
timestamp 1486834041
transform -1 0 50512 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1844_
timestamp 1486834041
transform 1 0 51856 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1845_
timestamp 1486834041
transform 1 0 50288 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1846_
timestamp 1486834041
transform -1 0 55888 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1847_
timestamp 1486834041
transform 1 0 50176 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1848_
timestamp 1486834041
transform 1 0 53312 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1849_
timestamp 1486834041
transform 1 0 50176 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1850_
timestamp 1486834041
transform 1 0 53200 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1851_
timestamp 1486834041
transform -1 0 54656 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1852_
timestamp 1486834041
transform 1 0 53536 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1853_
timestamp 1486834041
transform 1 0 51856 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1854_
timestamp 1486834041
transform 1 0 53536 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1855_
timestamp 1486834041
transform 1 0 50960 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1856_
timestamp 1486834041
transform 1 0 54096 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1857_
timestamp 1486834041
transform 1 0 48832 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1858_
timestamp 1486834041
transform 1 0 52976 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1859_
timestamp 1486834041
transform 1 0 49280 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1860_
timestamp 1486834041
transform 1 0 53312 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1861_
timestamp 1486834041
transform 1 0 47040 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1862_
timestamp 1486834041
transform 1 0 47152 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1863_
timestamp 1486834041
transform -1 0 50176 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1864_
timestamp 1486834041
transform 1 0 47936 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1865_
timestamp 1486834041
transform 1 0 53088 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1866_
timestamp 1486834041
transform 1 0 48496 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1867_
timestamp 1486834041
transform 1 0 48496 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1868_
timestamp 1486834041
transform 1 0 48496 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1869_
timestamp 1486834041
transform 1 0 48720 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1870_
timestamp 1486834041
transform 1 0 48496 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1871_
timestamp 1486834041
transform 1 0 52752 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1872_
timestamp 1486834041
transform 1 0 52080 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1873_
timestamp 1486834041
transform 1 0 54320 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1874_
timestamp 1486834041
transform 1 0 51072 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1875_
timestamp 1486834041
transform 1 0 50736 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1876_
timestamp 1486834041
transform 1 0 52864 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1877_
timestamp 1486834041
transform 1 0 53312 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1878_
timestamp 1486834041
transform -1 0 56336 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1879_
timestamp 1486834041
transform 1 0 51856 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1880_
timestamp 1486834041
transform 1 0 46256 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1881_
timestamp 1486834041
transform 1 0 48048 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1882_
timestamp 1486834041
transform 1 0 46256 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1883_
timestamp 1486834041
transform 1 0 53872 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1884_
timestamp 1486834041
transform 1 0 48160 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1885_
timestamp 1486834041
transform -1 0 56560 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1886_
timestamp 1486834041
transform 1 0 48944 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1887_
timestamp 1486834041
transform 1 0 50624 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1888_
timestamp 1486834041
transform 1 0 48832 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1889_
timestamp 1486834041
transform 1 0 52080 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1890_
timestamp 1486834041
transform 1 0 48384 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1891_
timestamp 1486834041
transform -1 0 55776 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1892_
timestamp 1486834041
transform 1 0 52752 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1893_
timestamp 1486834041
transform -1 0 55776 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1894_
timestamp 1486834041
transform 1 0 51856 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1895_
timestamp 1486834041
transform 1 0 49392 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1896_
timestamp 1486834041
transform 1 0 49392 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1897_
timestamp 1486834041
transform -1 0 54432 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1898_
timestamp 1486834041
transform -1 0 53872 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1899_
timestamp 1486834041
transform 1 0 45472 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1900_
timestamp 1486834041
transform 1 0 48496 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1901_
timestamp 1486834041
transform 1 0 50064 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1902_
timestamp 1486834041
transform 1 0 40432 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1903_
timestamp 1486834041
transform 1 0 44016 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1904_
timestamp 1486834041
transform 1 0 40320 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1905_
timestamp 1486834041
transform -1 0 46256 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1906_
timestamp 1486834041
transform 1 0 40096 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1907_
timestamp 1486834041
transform -1 0 45136 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1908_
timestamp 1486834041
transform 1 0 40208 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1909_
timestamp 1486834041
transform 1 0 43008 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1910_
timestamp 1486834041
transform -1 0 48608 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1911_
timestamp 1486834041
transform -1 0 48496 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1912_
timestamp 1486834041
transform -1 0 46256 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1913_
timestamp 1486834041
transform 1 0 43120 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1914_
timestamp 1486834041
transform 1 0 46704 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1915_
timestamp 1486834041
transform 1 0 45472 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1916_
timestamp 1486834041
transform -1 0 45808 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1917_
timestamp 1486834041
transform 1 0 43120 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1918_
timestamp 1486834041
transform 1 0 44576 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1919_
timestamp 1486834041
transform 1 0 40432 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1920_
timestamp 1486834041
transform 1 0 46816 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1921_
timestamp 1486834041
transform 1 0 38864 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1922_
timestamp 1486834041
transform -1 0 42336 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1923_
timestamp 1486834041
transform 1 0 37856 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1924_
timestamp 1486834041
transform 1 0 37296 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1925_
timestamp 1486834041
transform 1 0 35952 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1926_
timestamp 1486834041
transform 1 0 35056 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1927_
timestamp 1486834041
transform 1 0 36736 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1928_
timestamp 1486834041
transform -1 0 38416 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1929_
timestamp 1486834041
transform -1 0 34496 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1930_
timestamp 1486834041
transform 1 0 37632 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1931_
timestamp 1486834041
transform -1 0 35056 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1932_
timestamp 1486834041
transform 1 0 37408 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1933_
timestamp 1486834041
transform 1 0 32368 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1934_
timestamp 1486834041
transform 1 0 35056 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1935_
timestamp 1486834041
transform 1 0 32032 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1936_
timestamp 1486834041
transform 1 0 36176 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1937_
timestamp 1486834041
transform 1 0 40096 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1938_
timestamp 1486834041
transform 1 0 37184 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1939_
timestamp 1486834041
transform 1 0 42336 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1940_
timestamp 1486834041
transform 1 0 32816 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1941_
timestamp 1486834041
transform -1 0 34496 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1942_
timestamp 1486834041
transform -1 0 36736 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1943_
timestamp 1486834041
transform -1 0 34496 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1944_
timestamp 1486834041
transform 1 0 32816 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1945_
timestamp 1486834041
transform 1 0 30016 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1946_
timestamp 1486834041
transform 1 0 33152 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1947_
timestamp 1486834041
transform 1 0 30576 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1948_
timestamp 1486834041
transform -1 0 34496 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1949_
timestamp 1486834041
transform -1 0 34496 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1950_
timestamp 1486834041
transform -1 0 36736 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1951_
timestamp 1486834041
transform 1 0 29904 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1952_
timestamp 1486834041
transform -1 0 32704 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1953_
timestamp 1486834041
transform -1 0 34384 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1954_
timestamp 1486834041
transform 1 0 32704 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1955_
timestamp 1486834041
transform -1 0 34944 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1956_
timestamp 1486834041
transform 1 0 40096 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1957_
timestamp 1486834041
transform 1 0 36736 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1958_
timestamp 1486834041
transform 1 0 41440 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1959_
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1960_
timestamp 1486834041
transform 1 0 8848 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1961_
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1962_
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1963_
timestamp 1486834041
transform -1 0 3136 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1964_
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1965_
timestamp 1486834041
transform 1 0 1008 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1966_
timestamp 1486834041
transform -1 0 3136 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1967_
timestamp 1486834041
transform -1 0 7056 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1968_
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1969_
timestamp 1486834041
transform 1 0 10192 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1970_
timestamp 1486834041
transform 1 0 11872 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1971_
timestamp 1486834041
transform 1 0 10192 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1972_
timestamp 1486834041
transform -1 0 15680 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1973_
timestamp 1486834041
transform -1 0 14896 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1974_
timestamp 1486834041
transform 1 0 11872 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1975_
timestamp 1486834041
transform 1 0 10192 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1976_
timestamp 1486834041
transform 1 0 10192 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1977_
timestamp 1486834041
transform 1 0 23184 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1978_
timestamp 1486834041
transform 1 0 20944 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1979_
timestamp 1486834041
transform 1 0 18032 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1980_
timestamp 1486834041
transform -1 0 30576 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1981_
timestamp 1486834041
transform 1 0 28672 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1982_
timestamp 1486834041
transform 1 0 28224 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1983_
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1984_
timestamp 1486834041
transform 1 0 21392 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1985_
timestamp 1486834041
transform 1 0 20496 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1986_
timestamp 1486834041
transform 1 0 21392 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1987_
timestamp 1486834041
transform 1 0 21392 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1988_
timestamp 1486834041
transform -1 0 27776 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1989_
timestamp 1486834041
transform 1 0 42336 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1990_
timestamp 1486834041
transform 1 0 40992 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1991_
timestamp 1486834041
transform 1 0 9408 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1992_
timestamp 1486834041
transform -1 0 14896 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1993_
timestamp 1486834041
transform -1 0 42336 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1994_
timestamp 1486834041
transform 1 0 36736 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1995_
timestamp 1486834041
transform 1 0 33712 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1996_
timestamp 1486834041
transform 1 0 36176 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1997_
timestamp 1486834041
transform 1 0 10192 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1998_
timestamp 1486834041
transform 1 0 12656 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1999_
timestamp 1486834041
transform 1 0 14112 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2000_
timestamp 1486834041
transform 1 0 28560 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2001_
timestamp 1486834041
transform -1 0 34496 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2002_
timestamp 1486834041
transform -1 0 32816 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2003_
timestamp 1486834041
transform 1 0 35056 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2004_
timestamp 1486834041
transform -1 0 38416 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2005_
timestamp 1486834041
transform 1 0 36176 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2006_
timestamp 1486834041
transform 1 0 25872 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2007_
timestamp 1486834041
transform 1 0 25872 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2008_
timestamp 1486834041
transform 1 0 28448 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2009_
timestamp 1486834041
transform 1 0 18256 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2010_
timestamp 1486834041
transform 1 0 18032 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2011_
timestamp 1486834041
transform 1 0 18144 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2012_
timestamp 1486834041
transform 1 0 17360 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2013_
timestamp 1486834041
transform 1 0 18368 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2014_
timestamp 1486834041
transform 1 0 20720 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2015_
timestamp 1486834041
transform 1 0 18368 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2016_
timestamp 1486834041
transform 1 0 17472 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2017_
timestamp 1486834041
transform -1 0 26656 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2018_
timestamp 1486834041
transform 1 0 21168 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2019_
timestamp 1486834041
transform 1 0 20608 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2020_
timestamp 1486834041
transform 1 0 21952 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2021_
timestamp 1486834041
transform 1 0 24192 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2022_
timestamp 1486834041
transform -1 0 26320 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2023_
timestamp 1486834041
transform 1 0 21168 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2024_
timestamp 1486834041
transform 1 0 21392 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2025_
timestamp 1486834041
transform 1 0 32256 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2026_
timestamp 1486834041
transform 1 0 29792 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2027_
timestamp 1486834041
transform 1 0 32704 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2028_
timestamp 1486834041
transform -1 0 34496 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2029_
timestamp 1486834041
transform 1 0 36288 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2030_
timestamp 1486834041
transform 1 0 35840 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2031_
timestamp 1486834041
transform 1 0 36960 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2032_
timestamp 1486834041
transform 1 0 37856 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2033_
timestamp 1486834041
transform 1 0 32256 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2034_
timestamp 1486834041
transform 1 0 28336 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2035_
timestamp 1486834041
transform 1 0 32256 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2036_
timestamp 1486834041
transform 1 0 29232 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2037_
timestamp 1486834041
transform 1 0 29792 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2038_
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2039_
timestamp 1486834041
transform 1 0 36512 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2040_
timestamp 1486834041
transform 1 0 36400 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2041_
timestamp 1486834041
transform -1 0 42896 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2042_
timestamp 1486834041
transform 1 0 22848 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2043_
timestamp 1486834041
transform 1 0 28000 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2044_
timestamp 1486834041
transform 1 0 28336 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2045_
timestamp 1486834041
transform -1 0 7616 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2046_
timestamp 1486834041
transform -1 0 4480 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2047_
timestamp 1486834041
transform -1 0 14560 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2048_
timestamp 1486834041
transform -1 0 4816 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2049_
timestamp 1486834041
transform 1 0 1008 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2050_
timestamp 1486834041
transform -1 0 3136 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2051_
timestamp 1486834041
transform -1 0 13328 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2052_
timestamp 1486834041
transform -1 0 10752 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2053_
timestamp 1486834041
transform 1 0 7728 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2054_
timestamp 1486834041
transform 1 0 9968 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2055_
timestamp 1486834041
transform -1 0 10192 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2056_
timestamp 1486834041
transform 1 0 14112 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2057_
timestamp 1486834041
transform 1 0 14112 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2058_
timestamp 1486834041
transform 1 0 14112 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2059_
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2060_
timestamp 1486834041
transform 1 0 1456 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2061_
timestamp 1486834041
transform -1 0 3136 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2062_
timestamp 1486834041
transform 1 0 12880 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2063_
timestamp 1486834041
transform 1 0 14112 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2064_
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2065_
timestamp 1486834041
transform 1 0 2688 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2066_
timestamp 1486834041
transform 1 0 2352 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2067_
timestamp 1486834041
transform -1 0 3136 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2068_
timestamp 1486834041
transform 1 0 1792 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2069_
timestamp 1486834041
transform 1 0 13776 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2070_
timestamp 1486834041
transform 1 0 14000 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2071_
timestamp 1486834041
transform 1 0 14112 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2072_
timestamp 1486834041
transform -1 0 18816 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2073_
timestamp 1486834041
transform 1 0 44576 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2074_
timestamp 1486834041
transform 1 0 46256 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2075_
timestamp 1486834041
transform -1 0 46256 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2076_
timestamp 1486834041
transform 1 0 44688 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2077_
timestamp 1486834041
transform 1 0 33488 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2078_
timestamp 1486834041
transform -1 0 37072 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2079_
timestamp 1486834041
transform 1 0 41216 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2080_
timestamp 1486834041
transform 1 0 43680 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2081_
timestamp 1486834041
transform -1 0 50176 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2082_
timestamp 1486834041
transform -1 0 49504 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2083_
timestamp 1486834041
transform 1 0 45472 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2084_
timestamp 1486834041
transform 1 0 45360 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2085_
timestamp 1486834041
transform 1 0 43344 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2086_
timestamp 1486834041
transform -1 0 49616 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2087_
timestamp 1486834041
transform 1 0 33488 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2088_
timestamp 1486834041
transform 1 0 34720 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2089_
timestamp 1486834041
transform -1 0 46256 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2090_
timestamp 1486834041
transform 1 0 44352 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2091_
timestamp 1486834041
transform -1 0 53424 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2092_
timestamp 1486834041
transform -1 0 51520 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2093_
timestamp 1486834041
transform 1 0 44240 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2094_
timestamp 1486834041
transform 1 0 44800 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2095_
timestamp 1486834041
transform 1 0 40096 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2096_
timestamp 1486834041
transform 1 0 40880 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2097_
timestamp 1486834041
transform 1 0 21952 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2098_
timestamp 1486834041
transform 1 0 25312 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2099_
timestamp 1486834041
transform -1 0 43344 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2100_
timestamp 1486834041
transform 1 0 41440 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2101_
timestamp 1486834041
transform -1 0 50176 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2102_
timestamp 1486834041
transform 1 0 44688 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2103_
timestamp 1486834041
transform 1 0 44688 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2104_
timestamp 1486834041
transform 1 0 46256 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2105_
timestamp 1486834041
transform -1 0 42336 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2106_
timestamp 1486834041
transform -1 0 43680 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2107_
timestamp 1486834041
transform 1 0 22176 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2108_
timestamp 1486834041
transform 1 0 25872 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2109_
timestamp 1486834041
transform 1 0 43680 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2110_
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2111_
timestamp 1486834041
transform 1 0 46256 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2112_
timestamp 1486834041
transform 1 0 44016 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2113_
timestamp 1486834041
transform 1 0 37072 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2114_
timestamp 1486834041
transform -1 0 42336 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2115_
timestamp 1486834041
transform 1 0 37632 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2116_
timestamp 1486834041
transform 1 0 40096 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2117_
timestamp 1486834041
transform 1 0 19712 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2118_
timestamp 1486834041
transform 1 0 21952 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2119_
timestamp 1486834041
transform 1 0 38416 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2120_
timestamp 1486834041
transform 1 0 40656 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2121_
timestamp 1486834041
transform -1 0 52640 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2122_
timestamp 1486834041
transform 1 0 45808 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2123_
timestamp 1486834041
transform 1 0 37072 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2124_
timestamp 1486834041
transform 1 0 39312 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2125_
timestamp 1486834041
transform 1 0 36848 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2126_
timestamp 1486834041
transform 1 0 38864 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2127_
timestamp 1486834041
transform 1 0 21840 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2128_
timestamp 1486834041
transform 1 0 21840 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2129_
timestamp 1486834041
transform 1 0 40768 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2130_
timestamp 1486834041
transform 1 0 41328 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2131_
timestamp 1486834041
transform -1 0 47712 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2132_
timestamp 1486834041
transform 1 0 44912 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2133_
timestamp 1486834041
transform 1 0 36736 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2134_
timestamp 1486834041
transform 1 0 36960 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2135_
timestamp 1486834041
transform -1 0 34496 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2136_
timestamp 1486834041
transform 1 0 32592 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2137_
timestamp 1486834041
transform 1 0 23632 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2138_
timestamp 1486834041
transform 1 0 25872 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2139_
timestamp 1486834041
transform 1 0 34720 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2140_
timestamp 1486834041
transform 1 0 36176 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2141_
timestamp 1486834041
transform -1 0 43792 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2142_
timestamp 1486834041
transform 1 0 40320 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2143_
timestamp 1486834041
transform 1 0 34496 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2144_
timestamp 1486834041
transform 1 0 34496 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2145_
timestamp 1486834041
transform 1 0 31024 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2146_
timestamp 1486834041
transform -1 0 35504 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2147_
timestamp 1486834041
transform 1 0 23632 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2148_
timestamp 1486834041
transform 1 0 25872 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2149_
timestamp 1486834041
transform 1 0 34496 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2150_
timestamp 1486834041
transform 1 0 36736 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2151_
timestamp 1486834041
transform 1 0 41104 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2152_
timestamp 1486834041
transform -1 0 44800 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2153_
timestamp 1486834041
transform 1 0 13776 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2154_
timestamp 1486834041
transform 1 0 12768 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2155_
timestamp 1486834041
transform 1 0 5824 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2156_
timestamp 1486834041
transform 1 0 5488 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2157_
timestamp 1486834041
transform -1 0 19712 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2158_
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2159_
timestamp 1486834041
transform -1 0 10976 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2160_
timestamp 1486834041
transform 1 0 7280 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2161_
timestamp 1486834041
transform 1 0 40656 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2162_
timestamp 1486834041
transform -1 0 45136 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2163_
timestamp 1486834041
transform 1 0 44576 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2164_
timestamp 1486834041
transform 1 0 45136 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2165_
timestamp 1486834041
transform 1 0 16912 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2166_
timestamp 1486834041
transform 1 0 17248 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2167_
timestamp 1486834041
transform 1 0 26880 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2168_
timestamp 1486834041
transform 1 0 28560 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2169_
timestamp 1486834041
transform -1 0 46816 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2170_
timestamp 1486834041
transform 1 0 44576 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2171_
timestamp 1486834041
transform 1 0 44016 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2172_
timestamp 1486834041
transform 1 0 42336 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2173_
timestamp 1486834041
transform 1 0 21952 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2174_
timestamp 1486834041
transform 1 0 21952 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2175_
timestamp 1486834041
transform 1 0 25760 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2176_
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2177_
timestamp 1486834041
transform 1 0 41552 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2178_
timestamp 1486834041
transform -1 0 46256 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2179_
timestamp 1486834041
transform -1 0 45920 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2180_
timestamp 1486834041
transform 1 0 44016 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2181_
timestamp 1486834041
transform 1 0 22736 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2182_
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2183_
timestamp 1486834041
transform 1 0 21392 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2184_
timestamp 1486834041
transform -1 0 26656 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2185_
timestamp 1486834041
transform 1 0 34496 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2186_
timestamp 1486834041
transform 1 0 34832 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2187_
timestamp 1486834041
transform -1 0 38304 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2188_
timestamp 1486834041
transform 1 0 32816 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2189_
timestamp 1486834041
transform 1 0 21952 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2190_
timestamp 1486834041
transform 1 0 20720 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2191_
timestamp 1486834041
transform 1 0 18032 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2192_
timestamp 1486834041
transform 1 0 17472 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2193_
timestamp 1486834041
transform 1 0 42448 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2194_
timestamp 1486834041
transform -1 0 46256 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2195_
timestamp 1486834041
transform -1 0 34496 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2196_
timestamp 1486834041
transform 1 0 32144 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2197_
timestamp 1486834041
transform 1 0 25760 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2198_
timestamp 1486834041
transform 1 0 25872 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2199_
timestamp 1486834041
transform 1 0 40208 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2200_
timestamp 1486834041
transform 1 0 41552 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2201_
timestamp 1486834041
transform 1 0 41440 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2202_
timestamp 1486834041
transform -1 0 46256 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2203_
timestamp 1486834041
transform 1 0 23632 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2204_
timestamp 1486834041
transform 1 0 25760 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2205_
timestamp 1486834041
transform 1 0 25648 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2206_
timestamp 1486834041
transform 1 0 23632 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2207_
timestamp 1486834041
transform -1 0 42000 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2208_
timestamp 1486834041
transform 1 0 40320 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2209_
timestamp 1486834041
transform 1 0 36176 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2210_
timestamp 1486834041
transform 1 0 36736 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2211_
timestamp 1486834041
transform 1 0 34496 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2212_
timestamp 1486834041
transform 1 0 34048 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2213_
timestamp 1486834041
transform 1 0 24528 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2214_
timestamp 1486834041
transform 1 0 24528 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2215_
timestamp 1486834041
transform -1 0 43232 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2216_
timestamp 1486834041
transform -1 0 45248 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2217_
timestamp 1486834041
transform 1 0 35840 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2218_
timestamp 1486834041
transform 1 0 36400 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2219_
timestamp 1486834041
transform 1 0 25872 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2220_
timestamp 1486834041
transform 1 0 28448 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2221_
timestamp 1486834041
transform -1 0 30576 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2222_
timestamp 1486834041
transform 1 0 28336 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2223_
timestamp 1486834041
transform -1 0 39200 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2224_
timestamp 1486834041
transform 1 0 37184 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2225_
timestamp 1486834041
transform 1 0 28336 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2226_
timestamp 1486834041
transform 1 0 25648 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2227_
timestamp 1486834041
transform 1 0 25872 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2228_
timestamp 1486834041
transform 1 0 24528 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2229_
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2230_
timestamp 1486834041
transform 1 0 17808 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2231_
timestamp 1486834041
transform 1 0 25088 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2232_
timestamp 1486834041
transform 1 0 21952 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2233_
timestamp 1486834041
transform 1 0 25872 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2234_
timestamp 1486834041
transform 1 0 27552 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2235_
timestamp 1486834041
transform 1 0 21504 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2236_
timestamp 1486834041
transform 1 0 23632 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2237_
timestamp 1486834041
transform 1 0 14112 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2238_
timestamp 1486834041
transform 1 0 15792 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2239_
timestamp 1486834041
transform 1 0 29344 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2240_
timestamp 1486834041
transform 1 0 27104 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2241_
timestamp 1486834041
transform -1 0 34496 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2242_
timestamp 1486834041
transform 1 0 29456 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2243_
timestamp 1486834041
transform 1 0 28336 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2244_
timestamp 1486834041
transform 1 0 24864 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2245_
timestamp 1486834041
transform 1 0 11872 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2246_
timestamp 1486834041
transform 1 0 10192 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2247_
timestamp 1486834041
transform 1 0 13552 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2248_
timestamp 1486834041
transform 1 0 14112 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2249_
timestamp 1486834041
transform 1 0 12432 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2250_
timestamp 1486834041
transform 1 0 13552 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2251_
timestamp 1486834041
transform 1 0 21392 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2252_
timestamp 1486834041
transform 1 0 21840 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2253_
timestamp 1486834041
transform 1 0 12992 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2254_
timestamp 1486834041
transform 1 0 11872 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2255_
timestamp 1486834041
transform 1 0 11872 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2256_
timestamp 1486834041
transform 1 0 12992 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2257_
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2258_
timestamp 1486834041
transform 1 0 6608 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2259_
timestamp 1486834041
transform 1 0 8400 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2260_
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2261_
timestamp 1486834041
transform 1 0 8624 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2262_
timestamp 1486834041
transform 1 0 8848 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2263_
timestamp 1486834041
transform 1 0 8512 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2264_
timestamp 1486834041
transform 1 0 10304 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2265_
timestamp 1486834041
transform 1 0 16576 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2266_
timestamp 1486834041
transform 1 0 18032 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2267_
timestamp 1486834041
transform 1 0 16576 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2268_
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2269_
timestamp 1486834041
transform 1 0 12992 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2270_
timestamp 1486834041
transform 1 0 12768 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2271_
timestamp 1486834041
transform 1 0 12992 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2272_
timestamp 1486834041
transform 1 0 14112 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2273_
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2274_
timestamp 1486834041
transform 1 0 1008 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2275_
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2276_
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2277_
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2278_
timestamp 1486834041
transform 1 0 1008 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2279_
timestamp 1486834041
transform 1 0 1120 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2280_
timestamp 1486834041
transform 1 0 1232 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2281_
timestamp 1486834041
transform 1 0 9744 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2282_
timestamp 1486834041
transform 1 0 6272 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2283_
timestamp 1486834041
transform 1 0 5264 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2284_
timestamp 1486834041
transform 1 0 9184 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2285_
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2286_
timestamp 1486834041
transform 1 0 896 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2287_
timestamp 1486834041
transform 1 0 896 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2288_
timestamp 1486834041
transform 1 0 896 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2289_
timestamp 1486834041
transform 1 0 8960 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2290_
timestamp 1486834041
transform 1 0 6272 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2291_
timestamp 1486834041
transform 1 0 9072 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2292_
timestamp 1486834041
transform -1 0 11872 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2293_
timestamp 1486834041
transform 1 0 22288 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2294_
timestamp 1486834041
transform 1 0 23520 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2295_
timestamp 1486834041
transform 1 0 23184 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2296_
timestamp 1486834041
transform 1 0 25760 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2297_
timestamp 1486834041
transform 1 0 18032 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2298_
timestamp 1486834041
transform 1 0 18368 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2299_
timestamp 1486834041
transform 1 0 19712 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2300_
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2301_
timestamp 1486834041
transform 1 0 16800 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2302_
timestamp 1486834041
transform 1 0 17024 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2303_
timestamp 1486834041
transform 1 0 18368 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2304_
timestamp 1486834041
transform -1 0 22736 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2305_
timestamp 1486834041
transform 1 0 6272 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2306_
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2307_
timestamp 1486834041
transform 1 0 7168 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2308_
timestamp 1486834041
transform 1 0 4928 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2309_
timestamp 1486834041
transform 1 0 6160 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2310_
timestamp 1486834041
transform 1 0 6608 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2311_
timestamp 1486834041
transform 1 0 6496 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2312_
timestamp 1486834041
transform 1 0 5936 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2313_
timestamp 1486834041
transform 1 0 10192 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2314_
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2315_
timestamp 1486834041
transform -1 0 19264 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2316_
timestamp 1486834041
transform 1 0 13664 0 1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2317_
timestamp 1486834041
transform 1 0 10976 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2318_
timestamp 1486834041
transform 1 0 8848 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2319_
timestamp 1486834041
transform 1 0 9968 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2320_
timestamp 1486834041
transform 1 0 9520 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2321_
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2322_
timestamp 1486834041
transform 1 0 2352 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2323_
timestamp 1486834041
transform -1 0 7616 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2324_
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2325_
timestamp 1486834041
transform 1 0 29904 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2326_
timestamp 1486834041
transform 1 0 29792 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2327_
timestamp 1486834041
transform 1 0 29792 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2328_
timestamp 1486834041
transform 1 0 32256 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2329_
timestamp 1486834041
transform 1 0 14112 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2330_
timestamp 1486834041
transform 1 0 17136 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2331_
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2332_
timestamp 1486834041
transform 1 0 17136 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2333_
timestamp 1486834041
transform 1 0 17248 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2334_
timestamp 1486834041
transform 1 0 17136 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2335_
timestamp 1486834041
transform 1 0 17360 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2336_
timestamp 1486834041
transform 1 0 17920 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2337_
timestamp 1486834041
transform 1 0 12768 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2338_
timestamp 1486834041
transform 1 0 12768 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2339_
timestamp 1486834041
transform 1 0 12992 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2340_
timestamp 1486834041
transform 1 0 12880 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2341_
timestamp 1486834041
transform 1 0 5712 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2342_
timestamp 1486834041
transform 1 0 6048 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2343_
timestamp 1486834041
transform 1 0 5824 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2344_
timestamp 1486834041
transform 1 0 7056 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2345_
timestamp 1486834041
transform 1 0 21504 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2346_
timestamp 1486834041
transform 1 0 21952 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2347_
timestamp 1486834041
transform -1 0 25088 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2348_
timestamp 1486834041
transform -1 0 26432 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2349_
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2350_
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2351_
timestamp 1486834041
transform 1 0 1008 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2352_
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2353_
timestamp 1486834041
transform 1 0 1232 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2354_
timestamp 1486834041
transform 1 0 1232 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2355_
timestamp 1486834041
transform -1 0 3248 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2356_
timestamp 1486834041
transform 1 0 1120 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2357_
timestamp 1486834041
transform 1 0 2800 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2358_
timestamp 1486834041
transform 1 0 4816 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2359_
timestamp 1486834041
transform -1 0 7616 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2360_
timestamp 1486834041
transform -1 0 7280 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2361_
timestamp 1486834041
transform 1 0 29680 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2362_
timestamp 1486834041
transform 1 0 29568 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2363_
timestamp 1486834041
transform 1 0 30576 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2364_
timestamp 1486834041
transform -1 0 35056 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2365_
timestamp 1486834041
transform 1 0 13776 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2366_
timestamp 1486834041
transform 1 0 13440 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2367_
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2368_
timestamp 1486834041
transform 1 0 14112 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2369_
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2370_
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2371_
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2372_
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2373_
timestamp 1486834041
transform 1 0 896 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2374_
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2375_
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2376_
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2377_
timestamp 1486834041
transform 1 0 3024 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2378_
timestamp 1486834041
transform 1 0 2352 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2379_
timestamp 1486834041
transform 1 0 3696 0 -1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2380_
timestamp 1486834041
transform 1 0 4032 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2381_
timestamp 1486834041
transform 1 0 6160 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2382_
timestamp 1486834041
transform 1 0 2352 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2383_
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2384_
timestamp 1486834041
transform 1 0 5040 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2385_
timestamp 1486834041
transform 1 0 17584 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2386_
timestamp 1486834041
transform 1 0 18032 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2387_
timestamp 1486834041
transform 1 0 30688 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2388_
timestamp 1486834041
transform -1 0 35168 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2389_
timestamp 1486834041
transform 1 0 32704 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2390_
timestamp 1486834041
transform 1 0 33712 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2391_
timestamp 1486834041
transform 1 0 39424 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2392_
timestamp 1486834041
transform -1 0 43680 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2393_
timestamp 1486834041
transform 1 0 40208 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2394_
timestamp 1486834041
transform 1 0 38416 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2395_
timestamp 1486834041
transform 1 0 29456 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2396_
timestamp 1486834041
transform 1 0 28672 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2397_
timestamp 1486834041
transform 1 0 13104 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2398_
timestamp 1486834041
transform 1 0 14112 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2399_
timestamp 1486834041
transform 1 0 39312 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2400_
timestamp 1486834041
transform 1 0 37632 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2401_
timestamp 1486834041
transform 1 0 37632 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2402_
timestamp 1486834041
transform 1 0 36400 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2403_
timestamp 1486834041
transform 1 0 32256 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2404_
timestamp 1486834041
transform 1 0 30800 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2405_
timestamp 1486834041
transform 1 0 14112 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2406_
timestamp 1486834041
transform 1 0 16688 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2407_
timestamp 1486834041
transform 1 0 28336 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2408_
timestamp 1486834041
transform 1 0 26432 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2409_
timestamp 1486834041
transform 1 0 33264 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2410_
timestamp 1486834041
transform -1 0 38416 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2411_
timestamp 1486834041
transform 1 0 32256 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2412_
timestamp 1486834041
transform 1 0 32256 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2413_
timestamp 1486834041
transform 1 0 25088 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2414_
timestamp 1486834041
transform 1 0 25536 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2415_
timestamp 1486834041
transform -1 0 30576 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2416_
timestamp 1486834041
transform 1 0 24864 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2417_
timestamp 1486834041
transform 1 0 37520 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2418_
timestamp 1486834041
transform 1 0 39312 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2419_
timestamp 1486834041
transform 1 0 40096 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2420_
timestamp 1486834041
transform 1 0 36736 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2421_
timestamp 1486834041
transform 1 0 38976 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _2422_
timestamp 1486834041
transform 1 0 40208 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2423_
timestamp 1486834041
transform -1 0 46256 0 -1 49392
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2424_
timestamp 1486834041
transform 1 0 47936 0 -1 18032
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2425_
timestamp 1486834041
transform 1 0 47936 0 -1 24304
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2426_
timestamp 1486834041
transform 1 0 45696 0 1 25872
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2427_
timestamp 1486834041
transform 1 0 45360 0 1 36848
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2428_
timestamp 1486834041
transform -1 0 49504 0 1 50960
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2429_
timestamp 1486834041
transform -1 0 50064 0 1 47824
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2430_
timestamp 1486834041
transform -1 0 46368 0 -1 52528
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2431_
timestamp 1486834041
transform -1 0 47712 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1486834041
transform -1 0 53872 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2433_
timestamp 1486834041
transform 1 0 47040 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2434_
timestamp 1486834041
transform -1 0 50288 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2435_
timestamp 1486834041
transform 1 0 53200 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2436_
timestamp 1486834041
transform 1 0 54880 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2437_
timestamp 1486834041
transform 1 0 46368 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2438_
timestamp 1486834041
transform 1 0 55552 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1486834041
transform 1 0 55776 0 -1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2440_
timestamp 1486834041
transform 1 0 55776 0 1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2441_
timestamp 1486834041
transform 1 0 52528 0 -1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2442_
timestamp 1486834041
transform 1 0 55776 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2443_
timestamp 1486834041
transform 1 0 55776 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2444_
timestamp 1486834041
transform 1 0 49616 0 -1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2445_
timestamp 1486834041
transform 1 0 55776 0 -1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2446_
timestamp 1486834041
transform 1 0 55776 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2447_
timestamp 1486834041
transform 1 0 27440 0 1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2448_
timestamp 1486834041
transform 1 0 29904 0 1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2449_
timestamp 1486834041
transform 1 0 55776 0 -1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2450_
timestamp 1486834041
transform 1 0 55776 0 1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2451_
timestamp 1486834041
transform -1 0 55776 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2452_
timestamp 1486834041
transform 1 0 47040 0 -1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2453_
timestamp 1486834041
transform -1 0 55552 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2454_
timestamp 1486834041
transform -1 0 54880 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2455_
timestamp 1486834041
transform -1 0 55552 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2456_
timestamp 1486834041
transform 1 0 1568 0 -1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2458_
timestamp 1486834041
transform 1 0 1568 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2459_
timestamp 1486834041
transform 1 0 2240 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2460_
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1486834041
transform -1 0 54880 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2462_
timestamp 1486834041
transform -1 0 40320 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2463_
timestamp 1486834041
transform 1 0 55552 0 1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2464_
timestamp 1486834041
transform 1 0 55776 0 -1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2465_
timestamp 1486834041
transform 1 0 54880 0 -1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2466_
timestamp 1486834041
transform 1 0 54768 0 -1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2467_
timestamp 1486834041
transform 1 0 55776 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2468_
timestamp 1486834041
transform -1 0 55888 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2469_
timestamp 1486834041
transform 1 0 55888 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2470_
timestamp 1486834041
transform 1 0 54656 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1486834041
transform -1 0 56448 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2472_
timestamp 1486834041
transform 1 0 54880 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2473_
timestamp 1486834041
transform 1 0 43120 0 1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2474_
timestamp 1486834041
transform -1 0 55440 0 1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2475_
timestamp 1486834041
transform 1 0 54880 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1486834041
transform 1 0 54432 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2477_
timestamp 1486834041
transform 1 0 54544 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2478_
timestamp 1486834041
transform 1 0 51856 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2479_
timestamp 1486834041
transform -1 0 54208 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2480_
timestamp 1486834041
transform -1 0 55216 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2481_
timestamp 1486834041
transform -1 0 53872 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2482_
timestamp 1486834041
transform -1 0 31472 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2483_
timestamp 1486834041
transform -1 0 56224 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2484_
timestamp 1486834041
transform 1 0 40544 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2485_
timestamp 1486834041
transform -1 0 54544 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2486_
timestamp 1486834041
transform -1 0 31360 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2487_
timestamp 1486834041
transform -1 0 41552 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2488_
timestamp 1486834041
transform -1 0 30464 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2489_
timestamp 1486834041
transform 1 0 31360 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1486834041
transform -1 0 54880 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2491_
timestamp 1486834041
transform -1 0 31360 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2492_
timestamp 1486834041
transform 1 0 36288 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2493_
timestamp 1486834041
transform 1 0 28448 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2494_
timestamp 1486834041
transform 1 0 27776 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2495_
timestamp 1486834041
transform 1 0 33600 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2496_
timestamp 1486834041
transform 1 0 51856 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2497_
timestamp 1486834041
transform -1 0 51408 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1486834041
transform -1 0 56448 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2499_
timestamp 1486834041
transform -1 0 49616 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2500_
timestamp 1486834041
transform -1 0 51744 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2501_
timestamp 1486834041
transform -1 0 51072 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2502_
timestamp 1486834041
transform -1 0 47712 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2503_
timestamp 1486834041
transform -1 0 47040 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2504_
timestamp 1486834041
transform -1 0 46592 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2505_
timestamp 1486834041
transform -1 0 45920 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2506_
timestamp 1486834041
transform -1 0 45696 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2507_
timestamp 1486834041
transform -1 0 45024 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2508_
timestamp 1486834041
transform -1 0 45248 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1486834041
transform -1 0 44352 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2510_
timestamp 1486834041
transform -1 0 45024 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2511_
timestamp 1486834041
transform 1 0 45696 0 1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2512_
timestamp 1486834041
transform 1 0 48608 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2513_
timestamp 1486834041
transform -1 0 51072 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2514_
timestamp 1486834041
transform -1 0 52416 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2515_
timestamp 1486834041
transform -1 0 54208 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2516_
timestamp 1486834041
transform -1 0 52528 0 1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2517_
timestamp 1486834041
transform -1 0 53760 0 1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2518_
timestamp 1486834041
transform 1 0 49952 0 1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2519_
timestamp 1486834041
transform -1 0 53760 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2520_
timestamp 1486834041
transform 1 0 32704 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2521_
timestamp 1486834041
transform -1 0 54320 0 1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2522_
timestamp 1486834041
transform -1 0 53984 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2523_
timestamp 1486834041
transform 1 0 31360 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2524_
timestamp 1486834041
transform 1 0 32256 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2525_
timestamp 1486834041
transform 1 0 31360 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2526_
timestamp 1486834041
transform -1 0 47264 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2527_
timestamp 1486834041
transform -1 0 52416 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2528_
timestamp 1486834041
transform 1 0 39200 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2529_
timestamp 1486834041
transform -1 0 56448 0 1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2530_
timestamp 1486834041
transform -1 0 56448 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2531_
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2532_
timestamp 1486834041
transform 1 0 9520 0 1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2533_
timestamp 1486834041
transform -1 0 23184 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2534_
timestamp 1486834041
transform 1 0 7616 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2535_
timestamp 1486834041
transform 1 0 4928 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2536_
timestamp 1486834041
transform -1 0 15456 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2537_
timestamp 1486834041
transform 1 0 3248 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2538_
timestamp 1486834041
transform 1 0 4256 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2539_
timestamp 1486834041
transform -1 0 3024 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2540_
timestamp 1486834041
transform -1 0 12432 0 1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2541_
timestamp 1486834041
transform 1 0 1008 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2542_
timestamp 1486834041
transform -1 0 22512 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2543_
timestamp 1486834041
transform -1 0 5488 0 1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2544_
timestamp 1486834041
transform 1 0 3136 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2545_
timestamp 1486834041
transform -1 0 20048 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2546_
timestamp 1486834041
transform -1 0 8064 0 -1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2547_
timestamp 1486834041
transform -1 0 19376 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2548_
timestamp 1486834041
transform -1 0 21728 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2549_
timestamp 1486834041
transform 1 0 1120 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2550_
timestamp 1486834041
transform -1 0 4592 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2551_
timestamp 1486834041
transform 1 0 6496 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2552_
timestamp 1486834041
transform -1 0 8176 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2553_
timestamp 1486834041
transform 1 0 8176 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2554_
timestamp 1486834041
transform 1 0 7840 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2555_
timestamp 1486834041
transform -1 0 9520 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2556_
timestamp 1486834041
transform 1 0 8960 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2557_
timestamp 1486834041
transform -1 0 10864 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2558_
timestamp 1486834041
transform -1 0 10304 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2559_
timestamp 1486834041
transform -1 0 11536 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2560_
timestamp 1486834041
transform -1 0 11648 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2561_
timestamp 1486834041
transform -1 0 12992 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2562_
timestamp 1486834041
transform -1 0 15680 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2563_
timestamp 1486834041
transform -1 0 7840 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2564_
timestamp 1486834041
transform -1 0 10192 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2565_
timestamp 1486834041
transform 1 0 10304 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2566_
timestamp 1486834041
transform -1 0 14336 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2567_
timestamp 1486834041
transform -1 0 15008 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2568_
timestamp 1486834041
transform 1 0 15008 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2569_
timestamp 1486834041
transform -1 0 16352 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2570_
timestamp 1486834041
transform -1 0 17696 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2571_
timestamp 1486834041
transform -1 0 19824 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2572_
timestamp 1486834041
transform -1 0 20272 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2573_
timestamp 1486834041
transform -1 0 20048 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2574_
timestamp 1486834041
transform 1 0 20048 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2575_
timestamp 1486834041
transform -1 0 21728 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2576_
timestamp 1486834041
transform -1 0 21392 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2577_
timestamp 1486834041
transform -1 0 22064 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2578_
timestamp 1486834041
transform -1 0 22960 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2579_
timestamp 1486834041
transform -1 0 23408 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2580_
timestamp 1486834041
transform -1 0 28784 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2581_
timestamp 1486834041
transform -1 0 22736 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2582_
timestamp 1486834041
transform -1 0 25872 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2583_
timestamp 1486834041
transform -1 0 24192 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2584_
timestamp 1486834041
transform -1 0 23184 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2585_
timestamp 1486834041
transform -1 0 25088 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2586_
timestamp 1486834041
transform -1 0 25536 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2587_
timestamp 1486834041
transform 1 0 2128 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2588_
timestamp 1486834041
transform -1 0 25760 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2589_
timestamp 1486834041
transform -1 0 25088 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2590_
timestamp 1486834041
transform -1 0 26656 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2591_
timestamp 1486834041
transform 1 0 25312 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2592_
timestamp 1486834041
transform 1 0 25088 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2593_
timestamp 1486834041
transform -1 0 28112 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2594_
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2595_
timestamp 1486834041
transform 1 0 29232 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2596_
timestamp 1486834041
transform 1 0 29904 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2597_
timestamp 1486834041
transform 1 0 28560 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2598_
timestamp 1486834041
transform 1 0 32256 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2599_
timestamp 1486834041
transform 1 0 28448 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2600_
timestamp 1486834041
transform 1 0 29120 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2601_
timestamp 1486834041
transform 1 0 34160 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2602_
timestamp 1486834041
transform -1 0 35504 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2603_
timestamp 1486834041
transform 1 0 33376 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2604_
timestamp 1486834041
transform 1 0 35168 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2605_
timestamp 1486834041
transform 1 0 35840 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2606_
timestamp 1486834041
transform 1 0 35280 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2607_
timestamp 1486834041
transform -1 0 36624 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2608_
timestamp 1486834041
transform 1 0 36624 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2609_
timestamp 1486834041
transform 1 0 37296 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2610_
timestamp 1486834041
transform 1 0 38416 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2611_
timestamp 1486834041
transform -1 0 38640 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2612_
timestamp 1486834041
transform 1 0 39088 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2613_
timestamp 1486834041
transform -1 0 39648 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2614_
timestamp 1486834041
transform 1 0 40096 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2615_
timestamp 1486834041
transform 1 0 37520 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2616_
timestamp 1486834041
transform 1 0 39088 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2617_
timestamp 1486834041
transform 1 0 38416 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2618_
timestamp 1486834041
transform 1 0 39088 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2619_
timestamp 1486834041
transform 1 0 42000 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2620_
timestamp 1486834041
transform 1 0 42784 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2621_
timestamp 1486834041
transform 1 0 42672 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2622_
timestamp 1486834041
transform 1 0 44128 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2623_
timestamp 1486834041
transform 1 0 44800 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2624_
timestamp 1486834041
transform -1 0 44688 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2625_
timestamp 1486834041
transform 1 0 44688 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1486834041
transform 1 0 46144 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2627_
timestamp 1486834041
transform 1 0 44688 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2628_
timestamp 1486834041
transform -1 0 46704 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2629_
timestamp 1486834041
transform 1 0 46704 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2630_
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2631_
timestamp 1486834041
transform 1 0 45360 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2632_
timestamp 1486834041
transform -1 0 49280 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2633_
timestamp 1486834041
transform 1 0 39536 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2634_
timestamp 1486834041
transform 1 0 46032 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2635_
timestamp 1486834041
transform 1 0 47936 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2636_
timestamp 1486834041
transform 1 0 8960 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2637_
timestamp 1486834041
transform -1 0 17248 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2638_
timestamp 1486834041
transform 1 0 11760 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2639_
timestamp 1486834041
transform 1 0 11088 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2640_
timestamp 1486834041
transform 1 0 9632 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2641_
timestamp 1486834041
transform 1 0 13216 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2642_
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2643_
timestamp 1486834041
transform 1 0 5488 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2644_
timestamp 1486834041
transform -1 0 13216 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2645_
timestamp 1486834041
transform 1 0 1568 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2646_
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2647_
timestamp 1486834041
transform 1 0 7952 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2648_
timestamp 1486834041
transform 1 0 7840 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2649_
timestamp 1486834041
transform -1 0 38080 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2650_
timestamp 1486834041
transform -1 0 10080 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2651_
timestamp 1486834041
transform -1 0 25088 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2652_
timestamp 1486834041
transform -1 0 17248 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2653_
timestamp 1486834041
transform -1 0 24192 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2654_
timestamp 1486834041
transform 1 0 7056 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2655_
timestamp 1486834041
transform -1 0 37072 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2656_
timestamp 1486834041
transform -1 0 56000 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2657_
timestamp 1486834041
transform -1 0 56448 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2658_
timestamp 1486834041
transform -1 0 55776 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2659_
timestamp 1486834041
transform -1 0 51632 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2660_
timestamp 1486834041
transform -1 0 56560 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2661_
timestamp 1486834041
transform -1 0 53088 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2662_
timestamp 1486834041
transform -1 0 48608 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2663_
timestamp 1486834041
transform -1 0 47264 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2664_
timestamp 1486834041
transform -1 0 47040 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2665_
timestamp 1486834041
transform -1 0 50960 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2666_
timestamp 1486834041
transform -1 0 2240 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2667_
timestamp 1486834041
transform -1 0 2240 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2668_
timestamp 1486834041
transform -1 0 51632 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2669_
timestamp 1486834041
transform -1 0 53312 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2670_
timestamp 1486834041
transform -1 0 56448 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2671_
timestamp 1486834041
transform -1 0 55776 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2672_
timestamp 1486834041
transform -1 0 52864 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2673_
timestamp 1486834041
transform -1 0 54656 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2674_
timestamp 1486834041
transform -1 0 49952 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2675_
timestamp 1486834041
transform -1 0 56448 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2676_
timestamp 1486834041
transform -1 0 56560 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2677_
timestamp 1486834041
transform -1 0 50064 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2678_
timestamp 1486834041
transform -1 0 55552 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2679_
timestamp 1486834041
transform -1 0 50960 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2680_
timestamp 1486834041
transform 1 0 1568 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2681_
timestamp 1486834041
transform 1 0 3360 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2682_
timestamp 1486834041
transform 1 0 7616 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2683_
timestamp 1486834041
transform 1 0 4816 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_1
timestamp 1486834041
transform 1 0 44688 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_2
timestamp 1486834041
transform 1 0 54208 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_3
timestamp 1486834041
transform -1 0 54768 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_4
timestamp 1486834041
transform 1 0 30576 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_5
timestamp 1486834041
transform -1 0 10416 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_6
timestamp 1486834041
transform -1 0 9856 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_7
timestamp 1486834041
transform -1 0 11088 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_8
timestamp 1486834041
transform -1 0 11200 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_9
timestamp 1486834041
transform -1 0 12544 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_10
timestamp 1486834041
transform -1 0 15232 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_11
timestamp 1486834041
transform -1 0 6720 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_12
timestamp 1486834041
transform -1 0 7728 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_13
timestamp 1486834041
transform -1 0 8400 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_14
timestamp 1486834041
transform -1 0 8064 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_15
timestamp 1486834041
transform -1 0 9072 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_16
timestamp 1486834041
transform -1 0 9184 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_17
timestamp 1486834041
transform -1 0 19600 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_18
timestamp 1486834041
transform -1 0 20272 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_19
timestamp 1486834041
transform -1 0 21280 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_20
timestamp 1486834041
transform -1 0 20944 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_21
timestamp 1486834041
transform -1 0 21616 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_22
timestamp 1486834041
transform -1 0 22512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_23
timestamp 1486834041
transform -1 0 14560 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_24
timestamp 1486834041
transform -1 0 15232 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_25
timestamp 1486834041
transform -1 0 15904 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_26
timestamp 1486834041
transform -1 0 17248 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_27
timestamp 1486834041
transform -1 0 19376 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_28
timestamp 1486834041
transform -1 0 19824 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_29
timestamp 1486834041
transform -1 0 44912 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_30
timestamp 1486834041
transform -1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_31
timestamp 1486834041
transform -1 0 44912 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_32
timestamp 1486834041
transform -1 0 46256 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_33
timestamp 1486834041
transform -1 0 46928 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_34
timestamp 1486834041
transform -1 0 48160 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_35
timestamp 1486834041
transform -1 0 42224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_36
timestamp 1486834041
transform -1 0 43008 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_37
timestamp 1486834041
transform -1 0 42896 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_38
timestamp 1486834041
transform -1 0 44352 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_39
timestamp 1486834041
transform 1 0 44800 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_40
timestamp 1486834041
transform -1 0 44240 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_41
timestamp 1486834041
transform -1 0 23520 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_42
timestamp 1486834041
transform -1 0 7056 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_43
timestamp 1486834041
transform -1 0 5488 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_44
timestamp 1486834041
transform -1 0 1792 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_45
timestamp 1486834041
transform 1 0 9408 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_46
timestamp 1486834041
transform 1 0 55776 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_47
timestamp 1486834041
transform -1 0 6944 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_48
timestamp 1486834041
transform 1 0 56224 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_49
timestamp 1486834041
transform -1 0 42560 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_50
timestamp 1486834041
transform 1 0 8064 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_51
timestamp 1486834041
transform 1 0 20048 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_52
timestamp 1486834041
transform -1 0 1456 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_53
timestamp 1486834041
transform 1 0 7616 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK
timestamp 1486834041
transform 1 0 46032 0 1 54096
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp 1486834041
transform -1 0 53536 0 -1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp 1486834041
transform 1 0 47936 0 -1 55664
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp 1486834041
transform -1 0 51632 0 1 27440
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp 1486834041
transform -1 0 53536 0 -1 43120
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp 1486834041
transform 1 0 47936 0 -1 36848
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_124
timestamp 1486834041
transform 1 0 14560 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134
timestamp 1486834041
transform 1 0 15680 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144
timestamp 1486834041
transform 1 0 16800 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168
timestamp 1486834041
transform 1 0 19488 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_242
timestamp 1486834041
transform 1 0 27776 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_267
timestamp 1486834041
transform 1 0 30576 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_271
timestamp 1486834041
transform 1 0 31024 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_338
timestamp 1486834041
transform 1 0 38528 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_384
timestamp 1486834041
transform 1 0 43680 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_390
timestamp 1486834041
transform 1 0 44352 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_392
timestamp 1486834041
transform 1 0 44576 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_401
timestamp 1486834041
transform 1 0 45584 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_405
timestamp 1486834041
transform 1 0 46032 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_450
timestamp 1486834041
transform 1 0 51072 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_466
timestamp 1486834041
transform 1 0 52864 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_474
timestamp 1486834041
transform 1 0 53760 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_494
timestamp 1486834041
transform 1 0 56000 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_498
timestamp 1486834041
transform 1 0 56448 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_4
timestamp 1486834041
transform 1 0 1120 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_59
timestamp 1486834041
transform 1 0 7280 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_63
timestamp 1486834041
transform 1 0 7728 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_135
timestamp 1486834041
transform 1 0 15792 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_148
timestamp 1486834041
transform 1 0 17248 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_188
timestamp 1486834041
transform 1 0 21728 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_244
timestamp 1486834041
transform 1 0 28000 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_303
timestamp 1486834041
transform 1 0 34608 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_349
timestamp 1486834041
transform 1 0 39760 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_366
timestamp 1486834041
transform 1 0 41664 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_368
timestamp 1486834041
transform 1 0 41888 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_371
timestamp 1486834041
transform 1 0 42224 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_375
timestamp 1486834041
transform 1 0 42672 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_418
timestamp 1486834041
transform 1 0 47488 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_440
timestamp 1486834041
transform 1 0 49952 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_472
timestamp 1486834041
transform 1 0 53536 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_488
timestamp 1486834041
transform 1 0 55328 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_22
timestamp 1486834041
transform 1 0 3136 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_41
timestamp 1486834041
transform 1 0 5264 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_64
timestamp 1486834041
transform 1 0 7840 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_91
timestamp 1486834041
transform 1 0 10864 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_113
timestamp 1486834041
transform 1 0 13328 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_140
timestamp 1486834041
transform 1 0 16352 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_165
timestamp 1486834041
transform 1 0 19152 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_234
timestamp 1486834041
transform 1 0 26880 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_238
timestamp 1486834041
transform 1 0 27328 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_341
timestamp 1486834041
transform 1 0 38864 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_435
timestamp 1486834041
transform 1 0 49392 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 51184 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_457
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_473
timestamp 1486834041
transform 1 0 53648 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_481
timestamp 1486834041
transform 1 0 54544 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_485
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_498
timestamp 1486834041
transform 1 0 56448 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_4
timestamp 1486834041
transform 1 0 1120 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_57
timestamp 1486834041
transform 1 0 7056 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_118
timestamp 1486834041
transform 1 0 13888 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_150
timestamp 1486834041
transform 1 0 17472 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_174
timestamp 1486834041
transform 1 0 20160 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_276
timestamp 1486834041
transform 1 0 31584 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_288
timestamp 1486834041
transform 1 0 32928 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_292
timestamp 1486834041
transform 1 0 33376 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_335
timestamp 1486834041
transform 1 0 38192 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_343
timestamp 1486834041
transform 1 0 39088 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_373
timestamp 1486834041
transform 1 0 42448 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_383
timestamp 1486834041
transform 1 0 43568 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_389
timestamp 1486834041
transform 1 0 44240 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_407
timestamp 1486834041
transform 1 0 46256 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1486834041
transform 1 0 47600 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_454
timestamp 1486834041
transform 1 0 51520 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_470
timestamp 1486834041
transform 1 0 53312 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_478
timestamp 1486834041
transform 1 0 54208 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_482
timestamp 1486834041
transform 1 0 54656 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_102
timestamp 1486834041
transform 1 0 12096 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_104
timestamp 1486834041
transform 1 0 12320 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_221
timestamp 1486834041
transform 1 0 25424 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_225
timestamp 1486834041
transform 1 0 25872 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_240
timestamp 1486834041
transform 1 0 27552 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_244
timestamp 1486834041
transform 1 0 28000 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_253
timestamp 1486834041
transform 1 0 29008 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_257
timestamp 1486834041
transform 1 0 29456 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_259
timestamp 1486834041
transform 1 0 29680 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_304
timestamp 1486834041
transform 1 0 34720 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_308
timestamp 1486834041
transform 1 0 35168 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_321
timestamp 1486834041
transform 1 0 36624 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_329
timestamp 1486834041
transform 1 0 37520 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_331
timestamp 1486834041
transform 1 0 37744 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_338
timestamp 1486834041
transform 1 0 38528 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_346
timestamp 1486834041
transform 1 0 39424 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1486834041
transform 1 0 44576 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_395
timestamp 1486834041
transform 1 0 44912 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_403
timestamp 1486834041
transform 1 0 45808 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_411
timestamp 1486834041
transform 1 0 46704 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_443
timestamp 1486834041
transform 1 0 50288 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_451
timestamp 1486834041
transform 1 0 51184 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_457
timestamp 1486834041
transform 1 0 51856 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_473
timestamp 1486834041
transform 1 0 53648 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_475
timestamp 1486834041
transform 1 0 53872 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_497
timestamp 1486834041
transform 1 0 56336 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_8
timestamp 1486834041
transform 1 0 1568 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_84
timestamp 1486834041
transform 1 0 10080 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_137
timestamp 1486834041
transform 1 0 16016 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_139
timestamp 1486834041
transform 1 0 16240 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_147
timestamp 1486834041
transform 1 0 17136 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_201
timestamp 1486834041
transform 1 0 23184 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_203
timestamp 1486834041
transform 1 0 23408 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_222
timestamp 1486834041
transform 1 0 25536 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_246
timestamp 1486834041
transform 1 0 28224 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_278
timestamp 1486834041
transform 1 0 31808 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_304
timestamp 1486834041
transform 1 0 34720 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_312
timestamp 1486834041
transform 1 0 35616 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_316
timestamp 1486834041
transform 1 0 36064 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_318
timestamp 1486834041
transform 1 0 36288 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_327
timestamp 1486834041
transform 1 0 37296 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_331
timestamp 1486834041
transform 1 0 37744 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_348
timestamp 1486834041
transform 1 0 39648 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_360
timestamp 1486834041
transform 1 0 40992 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_396
timestamp 1486834041
transform 1 0 45024 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_412
timestamp 1486834041
transform 1 0 46816 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_454
timestamp 1486834041
transform 1 0 51520 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_462
timestamp 1486834041
transform 1 0 52416 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_466
timestamp 1486834041
transform 1 0 52864 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_468
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_23
timestamp 1486834041
transform 1 0 3248 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_30
timestamp 1486834041
transform 1 0 4032 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_94
timestamp 1486834041
transform 1 0 11200 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_115
timestamp 1486834041
transform 1 0 13552 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_117
timestamp 1486834041
transform 1 0 13776 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_158
timestamp 1486834041
transform 1 0 18368 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_166
timestamp 1486834041
transform 1 0 19264 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_168
timestamp 1486834041
transform 1 0 19488 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_191
timestamp 1486834041
transform 1 0 22064 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_253
timestamp 1486834041
transform 1 0 29008 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_275
timestamp 1486834041
transform 1 0 31472 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_279
timestamp 1486834041
transform 1 0 31920 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_281
timestamp 1486834041
transform 1 0 32144 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_308
timestamp 1486834041
transform 1 0 35168 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_312
timestamp 1486834041
transform 1 0 35616 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 35840 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_327
timestamp 1486834041
transform 1 0 37296 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_334
timestamp 1486834041
transform 1 0 38080 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_344
timestamp 1486834041
transform 1 0 39200 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_402
timestamp 1486834041
transform 1 0 45696 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_434
timestamp 1486834041
transform 1 0 49280 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_450
timestamp 1486834041
transform 1 0 51072 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1486834041
transform 1 0 51520 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_487
timestamp 1486834041
transform 1 0 55216 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_494
timestamp 1486834041
transform 1 0 56000 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_498
timestamp 1486834041
transform 1 0 56448 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_200
timestamp 1486834041
transform 1 0 23072 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_218
timestamp 1486834041
transform 1 0 25088 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_220
timestamp 1486834041
transform 1 0 25312 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_259
timestamp 1486834041
transform 1 0 29680 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_321
timestamp 1486834041
transform 1 0 36624 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_329
timestamp 1486834041
transform 1 0 37520 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_414
timestamp 1486834041
transform 1 0 47040 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_418
timestamp 1486834041
transform 1 0 47488 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_438
timestamp 1486834041
transform 1 0 49728 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_459
timestamp 1486834041
transform 1 0 52080 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_463
timestamp 1486834041
transform 1 0 52528 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_4
timestamp 1486834041
transform 1 0 1120 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_129
timestamp 1486834041
transform 1 0 15120 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_133
timestamp 1486834041
transform 1 0 15568 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_167
timestamp 1486834041
transform 1 0 19376 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_209
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_255
timestamp 1486834041
transform 1 0 29232 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_259
timestamp 1486834041
transform 1 0 29680 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_281
timestamp 1486834041
transform 1 0 32144 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_325
timestamp 1486834041
transform 1 0 37072 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_329
timestamp 1486834041
transform 1 0 37520 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_363
timestamp 1486834041
transform 1 0 41328 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_384
timestamp 1486834041
transform 1 0 43680 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_447
timestamp 1486834041
transform 1 0 50736 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_497
timestamp 1486834041
transform 1 0 56336 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_2
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_4
timestamp 1486834041
transform 1 0 1120 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_37
timestamp 1486834041
transform 1 0 4816 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_199
timestamp 1486834041
transform 1 0 22960 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1486834041
transform 1 0 23856 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_220
timestamp 1486834041
transform 1 0 25312 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_254
timestamp 1486834041
transform 1 0 29120 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_258
timestamp 1486834041
transform 1 0 29568 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_314
timestamp 1486834041
transform 1 0 35840 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_318
timestamp 1486834041
transform 1 0 36288 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_339
timestamp 1486834041
transform 1 0 38640 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_347
timestamp 1486834041
transform 1 0 39536 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_349
timestamp 1486834041
transform 1 0 39760 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_391
timestamp 1486834041
transform 1 0 44464 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_412
timestamp 1486834041
transform 1 0 46816 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_430
timestamp 1486834041
transform 1 0 48832 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_474
timestamp 1486834041
transform 1 0 53760 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_14
timestamp 1486834041
transform 1 0 2240 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_73
timestamp 1486834041
transform 1 0 8848 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_128
timestamp 1486834041
transform 1 0 15008 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_161
timestamp 1486834041
transform 1 0 18704 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_169
timestamp 1486834041
transform 1 0 19600 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_173
timestamp 1486834041
transform 1 0 20048 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_197
timestamp 1486834041
transform 1 0 22736 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_201
timestamp 1486834041
transform 1 0 23184 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_203
timestamp 1486834041
transform 1 0 23408 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_224
timestamp 1486834041
transform 1 0 25760 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_240
timestamp 1486834041
transform 1 0 27552 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_244
timestamp 1486834041
transform 1 0 28000 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_402
timestamp 1486834041
transform 1 0 45696 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_404
timestamp 1486834041
transform 1 0 45920 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_437
timestamp 1486834041
transform 1 0 49616 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_439
timestamp 1486834041
transform 1 0 49840 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_457
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_459
timestamp 1486834041
transform 1 0 52080 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_492
timestamp 1486834041
transform 1 0 55776 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_130
timestamp 1486834041
transform 1 0 15232 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_178
timestamp 1486834041
transform 1 0 20608 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_186
timestamp 1486834041
transform 1 0 21504 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_228
timestamp 1486834041
transform 1 0 26208 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 31584 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_340
timestamp 1486834041
transform 1 0 38752 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_348
timestamp 1486834041
transform 1 0 39648 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_397
timestamp 1486834041
transform 1 0 45136 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_413
timestamp 1486834041
transform 1 0 46928 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_437
timestamp 1486834041
transform 1 0 49616 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_468
timestamp 1486834041
transform 1 0 53088 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_102
timestamp 1486834041
transform 1 0 12096 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1486834041
transform 1 0 12320 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_171
timestamp 1486834041
transform 1 0 19824 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_230
timestamp 1486834041
transform 1 0 26432 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_238
timestamp 1486834041
transform 1 0 27328 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_242
timestamp 1486834041
transform 1 0 27776 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_244
timestamp 1486834041
transform 1 0 28000 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_251
timestamp 1486834041
transform 1 0 28784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_253
timestamp 1486834041
transform 1 0 29008 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_306
timestamp 1486834041
transform 1 0 34944 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_310
timestamp 1486834041
transform 1 0 35392 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_327
timestamp 1486834041
transform 1 0 37296 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_331
timestamp 1486834041
transform 1 0 37744 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_352
timestamp 1486834041
transform 1 0 40096 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_360
timestamp 1486834041
transform 1 0 40992 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_382
timestamp 1486834041
transform 1 0 43456 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 43680 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_395
timestamp 1486834041
transform 1 0 44912 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_411
timestamp 1486834041
transform 1 0 46704 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1486834041
transform 1 0 47600 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_467
timestamp 1486834041
transform 1 0 52976 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_488
timestamp 1486834041
transform 1 0 55328 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_492
timestamp 1486834041
transform 1 0 55776 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_196
timestamp 1486834041
transform 1 0 22624 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_204
timestamp 1486834041
transform 1 0 23520 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_208
timestamp 1486834041
transform 1 0 23968 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_268
timestamp 1486834041
transform 1 0 30688 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_276
timestamp 1486834041
transform 1 0 31584 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_298
timestamp 1486834041
transform 1 0 34048 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_331
timestamp 1486834041
transform 1 0 37744 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_437
timestamp 1486834041
transform 1 0 49616 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_439
timestamp 1486834041
transform 1 0 49840 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_480
timestamp 1486834041
transform 1 0 54432 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_107
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_109
timestamp 1486834041
transform 1 0 12880 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_162
timestamp 1486834041
transform 1 0 18816 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_235
timestamp 1486834041
transform 1 0 26992 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_243
timestamp 1486834041
transform 1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_267
timestamp 1486834041
transform 1 0 30576 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_289
timestamp 1486834041
transform 1 0 33040 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_293
timestamp 1486834041
transform 1 0 33488 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_325
timestamp 1486834041
transform 1 0 37072 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_329
timestamp 1486834041
transform 1 0 37520 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_331
timestamp 1486834041
transform 1 0 37744 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_384
timestamp 1486834041
transform 1 0 43680 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_403
timestamp 1486834041
transform 1 0 45808 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_411
timestamp 1486834041
transform 1 0 46704 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_431
timestamp 1486834041
transform 1 0 48944 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_433
timestamp 1486834041
transform 1 0 49168 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_472
timestamp 1486834041
transform 1 0 53536 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_22
timestamp 1486834041
transform 1 0 3136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_204
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_208
timestamp 1486834041
transform 1 0 23968 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_232
timestamp 1486834041
transform 1 0 26656 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_254
timestamp 1486834041
transform 1 0 29120 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_270
timestamp 1486834041
transform 1 0 30912 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_278
timestamp 1486834041
transform 1 0 31808 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_302
timestamp 1486834041
transform 1 0 34496 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_344
timestamp 1486834041
transform 1 0 39200 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_348
timestamp 1486834041
transform 1 0 39648 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_434
timestamp 1486834041
transform 1 0 49280 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_498
timestamp 1486834041
transform 1 0 56448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_30
timestamp 1486834041
transform 1 0 4032 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1486834041
transform 1 0 4480 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_43
timestamp 1486834041
transform 1 0 5488 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_45
timestamp 1486834041
transform 1 0 5712 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_84
timestamp 1486834041
transform 1 0 10080 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_107
timestamp 1486834041
transform 1 0 12656 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_109
timestamp 1486834041
transform 1 0 12880 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_229
timestamp 1486834041
transform 1 0 26320 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_247
timestamp 1486834041
transform 1 0 28336 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_269
timestamp 1486834041
transform 1 0 30800 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_277
timestamp 1486834041
transform 1 0 31696 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_313
timestamp 1486834041
transform 1 0 35728 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_317
timestamp 1486834041
transform 1 0 36176 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_325
timestamp 1486834041
transform 1 0 37072 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_366
timestamp 1486834041
transform 1 0 41664 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_374
timestamp 1486834041
transform 1 0 42560 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_378
timestamp 1486834041
transform 1 0 43008 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_380
timestamp 1486834041
transform 1 0 43232 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_419
timestamp 1486834041
transform 1 0 47600 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_445
timestamp 1486834041
transform 1 0 50512 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_78
timestamp 1486834041
transform 1 0 9408 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_80
timestamp 1486834041
transform 1 0 9632 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_113
timestamp 1486834041
transform 1 0 13328 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_117
timestamp 1486834041
transform 1 0 13776 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_119
timestamp 1486834041
transform 1 0 14000 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_142
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_195
timestamp 1486834041
transform 1 0 22512 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_203
timestamp 1486834041
transform 1 0 23408 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_207
timestamp 1486834041
transform 1 0 23856 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_209
timestamp 1486834041
transform 1 0 24080 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_245
timestamp 1486834041
transform 1 0 28112 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_247
timestamp 1486834041
transform 1 0 28336 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_282
timestamp 1486834041
transform 1 0 32256 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_298
timestamp 1486834041
transform 1 0 34048 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_302
timestamp 1486834041
transform 1 0 34496 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_304
timestamp 1486834041
transform 1 0 34720 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_337
timestamp 1486834041
transform 1 0 38416 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_345
timestamp 1486834041
transform 1 0 39312 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_349
timestamp 1486834041
transform 1 0 39760 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_352
timestamp 1486834041
transform 1 0 40096 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_356
timestamp 1486834041
transform 1 0 40544 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_358
timestamp 1486834041
transform 1 0 40768 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_391
timestamp 1486834041
transform 1 0 44464 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_398
timestamp 1486834041
transform 1 0 45248 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1486834041
transform 1 0 47600 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_433
timestamp 1486834041
transform 1 0 49168 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_461
timestamp 1486834041
transform 1 0 52304 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_488
timestamp 1486834041
transform 1 0 55328 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_492
timestamp 1486834041
transform 1 0 55776 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1486834041
transform 1 0 4480 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_43
timestamp 1486834041
transform 1 0 5488 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_82
timestamp 1486834041
transform 1 0 9856 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_84
timestamp 1486834041
transform 1 0 10080 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_139
timestamp 1486834041
transform 1 0 16240 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_197
timestamp 1486834041
transform 1 0 22736 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_205
timestamp 1486834041
transform 1 0 23632 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_209
timestamp 1486834041
transform 1 0 24080 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_230
timestamp 1486834041
transform 1 0 26432 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_238
timestamp 1486834041
transform 1 0 27328 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_242
timestamp 1486834041
transform 1 0 27776 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_244
timestamp 1486834041
transform 1 0 28000 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_247
timestamp 1486834041
transform 1 0 28336 0 1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_263
timestamp 1486834041
transform 1 0 30128 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_271
timestamp 1486834041
transform 1 0 31024 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_275
timestamp 1486834041
transform 1 0 31472 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_277
timestamp 1486834041
transform 1 0 31696 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_310
timestamp 1486834041
transform 1 0 35392 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_314
timestamp 1486834041
transform 1 0 35840 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_317
timestamp 1486834041
transform 1 0 36176 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_325
timestamp 1486834041
transform 1 0 37072 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_327
timestamp 1486834041
transform 1 0 37296 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_387
timestamp 1486834041
transform 1 0 44016 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1486834041
transform 1 0 44240 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_410
timestamp 1486834041
transform 1 0 46592 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_421
timestamp 1486834041
transform 1 0 47824 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_477
timestamp 1486834041
transform 1 0 54096 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_498
timestamp 1486834041
transform 1 0 56448 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_68
timestamp 1486834041
transform 1 0 8288 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_142
timestamp 1486834041
transform 1 0 16576 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_150
timestamp 1486834041
transform 1 0 17472 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_152
timestamp 1486834041
transform 1 0 17696 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_205
timestamp 1486834041
transform 1 0 23632 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_209
timestamp 1486834041
transform 1 0 24080 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_228
timestamp 1486834041
transform 1 0 26208 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_250
timestamp 1486834041
transform 1 0 28672 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_258
timestamp 1486834041
transform 1 0 29568 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_302
timestamp 1486834041
transform 1 0 34496 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_344
timestamp 1486834041
transform 1 0 39200 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_348
timestamp 1486834041
transform 1 0 39648 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_352
timestamp 1486834041
transform 1 0 40096 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_422
timestamp 1486834041
transform 1 0 47936 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_489
timestamp 1486834041
transform 1 0 55440 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_492
timestamp 1486834041
transform 1 0 55776 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_2
timestamp 1486834041
transform 1 0 896 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_6
timestamp 1486834041
transform 1 0 1344 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_37
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_49
timestamp 1486834041
transform 1 0 6160 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_107
timestamp 1486834041
transform 1 0 12656 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_109
timestamp 1486834041
transform 1 0 12880 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_177
timestamp 1486834041
transform 1 0 20496 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_237
timestamp 1486834041
transform 1 0 27216 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_267
timestamp 1486834041
transform 1 0 30576 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_313
timestamp 1486834041
transform 1 0 35728 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_414
timestamp 1486834041
transform 1 0 47040 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_420
timestamp 1486834041
transform 1 0 47712 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_454
timestamp 1486834041
transform 1 0 51520 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_457
timestamp 1486834041
transform 1 0 51856 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_459
timestamp 1486834041
transform 1 0 52080 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_496
timestamp 1486834041
transform 1 0 56224 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_498
timestamp 1486834041
transform 1 0 56448 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1486834041
transform 1 0 896 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_67
timestamp 1486834041
transform 1 0 8176 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_69
timestamp 1486834041
transform 1 0 8400 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_97
timestamp 1486834041
transform 1 0 11536 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_99
timestamp 1486834041
transform 1 0 11760 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_152
timestamp 1486834041
transform 1 0 17696 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_185
timestamp 1486834041
transform 1 0 21392 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_201
timestamp 1486834041
transform 1 0 23184 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_209
timestamp 1486834041
transform 1 0 24080 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_232
timestamp 1486834041
transform 1 0 26656 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_240
timestamp 1486834041
transform 1 0 27552 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_242
timestamp 1486834041
transform 1 0 27776 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_310
timestamp 1486834041
transform 1 0 35392 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_314
timestamp 1486834041
transform 1 0 35840 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_316
timestamp 1486834041
transform 1 0 36064 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_349
timestamp 1486834041
transform 1 0 39760 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_389
timestamp 1486834041
transform 1 0 44240 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_418
timestamp 1486834041
transform 1 0 47488 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_492
timestamp 1486834041
transform 1 0 55776 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_14
timestamp 1486834041
transform 1 0 2240 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_37
timestamp 1486834041
transform 1 0 4816 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_70
timestamp 1486834041
transform 1 0 8512 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_72
timestamp 1486834041
transform 1 0 8736 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_159
timestamp 1486834041
transform 1 0 18480 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_217
timestamp 1486834041
transform 1 0 24976 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_313
timestamp 1486834041
transform 1 0 35728 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_349
timestamp 1486834041
transform 1 0 39760 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_383
timestamp 1486834041
transform 1 0 43568 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_407
timestamp 1486834041
transform 1 0 46256 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_409
timestamp 1486834041
transform 1 0 46480 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_454
timestamp 1486834041
transform 1 0 51520 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1486834041
transform 1 0 896 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_116
timestamp 1486834041
transform 1 0 13664 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_162
timestamp 1486834041
transform 1 0 18816 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_164
timestamp 1486834041
transform 1 0 19040 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_197
timestamp 1486834041
transform 1 0 22736 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_205
timestamp 1486834041
transform 1 0 23632 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_209
timestamp 1486834041
transform 1 0 24080 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_265
timestamp 1486834041
transform 1 0 30352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_342
timestamp 1486834041
transform 1 0 38976 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_352
timestamp 1486834041
transform 1 0 40096 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_383
timestamp 1486834041
transform 1 0 43568 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_387
timestamp 1486834041
transform 1 0 44016 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1486834041
transform 1 0 48608 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_492
timestamp 1486834041
transform 1 0 55776 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1486834041
transform 1 0 4480 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_104
timestamp 1486834041
transform 1 0 12320 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_107
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_161
timestamp 1486834041
transform 1 0 18704 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_169
timestamp 1486834041
transform 1 0 19600 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_173
timestamp 1486834041
transform 1 0 20048 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_177
timestamp 1486834041
transform 1 0 20496 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_231
timestamp 1486834041
transform 1 0 26544 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_239
timestamp 1486834041
transform 1 0 27440 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_243
timestamp 1486834041
transform 1 0 27888 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_267
timestamp 1486834041
transform 1 0 30576 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_308
timestamp 1486834041
transform 1 0 35168 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_312
timestamp 1486834041
transform 1 0 35616 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_314
timestamp 1486834041
transform 1 0 35840 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_317
timestamp 1486834041
transform 1 0 36176 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1486834041
transform 1 0 36624 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_381
timestamp 1486834041
transform 1 0 43344 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_387
timestamp 1486834041
transform 1 0 44016 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_433
timestamp 1486834041
transform 1 0 49168 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_498
timestamp 1486834041
transform 1 0 56448 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_54
timestamp 1486834041
transform 1 0 6720 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_142
timestamp 1486834041
transform 1 0 16576 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_279
timestamp 1486834041
transform 1 0 31920 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_334
timestamp 1486834041
transform 1 0 38080 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_338
timestamp 1486834041
transform 1 0 38528 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_380
timestamp 1486834041
transform 1 0 43232 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_401
timestamp 1486834041
transform 1 0 45584 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_405
timestamp 1486834041
transform 1 0 46032 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_407
timestamp 1486834041
transform 1 0 46256 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_422
timestamp 1486834041
transform 1 0 47936 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_426
timestamp 1486834041
transform 1 0 48384 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_455
timestamp 1486834041
transform 1 0 51632 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_468
timestamp 1486834041
transform 1 0 53088 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_492
timestamp 1486834041
transform 1 0 55776 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_14
timestamp 1486834041
transform 1 0 2240 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_43
timestamp 1486834041
transform 1 0 5488 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_51
timestamp 1486834041
transform 1 0 6384 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_154
timestamp 1486834041
transform 1 0 17920 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_197
timestamp 1486834041
transform 1 0 22736 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_238
timestamp 1486834041
transform 1 0 27328 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_242
timestamp 1486834041
transform 1 0 27776 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_244
timestamp 1486834041
transform 1 0 28000 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_279
timestamp 1486834041
transform 1 0 31920 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_281
timestamp 1486834041
transform 1 0 32144 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_306
timestamp 1486834041
transform 1 0 34944 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_314
timestamp 1486834041
transform 1 0 35840 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_349
timestamp 1486834041
transform 1 0 39760 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_380
timestamp 1486834041
transform 1 0 43232 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_384
timestamp 1486834041
transform 1 0 43680 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_387
timestamp 1486834041
transform 1 0 44016 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_395
timestamp 1486834041
transform 1 0 44912 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_449
timestamp 1486834041
transform 1 0 50960 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_457
timestamp 1486834041
transform 1 0 51856 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_459
timestamp 1486834041
transform 1 0 52080 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_498
timestamp 1486834041
transform 1 0 56448 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_69
timestamp 1486834041
transform 1 0 8400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_72
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_76
timestamp 1486834041
transform 1 0 9184 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_130
timestamp 1486834041
transform 1 0 15232 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_142
timestamp 1486834041
transform 1 0 16576 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_203
timestamp 1486834041
transform 1 0 23408 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_207
timestamp 1486834041
transform 1 0 23856 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_220
timestamp 1486834041
transform 1 0 25312 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_276
timestamp 1486834041
transform 1 0 31584 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_282
timestamp 1486834041
transform 1 0 32256 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_338
timestamp 1486834041
transform 1 0 38528 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_346
timestamp 1486834041
transform 1 0 39424 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_352
timestamp 1486834041
transform 1 0 40096 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_368
timestamp 1486834041
transform 1 0 41888 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_401
timestamp 1486834041
transform 1 0 45584 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_442
timestamp 1486834041
transform 1 0 50176 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_444
timestamp 1486834041
transform 1 0 50400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_498
timestamp 1486834041
transform 1 0 56448 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1486834041
transform 1 0 896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_33
timestamp 1486834041
transform 1 0 4368 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_57
timestamp 1486834041
transform 1 0 7056 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_59
timestamp 1486834041
transform 1 0 7280 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_92
timestamp 1486834041
transform 1 0 10976 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_100
timestamp 1486834041
transform 1 0 11872 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_104
timestamp 1486834041
transform 1 0 12320 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_127
timestamp 1486834041
transform 1 0 14896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_172
timestamp 1486834041
transform 1 0 19936 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_174
timestamp 1486834041
transform 1 0 20160 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_177
timestamp 1486834041
transform 1 0 20496 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_181
timestamp 1486834041
transform 1 0 20944 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_235
timestamp 1486834041
transform 1 0 26992 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_243
timestamp 1486834041
transform 1 0 27888 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_247
timestamp 1486834041
transform 1 0 28336 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_249
timestamp 1486834041
transform 1 0 28560 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_302
timestamp 1486834041
transform 1 0 34496 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_306
timestamp 1486834041
transform 1 0 34944 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_331
timestamp 1486834041
transform 1 0 37744 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_333
timestamp 1486834041
transform 1 0 37968 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_366
timestamp 1486834041
transform 1 0 41664 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_382
timestamp 1486834041
transform 1 0 43456 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_384
timestamp 1486834041
transform 1 0 43680 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_387
timestamp 1486834041
transform 1 0 44016 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_395
timestamp 1486834041
transform 1 0 44912 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_431
timestamp 1486834041
transform 1 0 48944 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_433
timestamp 1486834041
transform 1 0 49168 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_454
timestamp 1486834041
transform 1 0 51520 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_477
timestamp 1486834041
transform 1 0 54096 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_479
timestamp 1486834041
transform 1 0 54320 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_490
timestamp 1486834041
transform 1 0 55552 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_498
timestamp 1486834041
transform 1 0 56448 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_2
timestamp 1486834041
transform 1 0 896 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_87
timestamp 1486834041
transform 1 0 10416 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_91
timestamp 1486834041
transform 1 0 10864 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_112
timestamp 1486834041
transform 1 0 13216 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_116
timestamp 1486834041
transform 1 0 13664 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_118
timestamp 1486834041
transform 1 0 13888 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_139
timestamp 1486834041
transform 1 0 16240 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_174
timestamp 1486834041
transform 1 0 20160 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_220
timestamp 1486834041
transform 1 0 25312 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_253
timestamp 1486834041
transform 1 0 29008 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_277
timestamp 1486834041
transform 1 0 31696 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_279
timestamp 1486834041
transform 1 0 31920 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_302
timestamp 1486834041
transform 1 0 34496 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_412
timestamp 1486834041
transform 1 0 46816 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_486
timestamp 1486834041
transform 1 0 55104 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_498
timestamp 1486834041
transform 1 0 56448 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_86
timestamp 1486834041
transform 1 0 10304 0 1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_102
timestamp 1486834041
transform 1 0 12096 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_104
timestamp 1486834041
transform 1 0 12320 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_107
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_115
timestamp 1486834041
transform 1 0 13552 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_137
timestamp 1486834041
transform 1 0 16016 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_173
timestamp 1486834041
transform 1 0 20048 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_279
timestamp 1486834041
transform 1 0 31920 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_283
timestamp 1486834041
transform 1 0 32368 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_293
timestamp 1486834041
transform 1 0 33488 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_337
timestamp 1486834041
transform 1 0 38416 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_339
timestamp 1486834041
transform 1 0 38640 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_371
timestamp 1486834041
transform 1 0 42224 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_379
timestamp 1486834041
transform 1 0 43120 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_383
timestamp 1486834041
transform 1 0 43568 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_407
timestamp 1486834041
transform 1 0 46256 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_454
timestamp 1486834041
transform 1 0 51520 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_492
timestamp 1486834041
transform 1 0 55776 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1486834041
transform 1 0 896 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_23
timestamp 1486834041
transform 1 0 3248 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_27
timestamp 1486834041
transform 1 0 3696 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_37
timestamp 1486834041
transform 1 0 4816 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_69
timestamp 1486834041
transform 1 0 8400 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_72
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_125
timestamp 1486834041
transform 1 0 14672 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_133
timestamp 1486834041
transform 1 0 15568 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_137
timestamp 1486834041
transform 1 0 16016 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_139
timestamp 1486834041
transform 1 0 16240 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_174
timestamp 1486834041
transform 1 0 20160 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_176
timestamp 1486834041
transform 1 0 20384 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_221
timestamp 1486834041
transform 1 0 25424 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_223
timestamp 1486834041
transform 1 0 25648 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_244
timestamp 1486834041
transform 1 0 28000 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_268
timestamp 1486834041
transform 1 0 30688 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_272
timestamp 1486834041
transform 1 0 31136 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_274
timestamp 1486834041
transform 1 0 31360 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_282
timestamp 1486834041
transform 1 0 32256 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_352
timestamp 1486834041
transform 1 0 40096 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_418
timestamp 1486834041
transform 1 0 47488 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_462
timestamp 1486834041
transform 1 0 52416 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_489
timestamp 1486834041
transform 1 0 55440 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_498
timestamp 1486834041
transform 1 0 56448 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_57
timestamp 1486834041
transform 1 0 7056 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_89
timestamp 1486834041
transform 1 0 10640 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_116
timestamp 1486834041
transform 1 0 13664 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_132
timestamp 1486834041
transform 1 0 15456 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_140
timestamp 1486834041
transform 1 0 16352 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_142
timestamp 1486834041
transform 1 0 16576 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_177
timestamp 1486834041
transform 1 0 20496 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_219
timestamp 1486834041
transform 1 0 25200 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_223
timestamp 1486834041
transform 1 0 25648 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_247
timestamp 1486834041
transform 1 0 28336 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_327
timestamp 1486834041
transform 1 0 37296 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_349
timestamp 1486834041
transform 1 0 39760 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_351
timestamp 1486834041
transform 1 0 39984 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_384
timestamp 1486834041
transform 1 0 43680 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_387
timestamp 1486834041
transform 1 0 44016 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_395
timestamp 1486834041
transform 1 0 44912 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_431
timestamp 1486834041
transform 1 0 48944 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_467
timestamp 1486834041
transform 1 0 52976 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_469
timestamp 1486834041
transform 1 0 53200 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_490
timestamp 1486834041
transform 1 0 55552 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_498
timestamp 1486834041
transform 1 0 56448 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_22
timestamp 1486834041
transform 1 0 3136 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_60
timestamp 1486834041
transform 1 0 7392 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_92
timestamp 1486834041
transform 1 0 10976 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_96
timestamp 1486834041
transform 1 0 11424 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_98
timestamp 1486834041
transform 1 0 11648 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_142
timestamp 1486834041
transform 1 0 16576 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_228
timestamp 1486834041
transform 1 0 26208 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_262
timestamp 1486834041
transform 1 0 30016 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_270
timestamp 1486834041
transform 1 0 30912 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_352
timestamp 1486834041
transform 1 0 40096 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_413
timestamp 1486834041
transform 1 0 46928 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_488
timestamp 1486834041
transform 1 0 55328 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_498
timestamp 1486834041
transform 1 0 56448 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1486834041
transform 1 0 896 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_99
timestamp 1486834041
transform 1 0 11760 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_238
timestamp 1486834041
transform 1 0 27328 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_247
timestamp 1486834041
transform 1 0 28336 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_255
timestamp 1486834041
transform 1 0 29232 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_259
timestamp 1486834041
transform 1 0 29680 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_355
timestamp 1486834041
transform 1 0 40432 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_384
timestamp 1486834041
transform 1 0 43680 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_387
timestamp 1486834041
transform 1 0 44016 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1486834041
transform 1 0 44240 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_402
timestamp 1486834041
transform 1 0 45696 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_404
timestamp 1486834041
transform 1 0 45920 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_22
timestamp 1486834041
transform 1 0 3136 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_80
timestamp 1486834041
transform 1 0 9632 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_82
timestamp 1486834041
transform 1 0 9856 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_103
timestamp 1486834041
transform 1 0 12208 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_137
timestamp 1486834041
transform 1 0 16016 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_139
timestamp 1486834041
transform 1 0 16240 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_176
timestamp 1486834041
transform 1 0 20384 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_209
timestamp 1486834041
transform 1 0 24080 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_220
timestamp 1486834041
transform 1 0 25312 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_222
timestamp 1486834041
transform 1 0 25536 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_347
timestamp 1486834041
transform 1 0 39536 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_349
timestamp 1486834041
transform 1 0 39760 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_372
timestamp 1486834041
transform 1 0 42336 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_414
timestamp 1486834041
transform 1 0 47040 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_489
timestamp 1486834041
transform 1 0 55440 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_498
timestamp 1486834041
transform 1 0 56448 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1486834041
transform 1 0 4480 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_53
timestamp 1486834041
transform 1 0 6608 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_85
timestamp 1486834041
transform 1 0 10192 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_127
timestamp 1486834041
transform 1 0 14896 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_135
timestamp 1486834041
transform 1 0 15792 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_314
timestamp 1486834041
transform 1 0 35840 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_373
timestamp 1486834041
transform 1 0 42448 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_381
timestamp 1486834041
transform 1 0 43344 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_452
timestamp 1486834041
transform 1 0 51296 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_454
timestamp 1486834041
transform 1 0 51520 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_498
timestamp 1486834041
transform 1 0 56448 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_22
timestamp 1486834041
transform 1 0 3136 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_24
timestamp 1486834041
transform 1 0 3360 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_57
timestamp 1486834041
transform 1 0 7056 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_61
timestamp 1486834041
transform 1 0 7504 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_72
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_91
timestamp 1486834041
transform 1 0 10864 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_99
timestamp 1486834041
transform 1 0 11760 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_199
timestamp 1486834041
transform 1 0 22960 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_207
timestamp 1486834041
transform 1 0 23856 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_209
timestamp 1486834041
transform 1 0 24080 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_270
timestamp 1486834041
transform 1 0 30912 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_347
timestamp 1486834041
transform 1 0 39536 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_349
timestamp 1486834041
transform 1 0 39760 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_384
timestamp 1486834041
transform 1 0 43680 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_388
timestamp 1486834041
transform 1 0 44128 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1486834041
transform 1 0 47600 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_464
timestamp 1486834041
transform 1 0 52640 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_466
timestamp 1486834041
transform 1 0 52864 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_487
timestamp 1486834041
transform 1 0 55216 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_489
timestamp 1486834041
transform 1 0 55440 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_498
timestamp 1486834041
transform 1 0 56448 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_45
timestamp 1486834041
transform 1 0 5712 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_98
timestamp 1486834041
transform 1 0 11648 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_102
timestamp 1486834041
transform 1 0 12096 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_104
timestamp 1486834041
transform 1 0 12320 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_107
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_109
timestamp 1486834041
transform 1 0 12880 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_142
timestamp 1486834041
transform 1 0 16576 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_229
timestamp 1486834041
transform 1 0 26320 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_247
timestamp 1486834041
transform 1 0 28336 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_249
timestamp 1486834041
transform 1 0 28560 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_357
timestamp 1486834041
transform 1 0 40656 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_379
timestamp 1486834041
transform 1 0 43120 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_387
timestamp 1486834041
transform 1 0 44016 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_424
timestamp 1486834041
transform 1 0 48160 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_497
timestamp 1486834041
transform 1 0 56336 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_104
timestamp 1486834041
transform 1 0 12320 0 -1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_142
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_150
timestamp 1486834041
transform 1 0 17472 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_154
timestamp 1486834041
transform 1 0 17920 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_187
timestamp 1486834041
transform 1 0 21616 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_189
timestamp 1486834041
transform 1 0 21840 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_227
timestamp 1486834041
transform 1 0 26096 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_261
timestamp 1486834041
transform 1 0 29904 0 -1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_277
timestamp 1486834041
transform 1 0 31696 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_279
timestamp 1486834041
transform 1 0 31920 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_349
timestamp 1486834041
transform 1 0 39760 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_352
timestamp 1486834041
transform 1 0 40096 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_360
timestamp 1486834041
transform 1 0 40992 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1486834041
transform 1 0 47600 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_430
timestamp 1486834041
transform 1 0 48832 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_448
timestamp 1486834041
transform 1 0 50848 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_469
timestamp 1486834041
transform 1 0 53200 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_492
timestamp 1486834041
transform 1 0 55776 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_100
timestamp 1486834041
transform 1 0 11872 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_104
timestamp 1486834041
transform 1 0 12320 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_107
timestamp 1486834041
transform 1 0 12656 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_163
timestamp 1486834041
transform 1 0 18928 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_171
timestamp 1486834041
transform 1 0 19824 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_229
timestamp 1486834041
transform 1 0 26320 0 1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_247
timestamp 1486834041
transform 1 0 28336 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_249
timestamp 1486834041
transform 1 0 28560 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_311
timestamp 1486834041
transform 1 0 35504 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_347
timestamp 1486834041
transform 1 0 39536 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_351
timestamp 1486834041
transform 1 0 39984 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_479
timestamp 1486834041
transform 1 0 54320 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_496
timestamp 1486834041
transform 1 0 56224 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_498
timestamp 1486834041
transform 1 0 56448 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_104
timestamp 1486834041
transform 1 0 12320 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_162
timestamp 1486834041
transform 1 0 18816 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_166
timestamp 1486834041
transform 1 0 19264 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_199
timestamp 1486834041
transform 1 0 22960 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_207
timestamp 1486834041
transform 1 0 23856 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_209
timestamp 1486834041
transform 1 0 24080 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_228
timestamp 1486834041
transform 1 0 26208 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_262
timestamp 1486834041
transform 1 0 30016 0 -1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_278
timestamp 1486834041
transform 1 0 31808 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_302
timestamp 1486834041
transform 1 0 34496 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_306
timestamp 1486834041
transform 1 0 34944 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_327
timestamp 1486834041
transform 1 0 37296 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_329
timestamp 1486834041
transform 1 0 37520 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_372
timestamp 1486834041
transform 1 0 42336 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_380
timestamp 1486834041
transform 1 0 43232 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_422
timestamp 1486834041
transform 1 0 47936 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_467
timestamp 1486834041
transform 1 0 52976 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_488
timestamp 1486834041
transform 1 0 55328 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_492
timestamp 1486834041
transform 1 0 55776 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_107
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_115
timestamp 1486834041
transform 1 0 13552 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_117
timestamp 1486834041
transform 1 0 13776 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_150
timestamp 1486834041
transform 1 0 17472 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1486834041
transform 1 0 20160 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_182
timestamp 1486834041
transform 1 0 21056 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_190
timestamp 1486834041
transform 1 0 21952 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1486834041
transform 1 0 28000 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_247
timestamp 1486834041
transform 1 0 28336 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_255
timestamp 1486834041
transform 1 0 29232 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_311
timestamp 1486834041
transform 1 0 35504 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_317
timestamp 1486834041
transform 1 0 36176 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1486834041
transform 1 0 36624 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_330
timestamp 1486834041
transform 1 0 37632 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1486834041
transform 1 0 43680 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_387
timestamp 1486834041
transform 1 0 44016 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_452
timestamp 1486834041
transform 1 0 51296 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1486834041
transform 1 0 51520 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_495
timestamp 1486834041
transform 1 0 56112 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_68
timestamp 1486834041
transform 1 0 8288 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_72
timestamp 1486834041
transform 1 0 8736 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_80
timestamp 1486834041
transform 1 0 9632 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_134
timestamp 1486834041
transform 1 0 15680 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_138
timestamp 1486834041
transform 1 0 16128 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_176
timestamp 1486834041
transform 1 0 20384 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_212
timestamp 1486834041
transform 1 0 24416 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_268
timestamp 1486834041
transform 1 0 30688 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_276
timestamp 1486834041
transform 1 0 31584 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_334
timestamp 1486834041
transform 1 0 38080 0 -1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_472
timestamp 1486834041
transform 1 0 53536 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_498
timestamp 1486834041
transform 1 0 56448 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1486834041
transform 1 0 896 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_69
timestamp 1486834041
transform 1 0 8400 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_107
timestamp 1486834041
transform 1 0 12656 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_135
timestamp 1486834041
transform 1 0 15792 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_301
timestamp 1486834041
transform 1 0 34384 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_309
timestamp 1486834041
transform 1 0 35280 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_313
timestamp 1486834041
transform 1 0 35728 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_337
timestamp 1486834041
transform 1 0 38416 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_339
timestamp 1486834041
transform 1 0 38640 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_372
timestamp 1486834041
transform 1 0 42336 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_498
timestamp 1486834041
transform 1 0 56448 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_115
timestamp 1486834041
transform 1 0 13552 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_119
timestamp 1486834041
transform 1 0 14000 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_194
timestamp 1486834041
transform 1 0 22400 0 -1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_244
timestamp 1486834041
transform 1 0 28000 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_252
timestamp 1486834041
transform 1 0 28896 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_256
timestamp 1486834041
transform 1 0 29344 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_277
timestamp 1486834041
transform 1 0 31696 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_279
timestamp 1486834041
transform 1 0 31920 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_282
timestamp 1486834041
transform 1 0 32256 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1486834041
transform 1 0 32704 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_339
timestamp 1486834041
transform 1 0 38640 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_347
timestamp 1486834041
transform 1 0 39536 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_349
timestamp 1486834041
transform 1 0 39760 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_352
timestamp 1486834041
transform 1 0 40096 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_498
timestamp 1486834041
transform 1 0 56448 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_103
timestamp 1486834041
transform 1 0 12208 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_115
timestamp 1486834041
transform 1 0 13552 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_119
timestamp 1486834041
transform 1 0 14000 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_121
timestamp 1486834041
transform 1 0 14224 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_154
timestamp 1486834041
transform 1 0 17920 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_185
timestamp 1486834041
transform 1 0 21392 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_241
timestamp 1486834041
transform 1 0 27664 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_279
timestamp 1486834041
transform 1 0 31920 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_317
timestamp 1486834041
transform 1 0 36176 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_371
timestamp 1486834041
transform 1 0 42224 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_373
timestamp 1486834041
transform 1 0 42448 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_395
timestamp 1486834041
transform 1 0 44912 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_428
timestamp 1486834041
transform 1 0 48608 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_457
timestamp 1486834041
transform 1 0 51856 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_22
timestamp 1486834041
transform 1 0 3136 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_24
timestamp 1486834041
transform 1 0 3360 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_142
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_158
timestamp 1486834041
transform 1 0 18368 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_160
timestamp 1486834041
transform 1 0 18592 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_193
timestamp 1486834041
transform 1 0 22288 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_220
timestamp 1486834041
transform 1 0 25312 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_222
timestamp 1486834041
transform 1 0 25536 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_243
timestamp 1486834041
transform 1 0 27888 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_277
timestamp 1486834041
transform 1 0 31696 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_279
timestamp 1486834041
transform 1 0 31920 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_282
timestamp 1486834041
transform 1 0 32256 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_336
timestamp 1486834041
transform 1 0 38304 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_344
timestamp 1486834041
transform 1 0 39200 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_348
timestamp 1486834041
transform 1 0 39648 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_406
timestamp 1486834041
transform 1 0 46144 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_408
timestamp 1486834041
transform 1 0 46368 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_447
timestamp 1486834041
transform 1 0 50736 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_449
timestamp 1486834041
transform 1 0 50960 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_492
timestamp 1486834041
transform 1 0 55776 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_43
timestamp 1486834041
transform 1 0 5488 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_45
timestamp 1486834041
transform 1 0 5712 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_102
timestamp 1486834041
transform 1 0 12096 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_104
timestamp 1486834041
transform 1 0 12320 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_112
timestamp 1486834041
transform 1 0 13216 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_120
timestamp 1486834041
transform 1 0 14112 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_153
timestamp 1486834041
transform 1 0 17808 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_221
timestamp 1486834041
transform 1 0 25424 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1486834041
transform 1 0 28336 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_268
timestamp 1486834041
transform 1 0 30688 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_270
timestamp 1486834041
transform 1 0 30912 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_442
timestamp 1486834041
transform 1 0 50176 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_454
timestamp 1486834041
transform 1 0 51520 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_497
timestamp 1486834041
transform 1 0 56336 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_104
timestamp 1486834041
transform 1 0 12320 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_106
timestamp 1486834041
transform 1 0 12544 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_127
timestamp 1486834041
transform 1 0 14896 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_135
timestamp 1486834041
transform 1 0 15792 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_142
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_150
timestamp 1486834041
transform 1 0 17472 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_154
timestamp 1486834041
transform 1 0 17920 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_208
timestamp 1486834041
transform 1 0 23968 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_228
timestamp 1486834041
transform 1 0 26208 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_276
timestamp 1486834041
transform 1 0 31584 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_322
timestamp 1486834041
transform 1 0 36736 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_324
timestamp 1486834041
transform 1 0 36960 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_404
timestamp 1486834041
transform 1 0 45920 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_413
timestamp 1486834041
transform 1 0 46928 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_487
timestamp 1486834041
transform 1 0 55216 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_489
timestamp 1486834041
transform 1 0 55440 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_498
timestamp 1486834041
transform 1 0 56448 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_46
timestamp 1486834041
transform 1 0 5824 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_113
timestamp 1486834041
transform 1 0 13328 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_146
timestamp 1486834041
transform 1 0 17024 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_154
timestamp 1486834041
transform 1 0 17920 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_177
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_185
timestamp 1486834041
transform 1 0 21392 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_221
timestamp 1486834041
transform 1 0 25424 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_247
timestamp 1486834041
transform 1 0 28336 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_301
timestamp 1486834041
transform 1 0 34384 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_322
timestamp 1486834041
transform 1 0 36736 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_454
timestamp 1486834041
transform 1 0 51520 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_497
timestamp 1486834041
transform 1 0 56336 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_22
timestamp 1486834041
transform 1 0 3136 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_68
timestamp 1486834041
transform 1 0 8288 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_116
timestamp 1486834041
transform 1 0 13664 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_209
timestamp 1486834041
transform 1 0 24080 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_220
timestamp 1486834041
transform 1 0 25312 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_274
timestamp 1486834041
transform 1 0 31360 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_278
timestamp 1486834041
transform 1 0 31808 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_282
timestamp 1486834041
transform 1 0 32256 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_284
timestamp 1486834041
transform 1 0 32480 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_403
timestamp 1486834041
transform 1 0 45808 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_498
timestamp 1486834041
transform 1 0 56448 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_72
timestamp 1486834041
transform 1 0 8736 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_177
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_185
timestamp 1486834041
transform 1 0 21392 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_238
timestamp 1486834041
transform 1 0 27328 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_242
timestamp 1486834041
transform 1 0 27776 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_244
timestamp 1486834041
transform 1 0 28000 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_247
timestamp 1486834041
transform 1 0 28336 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_263
timestamp 1486834041
transform 1 0 30128 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_265
timestamp 1486834041
transform 1 0 30352 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_298
timestamp 1486834041
transform 1 0 34048 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_340
timestamp 1486834041
transform 1 0 38752 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_361
timestamp 1486834041
transform 1 0 41104 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_447
timestamp 1486834041
transform 1 0 50736 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_457
timestamp 1486834041
transform 1 0 51856 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_83
timestamp 1486834041
transform 1 0 9968 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_146
timestamp 1486834041
transform 1 0 17024 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_148
timestamp 1486834041
transform 1 0 17248 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_201
timestamp 1486834041
transform 1 0 23184 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_209
timestamp 1486834041
transform 1 0 24080 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_228
timestamp 1486834041
transform 1 0 26208 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_261
timestamp 1486834041
transform 1 0 29904 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_352
timestamp 1486834041
transform 1 0 40096 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1486834041
transform 1 0 40320 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1486834041
transform 1 0 47600 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_489
timestamp 1486834041
transform 1 0 55440 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_492
timestamp 1486834041
transform 1 0 55776 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_2
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_4
timestamp 1486834041
transform 1 0 1120 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1486834041
transform 1 0 4480 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_109
timestamp 1486834041
transform 1 0 12880 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_130
timestamp 1486834041
transform 1 0 15232 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_177
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_185
timestamp 1486834041
transform 1 0 21392 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_241
timestamp 1486834041
transform 1 0 27664 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_317
timestamp 1486834041
transform 1 0 36176 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_374
timestamp 1486834041
transform 1 0 42560 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_454
timestamp 1486834041
transform 1 0 51520 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_474
timestamp 1486834041
transform 1 0 53760 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_2
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_24
timestamp 1486834041
transform 1 0 3360 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_147
timestamp 1486834041
transform 1 0 17136 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_149
timestamp 1486834041
transform 1 0 17360 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_347
timestamp 1486834041
transform 1 0 39536 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_349
timestamp 1486834041
transform 1 0 39760 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_352
timestamp 1486834041
transform 1 0 40096 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1486834041
transform 1 0 40320 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_399
timestamp 1486834041
transform 1 0 45360 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_422
timestamp 1486834041
transform 1 0 47936 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_492
timestamp 1486834041
transform 1 0 55776 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_2
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_115
timestamp 1486834041
transform 1 0 13552 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_117
timestamp 1486834041
transform 1 0 13776 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_170
timestamp 1486834041
transform 1 0 19712 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_174
timestamp 1486834041
transform 1 0 20160 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_185
timestamp 1486834041
transform 1 0 21392 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_241
timestamp 1486834041
transform 1 0 27664 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_307
timestamp 1486834041
transform 1 0 35056 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_314
timestamp 1486834041
transform 1 0 35840 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_317
timestamp 1486834041
transform 1 0 36176 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_319
timestamp 1486834041
transform 1 0 36400 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_346
timestamp 1486834041
transform 1 0 39424 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_383
timestamp 1486834041
transform 1 0 43568 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_52
timestamp 1486834041
transform 1 0 6496 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_54
timestamp 1486834041
transform 1 0 6720 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_137
timestamp 1486834041
transform 1 0 16016 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_139
timestamp 1486834041
transform 1 0 16240 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_162
timestamp 1486834041
transform 1 0 18816 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_398
timestamp 1486834041
transform 1 0 45248 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_422
timestamp 1486834041
transform 1 0 47936 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_488
timestamp 1486834041
transform 1 0 55328 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_498
timestamp 1486834041
transform 1 0 56448 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_37
timestamp 1486834041
transform 1 0 4816 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_78
timestamp 1486834041
transform 1 0 9408 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_80
timestamp 1486834041
transform 1 0 9632 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_107
timestamp 1486834041
transform 1 0 12656 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_182
timestamp 1486834041
transform 1 0 21056 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_184
timestamp 1486834041
transform 1 0 21280 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_247
timestamp 1486834041
transform 1 0 28336 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_251
timestamp 1486834041
transform 1 0 28784 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_282
timestamp 1486834041
transform 1 0 32256 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_352
timestamp 1486834041
transform 1 0 40096 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_384
timestamp 1486834041
transform 1 0 43680 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_432
timestamp 1486834041
transform 1 0 49056 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_434
timestamp 1486834041
transform 1 0 49280 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_457
timestamp 1486834041
transform 1 0 51856 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_459
timestamp 1486834041
transform 1 0 52080 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_492
timestamp 1486834041
transform 1 0 55776 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_22
timestamp 1486834041
transform 1 0 3136 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_61
timestamp 1486834041
transform 1 0 7504 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_106
timestamp 1486834041
transform 1 0 12544 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_142
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_227
timestamp 1486834041
transform 1 0 26096 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_263
timestamp 1486834041
transform 1 0 30128 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_282
timestamp 1486834041
transform 1 0 32256 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_284
timestamp 1486834041
transform 1 0 32480 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_341
timestamp 1486834041
transform 1 0 38864 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_376
timestamp 1486834041
transform 1 0 42784 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_397
timestamp 1486834041
transform 1 0 45136 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_399
timestamp 1486834041
transform 1 0 45360 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_488
timestamp 1486834041
transform 1 0 55328 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_492
timestamp 1486834041
transform 1 0 55776 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_2
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_182
timestamp 1486834041
transform 1 0 21056 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_184
timestamp 1486834041
transform 1 0 21280 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_247
timestamp 1486834041
transform 1 0 28336 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_255
timestamp 1486834041
transform 1 0 29232 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_259
timestamp 1486834041
transform 1 0 29680 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_301
timestamp 1486834041
transform 1 0 34384 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_303
timestamp 1486834041
transform 1 0 34608 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_314
timestamp 1486834041
transform 1 0 35840 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_328
timestamp 1486834041
transform 1 0 37408 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1486834041
transform 1 0 896 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_47
timestamp 1486834041
transform 1 0 5936 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_49
timestamp 1486834041
transform 1 0 6160 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_108
timestamp 1486834041
transform 1 0 12768 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_130
timestamp 1486834041
transform 1 0 15232 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_263
timestamp 1486834041
transform 1 0 30128 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_342
timestamp 1486834041
transform 1 0 38976 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_417
timestamp 1486834041
transform 1 0 47376 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_419
timestamp 1486834041
transform 1 0 47600 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_433
timestamp 1486834041
transform 1 0 49168 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_481
timestamp 1486834041
transform 1 0 54544 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_483
timestamp 1486834041
transform 1 0 54768 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_492
timestamp 1486834041
transform 1 0 55776 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_71
timestamp 1486834041
transform 1 0 8624 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_199
timestamp 1486834041
transform 1 0 22960 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_201
timestamp 1486834041
transform 1 0 23184 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_234
timestamp 1486834041
transform 1 0 26880 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_242
timestamp 1486834041
transform 1 0 27776 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_244
timestamp 1486834041
transform 1 0 28000 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_247
timestamp 1486834041
transform 1 0 28336 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_255
timestamp 1486834041
transform 1 0 29232 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_314
timestamp 1486834041
transform 1 0 35840 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_361
timestamp 1486834041
transform 1 0 41104 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_363
timestamp 1486834041
transform 1 0 41328 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_384
timestamp 1486834041
transform 1 0 43680 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_439
timestamp 1486834041
transform 1 0 49840 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_446
timestamp 1486834041
transform 1 0 50624 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_463
timestamp 1486834041
transform 1 0 52528 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_485
timestamp 1486834041
transform 1 0 54992 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_498
timestamp 1486834041
transform 1 0 56448 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_22
timestamp 1486834041
transform 1 0 3136 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_92
timestamp 1486834041
transform 1 0 10976 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_142
timestamp 1486834041
transform 1 0 16576 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_144
timestamp 1486834041
transform 1 0 16800 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_177
timestamp 1486834041
transform 1 0 20496 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_244
timestamp 1486834041
transform 1 0 28000 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_302
timestamp 1486834041
transform 1 0 34496 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_372
timestamp 1486834041
transform 1 0 42336 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_422
timestamp 1486834041
transform 1 0 47936 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_424
timestamp 1486834041
transform 1 0 48160 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_440
timestamp 1486834041
transform 1 0 49952 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_461
timestamp 1486834041
transform 1 0 52304 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_463
timestamp 1486834041
transform 1 0 52528 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_476
timestamp 1486834041
transform 1 0 53984 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_483
timestamp 1486834041
transform 1 0 54768 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_492
timestamp 1486834041
transform 1 0 55776 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_37
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_39
timestamp 1486834041
transform 1 0 5040 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_206
timestamp 1486834041
transform 1 0 23744 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1486834041
transform 1 0 28336 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_285
timestamp 1486834041
transform 1 0 32592 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_314
timestamp 1486834041
transform 1 0 35840 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_323
timestamp 1486834041
transform 1 0 36848 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_347
timestamp 1486834041
transform 1 0 39536 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_405
timestamp 1486834041
transform 1 0 46032 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_475
timestamp 1486834041
transform 1 0 53872 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_477
timestamp 1486834041
transform 1 0 54096 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_492
timestamp 1486834041
transform 1 0 55776 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_22
timestamp 1486834041
transform 1 0 3136 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_188
timestamp 1486834041
transform 1 0 21728 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_214
timestamp 1486834041
transform 1 0 24640 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_247
timestamp 1486834041
transform 1 0 28336 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_249
timestamp 1486834041
transform 1 0 28560 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_327
timestamp 1486834041
transform 1 0 37296 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_329
timestamp 1486834041
transform 1 0 37520 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_372
timestamp 1486834041
transform 1 0 42336 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_422
timestamp 1486834041
transform 1 0 47936 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_431
timestamp 1486834041
transform 1 0 48944 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_470
timestamp 1486834041
transform 1 0 53312 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_492
timestamp 1486834041
transform 1 0 55776 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_22
timestamp 1486834041
transform 1 0 3136 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_39
timestamp 1486834041
transform 1 0 5040 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_130
timestamp 1486834041
transform 1 0 15232 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_132
timestamp 1486834041
transform 1 0 15456 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_167
timestamp 1486834041
transform 1 0 19376 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_195
timestamp 1486834041
transform 1 0 22512 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_197
timestamp 1486834041
transform 1 0 22736 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_242
timestamp 1486834041
transform 1 0 27776 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_244
timestamp 1486834041
transform 1 0 28000 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_267
timestamp 1486834041
transform 1 0 30576 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_313
timestamp 1486834041
transform 1 0 35728 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_317
timestamp 1486834041
transform 1 0 36176 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_356
timestamp 1486834041
transform 1 0 40544 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_358
timestamp 1486834041
transform 1 0 40768 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_401
timestamp 1486834041
transform 1 0 45584 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_423
timestamp 1486834041
transform 1 0 48048 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_431
timestamp 1486834041
transform 1 0 48944 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_438
timestamp 1486834041
transform 1 0 49728 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_440
timestamp 1486834041
transform 1 0 49952 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_453
timestamp 1486834041
transform 1 0 51408 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_475
timestamp 1486834041
transform 1 0 53872 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_477
timestamp 1486834041
transform 1 0 54096 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_490
timestamp 1486834041
transform 1 0 55552 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_492
timestamp 1486834041
transform 1 0 55776 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_2
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1486834041
transform 1 0 8400 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_75
timestamp 1486834041
transform 1 0 9072 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_87
timestamp 1486834041
transform 1 0 10416 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_93
timestamp 1486834041
transform 1 0 11088 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_127
timestamp 1486834041
transform 1 0 14896 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_162
timestamp 1486834041
transform 1 0 18816 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_164
timestamp 1486834041
transform 1 0 19040 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_184
timestamp 1486834041
transform 1 0 21280 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_186
timestamp 1486834041
transform 1 0 21504 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_207
timestamp 1486834041
transform 1 0 23856 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1486834041
transform 1 0 24080 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_237
timestamp 1486834041
transform 1 0 27216 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_239
timestamp 1486834041
transform 1 0 27440 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_266
timestamp 1486834041
transform 1 0 30464 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_327
timestamp 1486834041
transform 1 0 37296 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_348
timestamp 1486834041
transform 1 0 39648 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_352
timestamp 1486834041
transform 1 0 40096 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1486834041
transform 1 0 40320 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_370
timestamp 1486834041
transform 1 0 42112 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_428
timestamp 1486834041
transform 1 0 48608 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_430
timestamp 1486834041
transform 1 0 48832 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_437
timestamp 1486834041
transform 1 0 49616 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_480
timestamp 1486834041
transform 1 0 54432 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_492
timestamp 1486834041
transform 1 0 55776 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_2
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_54
timestamp 1486834041
transform 1 0 6720 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_79
timestamp 1486834041
transform 1 0 9520 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_82
timestamp 1486834041
transform 1 0 9856 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_84
timestamp 1486834041
transform 1 0 10080 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_124
timestamp 1486834041
transform 1 0 14560 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_130
timestamp 1486834041
transform 1 0 15232 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_142
timestamp 1486834041
transform 1 0 16576 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_166
timestamp 1486834041
transform 1 0 19264 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_177
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_181
timestamp 1486834041
transform 1 0 20944 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_230
timestamp 1486834041
transform 1 0 26432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_232
timestamp 1486834041
transform 1 0 26656 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_267
timestamp 1486834041
transform 1 0 30576 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_300
timestamp 1486834041
transform 1 0 34272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_312
timestamp 1486834041
transform 1 0 35616 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_314
timestamp 1486834041
transform 1 0 35840 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_352
timestamp 1486834041
transform 1 0 40096 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_404
timestamp 1486834041
transform 1 0 45920 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_481
timestamp 1486834041
transform 1 0 54544 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_483
timestamp 1486834041
transform 1 0 54768 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_490
timestamp 1486834041
transform 1 0 55552 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_492
timestamp 1486834041
transform 1 0 55776 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_118
timestamp 1486834041
transform 1 0 13888 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_148
timestamp 1486834041
transform 1 0 17248 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_218
timestamp 1486834041
transform 1 0 25088 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_225
timestamp 1486834041
transform 1 0 25872 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_320
timestamp 1486834041
transform 1 0 36512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_349
timestamp 1486834041
transform 1 0 39760 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_358
timestamp 1486834041
transform 1 0 40768 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_402
timestamp 1486834041
transform 1 0 45696 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_416
timestamp 1486834041
transform 1 0 47264 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_478
timestamp 1486834041
transform 1 0 54208 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_480
timestamp 1486834041
transform 1 0 54432 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_487
timestamp 1486834041
transform 1 0 55216 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_489
timestamp 1486834041
transform 1 0 55440 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_498
timestamp 1486834041
transform 1 0 56448 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_2
timestamp 1486834041
transform 1 0 896 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_70
timestamp 1486834041
transform 1 0 8512 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_76
timestamp 1486834041
transform 1 0 9184 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_94
timestamp 1486834041
transform 1 0 11200 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_106
timestamp 1486834041
transform 1 0 12544 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_138
timestamp 1486834041
transform 1 0 16128 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_172
timestamp 1486834041
transform 1 0 19936 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_181
timestamp 1486834041
transform 1 0 20944 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_206
timestamp 1486834041
transform 1 0 23744 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_208
timestamp 1486834041
transform 1 0 23968 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_240
timestamp 1486834041
transform 1 0 27552 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_274
timestamp 1486834041
transform 1 0 31360 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_308
timestamp 1486834041
transform 1 0 35168 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_339
timestamp 1486834041
transform 1 0 38640 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_348
timestamp 1486834041
transform 1 0 39648 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_376
timestamp 1486834041
transform 1 0 42784 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_440
timestamp 1486834041
transform 1 0 49952 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_474
timestamp 1486834041
transform 1 0 53760 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_498
timestamp 1486834041
transform 1 0 56448 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output1
timestamp 1486834041
transform -1 0 24752 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output2
timestamp 1486834041
transform 1 0 46368 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output3
timestamp 1486834041
transform 1 0 48720 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output4
timestamp 1486834041
transform 1 0 55888 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output5
timestamp 1486834041
transform 1 0 48496 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output6
timestamp 1486834041
transform 1 0 55888 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output7
timestamp 1486834041
transform 1 0 55888 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output8
timestamp 1486834041
transform 1 0 55888 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output9
timestamp 1486834041
transform 1 0 55888 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output10
timestamp 1486834041
transform 1 0 55888 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output11
timestamp 1486834041
transform 1 0 55888 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output12
timestamp 1486834041
transform 1 0 55888 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output13
timestamp 1486834041
transform 1 0 55776 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output14
timestamp 1486834041
transform 1 0 55888 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output15
timestamp 1486834041
transform 1 0 55888 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output16
timestamp 1486834041
transform 1 0 55888 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output17
timestamp 1486834041
transform 1 0 55888 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output18
timestamp 1486834041
transform 1 0 55888 0 1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output19
timestamp 1486834041
transform 1 0 55888 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output20
timestamp 1486834041
transform 1 0 55888 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output21
timestamp 1486834041
transform 1 0 55888 0 -1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output22
timestamp 1486834041
transform 1 0 43120 0 1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output23
timestamp 1486834041
transform 1 0 30688 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output24
timestamp 1486834041
transform 1 0 27552 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output25
timestamp 1486834041
transform 1 0 55888 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output26
timestamp 1486834041
transform 1 0 53872 0 1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output27
timestamp 1486834041
transform 1 0 41216 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output28
timestamp 1486834041
transform 1 0 36512 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output29
timestamp 1486834041
transform 1 0 54880 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output30
timestamp 1486834041
transform 1 0 44016 0 1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output31
timestamp 1486834041
transform 1 0 48944 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output32
timestamp 1486834041
transform 1 0 47040 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output33
timestamp 1486834041
transform 1 0 31360 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output34
timestamp 1486834041
transform 1 0 55888 0 -1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output35
timestamp 1486834041
transform 1 0 55888 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output36
timestamp 1486834041
transform 1 0 53872 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output37
timestamp 1486834041
transform 1 0 54880 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output38
timestamp 1486834041
transform 1 0 55888 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output39
timestamp 1486834041
transform 1 0 55888 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output40
timestamp 1486834041
transform 1 0 54880 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output41
timestamp 1486834041
transform 1 0 55888 0 -1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output42
timestamp 1486834041
transform 1 0 55888 0 1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output43
timestamp 1486834041
transform 1 0 55888 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output44
timestamp 1486834041
transform 1 0 55888 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output45
timestamp 1486834041
transform 1 0 51856 0 1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output46
timestamp 1486834041
transform 1 0 55888 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output47
timestamp 1486834041
transform 1 0 55104 0 1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output48
timestamp 1486834041
transform 1 0 50960 0 1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output49
timestamp 1486834041
transform 1 0 55888 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output50
timestamp 1486834041
transform 1 0 26768 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output51
timestamp 1486834041
transform 1 0 53760 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output52
timestamp 1486834041
transform 1 0 36288 0 1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output53
timestamp 1486834041
transform 1 0 29344 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output54
timestamp 1486834041
transform 1 0 49728 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output55
timestamp 1486834041
transform 1 0 29120 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output56
timestamp 1486834041
transform 1 0 49056 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output57
timestamp 1486834041
transform 1 0 52416 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output58
timestamp 1486834041
transform 1 0 53200 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output59
timestamp 1486834041
transform 1 0 48272 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output60
timestamp 1486834041
transform 1 0 47040 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output61
timestamp 1486834041
transform 1 0 30016 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output62
timestamp 1486834041
transform 1 0 47936 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output63
timestamp 1486834041
transform 1 0 46368 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output64
timestamp 1486834041
transform 1 0 45696 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output65
timestamp 1486834041
transform 1 0 45024 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output66
timestamp 1486834041
transform 1 0 43008 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output67
timestamp 1486834041
transform 1 0 42336 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output68
timestamp 1486834041
transform 1 0 41664 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output69
timestamp 1486834041
transform 1 0 41216 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output70
timestamp 1486834041
transform 1 0 40992 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output71
timestamp 1486834041
transform 1 0 41664 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output72
timestamp 1486834041
transform 1 0 52640 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output73
timestamp 1486834041
transform 1 0 39872 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output74
timestamp 1486834041
transform 1 0 40992 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output75
timestamp 1486834041
transform 1 0 27440 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output76
timestamp 1486834041
transform 1 0 26768 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output77
timestamp 1486834041
transform 1 0 53200 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output78
timestamp 1486834041
transform 1 0 50064 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output79
timestamp 1486834041
transform 1 0 25984 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output80
timestamp 1486834041
transform 1 0 27440 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output81
timestamp 1486834041
transform 1 0 26656 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output82
timestamp 1486834041
transform -1 0 53088 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output83
timestamp 1486834041
transform 1 0 47264 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output84
timestamp 1486834041
transform 1 0 46592 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output85
timestamp 1486834041
transform 1 0 45024 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output86
timestamp 1486834041
transform 1 0 45696 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output87
timestamp 1486834041
transform 1 0 43680 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output88
timestamp 1486834041
transform 1 0 43008 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output89
timestamp 1486834041
transform 1 0 41888 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output90
timestamp 1486834041
transform 1 0 40544 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output91
timestamp 1486834041
transform 1 0 40320 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output92
timestamp 1486834041
transform 1 0 42448 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output93
timestamp 1486834041
transform -1 0 53760 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output94
timestamp 1486834041
transform 1 0 34272 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output95
timestamp 1486834041
transform 1 0 32928 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output96
timestamp 1486834041
transform 1 0 26096 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output97
timestamp 1486834041
transform 1 0 31584 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output98
timestamp 1486834041
transform 1 0 30464 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output99
timestamp 1486834041
transform -1 0 53200 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output100
timestamp 1486834041
transform -1 0 52528 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output101
timestamp 1486834041
transform 1 0 49280 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output102
timestamp 1486834041
transform -1 0 23632 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output103
timestamp 1486834041
transform -1 0 22288 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output104
timestamp 1486834041
transform -1 0 21840 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 24080 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output106
timestamp 1486834041
transform -1 0 21168 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output107
timestamp 1486834041
transform -1 0 7056 0 -1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output108
timestamp 1486834041
transform -1 0 5488 0 1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output109
timestamp 1486834041
transform -1 0 7616 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output110
timestamp 1486834041
transform 1 0 1008 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output111
timestamp 1486834041
transform 1 0 1680 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output112
timestamp 1486834041
transform 1 0 3360 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output113
timestamp 1486834041
transform 1 0 1680 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output114
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output115
timestamp 1486834041
transform -1 0 13328 0 1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output116
timestamp 1486834041
transform -1 0 9408 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output117
timestamp 1486834041
transform 1 0 3248 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output118
timestamp 1486834041
transform -1 0 13664 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output119
timestamp 1486834041
transform -1 0 12992 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output120
timestamp 1486834041
transform 1 0 7392 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output121
timestamp 1486834041
transform 1 0 1008 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output122
timestamp 1486834041
transform 1 0 6720 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output123
timestamp 1486834041
transform 1 0 5152 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output124
timestamp 1486834041
transform 1 0 5824 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output125
timestamp 1486834041
transform 1 0 6496 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output126
timestamp 1486834041
transform 1 0 7168 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output127
timestamp 1486834041
transform 1 0 15680 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output128
timestamp 1486834041
transform 1 0 11648 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output129
timestamp 1486834041
transform 1 0 1680 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output130
timestamp 1486834041
transform -1 0 23856 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output131
timestamp 1486834041
transform -1 0 25088 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output132
timestamp 1486834041
transform 1 0 2464 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output133
timestamp 1486834041
transform -1 0 25424 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output134
timestamp 1486834041
transform 1 0 1792 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output135
timestamp 1486834041
transform 1 0 6832 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output136
timestamp 1486834041
transform 1 0 3136 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output137
timestamp 1486834041
transform 1 0 3808 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output138
timestamp 1486834041
transform 1 0 9632 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output139
timestamp 1486834041
transform 1 0 20384 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output140
timestamp 1486834041
transform 1 0 18704 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output141
timestamp 1486834041
transform 1 0 18368 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output142
timestamp 1486834041
transform 1 0 19040 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output143
timestamp 1486834041
transform 1 0 22176 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output144
timestamp 1486834041
transform 1 0 22848 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output145
timestamp 1486834041
transform 1 0 15904 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output146
timestamp 1486834041
transform 1 0 10304 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output147
timestamp 1486834041
transform 1 0 11424 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output148
timestamp 1486834041
transform 1 0 12992 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output149
timestamp 1486834041
transform 1 0 16352 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output150
timestamp 1486834041
transform 1 0 17360 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output151
timestamp 1486834041
transform -1 0 20944 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output152
timestamp 1486834041
transform 1 0 18032 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output153
timestamp 1486834041
transform 1 0 17696 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output154
timestamp 1486834041
transform 1 0 21840 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output155
timestamp 1486834041
transform 1 0 20160 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output156
timestamp 1486834041
transform 1 0 20832 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output157
timestamp 1486834041
transform 1 0 21504 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output158
timestamp 1486834041
transform 1 0 22176 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output159
timestamp 1486834041
transform 1 0 22848 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output160
timestamp 1486834041
transform 1 0 23968 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output161
timestamp 1486834041
transform 1 0 24640 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output162
timestamp 1486834041
transform -1 0 29008 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output163
timestamp 1486834041
transform 1 0 25984 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output164
timestamp 1486834041
transform 1 0 26656 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output165
timestamp 1486834041
transform 1 0 27888 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output166
timestamp 1486834041
transform -1 0 30464 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output167
timestamp 1486834041
transform -1 0 34272 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output168
timestamp 1486834041
transform -1 0 34944 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output169
timestamp 1486834041
transform -1 0 34608 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output170
timestamp 1486834041
transform -1 0 35840 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output171
timestamp 1486834041
transform -1 0 36512 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output172
timestamp 1486834041
transform -1 0 37184 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output173
timestamp 1486834041
transform -1 0 34720 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output174
timestamp 1486834041
transform -1 0 37856 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output175
timestamp 1486834041
transform -1 0 38864 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output176
timestamp 1486834041
transform -1 0 40992 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output177
timestamp 1486834041
transform -1 0 41664 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output178
timestamp 1486834041
transform -1 0 43680 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output179
timestamp 1486834041
transform 1 0 39200 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output180
timestamp 1486834041
transform -1 0 45584 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output181
timestamp 1486834041
transform -1 0 36848 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output182
timestamp 1486834041
transform -1 0 38528 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output183
timestamp 1486834041
transform -1 0 37744 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output184
timestamp 1486834041
transform -1 0 35952 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output185
timestamp 1486834041
transform -1 0 37520 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output186
timestamp 1486834041
transform -1 0 38416 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output187
timestamp 1486834041
transform -1 0 39648 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output188
timestamp 1486834041
transform -1 0 37744 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output189
timestamp 1486834041
transform -1 0 40320 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output190
timestamp 1486834041
transform -1 0 46144 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output191
timestamp 1486834041
transform -1 0 48720 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output192
timestamp 1486834041
transform -1 0 49392 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output193
timestamp 1486834041
transform -1 0 48048 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output194
timestamp 1486834041
transform -1 0 47600 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output195
timestamp 1486834041
transform -1 0 51072 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output196
timestamp 1486834041
transform -1 0 49952 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output197
timestamp 1486834041
transform -1 0 47264 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output198
timestamp 1486834041
transform -1 0 44128 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output199
timestamp 1486834041
transform -1 0 47936 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output200
timestamp 1486834041
transform -1 0 48832 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output201
timestamp 1486834041
transform -1 0 43568 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output202
timestamp 1486834041
transform -1 0 47488 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output203
timestamp 1486834041
transform -1 0 49504 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output204
timestamp 1486834041
transform -1 0 50176 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output205
timestamp 1486834041
transform -1 0 46032 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output206
timestamp 1486834041
transform -1 0 51744 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output207
timestamp 1486834041
transform -1 0 15792 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output208
timestamp 1486834041
transform -1 0 15680 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output209
timestamp 1486834041
transform -1 0 15120 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output210
timestamp 1486834041
transform -1 0 12096 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output211
timestamp 1486834041
transform -1 0 16800 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output212
timestamp 1486834041
transform -1 0 14448 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output213
timestamp 1486834041
transform -1 0 8288 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output214
timestamp 1486834041
transform -1 0 13328 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output215
timestamp 1486834041
transform -1 0 7840 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output216
timestamp 1486834041
transform -1 0 8512 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output217
timestamp 1486834041
transform -1 0 11424 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output218
timestamp 1486834041
transform -1 0 13328 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output219
timestamp 1486834041
transform -1 0 12096 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output220
timestamp 1486834041
transform -1 0 11424 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output221
timestamp 1486834041
transform -1 0 4592 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output222
timestamp 1486834041
transform -1 0 3920 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output223
timestamp 1486834041
transform -1 0 6832 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output224
timestamp 1486834041
transform -1 0 9408 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output225
timestamp 1486834041
transform -1 0 8400 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output226
timestamp 1486834041
transform -1 0 16352 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output227
timestamp 1486834041
transform -1 0 1568 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output228
timestamp 1486834041
transform -1 0 1568 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output229
timestamp 1486834041
transform -1 0 1568 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output230
timestamp 1486834041
transform -1 0 3920 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output231
timestamp 1486834041
transform -1 0 7616 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output232
timestamp 1486834041
transform -1 0 6160 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output233
timestamp 1486834041
transform -1 0 1568 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output234
timestamp 1486834041
transform -1 0 2240 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output235
timestamp 1486834041
transform -1 0 1568 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output236
timestamp 1486834041
transform -1 0 5488 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output237
timestamp 1486834041
transform -1 0 4480 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output238
timestamp 1486834041
transform -1 0 3808 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output239
timestamp 1486834041
transform -1 0 2128 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output240
timestamp 1486834041
transform -1 0 14000 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output241
timestamp 1486834041
transform -1 0 10080 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output242
timestamp 1486834041
transform -1 0 4144 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output243
timestamp 1486834041
transform -1 0 8512 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output244
timestamp 1486834041
transform -1 0 9408 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output245
timestamp 1486834041
transform -1 0 9856 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output246
timestamp 1486834041
transform -1 0 2576 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output247
timestamp 1486834041
transform -1 0 8848 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output248
timestamp 1486834041
transform -1 0 9408 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output249
timestamp 1486834041
transform -1 0 1904 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output250
timestamp 1486834041
transform -1 0 4592 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output251
timestamp 1486834041
transform -1 0 3920 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output252
timestamp 1486834041
transform -1 0 4032 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output253
timestamp 1486834041
transform -1 0 4144 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output254
timestamp 1486834041
transform -1 0 4816 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_71
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_72
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_73
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_74
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_75
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_76
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_77
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_78
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_79
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_80
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_81
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_82
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_83
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_84
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_85
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_86
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_87
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 56784 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_88
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 56784 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_89
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 56784 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_90
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 56784 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_91
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 56784 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_92
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 56784 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_93
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 56784 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_94
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 56784 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_95
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 56784 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_96
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 56784 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_97
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 56784 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_98
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 56784 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_99
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 56784 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_100
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 56784 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_101
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 56784 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_102
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 56784 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_103
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 56784 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_104
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 56784 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_105
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 56784 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_106
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 56784 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_107
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 56784 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_108
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 56784 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_109
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 56784 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_110
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 56784 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_111
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 56784 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_112
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 56784 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_113
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 56784 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_114
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 56784 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_115
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 56784 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_116
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 56784 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_117
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 56784 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_118
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 56784 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_119
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 56784 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_120
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 56784 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_121
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 56784 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_122
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 56784 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_123
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 56784 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_124
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 56784 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_125
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 56784 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_126
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 56784 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_127
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 56784 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_128
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 56784 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_129
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 56784 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_130
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 56784 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_131
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 56784 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_132
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 56784 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_133
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 56784 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_134
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 56784 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_135
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 56784 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_136
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 56784 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_137
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 56784 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_138
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 56784 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_139
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 56784 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_140
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 56784 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_141
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 56784 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_157
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_158
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_159
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_160
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_161
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_162
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_164
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_165
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_166
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_167
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_168
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_169
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_171
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_172
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_173
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_174
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_175
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_176
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_178
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_179
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_180
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_181
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_182
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_183
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_185
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_186
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_187
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_188
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_189
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_190
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_192
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_193
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_194
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_195
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_196
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_197
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_199
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_200
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_201
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_202
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_203
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_204
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_206
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_207
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_208
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_209
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_210
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_211
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_213
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_214
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_215
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_216
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_217
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_218
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_220
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_221
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_222
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_223
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_224
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_225
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_227
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_228
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_229
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_230
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_231
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_232
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_234
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_235
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_236
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_237
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_238
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_239
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_241
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_242
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_243
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_244
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_245
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_246
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_248
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_249
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_250
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_251
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_252
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_253
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_255
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_256
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_257
timestamp 1486834041
transform 1 0 32032 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_258
timestamp 1486834041
transform 1 0 39872 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_259
timestamp 1486834041
transform 1 0 47712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_260
timestamp 1486834041
transform 1 0 55552 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_262
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_263
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_264
timestamp 1486834041
transform 1 0 28112 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_265
timestamp 1486834041
transform 1 0 35952 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_266
timestamp 1486834041
transform 1 0 43792 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_267
timestamp 1486834041
transform 1 0 51632 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_269
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_270
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_271
timestamp 1486834041
transform 1 0 32032 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_272
timestamp 1486834041
transform 1 0 39872 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_273
timestamp 1486834041
transform 1 0 47712 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_274
timestamp 1486834041
transform 1 0 55552 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_276
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_277
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_278
timestamp 1486834041
transform 1 0 28112 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_279
timestamp 1486834041
transform 1 0 35952 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_280
timestamp 1486834041
transform 1 0 43792 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_281
timestamp 1486834041
transform 1 0 51632 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_283
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_284
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_285
timestamp 1486834041
transform 1 0 32032 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_286
timestamp 1486834041
transform 1 0 39872 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_287
timestamp 1486834041
transform 1 0 47712 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_288
timestamp 1486834041
transform 1 0 55552 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_290
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_291
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_292
timestamp 1486834041
transform 1 0 28112 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_293
timestamp 1486834041
transform 1 0 35952 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_294
timestamp 1486834041
transform 1 0 43792 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_295
timestamp 1486834041
transform 1 0 51632 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_297
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_298
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_299
timestamp 1486834041
transform 1 0 32032 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_300
timestamp 1486834041
transform 1 0 39872 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_301
timestamp 1486834041
transform 1 0 47712 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_302
timestamp 1486834041
transform 1 0 55552 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_304
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_305
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_306
timestamp 1486834041
transform 1 0 28112 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_307
timestamp 1486834041
transform 1 0 35952 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_308
timestamp 1486834041
transform 1 0 43792 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_309
timestamp 1486834041
transform 1 0 51632 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_311
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_312
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_313
timestamp 1486834041
transform 1 0 32032 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_314
timestamp 1486834041
transform 1 0 39872 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_315
timestamp 1486834041
transform 1 0 47712 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_316
timestamp 1486834041
transform 1 0 55552 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_318
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_319
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_320
timestamp 1486834041
transform 1 0 28112 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_321
timestamp 1486834041
transform 1 0 35952 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_322
timestamp 1486834041
transform 1 0 43792 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_323
timestamp 1486834041
transform 1 0 51632 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_325
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_326
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_327
timestamp 1486834041
transform 1 0 32032 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_328
timestamp 1486834041
transform 1 0 39872 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_329
timestamp 1486834041
transform 1 0 47712 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_330
timestamp 1486834041
transform 1 0 55552 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_332
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_333
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_334
timestamp 1486834041
transform 1 0 28112 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_335
timestamp 1486834041
transform 1 0 35952 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_336
timestamp 1486834041
transform 1 0 43792 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_337
timestamp 1486834041
transform 1 0 51632 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_339
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_340
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_341
timestamp 1486834041
transform 1 0 32032 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_342
timestamp 1486834041
transform 1 0 39872 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_343
timestamp 1486834041
transform 1 0 47712 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_344
timestamp 1486834041
transform 1 0 55552 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_346
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_347
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_348
timestamp 1486834041
transform 1 0 28112 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_349
timestamp 1486834041
transform 1 0 35952 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_350
timestamp 1486834041
transform 1 0 43792 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_351
timestamp 1486834041
transform 1 0 51632 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_353
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_354
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_355
timestamp 1486834041
transform 1 0 32032 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_356
timestamp 1486834041
transform 1 0 39872 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_357
timestamp 1486834041
transform 1 0 47712 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_358
timestamp 1486834041
transform 1 0 55552 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_360
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_361
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_362
timestamp 1486834041
transform 1 0 28112 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_363
timestamp 1486834041
transform 1 0 35952 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_364
timestamp 1486834041
transform 1 0 43792 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_365
timestamp 1486834041
transform 1 0 51632 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_367
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_368
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_369
timestamp 1486834041
transform 1 0 32032 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_370
timestamp 1486834041
transform 1 0 39872 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_371
timestamp 1486834041
transform 1 0 47712 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_372
timestamp 1486834041
transform 1 0 55552 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_374
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_375
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_376
timestamp 1486834041
transform 1 0 28112 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_377
timestamp 1486834041
transform 1 0 35952 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_378
timestamp 1486834041
transform 1 0 43792 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_379
timestamp 1486834041
transform 1 0 51632 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_381
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_382
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_383
timestamp 1486834041
transform 1 0 32032 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_384
timestamp 1486834041
transform 1 0 39872 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_385
timestamp 1486834041
transform 1 0 47712 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_386
timestamp 1486834041
transform 1 0 55552 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_388
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_389
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_390
timestamp 1486834041
transform 1 0 28112 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_391
timestamp 1486834041
transform 1 0 35952 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_392
timestamp 1486834041
transform 1 0 43792 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_393
timestamp 1486834041
transform 1 0 51632 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_395
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_396
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_397
timestamp 1486834041
transform 1 0 32032 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_398
timestamp 1486834041
transform 1 0 39872 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_399
timestamp 1486834041
transform 1 0 47712 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_400
timestamp 1486834041
transform 1 0 55552 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_402
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_403
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_404
timestamp 1486834041
transform 1 0 28112 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_405
timestamp 1486834041
transform 1 0 35952 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_406
timestamp 1486834041
transform 1 0 43792 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_407
timestamp 1486834041
transform 1 0 51632 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_409
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_410
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_411
timestamp 1486834041
transform 1 0 32032 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_412
timestamp 1486834041
transform 1 0 39872 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_413
timestamp 1486834041
transform 1 0 47712 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_414
timestamp 1486834041
transform 1 0 55552 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_416
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_417
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_418
timestamp 1486834041
transform 1 0 28112 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_419
timestamp 1486834041
transform 1 0 35952 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_420
timestamp 1486834041
transform 1 0 43792 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_421
timestamp 1486834041
transform 1 0 51632 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_423
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_424
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_425
timestamp 1486834041
transform 1 0 32032 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_426
timestamp 1486834041
transform 1 0 39872 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_427
timestamp 1486834041
transform 1 0 47712 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_428
timestamp 1486834041
transform 1 0 55552 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_430
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_431
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_432
timestamp 1486834041
transform 1 0 28112 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_433
timestamp 1486834041
transform 1 0 35952 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_434
timestamp 1486834041
transform 1 0 43792 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_435
timestamp 1486834041
transform 1 0 51632 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_437
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_438
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_439
timestamp 1486834041
transform 1 0 32032 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_440
timestamp 1486834041
transform 1 0 39872 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_441
timestamp 1486834041
transform 1 0 47712 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_442
timestamp 1486834041
transform 1 0 55552 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_444
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_445
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_446
timestamp 1486834041
transform 1 0 28112 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_447
timestamp 1486834041
transform 1 0 35952 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_448
timestamp 1486834041
transform 1 0 43792 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_449
timestamp 1486834041
transform 1 0 51632 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_451
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_452
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_453
timestamp 1486834041
transform 1 0 32032 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_454
timestamp 1486834041
transform 1 0 39872 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_455
timestamp 1486834041
transform 1 0 47712 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_456
timestamp 1486834041
transform 1 0 55552 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_458
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_459
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_460
timestamp 1486834041
transform 1 0 28112 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_461
timestamp 1486834041
transform 1 0 35952 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_462
timestamp 1486834041
transform 1 0 43792 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_463
timestamp 1486834041
transform 1 0 51632 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_465
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_466
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_467
timestamp 1486834041
transform 1 0 32032 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_468
timestamp 1486834041
transform 1 0 39872 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_469
timestamp 1486834041
transform 1 0 47712 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_470
timestamp 1486834041
transform 1 0 55552 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_472
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_473
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_474
timestamp 1486834041
transform 1 0 28112 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_475
timestamp 1486834041
transform 1 0 35952 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_476
timestamp 1486834041
transform 1 0 43792 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_477
timestamp 1486834041
transform 1 0 51632 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_479
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_480
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_481
timestamp 1486834041
transform 1 0 32032 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_482
timestamp 1486834041
transform 1 0 39872 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_483
timestamp 1486834041
transform 1 0 47712 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_484
timestamp 1486834041
transform 1 0 55552 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_486
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_487
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_488
timestamp 1486834041
transform 1 0 28112 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_489
timestamp 1486834041
transform 1 0 35952 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_490
timestamp 1486834041
transform 1 0 43792 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_491
timestamp 1486834041
transform 1 0 51632 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_493
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_494
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_495
timestamp 1486834041
transform 1 0 32032 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_496
timestamp 1486834041
transform 1 0 39872 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_497
timestamp 1486834041
transform 1 0 47712 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_498
timestamp 1486834041
transform 1 0 55552 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_500
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_501
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_502
timestamp 1486834041
transform 1 0 28112 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_503
timestamp 1486834041
transform 1 0 35952 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_504
timestamp 1486834041
transform 1 0 43792 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_505
timestamp 1486834041
transform 1 0 51632 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_507
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_508
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_509
timestamp 1486834041
transform 1 0 32032 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_510
timestamp 1486834041
transform 1 0 39872 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_511
timestamp 1486834041
transform 1 0 47712 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_512
timestamp 1486834041
transform 1 0 55552 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_514
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_515
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_516
timestamp 1486834041
transform 1 0 28112 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_517
timestamp 1486834041
transform 1 0 35952 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_518
timestamp 1486834041
transform 1 0 43792 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_519
timestamp 1486834041
transform 1 0 51632 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_521
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_522
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_523
timestamp 1486834041
transform 1 0 32032 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_524
timestamp 1486834041
transform 1 0 39872 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_525
timestamp 1486834041
transform 1 0 47712 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_526
timestamp 1486834041
transform 1 0 55552 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_528
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_529
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_530
timestamp 1486834041
transform 1 0 28112 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_531
timestamp 1486834041
transform 1 0 35952 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_532
timestamp 1486834041
transform 1 0 43792 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_533
timestamp 1486834041
transform 1 0 51632 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_535
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_536
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_537
timestamp 1486834041
transform 1 0 32032 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_538
timestamp 1486834041
transform 1 0 39872 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_539
timestamp 1486834041
transform 1 0 47712 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_540
timestamp 1486834041
transform 1 0 55552 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_542
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_543
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_544
timestamp 1486834041
transform 1 0 28112 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_545
timestamp 1486834041
transform 1 0 35952 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_546
timestamp 1486834041
transform 1 0 43792 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_547
timestamp 1486834041
transform 1 0 51632 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_549
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_550
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_551
timestamp 1486834041
transform 1 0 32032 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_552
timestamp 1486834041
transform 1 0 39872 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_553
timestamp 1486834041
transform 1 0 47712 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_554
timestamp 1486834041
transform 1 0 55552 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_556
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_557
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_558
timestamp 1486834041
transform 1 0 28112 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_559
timestamp 1486834041
transform 1 0 35952 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_560
timestamp 1486834041
transform 1 0 43792 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_561
timestamp 1486834041
transform 1 0 51632 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_563
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_564
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_565
timestamp 1486834041
transform 1 0 32032 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_566
timestamp 1486834041
transform 1 0 39872 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_567
timestamp 1486834041
transform 1 0 47712 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_568
timestamp 1486834041
transform 1 0 55552 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_570
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_571
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_572
timestamp 1486834041
transform 1 0 28112 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_573
timestamp 1486834041
transform 1 0 35952 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_574
timestamp 1486834041
transform 1 0 43792 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_575
timestamp 1486834041
transform 1 0 51632 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_577
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_578
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_579
timestamp 1486834041
transform 1 0 32032 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_580
timestamp 1486834041
transform 1 0 39872 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_581
timestamp 1486834041
transform 1 0 47712 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_582
timestamp 1486834041
transform 1 0 55552 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_584
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_585
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_586
timestamp 1486834041
transform 1 0 28112 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_587
timestamp 1486834041
transform 1 0 35952 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_588
timestamp 1486834041
transform 1 0 43792 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_589
timestamp 1486834041
transform 1 0 51632 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_591
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_592
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_593
timestamp 1486834041
transform 1 0 32032 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_594
timestamp 1486834041
transform 1 0 39872 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_595
timestamp 1486834041
transform 1 0 47712 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_596
timestamp 1486834041
transform 1 0 55552 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_598
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_599
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_600
timestamp 1486834041
transform 1 0 28112 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_601
timestamp 1486834041
transform 1 0 35952 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_602
timestamp 1486834041
transform 1 0 43792 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_603
timestamp 1486834041
transform 1 0 51632 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_605
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_606
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_607
timestamp 1486834041
transform 1 0 32032 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_608
timestamp 1486834041
transform 1 0 39872 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_609
timestamp 1486834041
transform 1 0 47712 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_610
timestamp 1486834041
transform 1 0 55552 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_612
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_613
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_614
timestamp 1486834041
transform 1 0 28112 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_615
timestamp 1486834041
transform 1 0 35952 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_616
timestamp 1486834041
transform 1 0 43792 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_617
timestamp 1486834041
transform 1 0 51632 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1486834041
transform 1 0 32032 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1486834041
transform 1 0 39872 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1486834041
transform 1 0 47712 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1486834041
transform 1 0 55552 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_625
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_626
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_627
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_628
timestamp 1486834041
transform 1 0 28112 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_629
timestamp 1486834041
transform 1 0 35952 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_630
timestamp 1486834041
transform 1 0 43792 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_631
timestamp 1486834041
transform 1 0 51632 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_632
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_633
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_634
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_635
timestamp 1486834041
transform 1 0 32032 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_636
timestamp 1486834041
transform 1 0 39872 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_637
timestamp 1486834041
transform 1 0 47712 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_638
timestamp 1486834041
transform 1 0 55552 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_639
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_640
timestamp 1486834041
transform 1 0 8288 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_641
timestamp 1486834041
transform 1 0 12096 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_642
timestamp 1486834041
transform 1 0 15904 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_643
timestamp 1486834041
transform 1 0 19712 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_644
timestamp 1486834041
transform 1 0 23520 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_645
timestamp 1486834041
transform 1 0 27328 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_646
timestamp 1486834041
transform 1 0 31136 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_647
timestamp 1486834041
transform 1 0 34944 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_648
timestamp 1486834041
transform 1 0 38752 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_649
timestamp 1486834041
transform 1 0 42560 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_650
timestamp 1486834041
transform 1 0 46368 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_651
timestamp 1486834041
transform 1 0 50176 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_652
timestamp 1486834041
transform 1 0 53984 0 1 55664
box -86 -86 310 870
<< labels >>
flabel metal2 s 23968 0 24080 112 0 FreeSans 448 0 0 0 Ci
port 0 nsew signal input
flabel metal2 s 23968 57344 24080 57456 0 FreeSans 448 0 0 0 Co
port 1 nsew signal output
flabel metal3 s 57344 21728 57456 21840 0 FreeSans 448 0 0 0 E1BEG[0]
port 2 nsew signal output
flabel metal3 s 57344 22176 57456 22288 0 FreeSans 448 0 0 0 E1BEG[1]
port 3 nsew signal output
flabel metal3 s 57344 22624 57456 22736 0 FreeSans 448 0 0 0 E1BEG[2]
port 4 nsew signal output
flabel metal3 s 57344 23072 57456 23184 0 FreeSans 448 0 0 0 E1BEG[3]
port 5 nsew signal output
flabel metal3 s 0 21728 112 21840 0 FreeSans 448 0 0 0 E1END[0]
port 6 nsew signal input
flabel metal3 s 0 22176 112 22288 0 FreeSans 448 0 0 0 E1END[1]
port 7 nsew signal input
flabel metal3 s 0 22624 112 22736 0 FreeSans 448 0 0 0 E1END[2]
port 8 nsew signal input
flabel metal3 s 0 23072 112 23184 0 FreeSans 448 0 0 0 E1END[3]
port 9 nsew signal input
flabel metal3 s 57344 23520 57456 23632 0 FreeSans 448 0 0 0 E2BEG[0]
port 10 nsew signal output
flabel metal3 s 57344 23968 57456 24080 0 FreeSans 448 0 0 0 E2BEG[1]
port 11 nsew signal output
flabel metal3 s 57344 24416 57456 24528 0 FreeSans 448 0 0 0 E2BEG[2]
port 12 nsew signal output
flabel metal3 s 57344 24864 57456 24976 0 FreeSans 448 0 0 0 E2BEG[3]
port 13 nsew signal output
flabel metal3 s 57344 25312 57456 25424 0 FreeSans 448 0 0 0 E2BEG[4]
port 14 nsew signal output
flabel metal3 s 57344 25760 57456 25872 0 FreeSans 448 0 0 0 E2BEG[5]
port 15 nsew signal output
flabel metal3 s 57344 26208 57456 26320 0 FreeSans 448 0 0 0 E2BEG[6]
port 16 nsew signal output
flabel metal3 s 57344 26656 57456 26768 0 FreeSans 448 0 0 0 E2BEG[7]
port 17 nsew signal output
flabel metal3 s 57344 27104 57456 27216 0 FreeSans 448 0 0 0 E2BEGb[0]
port 18 nsew signal output
flabel metal3 s 57344 27552 57456 27664 0 FreeSans 448 0 0 0 E2BEGb[1]
port 19 nsew signal output
flabel metal3 s 57344 28000 57456 28112 0 FreeSans 448 0 0 0 E2BEGb[2]
port 20 nsew signal output
flabel metal3 s 57344 28448 57456 28560 0 FreeSans 448 0 0 0 E2BEGb[3]
port 21 nsew signal output
flabel metal3 s 57344 28896 57456 29008 0 FreeSans 448 0 0 0 E2BEGb[4]
port 22 nsew signal output
flabel metal3 s 57344 29344 57456 29456 0 FreeSans 448 0 0 0 E2BEGb[5]
port 23 nsew signal output
flabel metal3 s 57344 29792 57456 29904 0 FreeSans 448 0 0 0 E2BEGb[6]
port 24 nsew signal output
flabel metal3 s 57344 30240 57456 30352 0 FreeSans 448 0 0 0 E2BEGb[7]
port 25 nsew signal output
flabel metal3 s 0 27104 112 27216 0 FreeSans 448 0 0 0 E2END[0]
port 26 nsew signal input
flabel metal3 s 0 27552 112 27664 0 FreeSans 448 0 0 0 E2END[1]
port 27 nsew signal input
flabel metal3 s 0 28000 112 28112 0 FreeSans 448 0 0 0 E2END[2]
port 28 nsew signal input
flabel metal3 s 0 28448 112 28560 0 FreeSans 448 0 0 0 E2END[3]
port 29 nsew signal input
flabel metal3 s 0 28896 112 29008 0 FreeSans 448 0 0 0 E2END[4]
port 30 nsew signal input
flabel metal3 s 0 29344 112 29456 0 FreeSans 448 0 0 0 E2END[5]
port 31 nsew signal input
flabel metal3 s 0 29792 112 29904 0 FreeSans 448 0 0 0 E2END[6]
port 32 nsew signal input
flabel metal3 s 0 30240 112 30352 0 FreeSans 448 0 0 0 E2END[7]
port 33 nsew signal input
flabel metal3 s 0 23520 112 23632 0 FreeSans 448 0 0 0 E2MID[0]
port 34 nsew signal input
flabel metal3 s 0 23968 112 24080 0 FreeSans 448 0 0 0 E2MID[1]
port 35 nsew signal input
flabel metal3 s 0 24416 112 24528 0 FreeSans 448 0 0 0 E2MID[2]
port 36 nsew signal input
flabel metal3 s 0 24864 112 24976 0 FreeSans 448 0 0 0 E2MID[3]
port 37 nsew signal input
flabel metal3 s 0 25312 112 25424 0 FreeSans 448 0 0 0 E2MID[4]
port 38 nsew signal input
flabel metal3 s 0 25760 112 25872 0 FreeSans 448 0 0 0 E2MID[5]
port 39 nsew signal input
flabel metal3 s 0 26208 112 26320 0 FreeSans 448 0 0 0 E2MID[6]
port 40 nsew signal input
flabel metal3 s 0 26656 112 26768 0 FreeSans 448 0 0 0 E2MID[7]
port 41 nsew signal input
flabel metal3 s 57344 37856 57456 37968 0 FreeSans 448 0 0 0 E6BEG[0]
port 42 nsew signal output
flabel metal3 s 57344 42336 57456 42448 0 FreeSans 448 0 0 0 E6BEG[10]
port 43 nsew signal output
flabel metal3 s 57344 42784 57456 42896 0 FreeSans 448 0 0 0 E6BEG[11]
port 44 nsew signal output
flabel metal3 s 57344 38304 57456 38416 0 FreeSans 448 0 0 0 E6BEG[1]
port 45 nsew signal output
flabel metal3 s 57344 38752 57456 38864 0 FreeSans 448 0 0 0 E6BEG[2]
port 46 nsew signal output
flabel metal3 s 57344 39200 57456 39312 0 FreeSans 448 0 0 0 E6BEG[3]
port 47 nsew signal output
flabel metal3 s 57344 39648 57456 39760 0 FreeSans 448 0 0 0 E6BEG[4]
port 48 nsew signal output
flabel metal3 s 57344 40096 57456 40208 0 FreeSans 448 0 0 0 E6BEG[5]
port 49 nsew signal output
flabel metal3 s 57344 40544 57456 40656 0 FreeSans 448 0 0 0 E6BEG[6]
port 50 nsew signal output
flabel metal3 s 57344 40992 57456 41104 0 FreeSans 448 0 0 0 E6BEG[7]
port 51 nsew signal output
flabel metal3 s 57344 41440 57456 41552 0 FreeSans 448 0 0 0 E6BEG[8]
port 52 nsew signal output
flabel metal3 s 57344 41888 57456 42000 0 FreeSans 448 0 0 0 E6BEG[9]
port 53 nsew signal output
flabel metal3 s 0 37856 112 37968 0 FreeSans 448 0 0 0 E6END[0]
port 54 nsew signal input
flabel metal3 s 0 42336 112 42448 0 FreeSans 448 0 0 0 E6END[10]
port 55 nsew signal input
flabel metal3 s 0 42784 112 42896 0 FreeSans 448 0 0 0 E6END[11]
port 56 nsew signal input
flabel metal3 s 0 38304 112 38416 0 FreeSans 448 0 0 0 E6END[1]
port 57 nsew signal input
flabel metal3 s 0 38752 112 38864 0 FreeSans 448 0 0 0 E6END[2]
port 58 nsew signal input
flabel metal3 s 0 39200 112 39312 0 FreeSans 448 0 0 0 E6END[3]
port 59 nsew signal input
flabel metal3 s 0 39648 112 39760 0 FreeSans 448 0 0 0 E6END[4]
port 60 nsew signal input
flabel metal3 s 0 40096 112 40208 0 FreeSans 448 0 0 0 E6END[5]
port 61 nsew signal input
flabel metal3 s 0 40544 112 40656 0 FreeSans 448 0 0 0 E6END[6]
port 62 nsew signal input
flabel metal3 s 0 40992 112 41104 0 FreeSans 448 0 0 0 E6END[7]
port 63 nsew signal input
flabel metal3 s 0 41440 112 41552 0 FreeSans 448 0 0 0 E6END[8]
port 64 nsew signal input
flabel metal3 s 0 41888 112 42000 0 FreeSans 448 0 0 0 E6END[9]
port 65 nsew signal input
flabel metal3 s 57344 30688 57456 30800 0 FreeSans 448 0 0 0 EE4BEG[0]
port 66 nsew signal output
flabel metal3 s 57344 35168 57456 35280 0 FreeSans 448 0 0 0 EE4BEG[10]
port 67 nsew signal output
flabel metal3 s 57344 35616 57456 35728 0 FreeSans 448 0 0 0 EE4BEG[11]
port 68 nsew signal output
flabel metal3 s 57344 36064 57456 36176 0 FreeSans 448 0 0 0 EE4BEG[12]
port 69 nsew signal output
flabel metal3 s 57344 36512 57456 36624 0 FreeSans 448 0 0 0 EE4BEG[13]
port 70 nsew signal output
flabel metal3 s 57344 36960 57456 37072 0 FreeSans 448 0 0 0 EE4BEG[14]
port 71 nsew signal output
flabel metal3 s 57344 37408 57456 37520 0 FreeSans 448 0 0 0 EE4BEG[15]
port 72 nsew signal output
flabel metal3 s 57344 31136 57456 31248 0 FreeSans 448 0 0 0 EE4BEG[1]
port 73 nsew signal output
flabel metal3 s 57344 31584 57456 31696 0 FreeSans 448 0 0 0 EE4BEG[2]
port 74 nsew signal output
flabel metal3 s 57344 32032 57456 32144 0 FreeSans 448 0 0 0 EE4BEG[3]
port 75 nsew signal output
flabel metal3 s 57344 32480 57456 32592 0 FreeSans 448 0 0 0 EE4BEG[4]
port 76 nsew signal output
flabel metal3 s 57344 32928 57456 33040 0 FreeSans 448 0 0 0 EE4BEG[5]
port 77 nsew signal output
flabel metal3 s 57344 33376 57456 33488 0 FreeSans 448 0 0 0 EE4BEG[6]
port 78 nsew signal output
flabel metal3 s 57344 33824 57456 33936 0 FreeSans 448 0 0 0 EE4BEG[7]
port 79 nsew signal output
flabel metal3 s 57344 34272 57456 34384 0 FreeSans 448 0 0 0 EE4BEG[8]
port 80 nsew signal output
flabel metal3 s 57344 34720 57456 34832 0 FreeSans 448 0 0 0 EE4BEG[9]
port 81 nsew signal output
flabel metal3 s 0 30688 112 30800 0 FreeSans 448 0 0 0 EE4END[0]
port 82 nsew signal input
flabel metal3 s 0 35168 112 35280 0 FreeSans 448 0 0 0 EE4END[10]
port 83 nsew signal input
flabel metal3 s 0 35616 112 35728 0 FreeSans 448 0 0 0 EE4END[11]
port 84 nsew signal input
flabel metal3 s 0 36064 112 36176 0 FreeSans 448 0 0 0 EE4END[12]
port 85 nsew signal input
flabel metal3 s 0 36512 112 36624 0 FreeSans 448 0 0 0 EE4END[13]
port 86 nsew signal input
flabel metal3 s 0 36960 112 37072 0 FreeSans 448 0 0 0 EE4END[14]
port 87 nsew signal input
flabel metal3 s 0 37408 112 37520 0 FreeSans 448 0 0 0 EE4END[15]
port 88 nsew signal input
flabel metal3 s 0 31136 112 31248 0 FreeSans 448 0 0 0 EE4END[1]
port 89 nsew signal input
flabel metal3 s 0 31584 112 31696 0 FreeSans 448 0 0 0 EE4END[2]
port 90 nsew signal input
flabel metal3 s 0 32032 112 32144 0 FreeSans 448 0 0 0 EE4END[3]
port 91 nsew signal input
flabel metal3 s 0 32480 112 32592 0 FreeSans 448 0 0 0 EE4END[4]
port 92 nsew signal input
flabel metal3 s 0 32928 112 33040 0 FreeSans 448 0 0 0 EE4END[5]
port 93 nsew signal input
flabel metal3 s 0 33376 112 33488 0 FreeSans 448 0 0 0 EE4END[6]
port 94 nsew signal input
flabel metal3 s 0 33824 112 33936 0 FreeSans 448 0 0 0 EE4END[7]
port 95 nsew signal input
flabel metal3 s 0 34272 112 34384 0 FreeSans 448 0 0 0 EE4END[8]
port 96 nsew signal input
flabel metal3 s 0 34720 112 34832 0 FreeSans 448 0 0 0 EE4END[9]
port 97 nsew signal input
flabel metal3 s 0 43232 112 43344 0 FreeSans 448 0 0 0 FrameData[0]
port 98 nsew signal input
flabel metal3 s 0 47712 112 47824 0 FreeSans 448 0 0 0 FrameData[10]
port 99 nsew signal input
flabel metal3 s 0 48160 112 48272 0 FreeSans 448 0 0 0 FrameData[11]
port 100 nsew signal input
flabel metal3 s 0 48608 112 48720 0 FreeSans 448 0 0 0 FrameData[12]
port 101 nsew signal input
flabel metal3 s 0 49056 112 49168 0 FreeSans 448 0 0 0 FrameData[13]
port 102 nsew signal input
flabel metal3 s 0 49504 112 49616 0 FreeSans 448 0 0 0 FrameData[14]
port 103 nsew signal input
flabel metal3 s 0 49952 112 50064 0 FreeSans 448 0 0 0 FrameData[15]
port 104 nsew signal input
flabel metal3 s 0 50400 112 50512 0 FreeSans 448 0 0 0 FrameData[16]
port 105 nsew signal input
flabel metal3 s 0 50848 112 50960 0 FreeSans 448 0 0 0 FrameData[17]
port 106 nsew signal input
flabel metal3 s 0 51296 112 51408 0 FreeSans 448 0 0 0 FrameData[18]
port 107 nsew signal input
flabel metal3 s 0 51744 112 51856 0 FreeSans 448 0 0 0 FrameData[19]
port 108 nsew signal input
flabel metal3 s 0 43680 112 43792 0 FreeSans 448 0 0 0 FrameData[1]
port 109 nsew signal input
flabel metal3 s 0 52192 112 52304 0 FreeSans 448 0 0 0 FrameData[20]
port 110 nsew signal input
flabel metal3 s 0 52640 112 52752 0 FreeSans 448 0 0 0 FrameData[21]
port 111 nsew signal input
flabel metal3 s 0 53088 112 53200 0 FreeSans 448 0 0 0 FrameData[22]
port 112 nsew signal input
flabel metal3 s 0 53536 112 53648 0 FreeSans 448 0 0 0 FrameData[23]
port 113 nsew signal input
flabel metal3 s 0 53984 112 54096 0 FreeSans 448 0 0 0 FrameData[24]
port 114 nsew signal input
flabel metal3 s 0 54432 112 54544 0 FreeSans 448 0 0 0 FrameData[25]
port 115 nsew signal input
flabel metal3 s 0 54880 112 54992 0 FreeSans 448 0 0 0 FrameData[26]
port 116 nsew signal input
flabel metal3 s 0 55328 112 55440 0 FreeSans 448 0 0 0 FrameData[27]
port 117 nsew signal input
flabel metal3 s 0 55776 112 55888 0 FreeSans 448 0 0 0 FrameData[28]
port 118 nsew signal input
flabel metal3 s 0 56224 112 56336 0 FreeSans 448 0 0 0 FrameData[29]
port 119 nsew signal input
flabel metal3 s 0 44128 112 44240 0 FreeSans 448 0 0 0 FrameData[2]
port 120 nsew signal input
flabel metal3 s 0 56672 112 56784 0 FreeSans 448 0 0 0 FrameData[30]
port 121 nsew signal input
flabel metal3 s 0 57120 112 57232 0 FreeSans 448 0 0 0 FrameData[31]
port 122 nsew signal input
flabel metal3 s 0 44576 112 44688 0 FreeSans 448 0 0 0 FrameData[3]
port 123 nsew signal input
flabel metal3 s 0 45024 112 45136 0 FreeSans 448 0 0 0 FrameData[4]
port 124 nsew signal input
flabel metal3 s 0 45472 112 45584 0 FreeSans 448 0 0 0 FrameData[5]
port 125 nsew signal input
flabel metal3 s 0 45920 112 46032 0 FreeSans 448 0 0 0 FrameData[6]
port 126 nsew signal input
flabel metal3 s 0 46368 112 46480 0 FreeSans 448 0 0 0 FrameData[7]
port 127 nsew signal input
flabel metal3 s 0 46816 112 46928 0 FreeSans 448 0 0 0 FrameData[8]
port 128 nsew signal input
flabel metal3 s 0 47264 112 47376 0 FreeSans 448 0 0 0 FrameData[9]
port 129 nsew signal input
flabel metal3 s 57344 43232 57456 43344 0 FreeSans 448 0 0 0 FrameData_O[0]
port 130 nsew signal output
flabel metal3 s 57344 47712 57456 47824 0 FreeSans 448 0 0 0 FrameData_O[10]
port 131 nsew signal output
flabel metal3 s 57344 48160 57456 48272 0 FreeSans 448 0 0 0 FrameData_O[11]
port 132 nsew signal output
flabel metal3 s 57344 48608 57456 48720 0 FreeSans 448 0 0 0 FrameData_O[12]
port 133 nsew signal output
flabel metal3 s 57344 49056 57456 49168 0 FreeSans 448 0 0 0 FrameData_O[13]
port 134 nsew signal output
flabel metal3 s 57344 49504 57456 49616 0 FreeSans 448 0 0 0 FrameData_O[14]
port 135 nsew signal output
flabel metal3 s 57344 49952 57456 50064 0 FreeSans 448 0 0 0 FrameData_O[15]
port 136 nsew signal output
flabel metal3 s 57344 50400 57456 50512 0 FreeSans 448 0 0 0 FrameData_O[16]
port 137 nsew signal output
flabel metal3 s 57344 50848 57456 50960 0 FreeSans 448 0 0 0 FrameData_O[17]
port 138 nsew signal output
flabel metal3 s 57344 51296 57456 51408 0 FreeSans 448 0 0 0 FrameData_O[18]
port 139 nsew signal output
flabel metal3 s 57344 51744 57456 51856 0 FreeSans 448 0 0 0 FrameData_O[19]
port 140 nsew signal output
flabel metal3 s 57344 43680 57456 43792 0 FreeSans 448 0 0 0 FrameData_O[1]
port 141 nsew signal output
flabel metal3 s 57344 52192 57456 52304 0 FreeSans 448 0 0 0 FrameData_O[20]
port 142 nsew signal output
flabel metal3 s 57344 52640 57456 52752 0 FreeSans 448 0 0 0 FrameData_O[21]
port 143 nsew signal output
flabel metal3 s 57344 53088 57456 53200 0 FreeSans 448 0 0 0 FrameData_O[22]
port 144 nsew signal output
flabel metal3 s 57344 53536 57456 53648 0 FreeSans 448 0 0 0 FrameData_O[23]
port 145 nsew signal output
flabel metal3 s 57344 53984 57456 54096 0 FreeSans 448 0 0 0 FrameData_O[24]
port 146 nsew signal output
flabel metal3 s 57344 54432 57456 54544 0 FreeSans 448 0 0 0 FrameData_O[25]
port 147 nsew signal output
flabel metal3 s 57344 54880 57456 54992 0 FreeSans 448 0 0 0 FrameData_O[26]
port 148 nsew signal output
flabel metal3 s 57344 55328 57456 55440 0 FreeSans 448 0 0 0 FrameData_O[27]
port 149 nsew signal output
flabel metal3 s 57344 55776 57456 55888 0 FreeSans 448 0 0 0 FrameData_O[28]
port 150 nsew signal output
flabel metal3 s 57344 56224 57456 56336 0 FreeSans 448 0 0 0 FrameData_O[29]
port 151 nsew signal output
flabel metal3 s 57344 44128 57456 44240 0 FreeSans 448 0 0 0 FrameData_O[2]
port 152 nsew signal output
flabel metal3 s 57344 56672 57456 56784 0 FreeSans 448 0 0 0 FrameData_O[30]
port 153 nsew signal output
flabel metal3 s 57344 57120 57456 57232 0 FreeSans 448 0 0 0 FrameData_O[31]
port 154 nsew signal output
flabel metal3 s 57344 44576 57456 44688 0 FreeSans 448 0 0 0 FrameData_O[3]
port 155 nsew signal output
flabel metal3 s 57344 45024 57456 45136 0 FreeSans 448 0 0 0 FrameData_O[4]
port 156 nsew signal output
flabel metal3 s 57344 45472 57456 45584 0 FreeSans 448 0 0 0 FrameData_O[5]
port 157 nsew signal output
flabel metal3 s 57344 45920 57456 46032 0 FreeSans 448 0 0 0 FrameData_O[6]
port 158 nsew signal output
flabel metal3 s 57344 46368 57456 46480 0 FreeSans 448 0 0 0 FrameData_O[7]
port 159 nsew signal output
flabel metal3 s 57344 46816 57456 46928 0 FreeSans 448 0 0 0 FrameData_O[8]
port 160 nsew signal output
flabel metal3 s 57344 47264 57456 47376 0 FreeSans 448 0 0 0 FrameData_O[9]
port 161 nsew signal output
flabel metal2 s 48160 0 48272 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 162 nsew signal input
flabel metal2 s 52640 0 52752 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 163 nsew signal input
flabel metal2 s 53088 0 53200 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 164 nsew signal input
flabel metal2 s 53536 0 53648 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 165 nsew signal input
flabel metal2 s 53984 0 54096 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 166 nsew signal input
flabel metal2 s 54432 0 54544 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 167 nsew signal input
flabel metal2 s 54880 0 54992 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 168 nsew signal input
flabel metal2 s 55328 0 55440 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 169 nsew signal input
flabel metal2 s 55776 0 55888 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 170 nsew signal input
flabel metal2 s 56224 0 56336 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 171 nsew signal input
flabel metal2 s 56672 0 56784 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 172 nsew signal input
flabel metal2 s 48608 0 48720 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 173 nsew signal input
flabel metal2 s 49056 0 49168 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 174 nsew signal input
flabel metal2 s 49504 0 49616 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 175 nsew signal input
flabel metal2 s 49952 0 50064 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 176 nsew signal input
flabel metal2 s 50400 0 50512 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 177 nsew signal input
flabel metal2 s 50848 0 50960 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 178 nsew signal input
flabel metal2 s 51296 0 51408 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 179 nsew signal input
flabel metal2 s 51744 0 51856 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 180 nsew signal input
flabel metal2 s 52192 0 52304 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 181 nsew signal input
flabel metal2 s 48160 57344 48272 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 182 nsew signal output
flabel metal2 s 52640 57344 52752 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 183 nsew signal output
flabel metal2 s 53088 57344 53200 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 184 nsew signal output
flabel metal2 s 53536 57344 53648 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 185 nsew signal output
flabel metal2 s 53984 57344 54096 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 186 nsew signal output
flabel metal2 s 54432 57344 54544 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 187 nsew signal output
flabel metal2 s 54880 57344 54992 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 188 nsew signal output
flabel metal2 s 55328 57344 55440 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 189 nsew signal output
flabel metal2 s 55776 57344 55888 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 190 nsew signal output
flabel metal2 s 56224 57344 56336 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 191 nsew signal output
flabel metal2 s 56672 57344 56784 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 192 nsew signal output
flabel metal2 s 48608 57344 48720 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 193 nsew signal output
flabel metal2 s 49056 57344 49168 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 194 nsew signal output
flabel metal2 s 49504 57344 49616 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 195 nsew signal output
flabel metal2 s 49952 57344 50064 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 196 nsew signal output
flabel metal2 s 50400 57344 50512 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 197 nsew signal output
flabel metal2 s 50848 57344 50960 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 198 nsew signal output
flabel metal2 s 51296 57344 51408 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 199 nsew signal output
flabel metal2 s 51744 57344 51856 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 200 nsew signal output
flabel metal2 s 52192 57344 52304 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 201 nsew signal output
flabel metal2 s 672 57344 784 57456 0 FreeSans 448 0 0 0 N1BEG[0]
port 202 nsew signal output
flabel metal2 s 1120 57344 1232 57456 0 FreeSans 448 0 0 0 N1BEG[1]
port 203 nsew signal output
flabel metal2 s 1568 57344 1680 57456 0 FreeSans 448 0 0 0 N1BEG[2]
port 204 nsew signal output
flabel metal2 s 2016 57344 2128 57456 0 FreeSans 448 0 0 0 N1BEG[3]
port 205 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 N1END[0]
port 206 nsew signal input
flabel metal2 s 1120 0 1232 112 0 FreeSans 448 0 0 0 N1END[1]
port 207 nsew signal input
flabel metal2 s 1568 0 1680 112 0 FreeSans 448 0 0 0 N1END[2]
port 208 nsew signal input
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 N1END[3]
port 209 nsew signal input
flabel metal2 s 2464 57344 2576 57456 0 FreeSans 448 0 0 0 N2BEG[0]
port 210 nsew signal output
flabel metal2 s 2912 57344 3024 57456 0 FreeSans 448 0 0 0 N2BEG[1]
port 211 nsew signal output
flabel metal2 s 3360 57344 3472 57456 0 FreeSans 448 0 0 0 N2BEG[2]
port 212 nsew signal output
flabel metal2 s 3808 57344 3920 57456 0 FreeSans 448 0 0 0 N2BEG[3]
port 213 nsew signal output
flabel metal2 s 4256 57344 4368 57456 0 FreeSans 448 0 0 0 N2BEG[4]
port 214 nsew signal output
flabel metal2 s 4704 57344 4816 57456 0 FreeSans 448 0 0 0 N2BEG[5]
port 215 nsew signal output
flabel metal2 s 5152 57344 5264 57456 0 FreeSans 448 0 0 0 N2BEG[6]
port 216 nsew signal output
flabel metal2 s 5600 57344 5712 57456 0 FreeSans 448 0 0 0 N2BEG[7]
port 217 nsew signal output
flabel metal2 s 6048 57344 6160 57456 0 FreeSans 448 0 0 0 N2BEGb[0]
port 218 nsew signal output
flabel metal2 s 6496 57344 6608 57456 0 FreeSans 448 0 0 0 N2BEGb[1]
port 219 nsew signal output
flabel metal2 s 6944 57344 7056 57456 0 FreeSans 448 0 0 0 N2BEGb[2]
port 220 nsew signal output
flabel metal2 s 7392 57344 7504 57456 0 FreeSans 448 0 0 0 N2BEGb[3]
port 221 nsew signal output
flabel metal2 s 7840 57344 7952 57456 0 FreeSans 448 0 0 0 N2BEGb[4]
port 222 nsew signal output
flabel metal2 s 8288 57344 8400 57456 0 FreeSans 448 0 0 0 N2BEGb[5]
port 223 nsew signal output
flabel metal2 s 8736 57344 8848 57456 0 FreeSans 448 0 0 0 N2BEGb[6]
port 224 nsew signal output
flabel metal2 s 9184 57344 9296 57456 0 FreeSans 448 0 0 0 N2BEGb[7]
port 225 nsew signal output
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 N2END[0]
port 226 nsew signal input
flabel metal2 s 6496 0 6608 112 0 FreeSans 448 0 0 0 N2END[1]
port 227 nsew signal input
flabel metal2 s 6944 0 7056 112 0 FreeSans 448 0 0 0 N2END[2]
port 228 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 N2END[3]
port 229 nsew signal input
flabel metal2 s 7840 0 7952 112 0 FreeSans 448 0 0 0 N2END[4]
port 230 nsew signal input
flabel metal2 s 8288 0 8400 112 0 FreeSans 448 0 0 0 N2END[5]
port 231 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 N2END[6]
port 232 nsew signal input
flabel metal2 s 9184 0 9296 112 0 FreeSans 448 0 0 0 N2END[7]
port 233 nsew signal input
flabel metal2 s 2464 0 2576 112 0 FreeSans 448 0 0 0 N2MID[0]
port 234 nsew signal input
flabel metal2 s 2912 0 3024 112 0 FreeSans 448 0 0 0 N2MID[1]
port 235 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 N2MID[2]
port 236 nsew signal input
flabel metal2 s 3808 0 3920 112 0 FreeSans 448 0 0 0 N2MID[3]
port 237 nsew signal input
flabel metal2 s 4256 0 4368 112 0 FreeSans 448 0 0 0 N2MID[4]
port 238 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 N2MID[5]
port 239 nsew signal input
flabel metal2 s 5152 0 5264 112 0 FreeSans 448 0 0 0 N2MID[6]
port 240 nsew signal input
flabel metal2 s 5600 0 5712 112 0 FreeSans 448 0 0 0 N2MID[7]
port 241 nsew signal input
flabel metal2 s 9632 57344 9744 57456 0 FreeSans 448 0 0 0 N4BEG[0]
port 242 nsew signal output
flabel metal2 s 14112 57344 14224 57456 0 FreeSans 448 0 0 0 N4BEG[10]
port 243 nsew signal output
flabel metal2 s 14560 57344 14672 57456 0 FreeSans 448 0 0 0 N4BEG[11]
port 244 nsew signal output
flabel metal2 s 15008 57344 15120 57456 0 FreeSans 448 0 0 0 N4BEG[12]
port 245 nsew signal output
flabel metal2 s 15456 57344 15568 57456 0 FreeSans 448 0 0 0 N4BEG[13]
port 246 nsew signal output
flabel metal2 s 15904 57344 16016 57456 0 FreeSans 448 0 0 0 N4BEG[14]
port 247 nsew signal output
flabel metal2 s 16352 57344 16464 57456 0 FreeSans 448 0 0 0 N4BEG[15]
port 248 nsew signal output
flabel metal2 s 10080 57344 10192 57456 0 FreeSans 448 0 0 0 N4BEG[1]
port 249 nsew signal output
flabel metal2 s 10528 57344 10640 57456 0 FreeSans 448 0 0 0 N4BEG[2]
port 250 nsew signal output
flabel metal2 s 10976 57344 11088 57456 0 FreeSans 448 0 0 0 N4BEG[3]
port 251 nsew signal output
flabel metal2 s 11424 57344 11536 57456 0 FreeSans 448 0 0 0 N4BEG[4]
port 252 nsew signal output
flabel metal2 s 11872 57344 11984 57456 0 FreeSans 448 0 0 0 N4BEG[5]
port 253 nsew signal output
flabel metal2 s 12320 57344 12432 57456 0 FreeSans 448 0 0 0 N4BEG[6]
port 254 nsew signal output
flabel metal2 s 12768 57344 12880 57456 0 FreeSans 448 0 0 0 N4BEG[7]
port 255 nsew signal output
flabel metal2 s 13216 57344 13328 57456 0 FreeSans 448 0 0 0 N4BEG[8]
port 256 nsew signal output
flabel metal2 s 13664 57344 13776 57456 0 FreeSans 448 0 0 0 N4BEG[9]
port 257 nsew signal output
flabel metal2 s 9632 0 9744 112 0 FreeSans 448 0 0 0 N4END[0]
port 258 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 N4END[10]
port 259 nsew signal input
flabel metal2 s 14560 0 14672 112 0 FreeSans 448 0 0 0 N4END[11]
port 260 nsew signal input
flabel metal2 s 15008 0 15120 112 0 FreeSans 448 0 0 0 N4END[12]
port 261 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 N4END[13]
port 262 nsew signal input
flabel metal2 s 15904 0 16016 112 0 FreeSans 448 0 0 0 N4END[14]
port 263 nsew signal input
flabel metal2 s 16352 0 16464 112 0 FreeSans 448 0 0 0 N4END[15]
port 264 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 N4END[1]
port 265 nsew signal input
flabel metal2 s 10528 0 10640 112 0 FreeSans 448 0 0 0 N4END[2]
port 266 nsew signal input
flabel metal2 s 10976 0 11088 112 0 FreeSans 448 0 0 0 N4END[3]
port 267 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 N4END[4]
port 268 nsew signal input
flabel metal2 s 11872 0 11984 112 0 FreeSans 448 0 0 0 N4END[5]
port 269 nsew signal input
flabel metal2 s 12320 0 12432 112 0 FreeSans 448 0 0 0 N4END[6]
port 270 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 N4END[7]
port 271 nsew signal input
flabel metal2 s 13216 0 13328 112 0 FreeSans 448 0 0 0 N4END[8]
port 272 nsew signal input
flabel metal2 s 13664 0 13776 112 0 FreeSans 448 0 0 0 N4END[9]
port 273 nsew signal input
flabel metal2 s 16800 57344 16912 57456 0 FreeSans 448 0 0 0 NN4BEG[0]
port 274 nsew signal output
flabel metal2 s 21280 57344 21392 57456 0 FreeSans 448 0 0 0 NN4BEG[10]
port 275 nsew signal output
flabel metal2 s 21728 57344 21840 57456 0 FreeSans 448 0 0 0 NN4BEG[11]
port 276 nsew signal output
flabel metal2 s 22176 57344 22288 57456 0 FreeSans 448 0 0 0 NN4BEG[12]
port 277 nsew signal output
flabel metal2 s 22624 57344 22736 57456 0 FreeSans 448 0 0 0 NN4BEG[13]
port 278 nsew signal output
flabel metal2 s 23072 57344 23184 57456 0 FreeSans 448 0 0 0 NN4BEG[14]
port 279 nsew signal output
flabel metal2 s 23520 57344 23632 57456 0 FreeSans 448 0 0 0 NN4BEG[15]
port 280 nsew signal output
flabel metal2 s 17248 57344 17360 57456 0 FreeSans 448 0 0 0 NN4BEG[1]
port 281 nsew signal output
flabel metal2 s 17696 57344 17808 57456 0 FreeSans 448 0 0 0 NN4BEG[2]
port 282 nsew signal output
flabel metal2 s 18144 57344 18256 57456 0 FreeSans 448 0 0 0 NN4BEG[3]
port 283 nsew signal output
flabel metal2 s 18592 57344 18704 57456 0 FreeSans 448 0 0 0 NN4BEG[4]
port 284 nsew signal output
flabel metal2 s 19040 57344 19152 57456 0 FreeSans 448 0 0 0 NN4BEG[5]
port 285 nsew signal output
flabel metal2 s 19488 57344 19600 57456 0 FreeSans 448 0 0 0 NN4BEG[6]
port 286 nsew signal output
flabel metal2 s 19936 57344 20048 57456 0 FreeSans 448 0 0 0 NN4BEG[7]
port 287 nsew signal output
flabel metal2 s 20384 57344 20496 57456 0 FreeSans 448 0 0 0 NN4BEG[8]
port 288 nsew signal output
flabel metal2 s 20832 57344 20944 57456 0 FreeSans 448 0 0 0 NN4BEG[9]
port 289 nsew signal output
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 NN4END[0]
port 290 nsew signal input
flabel metal2 s 21280 0 21392 112 0 FreeSans 448 0 0 0 NN4END[10]
port 291 nsew signal input
flabel metal2 s 21728 0 21840 112 0 FreeSans 448 0 0 0 NN4END[11]
port 292 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 NN4END[12]
port 293 nsew signal input
flabel metal2 s 22624 0 22736 112 0 FreeSans 448 0 0 0 NN4END[13]
port 294 nsew signal input
flabel metal2 s 23072 0 23184 112 0 FreeSans 448 0 0 0 NN4END[14]
port 295 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 NN4END[15]
port 296 nsew signal input
flabel metal2 s 17248 0 17360 112 0 FreeSans 448 0 0 0 NN4END[1]
port 297 nsew signal input
flabel metal2 s 17696 0 17808 112 0 FreeSans 448 0 0 0 NN4END[2]
port 298 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 NN4END[3]
port 299 nsew signal input
flabel metal2 s 18592 0 18704 112 0 FreeSans 448 0 0 0 NN4END[4]
port 300 nsew signal input
flabel metal2 s 19040 0 19152 112 0 FreeSans 448 0 0 0 NN4END[5]
port 301 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 NN4END[6]
port 302 nsew signal input
flabel metal2 s 19936 0 20048 112 0 FreeSans 448 0 0 0 NN4END[7]
port 303 nsew signal input
flabel metal2 s 20384 0 20496 112 0 FreeSans 448 0 0 0 NN4END[8]
port 304 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 NN4END[9]
port 305 nsew signal input
flabel metal2 s 24416 0 24528 112 0 FreeSans 448 0 0 0 S1BEG[0]
port 306 nsew signal output
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 S1BEG[1]
port 307 nsew signal output
flabel metal2 s 25312 0 25424 112 0 FreeSans 448 0 0 0 S1BEG[2]
port 308 nsew signal output
flabel metal2 s 25760 0 25872 112 0 FreeSans 448 0 0 0 S1BEG[3]
port 309 nsew signal output
flabel metal2 s 24416 57344 24528 57456 0 FreeSans 448 0 0 0 S1END[0]
port 310 nsew signal input
flabel metal2 s 24864 57344 24976 57456 0 FreeSans 448 0 0 0 S1END[1]
port 311 nsew signal input
flabel metal2 s 25312 57344 25424 57456 0 FreeSans 448 0 0 0 S1END[2]
port 312 nsew signal input
flabel metal2 s 25760 57344 25872 57456 0 FreeSans 448 0 0 0 S1END[3]
port 313 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 S2BEG[0]
port 314 nsew signal output
flabel metal2 s 26656 0 26768 112 0 FreeSans 448 0 0 0 S2BEG[1]
port 315 nsew signal output
flabel metal2 s 27104 0 27216 112 0 FreeSans 448 0 0 0 S2BEG[2]
port 316 nsew signal output
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 S2BEG[3]
port 317 nsew signal output
flabel metal2 s 28000 0 28112 112 0 FreeSans 448 0 0 0 S2BEG[4]
port 318 nsew signal output
flabel metal2 s 28448 0 28560 112 0 FreeSans 448 0 0 0 S2BEG[5]
port 319 nsew signal output
flabel metal2 s 28896 0 29008 112 0 FreeSans 448 0 0 0 S2BEG[6]
port 320 nsew signal output
flabel metal2 s 29344 0 29456 112 0 FreeSans 448 0 0 0 S2BEG[7]
port 321 nsew signal output
flabel metal2 s 29792 0 29904 112 0 FreeSans 448 0 0 0 S2BEGb[0]
port 322 nsew signal output
flabel metal2 s 30240 0 30352 112 0 FreeSans 448 0 0 0 S2BEGb[1]
port 323 nsew signal output
flabel metal2 s 30688 0 30800 112 0 FreeSans 448 0 0 0 S2BEGb[2]
port 324 nsew signal output
flabel metal2 s 31136 0 31248 112 0 FreeSans 448 0 0 0 S2BEGb[3]
port 325 nsew signal output
flabel metal2 s 31584 0 31696 112 0 FreeSans 448 0 0 0 S2BEGb[4]
port 326 nsew signal output
flabel metal2 s 32032 0 32144 112 0 FreeSans 448 0 0 0 S2BEGb[5]
port 327 nsew signal output
flabel metal2 s 32480 0 32592 112 0 FreeSans 448 0 0 0 S2BEGb[6]
port 328 nsew signal output
flabel metal2 s 32928 0 33040 112 0 FreeSans 448 0 0 0 S2BEGb[7]
port 329 nsew signal output
flabel metal2 s 29792 57344 29904 57456 0 FreeSans 448 0 0 0 S2END[0]
port 330 nsew signal input
flabel metal2 s 30240 57344 30352 57456 0 FreeSans 448 0 0 0 S2END[1]
port 331 nsew signal input
flabel metal2 s 30688 57344 30800 57456 0 FreeSans 448 0 0 0 S2END[2]
port 332 nsew signal input
flabel metal2 s 31136 57344 31248 57456 0 FreeSans 448 0 0 0 S2END[3]
port 333 nsew signal input
flabel metal2 s 31584 57344 31696 57456 0 FreeSans 448 0 0 0 S2END[4]
port 334 nsew signal input
flabel metal2 s 32032 57344 32144 57456 0 FreeSans 448 0 0 0 S2END[5]
port 335 nsew signal input
flabel metal2 s 32480 57344 32592 57456 0 FreeSans 448 0 0 0 S2END[6]
port 336 nsew signal input
flabel metal2 s 32928 57344 33040 57456 0 FreeSans 448 0 0 0 S2END[7]
port 337 nsew signal input
flabel metal2 s 26208 57344 26320 57456 0 FreeSans 448 0 0 0 S2MID[0]
port 338 nsew signal input
flabel metal2 s 26656 57344 26768 57456 0 FreeSans 448 0 0 0 S2MID[1]
port 339 nsew signal input
flabel metal2 s 27104 57344 27216 57456 0 FreeSans 448 0 0 0 S2MID[2]
port 340 nsew signal input
flabel metal2 s 27552 57344 27664 57456 0 FreeSans 448 0 0 0 S2MID[3]
port 341 nsew signal input
flabel metal2 s 28000 57344 28112 57456 0 FreeSans 448 0 0 0 S2MID[4]
port 342 nsew signal input
flabel metal2 s 28448 57344 28560 57456 0 FreeSans 448 0 0 0 S2MID[5]
port 343 nsew signal input
flabel metal2 s 28896 57344 29008 57456 0 FreeSans 448 0 0 0 S2MID[6]
port 344 nsew signal input
flabel metal2 s 29344 57344 29456 57456 0 FreeSans 448 0 0 0 S2MID[7]
port 345 nsew signal input
flabel metal2 s 33376 0 33488 112 0 FreeSans 448 0 0 0 S4BEG[0]
port 346 nsew signal output
flabel metal2 s 37856 0 37968 112 0 FreeSans 448 0 0 0 S4BEG[10]
port 347 nsew signal output
flabel metal2 s 38304 0 38416 112 0 FreeSans 448 0 0 0 S4BEG[11]
port 348 nsew signal output
flabel metal2 s 38752 0 38864 112 0 FreeSans 448 0 0 0 S4BEG[12]
port 349 nsew signal output
flabel metal2 s 39200 0 39312 112 0 FreeSans 448 0 0 0 S4BEG[13]
port 350 nsew signal output
flabel metal2 s 39648 0 39760 112 0 FreeSans 448 0 0 0 S4BEG[14]
port 351 nsew signal output
flabel metal2 s 40096 0 40208 112 0 FreeSans 448 0 0 0 S4BEG[15]
port 352 nsew signal output
flabel metal2 s 33824 0 33936 112 0 FreeSans 448 0 0 0 S4BEG[1]
port 353 nsew signal output
flabel metal2 s 34272 0 34384 112 0 FreeSans 448 0 0 0 S4BEG[2]
port 354 nsew signal output
flabel metal2 s 34720 0 34832 112 0 FreeSans 448 0 0 0 S4BEG[3]
port 355 nsew signal output
flabel metal2 s 35168 0 35280 112 0 FreeSans 448 0 0 0 S4BEG[4]
port 356 nsew signal output
flabel metal2 s 35616 0 35728 112 0 FreeSans 448 0 0 0 S4BEG[5]
port 357 nsew signal output
flabel metal2 s 36064 0 36176 112 0 FreeSans 448 0 0 0 S4BEG[6]
port 358 nsew signal output
flabel metal2 s 36512 0 36624 112 0 FreeSans 448 0 0 0 S4BEG[7]
port 359 nsew signal output
flabel metal2 s 36960 0 37072 112 0 FreeSans 448 0 0 0 S4BEG[8]
port 360 nsew signal output
flabel metal2 s 37408 0 37520 112 0 FreeSans 448 0 0 0 S4BEG[9]
port 361 nsew signal output
flabel metal2 s 33376 57344 33488 57456 0 FreeSans 448 0 0 0 S4END[0]
port 362 nsew signal input
flabel metal2 s 37856 57344 37968 57456 0 FreeSans 448 0 0 0 S4END[10]
port 363 nsew signal input
flabel metal2 s 38304 57344 38416 57456 0 FreeSans 448 0 0 0 S4END[11]
port 364 nsew signal input
flabel metal2 s 38752 57344 38864 57456 0 FreeSans 448 0 0 0 S4END[12]
port 365 nsew signal input
flabel metal2 s 39200 57344 39312 57456 0 FreeSans 448 0 0 0 S4END[13]
port 366 nsew signal input
flabel metal2 s 39648 57344 39760 57456 0 FreeSans 448 0 0 0 S4END[14]
port 367 nsew signal input
flabel metal2 s 40096 57344 40208 57456 0 FreeSans 448 0 0 0 S4END[15]
port 368 nsew signal input
flabel metal2 s 33824 57344 33936 57456 0 FreeSans 448 0 0 0 S4END[1]
port 369 nsew signal input
flabel metal2 s 34272 57344 34384 57456 0 FreeSans 448 0 0 0 S4END[2]
port 370 nsew signal input
flabel metal2 s 34720 57344 34832 57456 0 FreeSans 448 0 0 0 S4END[3]
port 371 nsew signal input
flabel metal2 s 35168 57344 35280 57456 0 FreeSans 448 0 0 0 S4END[4]
port 372 nsew signal input
flabel metal2 s 35616 57344 35728 57456 0 FreeSans 448 0 0 0 S4END[5]
port 373 nsew signal input
flabel metal2 s 36064 57344 36176 57456 0 FreeSans 448 0 0 0 S4END[6]
port 374 nsew signal input
flabel metal2 s 36512 57344 36624 57456 0 FreeSans 448 0 0 0 S4END[7]
port 375 nsew signal input
flabel metal2 s 36960 57344 37072 57456 0 FreeSans 448 0 0 0 S4END[8]
port 376 nsew signal input
flabel metal2 s 37408 57344 37520 57456 0 FreeSans 448 0 0 0 S4END[9]
port 377 nsew signal input
flabel metal2 s 40544 0 40656 112 0 FreeSans 448 0 0 0 SS4BEG[0]
port 378 nsew signal output
flabel metal2 s 45024 0 45136 112 0 FreeSans 448 0 0 0 SS4BEG[10]
port 379 nsew signal output
flabel metal2 s 45472 0 45584 112 0 FreeSans 448 0 0 0 SS4BEG[11]
port 380 nsew signal output
flabel metal2 s 45920 0 46032 112 0 FreeSans 448 0 0 0 SS4BEG[12]
port 381 nsew signal output
flabel metal2 s 46368 0 46480 112 0 FreeSans 448 0 0 0 SS4BEG[13]
port 382 nsew signal output
flabel metal2 s 46816 0 46928 112 0 FreeSans 448 0 0 0 SS4BEG[14]
port 383 nsew signal output
flabel metal2 s 47264 0 47376 112 0 FreeSans 448 0 0 0 SS4BEG[15]
port 384 nsew signal output
flabel metal2 s 40992 0 41104 112 0 FreeSans 448 0 0 0 SS4BEG[1]
port 385 nsew signal output
flabel metal2 s 41440 0 41552 112 0 FreeSans 448 0 0 0 SS4BEG[2]
port 386 nsew signal output
flabel metal2 s 41888 0 42000 112 0 FreeSans 448 0 0 0 SS4BEG[3]
port 387 nsew signal output
flabel metal2 s 42336 0 42448 112 0 FreeSans 448 0 0 0 SS4BEG[4]
port 388 nsew signal output
flabel metal2 s 42784 0 42896 112 0 FreeSans 448 0 0 0 SS4BEG[5]
port 389 nsew signal output
flabel metal2 s 43232 0 43344 112 0 FreeSans 448 0 0 0 SS4BEG[6]
port 390 nsew signal output
flabel metal2 s 43680 0 43792 112 0 FreeSans 448 0 0 0 SS4BEG[7]
port 391 nsew signal output
flabel metal2 s 44128 0 44240 112 0 FreeSans 448 0 0 0 SS4BEG[8]
port 392 nsew signal output
flabel metal2 s 44576 0 44688 112 0 FreeSans 448 0 0 0 SS4BEG[9]
port 393 nsew signal output
flabel metal2 s 40544 57344 40656 57456 0 FreeSans 448 0 0 0 SS4END[0]
port 394 nsew signal input
flabel metal2 s 45024 57344 45136 57456 0 FreeSans 448 0 0 0 SS4END[10]
port 395 nsew signal input
flabel metal2 s 45472 57344 45584 57456 0 FreeSans 448 0 0 0 SS4END[11]
port 396 nsew signal input
flabel metal2 s 45920 57344 46032 57456 0 FreeSans 448 0 0 0 SS4END[12]
port 397 nsew signal input
flabel metal2 s 46368 57344 46480 57456 0 FreeSans 448 0 0 0 SS4END[13]
port 398 nsew signal input
flabel metal2 s 46816 57344 46928 57456 0 FreeSans 448 0 0 0 SS4END[14]
port 399 nsew signal input
flabel metal2 s 47264 57344 47376 57456 0 FreeSans 448 0 0 0 SS4END[15]
port 400 nsew signal input
flabel metal2 s 40992 57344 41104 57456 0 FreeSans 448 0 0 0 SS4END[1]
port 401 nsew signal input
flabel metal2 s 41440 57344 41552 57456 0 FreeSans 448 0 0 0 SS4END[2]
port 402 nsew signal input
flabel metal2 s 41888 57344 42000 57456 0 FreeSans 448 0 0 0 SS4END[3]
port 403 nsew signal input
flabel metal2 s 42336 57344 42448 57456 0 FreeSans 448 0 0 0 SS4END[4]
port 404 nsew signal input
flabel metal2 s 42784 57344 42896 57456 0 FreeSans 448 0 0 0 SS4END[5]
port 405 nsew signal input
flabel metal2 s 43232 57344 43344 57456 0 FreeSans 448 0 0 0 SS4END[6]
port 406 nsew signal input
flabel metal2 s 43680 57344 43792 57456 0 FreeSans 448 0 0 0 SS4END[7]
port 407 nsew signal input
flabel metal2 s 44128 57344 44240 57456 0 FreeSans 448 0 0 0 SS4END[8]
port 408 nsew signal input
flabel metal2 s 44576 57344 44688 57456 0 FreeSans 448 0 0 0 SS4END[9]
port 409 nsew signal input
flabel metal2 s 47712 0 47824 112 0 FreeSans 448 0 0 0 UserCLK
port 410 nsew signal input
flabel metal2 s 47712 57344 47824 57456 0 FreeSans 448 0 0 0 UserCLKo
port 411 nsew signal output
flabel metal4 s 3776 0 4096 57456 0 FreeSans 1472 90 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 3776 57400 4096 57456 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 23776 0 24096 57456 0 FreeSans 1472 90 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 23776 57400 24096 57456 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 43776 0 44096 57456 0 FreeSans 1472 90 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 43776 57400 44096 57456 0 FreeSans 368 0 0 0 VDD
port 412 nsew power bidirectional
flabel metal4 s 4436 0 4756 57456 0 FreeSans 1472 90 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 4436 57400 4756 57456 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 24436 0 24756 57456 0 FreeSans 1472 90 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 24436 57400 24756 57456 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 44436 0 44756 57456 0 FreeSans 1472 90 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal4 s 44436 57400 44756 57456 0 FreeSans 368 0 0 0 VSS
port 413 nsew ground bidirectional
flabel metal3 s 0 224 112 336 0 FreeSans 448 0 0 0 W1BEG[0]
port 414 nsew signal output
flabel metal3 s 0 672 112 784 0 FreeSans 448 0 0 0 W1BEG[1]
port 415 nsew signal output
flabel metal3 s 0 1120 112 1232 0 FreeSans 448 0 0 0 W1BEG[2]
port 416 nsew signal output
flabel metal3 s 0 1568 112 1680 0 FreeSans 448 0 0 0 W1BEG[3]
port 417 nsew signal output
flabel metal3 s 57344 224 57456 336 0 FreeSans 448 0 0 0 W1END[0]
port 418 nsew signal input
flabel metal3 s 57344 672 57456 784 0 FreeSans 448 0 0 0 W1END[1]
port 419 nsew signal input
flabel metal3 s 57344 1120 57456 1232 0 FreeSans 448 0 0 0 W1END[2]
port 420 nsew signal input
flabel metal3 s 57344 1568 57456 1680 0 FreeSans 448 0 0 0 W1END[3]
port 421 nsew signal input
flabel metal3 s 0 2016 112 2128 0 FreeSans 448 0 0 0 W2BEG[0]
port 422 nsew signal output
flabel metal3 s 0 2464 112 2576 0 FreeSans 448 0 0 0 W2BEG[1]
port 423 nsew signal output
flabel metal3 s 0 2912 112 3024 0 FreeSans 448 0 0 0 W2BEG[2]
port 424 nsew signal output
flabel metal3 s 0 3360 112 3472 0 FreeSans 448 0 0 0 W2BEG[3]
port 425 nsew signal output
flabel metal3 s 0 3808 112 3920 0 FreeSans 448 0 0 0 W2BEG[4]
port 426 nsew signal output
flabel metal3 s 0 4256 112 4368 0 FreeSans 448 0 0 0 W2BEG[5]
port 427 nsew signal output
flabel metal3 s 0 4704 112 4816 0 FreeSans 448 0 0 0 W2BEG[6]
port 428 nsew signal output
flabel metal3 s 0 5152 112 5264 0 FreeSans 448 0 0 0 W2BEG[7]
port 429 nsew signal output
flabel metal3 s 0 5600 112 5712 0 FreeSans 448 0 0 0 W2BEGb[0]
port 430 nsew signal output
flabel metal3 s 0 6048 112 6160 0 FreeSans 448 0 0 0 W2BEGb[1]
port 431 nsew signal output
flabel metal3 s 0 6496 112 6608 0 FreeSans 448 0 0 0 W2BEGb[2]
port 432 nsew signal output
flabel metal3 s 0 6944 112 7056 0 FreeSans 448 0 0 0 W2BEGb[3]
port 433 nsew signal output
flabel metal3 s 0 7392 112 7504 0 FreeSans 448 0 0 0 W2BEGb[4]
port 434 nsew signal output
flabel metal3 s 0 7840 112 7952 0 FreeSans 448 0 0 0 W2BEGb[5]
port 435 nsew signal output
flabel metal3 s 0 8288 112 8400 0 FreeSans 448 0 0 0 W2BEGb[6]
port 436 nsew signal output
flabel metal3 s 0 8736 112 8848 0 FreeSans 448 0 0 0 W2BEGb[7]
port 437 nsew signal output
flabel metal3 s 57344 5600 57456 5712 0 FreeSans 448 0 0 0 W2END[0]
port 438 nsew signal input
flabel metal3 s 57344 6048 57456 6160 0 FreeSans 448 0 0 0 W2END[1]
port 439 nsew signal input
flabel metal3 s 57344 6496 57456 6608 0 FreeSans 448 0 0 0 W2END[2]
port 440 nsew signal input
flabel metal3 s 57344 6944 57456 7056 0 FreeSans 448 0 0 0 W2END[3]
port 441 nsew signal input
flabel metal3 s 57344 7392 57456 7504 0 FreeSans 448 0 0 0 W2END[4]
port 442 nsew signal input
flabel metal3 s 57344 7840 57456 7952 0 FreeSans 448 0 0 0 W2END[5]
port 443 nsew signal input
flabel metal3 s 57344 8288 57456 8400 0 FreeSans 448 0 0 0 W2END[6]
port 444 nsew signal input
flabel metal3 s 57344 8736 57456 8848 0 FreeSans 448 0 0 0 W2END[7]
port 445 nsew signal input
flabel metal3 s 57344 2016 57456 2128 0 FreeSans 448 0 0 0 W2MID[0]
port 446 nsew signal input
flabel metal3 s 57344 2464 57456 2576 0 FreeSans 448 0 0 0 W2MID[1]
port 447 nsew signal input
flabel metal3 s 57344 2912 57456 3024 0 FreeSans 448 0 0 0 W2MID[2]
port 448 nsew signal input
flabel metal3 s 57344 3360 57456 3472 0 FreeSans 448 0 0 0 W2MID[3]
port 449 nsew signal input
flabel metal3 s 57344 3808 57456 3920 0 FreeSans 448 0 0 0 W2MID[4]
port 450 nsew signal input
flabel metal3 s 57344 4256 57456 4368 0 FreeSans 448 0 0 0 W2MID[5]
port 451 nsew signal input
flabel metal3 s 57344 4704 57456 4816 0 FreeSans 448 0 0 0 W2MID[6]
port 452 nsew signal input
flabel metal3 s 57344 5152 57456 5264 0 FreeSans 448 0 0 0 W2MID[7]
port 453 nsew signal input
flabel metal3 s 0 16352 112 16464 0 FreeSans 448 0 0 0 W6BEG[0]
port 454 nsew signal output
flabel metal3 s 0 20832 112 20944 0 FreeSans 448 0 0 0 W6BEG[10]
port 455 nsew signal output
flabel metal3 s 0 21280 112 21392 0 FreeSans 448 0 0 0 W6BEG[11]
port 456 nsew signal output
flabel metal3 s 0 16800 112 16912 0 FreeSans 448 0 0 0 W6BEG[1]
port 457 nsew signal output
flabel metal3 s 0 17248 112 17360 0 FreeSans 448 0 0 0 W6BEG[2]
port 458 nsew signal output
flabel metal3 s 0 17696 112 17808 0 FreeSans 448 0 0 0 W6BEG[3]
port 459 nsew signal output
flabel metal3 s 0 18144 112 18256 0 FreeSans 448 0 0 0 W6BEG[4]
port 460 nsew signal output
flabel metal3 s 0 18592 112 18704 0 FreeSans 448 0 0 0 W6BEG[5]
port 461 nsew signal output
flabel metal3 s 0 19040 112 19152 0 FreeSans 448 0 0 0 W6BEG[6]
port 462 nsew signal output
flabel metal3 s 0 19488 112 19600 0 FreeSans 448 0 0 0 W6BEG[7]
port 463 nsew signal output
flabel metal3 s 0 19936 112 20048 0 FreeSans 448 0 0 0 W6BEG[8]
port 464 nsew signal output
flabel metal3 s 0 20384 112 20496 0 FreeSans 448 0 0 0 W6BEG[9]
port 465 nsew signal output
flabel metal3 s 57344 16352 57456 16464 0 FreeSans 448 0 0 0 W6END[0]
port 466 nsew signal input
flabel metal3 s 57344 20832 57456 20944 0 FreeSans 448 0 0 0 W6END[10]
port 467 nsew signal input
flabel metal3 s 57344 21280 57456 21392 0 FreeSans 448 0 0 0 W6END[11]
port 468 nsew signal input
flabel metal3 s 57344 16800 57456 16912 0 FreeSans 448 0 0 0 W6END[1]
port 469 nsew signal input
flabel metal3 s 57344 17248 57456 17360 0 FreeSans 448 0 0 0 W6END[2]
port 470 nsew signal input
flabel metal3 s 57344 17696 57456 17808 0 FreeSans 448 0 0 0 W6END[3]
port 471 nsew signal input
flabel metal3 s 57344 18144 57456 18256 0 FreeSans 448 0 0 0 W6END[4]
port 472 nsew signal input
flabel metal3 s 57344 18592 57456 18704 0 FreeSans 448 0 0 0 W6END[5]
port 473 nsew signal input
flabel metal3 s 57344 19040 57456 19152 0 FreeSans 448 0 0 0 W6END[6]
port 474 nsew signal input
flabel metal3 s 57344 19488 57456 19600 0 FreeSans 448 0 0 0 W6END[7]
port 475 nsew signal input
flabel metal3 s 57344 19936 57456 20048 0 FreeSans 448 0 0 0 W6END[8]
port 476 nsew signal input
flabel metal3 s 57344 20384 57456 20496 0 FreeSans 448 0 0 0 W6END[9]
port 477 nsew signal input
flabel metal3 s 0 9184 112 9296 0 FreeSans 448 0 0 0 WW4BEG[0]
port 478 nsew signal output
flabel metal3 s 0 13664 112 13776 0 FreeSans 448 0 0 0 WW4BEG[10]
port 479 nsew signal output
flabel metal3 s 0 14112 112 14224 0 FreeSans 448 0 0 0 WW4BEG[11]
port 480 nsew signal output
flabel metal3 s 0 14560 112 14672 0 FreeSans 448 0 0 0 WW4BEG[12]
port 481 nsew signal output
flabel metal3 s 0 15008 112 15120 0 FreeSans 448 0 0 0 WW4BEG[13]
port 482 nsew signal output
flabel metal3 s 0 15456 112 15568 0 FreeSans 448 0 0 0 WW4BEG[14]
port 483 nsew signal output
flabel metal3 s 0 15904 112 16016 0 FreeSans 448 0 0 0 WW4BEG[15]
port 484 nsew signal output
flabel metal3 s 0 9632 112 9744 0 FreeSans 448 0 0 0 WW4BEG[1]
port 485 nsew signal output
flabel metal3 s 0 10080 112 10192 0 FreeSans 448 0 0 0 WW4BEG[2]
port 486 nsew signal output
flabel metal3 s 0 10528 112 10640 0 FreeSans 448 0 0 0 WW4BEG[3]
port 487 nsew signal output
flabel metal3 s 0 10976 112 11088 0 FreeSans 448 0 0 0 WW4BEG[4]
port 488 nsew signal output
flabel metal3 s 0 11424 112 11536 0 FreeSans 448 0 0 0 WW4BEG[5]
port 489 nsew signal output
flabel metal3 s 0 11872 112 11984 0 FreeSans 448 0 0 0 WW4BEG[6]
port 490 nsew signal output
flabel metal3 s 0 12320 112 12432 0 FreeSans 448 0 0 0 WW4BEG[7]
port 491 nsew signal output
flabel metal3 s 0 12768 112 12880 0 FreeSans 448 0 0 0 WW4BEG[8]
port 492 nsew signal output
flabel metal3 s 0 13216 112 13328 0 FreeSans 448 0 0 0 WW4BEG[9]
port 493 nsew signal output
flabel metal3 s 57344 9184 57456 9296 0 FreeSans 448 0 0 0 WW4END[0]
port 494 nsew signal input
flabel metal3 s 57344 13664 57456 13776 0 FreeSans 448 0 0 0 WW4END[10]
port 495 nsew signal input
flabel metal3 s 57344 14112 57456 14224 0 FreeSans 448 0 0 0 WW4END[11]
port 496 nsew signal input
flabel metal3 s 57344 14560 57456 14672 0 FreeSans 448 0 0 0 WW4END[12]
port 497 nsew signal input
flabel metal3 s 57344 15008 57456 15120 0 FreeSans 448 0 0 0 WW4END[13]
port 498 nsew signal input
flabel metal3 s 57344 15456 57456 15568 0 FreeSans 448 0 0 0 WW4END[14]
port 499 nsew signal input
flabel metal3 s 57344 15904 57456 16016 0 FreeSans 448 0 0 0 WW4END[15]
port 500 nsew signal input
flabel metal3 s 57344 9632 57456 9744 0 FreeSans 448 0 0 0 WW4END[1]
port 501 nsew signal input
flabel metal3 s 57344 10080 57456 10192 0 FreeSans 448 0 0 0 WW4END[2]
port 502 nsew signal input
flabel metal3 s 57344 10528 57456 10640 0 FreeSans 448 0 0 0 WW4END[3]
port 503 nsew signal input
flabel metal3 s 57344 10976 57456 11088 0 FreeSans 448 0 0 0 WW4END[4]
port 504 nsew signal input
flabel metal3 s 57344 11424 57456 11536 0 FreeSans 448 0 0 0 WW4END[5]
port 505 nsew signal input
flabel metal3 s 57344 11872 57456 11984 0 FreeSans 448 0 0 0 WW4END[6]
port 506 nsew signal input
flabel metal3 s 57344 12320 57456 12432 0 FreeSans 448 0 0 0 WW4END[7]
port 507 nsew signal input
flabel metal3 s 57344 12768 57456 12880 0 FreeSans 448 0 0 0 WW4END[8]
port 508 nsew signal input
flabel metal3 s 57344 13216 57456 13328 0 FreeSans 448 0 0 0 WW4END[9]
port 509 nsew signal input
rlabel metal1 28728 56448 28728 56448 0 VDD
rlabel metal1 28728 55664 28728 55664 0 VSS
rlabel metal3 16968 15176 16968 15176 0 A
rlabel metal2 3192 39928 3192 39928 0 B
rlabel metal2 19040 23128 19040 23128 0 C
rlabel metal2 49000 9856 49000 9856 0 Ci
rlabel metal2 24248 56280 24248 56280 0 Co
rlabel metal3 2520 47096 2520 47096 0 D
rlabel metal2 21672 42672 21672 42672 0 E
rlabel metal3 56406 21784 56406 21784 0 E1BEG[0]
rlabel metal2 50568 20832 50568 20832 0 E1BEG[1]
rlabel metal3 57330 22680 57330 22680 0 E1BEG[2]
rlabel metal2 49000 21504 49000 21504 0 E1BEG[3]
rlabel metal2 26152 31136 26152 31136 0 E1END[0]
rlabel metal3 406 22232 406 22232 0 E1END[1]
rlabel metal3 1414 22680 1414 22680 0 E1END[2]
rlabel metal2 23464 49616 23464 49616 0 E1END[3]
rlabel metal3 56882 23576 56882 23576 0 E2BEG[0]
rlabel metal3 57106 24024 57106 24024 0 E2BEG[1]
rlabel metal3 56938 24472 56938 24472 0 E2BEG[2]
rlabel metal3 57106 24920 57106 24920 0 E2BEG[3]
rlabel metal3 57330 25368 57330 25368 0 E2BEG[4]
rlabel metal3 56546 25816 56546 25816 0 E2BEG[5]
rlabel metal3 57162 26264 57162 26264 0 E2BEG[6]
rlabel metal2 56280 22680 56280 22680 0 E2BEG[7]
rlabel metal3 56728 17864 56728 17864 0 E2BEGb[0]
rlabel metal3 56784 19432 56784 19432 0 E2BEGb[1]
rlabel metal3 56000 21000 56000 21000 0 E2BEGb[2]
rlabel metal2 56448 24584 56448 24584 0 E2BEGb[3]
rlabel metal2 56392 28336 56392 28336 0 E2BEGb[4]
rlabel metal3 56882 29400 56882 29400 0 E2BEGb[5]
rlabel metal3 56994 29848 56994 29848 0 E2BEGb[6]
rlabel metal3 57106 30296 57106 30296 0 E2BEGb[7]
rlabel metal3 22232 26488 22232 26488 0 E2END[0]
rlabel metal2 16800 13720 16800 13720 0 E2END[1]
rlabel metal2 2520 21000 2520 21000 0 E2END[2]
rlabel metal2 21448 29232 21448 29232 0 E2END[3]
rlabel metal3 1358 28952 1358 28952 0 E2END[4]
rlabel metal2 3192 45192 3192 45192 0 E2END[5]
rlabel metal2 3696 38808 3696 38808 0 E2END[6]
rlabel metal2 16184 34608 16184 34608 0 E2END[7]
rlabel metal2 21336 19376 21336 19376 0 E2MID[0]
rlabel metal3 43568 5096 43568 5096 0 E2MID[1]
rlabel metal2 52136 25200 52136 25200 0 E2MID[2]
rlabel metal2 55944 23296 55944 23296 0 E2MID[3]
rlabel metal2 25704 2968 25704 2968 0 E2MID[4]
rlabel metal4 21896 26040 21896 26040 0 E2MID[5]
rlabel metal3 22120 42504 22120 42504 0 E2MID[6]
rlabel metal2 16520 26936 16520 26936 0 E2MID[7]
rlabel metal2 43512 40152 43512 40152 0 E6BEG[0]
rlabel metal4 38976 49770 38976 49770 0 E6BEG[10]
rlabel metal4 48776 33040 48776 33040 0 E6BEG[11]
rlabel metal2 56672 48104 56672 48104 0 E6BEG[1]
rlabel metal3 56658 38808 56658 38808 0 E6BEG[2]
rlabel metal4 45976 39144 45976 39144 0 E6BEG[3]
rlabel metal3 38752 35112 38752 35112 0 E6BEG[4]
rlabel metal3 55426 40152 55426 40152 0 E6BEG[5]
rlabel metal2 44520 37184 44520 37184 0 E6BEG[6]
rlabel metal2 49448 31640 49448 31640 0 E6BEG[7]
rlabel metal3 48888 33432 48888 33432 0 E6BEG[8]
rlabel metal2 49784 40320 49784 40320 0 E6BEG[9]
rlabel metal3 1078 37912 1078 37912 0 E6END[0]
rlabel metal3 1246 42392 1246 42392 0 E6END[10]
rlabel metal3 574 42840 574 42840 0 E6END[11]
rlabel metal3 182 38360 182 38360 0 E6END[1]
rlabel metal4 21000 43624 21000 43624 0 E6END[2]
rlabel metal3 24248 39312 24248 39312 0 E6END[3]
rlabel metal3 21000 39872 21000 39872 0 E6END[4]
rlabel metal3 910 40152 910 40152 0 E6END[5]
rlabel metal4 21000 41608 21000 41608 0 E6END[6]
rlabel metal3 910 41048 910 41048 0 E6END[7]
rlabel metal3 574 41496 574 41496 0 E6END[8]
rlabel metal3 910 41944 910 41944 0 E6END[9]
rlabel metal3 57330 30744 57330 30744 0 EE4BEG[0]
rlabel metal3 57330 35224 57330 35224 0 EE4BEG[10]
rlabel metal2 54264 49112 54264 49112 0 EE4BEG[11]
rlabel metal3 56938 36120 56938 36120 0 EE4BEG[12]
rlabel metal3 57162 36568 57162 36568 0 EE4BEG[13]
rlabel metal3 57330 37016 57330 37016 0 EE4BEG[14]
rlabel metal3 56322 37464 56322 37464 0 EE4BEG[15]
rlabel metal3 57162 31192 57162 31192 0 EE4BEG[1]
rlabel metal2 57232 41384 57232 41384 0 EE4BEG[2]
rlabel metal3 56728 47544 56728 47544 0 EE4BEG[3]
rlabel metal2 56504 47992 56504 47992 0 EE4BEG[4]
rlabel metal2 52304 32312 52304 32312 0 EE4BEG[5]
rlabel metal3 55818 33432 55818 33432 0 EE4BEG[6]
rlabel metal3 56056 39480 56056 39480 0 EE4BEG[7]
rlabel metal3 54586 34328 54586 34328 0 EE4BEG[8]
rlabel metal3 57274 34776 57274 34776 0 EE4BEG[9]
rlabel metal2 20216 16352 20216 16352 0 EE4END[0]
rlabel metal4 50344 25368 50344 25368 0 EE4END[10]
rlabel metal4 22456 35504 22456 35504 0 EE4END[11]
rlabel metal2 41384 35280 41384 35280 0 EE4END[12]
rlabel metal3 41384 35952 41384 35952 0 EE4END[13]
rlabel metal3 19208 38024 19208 38024 0 EE4END[14]
rlabel metal4 33656 36568 33656 36568 0 EE4END[15]
rlabel metal4 24248 17080 24248 17080 0 EE4END[1]
rlabel metal3 18424 31920 18424 31920 0 EE4END[2]
rlabel metal3 462 32088 462 32088 0 EE4END[3]
rlabel metal3 21336 31472 21336 31472 0 EE4END[4]
rlabel metal3 350 32984 350 32984 0 EE4END[5]
rlabel metal3 39088 26712 39088 26712 0 EE4END[6]
rlabel metal3 41160 34608 41160 34608 0 EE4END[7]
rlabel metal2 55384 23464 55384 23464 0 EE4END[8]
rlabel metal4 40152 34720 40152 34720 0 EE4END[9]
rlabel metal2 15232 23576 15232 23576 0 F
rlabel metal2 51016 25536 51016 25536 0 FrameData[0]
rlabel metal3 21000 42392 21000 42392 0 FrameData[10]
rlabel metal2 2296 2688 2296 2688 0 FrameData[11]
rlabel metal2 1624 47768 1624 47768 0 FrameData[12]
rlabel via3 26152 48104 26152 48104 0 FrameData[13]
rlabel metal3 54264 15176 54264 15176 0 FrameData[14]
rlabel metal3 52920 16296 52920 16296 0 FrameData[15]
rlabel metal2 54712 17864 54712 17864 0 FrameData[16]
rlabel metal2 26152 16408 26152 16408 0 FrameData[17]
rlabel metal2 52472 19880 52472 19880 0 FrameData[18]
rlabel metal2 53816 21504 53816 21504 0 FrameData[19]
rlabel metal2 54040 26488 54040 26488 0 FrameData[1]
rlabel metal2 52584 24248 52584 24248 0 FrameData[20]
rlabel metal2 50680 24640 50680 24640 0 FrameData[21]
rlabel metal2 51800 23968 51800 23968 0 FrameData[22]
rlabel metal2 3192 21000 3192 21000 0 FrameData[23]
rlabel metal3 54488 21784 54488 21784 0 FrameData[24]
rlabel via3 52024 18987 52024 18987 0 FrameData[25]
rlabel metal2 18424 22624 18424 22624 0 FrameData[26]
rlabel metal4 3192 18480 3192 18480 0 FrameData[27]
rlabel metal3 54544 19320 54544 19320 0 FrameData[28]
rlabel metal3 52304 21784 52304 21784 0 FrameData[29]
rlabel metal3 966 44184 966 44184 0 FrameData[2]
rlabel metal2 3304 2744 3304 2744 0 FrameData[30]
rlabel metal4 2408 46350 2408 46350 0 FrameData[31]
rlabel metal3 18536 40264 18536 40264 0 FrameData[3]
rlabel metal3 1190 45080 1190 45080 0 FrameData[4]
rlabel metal3 52976 24584 52976 24584 0 FrameData[5]
rlabel metal3 630 45976 630 45976 0 FrameData[6]
rlabel metal3 238 46424 238 46424 0 FrameData[7]
rlabel metal3 40768 2632 40768 2632 0 FrameData[8]
rlabel metal2 40992 1064 40992 1064 0 FrameData[9]
rlabel metal3 56434 43288 56434 43288 0 FrameData_O[0]
rlabel metal3 57218 47768 57218 47768 0 FrameData_O[10]
rlabel metal3 56826 48216 56826 48216 0 FrameData_O[11]
rlabel metal3 49224 40656 49224 40656 0 FrameData_O[12]
rlabel metal2 50288 52920 50288 52920 0 FrameData_O[13]
rlabel metal2 39032 42000 39032 42000 0 FrameData_O[14]
rlabel metal2 50008 50204 50008 50204 0 FrameData_O[15]
rlabel metal3 55986 50456 55986 50456 0 FrameData_O[16]
rlabel metal3 56378 50904 56378 50904 0 FrameData_O[17]
rlabel metal2 48776 52472 48776 52472 0 FrameData_O[18]
rlabel metal2 47544 52024 47544 52024 0 FrameData_O[19]
rlabel metal3 56392 24248 56392 24248 0 FrameData_O[1]
rlabel metal2 48552 53088 48552 53088 0 FrameData_O[20]
rlabel metal2 46872 52136 46872 52136 0 FrameData_O[21]
rlabel metal2 46200 53480 46200 53480 0 FrameData_O[22]
rlabel metal2 45528 53592 45528 53592 0 FrameData_O[23]
rlabel metal2 49000 54936 49000 54936 0 FrameData_O[24]
rlabel metal2 46648 51744 46648 51744 0 FrameData_O[25]
rlabel metal2 42168 54992 42168 54992 0 FrameData_O[26]
rlabel metal2 42000 49000 42000 49000 0 FrameData_O[27]
rlabel metal3 43680 49224 43680 49224 0 FrameData_O[28]
rlabel metal2 49224 54768 49224 54768 0 FrameData_O[29]
rlabel metal3 56770 44184 56770 44184 0 FrameData_O[2]
rlabel metal2 40432 50792 40432 50792 0 FrameData_O[30]
rlabel metal3 50400 48720 50400 48720 0 FrameData_O[31]
rlabel metal3 29008 45416 29008 45416 0 FrameData_O[3]
rlabel metal4 40040 45976 40040 45976 0 FrameData_O[4]
rlabel metal3 55594 45528 55594 45528 0 FrameData_O[5]
rlabel metal3 56378 45976 56378 45976 0 FrameData_O[6]
rlabel metal4 26488 53144 26488 53144 0 FrameData_O[7]
rlabel metal3 39704 48272 39704 48272 0 FrameData_O[8]
rlabel metal3 32536 49112 32536 49112 0 FrameData_O[9]
rlabel metal3 18088 16744 18088 16744 0 FrameStrobe[0]
rlabel metal2 52640 840 52640 840 0 FrameStrobe[10]
rlabel metal2 2744 2632 2744 2632 0 FrameStrobe[11]
rlabel metal2 30072 1680 30072 1680 0 FrameStrobe[12]
rlabel metal2 21616 48216 21616 48216 0 FrameStrobe[13]
rlabel metal2 54488 742 54488 742 0 FrameStrobe[14]
rlabel metal2 40880 42616 40880 42616 0 FrameStrobe[15]
rlabel metal2 55384 686 55384 686 0 FrameStrobe[16]
rlabel metal2 53928 22960 53928 22960 0 FrameStrobe[17]
rlabel metal2 50456 24864 50456 24864 0 FrameStrobe[18]
rlabel metal2 56896 2408 56896 2408 0 FrameStrobe[19]
rlabel metal2 48664 406 48664 406 0 FrameStrobe[1]
rlabel metal2 49056 1960 49056 1960 0 FrameStrobe[2]
rlabel metal2 49560 1582 49560 1582 0 FrameStrobe[3]
rlabel metal2 50008 350 50008 350 0 FrameStrobe[4]
rlabel metal3 51632 23016 51632 23016 0 FrameStrobe[5]
rlabel metal2 50904 574 50904 574 0 FrameStrobe[6]
rlabel metal2 26264 25088 26264 25088 0 FrameStrobe[7]
rlabel metal2 51800 406 51800 406 0 FrameStrobe[8]
rlabel metal2 52752 25480 52752 25480 0 FrameStrobe[9]
rlabel metal2 48216 56714 48216 56714 0 FrameStrobe_O[0]
rlabel metal2 47768 56056 47768 56056 0 FrameStrobe_O[10]
rlabel metal2 47096 56280 47096 56280 0 FrameStrobe_O[11]
rlabel metal3 47992 54992 47992 54992 0 FrameStrobe_O[12]
rlabel metal2 46200 56616 46200 56616 0 FrameStrobe_O[13]
rlabel metal2 44184 56168 44184 56168 0 FrameStrobe_O[14]
rlabel metal2 43512 56448 43512 56448 0 FrameStrobe_O[15]
rlabel metal2 55384 57330 55384 57330 0 FrameStrobe_O[16]
rlabel metal4 50120 53760 50120 53760 0 FrameStrobe_O[17]
rlabel metal2 40824 55720 40824 55720 0 FrameStrobe_O[18]
rlabel metal3 43624 48888 43624 48888 0 FrameStrobe_O[19]
rlabel metal2 48664 57050 48664 57050 0 FrameStrobe_O[1]
rlabel metal2 33992 53424 33992 53424 0 FrameStrobe_O[2]
rlabel metal2 49560 57106 49560 57106 0 FrameStrobe_O[3]
rlabel metal2 44184 49056 44184 49056 0 FrameStrobe_O[4]
rlabel metal2 32312 52976 32312 52976 0 FrameStrobe_O[5]
rlabel metal2 41832 55496 41832 55496 0 FrameStrobe_O[6]
rlabel metal2 52696 54936 52696 54936 0 FrameStrobe_O[7]
rlabel metal2 51912 54376 51912 54376 0 FrameStrobe_O[8]
rlabel metal2 49784 56224 49784 56224 0 FrameStrobe_O[9]
rlabel metal2 22904 15960 22904 15960 0 G
rlabel metal3 20328 25480 20328 25480 0 H
rlabel metal2 50960 17528 50960 17528 0 Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 48776 8792 48776 8792 0 Inst_LA_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal3 48496 15512 48496 15512 0 Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 49784 16800 49784 16800 0 Inst_LA_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal2 53592 12376 53592 12376 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal2 50960 12376 50960 12376 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal2 51184 9912 51184 9912 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 49560 8624 49560 8624 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal3 51240 12712 51240 12712 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 52808 11088 52808 11088 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal2 52472 11704 52472 11704 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal3 52136 11592 52136 11592 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 55048 9240 55048 9240 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 54488 9296 54488 9296 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 55160 5432 55160 5432 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 55888 4536 55888 4536 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 55272 5824 55272 5824 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal2 54544 4984 54544 4984 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 53256 6496 53256 6496 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal3 52136 6104 52136 6104 0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 51016 24360 51016 24360 0 Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 47992 13832 47992 13832 0 Inst_LB_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal2 51240 24808 51240 24808 0 Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal3 54152 23240 54152 23240 0 Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal2 52920 17080 52920 17080 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal3 53816 17080 53816 17080 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal2 52024 18707 52024 18707 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 56000 21560 56000 21560 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal2 54712 16296 54712 16296 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 55272 21280 55272 21280 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal3 52192 18648 52192 18648 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal3 51632 20216 51632 20216 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal3 52696 14728 52696 14728 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 55384 16576 55384 16576 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal3 51912 16072 51912 16072 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 55832 17976 55832 17976 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal3 51352 15512 51352 15512 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal3 53928 19320 53928 19320 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 55104 21336 55104 21336 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 52752 20888 52752 20888 0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 48776 26628 48776 26628 0 Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 49168 29176 49168 29176 0 Inst_LC_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal2 49000 26768 49000 26768 0 Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 48216 26096 48216 26096 0 Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal2 52472 26432 52472 26432 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal3 53928 28112 53928 28112 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal2 52864 31976 52864 31976 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 56112 31192 56112 31192 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal3 51240 30184 51240 30184 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 54880 30184 54880 30184 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal3 51688 30296 51688 30296 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal2 55384 31864 55384 31864 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 52136 25760 52136 25760 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 55272 26600 55272 26600 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 52080 26488 52080 26488 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 54656 23352 54656 23352 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal3 52920 27160 52920 27160 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal2 55048 23800 55048 23800 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 53816 31584 53816 31584 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 55496 30632 55496 30632 0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal3 48664 38248 48664 38248 0 Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 49952 32424 49952 32424 0 Inst_LD_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal2 48216 35952 48216 35952 0 Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 48272 39032 48272 39032 0 Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal3 50792 33936 50792 33936 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal2 55048 34048 55048 34048 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal2 53648 36456 53648 36456 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal3 52920 39368 52920 39368 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal2 55048 40264 55048 40264 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 55328 35896 55328 35896 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal2 54600 39984 54600 39984 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal2 53592 39984 53592 39984 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 52024 39592 52024 39592 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 50512 38248 50512 38248 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal3 51464 38808 51464 38808 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 50792 37464 50792 37464 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 50344 34552 50344 34552 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal2 54544 34328 54544 34328 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 54096 36680 54096 36680 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 54936 36064 54936 36064 0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 48888 50680 48888 50680 0 Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 50456 42639 50456 42639 0 Inst_LE_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal3 48272 50680 48272 50680 0 Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 52024 51632 52024 51632 0 Inst_LE_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal3 56112 43400 56112 43400 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal2 50120 45136 50120 45136 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal3 53592 46648 53592 46648 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 53480 47712 53480 47712 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal2 51352 47096 51352 47096 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 51296 47544 51296 47544 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal2 52416 46088 52416 46088 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal2 51968 47432 51968 47432 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal3 54208 42168 54208 42168 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 50904 45360 50904 45360 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 52640 51352 52640 51352 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 50904 47656 50904 47656 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 54040 43008 54040 43008 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal3 50568 45864 50568 45864 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 53872 45304 53872 45304 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 54432 47432 54432 47432 0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 46592 46424 46592 46424 0 Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal3 42168 41832 42168 41832 0 Inst_LF_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal3 48440 47432 48440 47432 0 Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 48776 48048 48776 48048 0 Inst_LF_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal2 42392 44576 42392 44576 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal3 46592 45304 46592 45304 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal3 43568 40488 43568 40488 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 45136 42952 45136 42952 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal3 49224 43400 49224 43400 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal3 48328 43512 48328 43512 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal3 43344 41384 43344 41384 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal3 45528 42840 45528 42840 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 43064 45192 43064 45192 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 43176 43456 43176 43456 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 42616 45528 42616 45528 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal2 43624 45416 43624 45416 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 42056 45080 42056 45080 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal3 45864 45640 45864 45640 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal2 47208 42280 47208 42280 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 46592 41160 46592 41160 0 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 41104 53480 41104 53480 0 Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal2 39144 45528 39144 45528 0 Inst_LG_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal2 42056 52808 42056 52808 0 Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal2 45304 53088 45304 53088 0 Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal2 40824 48888 40824 48888 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal3 39984 50568 39984 50568 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal3 32592 53144 32592 53144 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 39368 53200 39368 53200 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal2 34328 53200 34328 53200 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal2 37072 53032 37072 53032 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal2 33992 54880 33992 54880 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal2 38080 52920 38080 52920 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 39816 47544 39816 47544 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 38696 50848 38696 50848 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 37912 47880 37912 47880 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal3 36736 50680 36736 50680 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 38696 48496 38696 48496 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal3 36848 50008 36848 50008 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal3 31808 52136 31808 52136 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 39592 52640 39592 52640 0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 43176 50176 43176 50176 0 Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
rlabel metal3 42560 44408 42560 44408 0 Inst_LH_LUT4c_frame_config_dffesr.c_I0mux
rlabel metal2 42056 48160 42056 48160 0 Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
rlabel metal3 44520 50008 44520 50008 0 Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
rlabel metal3 35840 43624 35840 43624 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
rlabel metal3 32200 45640 32200 45640 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
rlabel metal2 34776 49812 34776 49812 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
rlabel metal2 31864 47712 31864 47712 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
rlabel metal2 31416 49448 31416 49448 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
rlabel metal3 31920 47656 31920 47656 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
rlabel metal2 34608 51576 34608 51576 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
rlabel metal3 31640 49784 31640 49784 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
rlabel metal2 34776 46368 34776 46368 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
rlabel metal2 32480 44072 32480 44072 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
rlabel metal2 37352 44688 37352 44688 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
rlabel metal3 31696 44520 31696 44520 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
rlabel metal2 35056 46872 35056 46872 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
rlabel metal3 32200 44296 32200 44296 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
rlabel metal3 32200 48776 32200 48776 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
rlabel metal2 29848 50064 29848 50064 0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
rlabel metal2 40712 13216 40712 13216 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 41720 12656 41720 12656 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 39592 33824 39592 33824 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 40824 34160 40824 34160 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 34216 13440 34216 13440 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 32760 13048 32760 13048 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 16856 15288 16856 15288 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 18592 14728 18592 14728 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 30016 17080 30016 17080 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 28392 16968 28392 16968 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 35168 34328 35168 34328 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 36400 34888 36400 34888 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 42168 29904 42168 29904 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 34216 32200 34216 32200 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 34888 32816 34888 32816 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 26992 39592 26992 39592 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 28056 39872 28056 39872 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 28672 11480 28672 11480 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 27216 11368 27216 11368 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 39424 26040 39424 26040 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 41888 25592 41888 25592 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 42336 26152 42336 26152 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 40600 20720 40600 20720 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 40600 30464 40600 30464 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 40880 19768 40880 19768 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 41608 21224 41608 21224 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 33880 23184 33880 23184 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
rlabel metal3 31640 23128 31640 23128 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q
rlabel metal3 15456 32536 15456 32536 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 16072 32144 16072 32144 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 41720 6384 41720 6384 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 40096 6664 40096 6664 0 Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 17192 22064 17192 22064 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
rlabel metal2 17136 26488 17136 26488 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
rlabel metal3 47152 22456 47152 22456 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q
rlabel metal2 47208 17976 47208 17976 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q
rlabel metal3 48104 11480 48104 11480 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q
rlabel metal2 47376 13160 47376 13160 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q
rlabel metal2 45360 19992 45360 19992 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q
rlabel metal2 46760 20664 46760 20664 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q
rlabel metal2 35448 15568 35448 15568 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
rlabel metal2 36680 13832 36680 13832 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q
rlabel metal2 43568 15176 43568 15176 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
rlabel metal2 46760 16184 46760 16184 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q
rlabel metal2 46536 8736 46536 8736 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q
rlabel metal2 51408 21448 51408 21448 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q
rlabel metal3 48664 20720 48664 20720 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q
rlabel metal2 47208 30408 47208 30408 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q
rlabel metal2 46760 29512 46760 29512 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
rlabel metal2 41832 31752 41832 31752 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q
rlabel metal2 42840 31472 42840 31472 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q
rlabel metal3 25424 31752 25424 31752 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
rlabel metal2 27944 31080 27944 31080 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q
rlabel metal2 44072 8680 44072 8680 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
rlabel metal2 43456 8232 43456 8232 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
rlabel metal2 48216 7840 48216 7840 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q
rlabel metal3 46816 26936 46816 26936 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
rlabel metal2 46704 26824 46704 26824 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q
rlabel metal2 44352 18648 44352 18648 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q
rlabel metal2 46648 18536 46648 18536 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q
rlabel metal2 22232 3136 22232 3136 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q
rlabel metal3 35392 2184 35392 2184 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q
rlabel metal2 43176 12264 43176 12264 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
rlabel metal2 45640 13384 45640 13384 0 Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q
rlabel metal2 38472 9128 38472 9128 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
rlabel metal3 38024 8344 38024 8344 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
rlabel metal3 2800 4536 2800 4536 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q
rlabel metal2 1176 4928 1176 4928 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
rlabel metal2 11368 2772 11368 2772 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
rlabel metal2 8792 1456 8792 1456 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q
rlabel metal2 10472 36736 10472 36736 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q
rlabel metal2 11704 35672 11704 35672 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
rlabel metal2 8232 33600 8232 33600 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q
rlabel metal2 17192 43568 17192 43568 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q
rlabel metal2 18312 42672 18312 42672 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
rlabel metal3 16744 41272 16744 41272 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q
rlabel metal3 39984 11480 39984 11480 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q
rlabel metal3 2856 20832 2856 20832 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
rlabel metal2 3584 20776 3584 20776 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
rlabel metal2 1176 17136 1176 17136 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q
rlabel metal2 15512 19208 15512 19208 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q
rlabel metal3 16464 19432 16464 19432 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
rlabel metal2 16856 21168 16856 21168 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q
rlabel metal2 5432 18200 5432 18200 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q
rlabel metal3 5432 18424 5432 18424 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
rlabel metal3 1624 15736 1624 15736 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q
rlabel metal2 3304 17696 3304 17696 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
rlabel metal3 26824 21560 26824 21560 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q
rlabel metal2 17080 25088 17080 25088 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q
rlabel metal2 17304 23408 17304 23408 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
rlabel metal2 29904 21560 29904 21560 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
rlabel metal2 30408 19880 30408 19880 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q
rlabel metal2 5600 1400 5600 1400 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q
rlabel metal2 2464 5096 2464 5096 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
rlabel metal3 11536 1176 11536 1176 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
rlabel metal2 2856 4088 2856 4088 0 Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q
rlabel metal2 29736 38360 29736 38360 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
rlabel metal2 30408 39312 30408 39312 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q
rlabel metal2 25032 12432 25032 12432 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q
rlabel metal3 23520 12152 23520 12152 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
rlabel metal2 23352 10752 23352 10752 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
rlabel metal2 23912 10304 23912 10304 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q
rlabel metal2 26152 14840 26152 14840 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q
rlabel metal2 24360 14000 24360 14000 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
rlabel metal3 23520 23128 23520 23128 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
rlabel metal2 25032 23184 25032 23184 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q
rlabel metal2 33656 15568 33656 15568 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
rlabel metal3 32032 15288 32032 15288 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q
rlabel metal2 20216 42056 20216 42056 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q
rlabel metal2 34608 21784 34608 21784 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
rlabel metal2 33208 22932 33208 22932 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q
rlabel metal2 38136 21840 38136 21840 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
rlabel metal2 37800 21280 37800 21280 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q
rlabel metal3 39872 12152 39872 12152 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q
rlabel metal2 39816 11424 39816 11424 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
rlabel metal2 34216 18872 34216 18872 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
rlabel metal3 31920 18424 31920 18424 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
rlabel metal2 34216 17136 34216 17136 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
rlabel metal2 31136 4312 31136 4312 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q
rlabel metal2 22120 39984 22120 39984 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
rlabel metal2 31808 2184 31808 2184 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
rlabel metal2 33096 1736 33096 1736 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q
rlabel metal2 20104 39928 20104 39928 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q
rlabel metal3 20720 41272 20720 41272 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
rlabel metal2 21112 46648 21112 46648 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q
rlabel metal2 22680 50288 22680 50288 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
rlabel metal3 22848 47544 22848 47544 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q
rlabel metal2 19432 45192 19432 45192 0 Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
rlabel metal2 14392 15232 14392 15232 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
rlabel metal2 13104 15288 13104 15288 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q
rlabel metal3 23856 31864 23856 31864 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q
rlabel metal3 25088 46872 25088 46872 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q
rlabel metal2 23352 47824 23352 47824 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
rlabel metal2 25816 50904 25816 50904 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q
rlabel metal2 43848 22680 43848 22680 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q
rlabel metal2 42896 21784 42896 21784 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
rlabel metal3 11760 22344 11760 22344 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
rlabel metal2 13272 22680 13272 22680 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q
rlabel metal2 40320 23576 40320 23576 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q
rlabel metal2 38696 24192 38696 24192 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
rlabel metal3 25424 37240 25424 37240 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
rlabel metal2 36792 24080 36792 24080 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
rlabel metal2 38136 24192 38136 24192 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q
rlabel metal3 13496 38248 13496 38248 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
rlabel metal2 15848 38976 15848 38976 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
rlabel metal2 15064 37912 15064 37912 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q
rlabel metal2 31304 41160 31304 41160 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q
rlabel metal2 32312 42224 32312 42224 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
rlabel metal2 30856 43008 30856 43008 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q
rlabel metal2 37016 33376 37016 33376 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
rlabel metal2 36792 32088 36792 32088 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
rlabel metal2 24584 37576 24584 37576 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
rlabel metal2 39256 31640 39256 31640 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
rlabel metal2 27888 40152 27888 40152 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q
rlabel metal2 19992 37744 19992 37744 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q
rlabel metal2 29456 51352 29456 51352 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q
rlabel metal2 30632 51632 30632 51632 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
rlabel metal2 30184 54208 30184 54208 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q
rlabel metal2 24584 31472 24584 31472 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
rlabel metal2 25704 30632 25704 30632 0 Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
rlabel metal2 11144 44044 11144 44044 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q
rlabel metal3 10752 44968 10752 44968 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q
rlabel metal2 2912 11592 2912 11592 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q
rlabel metal3 3696 17640 3696 17640 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
rlabel metal2 1176 40712 1176 40712 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
rlabel metal2 2968 37912 2968 37912 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q
rlabel metal2 2912 23352 2912 23352 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q
rlabel metal3 1344 19768 1344 19768 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
rlabel metal2 4312 24528 4312 24528 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
rlabel metal2 2856 21056 2856 21056 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q
rlabel metal2 13160 21672 13160 21672 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q
rlabel metal2 13888 21000 13888 21000 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
rlabel metal2 13272 33432 13272 33432 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q
rlabel metal2 14392 33712 14392 33712 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
rlabel metal3 13216 29624 13216 29624 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q
rlabel metal3 14224 30408 14224 30408 0 Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
rlabel metal2 5712 2968 5712 2968 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 4312 6496 4312 6496 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q
rlabel metal4 3304 45360 3304 45360 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 2856 45752 2856 45752 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 4760 46088 4760 46088 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 2856 49392 2856 49392 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 2856 37464 2856 37464 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 2856 36064 2856 36064 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 2856 33656 2856 33656 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 5544 33264 5544 33264 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 5768 52920 5768 52920 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 7672 53032 7672 53032 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 32424 31472 32424 31472 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 5544 52696 5544 52696 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 5992 52696 5992 52696 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 6776 23800 6776 23800 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 5432 22848 5432 22848 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 6832 23352 6832 23352 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q
rlabel metal3 7448 25592 7448 25592 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 20496 22344 20496 22344 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 20048 21784 20048 21784 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 32704 20216 32704 20216 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 33880 20664 33880 20664 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 32760 30464 32760 30464 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 34608 10360 34608 10360 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 35840 11368 35840 11368 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 35560 29400 35560 29400 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 33096 28448 33096 28448 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 16520 6608 16520 6608 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 15400 3164 15400 3164 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 16240 2072 16240 2072 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 16688 2856 16688 2856 0 Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 34888 5824 34888 5824 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q
rlabel metal3 35112 6104 35112 6104 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 15624 49000 15624 49000 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 16632 47040 16632 47040 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 16800 50344 16800 50344 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 16296 43400 16296 43400 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 8792 32368 8792 32368 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 9240 33040 9240 33040 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 8512 30184 8512 30184 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 9016 29848 9016 29848 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 23464 51072 23464 51072 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 25256 52192 25256 52192 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 17192 30576 17192 30576 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 23128 53200 23128 53200 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 25032 53984 25032 53984 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 3920 27832 3920 27832 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 4536 27048 4536 27048 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 3528 27328 3528 27328 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 3304 29064 3304 29064 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 3024 7672 3024 7672 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 3248 8008 3248 8008 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
rlabel metal3 840 7224 840 7224 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 3080 7448 3080 7448 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19992 30968 19992 30968 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 5488 2072 5488 2072 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 8120 5656 8120 5656 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 17472 28840 17472 28840 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q
rlabel metal3 20160 27832 20160 27832 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
rlabel metal3 20440 7448 20440 7448 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 20048 8232 20048 8232 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 19320 5600 19320 5600 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 21784 4200 21784 4200 0 Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 25592 6664 25592 6664 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 27608 3304 27608 3304 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q
rlabel metal3 10192 49000 10192 49000 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 10584 47880 10584 47880 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 9128 45864 9128 45864 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 8680 46592 8680 46592 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 9408 41160 9408 41160 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
rlabel metal3 9464 41272 9464 41272 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 8512 39816 8512 39816 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 7896 39144 7896 39144 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 17192 51408 17192 51408 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 18536 53312 18536 53312 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 21000 25536 21000 25536 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
rlabel metal3 16576 52136 16576 52136 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 15624 54040 15624 54040 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 12936 24808 12936 24808 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 11704 25704 11704 25704 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 11928 29064 11928 29064 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 11256 28672 11256 28672 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 6832 9240 6832 9240 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 7000 10024 7000 10024 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 5712 5320 5712 5320 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 7896 8960 7896 8960 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 22792 26096 22792 26096 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 32424 8680 32424 8680 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 32872 7728 32872 7728 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 20888 26320 20888 26320 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 21336 23856 21336 23856 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 19544 11536 19544 11536 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 21112 13216 21112 13216 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 21000 12600 21000 12600 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 19656 11704 19656 11704 0 Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 13160 5712 13160 5712 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 13608 2408 13608 2408 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 2968 49168 2968 49168 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
rlabel metal3 2576 48216 2576 48216 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
rlabel metal3 18536 42616 18536 42616 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 2856 54096 2856 54096 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q
rlabel via2 2856 41048 2856 41048 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 2632 41440 2632 41440 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 3080 43176 3080 43176 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 3192 42840 3192 42840 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 13104 51352 13104 51352 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 11816 51352 11816 51352 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 21112 34104 21112 34104 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 9856 52696 9856 52696 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 11144 52416 11144 52416 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 2856 32032 2856 32032 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
rlabel metal4 4312 32312 4312 32312 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 3248 32424 3248 32424 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q
rlabel metal3 4928 29400 4928 29400 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 10584 13048 10584 13048 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 9352 11872 9352 11872 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
rlabel metal3 12544 9912 12544 9912 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 9632 9912 9632 9912 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 20272 38136 20272 38136 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
rlabel metal3 24640 5880 24640 5880 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 26152 7896 26152 7896 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
rlabel metal3 19656 33992 19656 33992 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 18984 33768 18984 33768 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 16744 10696 16744 10696 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
rlabel metal3 15736 9016 15736 9016 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
rlabel metal3 14392 10808 14392 10808 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 16744 12292 16744 12292 0 Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 27048 22848 27048 22848 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
rlabel metal3 24920 23912 24920 23912 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 32536 35392 32536 35392 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 33768 35840 33768 35840 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 31304 34776 31304 34776 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 26824 34384 26824 34384 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 16184 43008 16184 43008 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q
rlabel metal3 13496 41944 13496 41944 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q
rlabel metal3 15400 13160 15400 13160 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 16296 14000 16296 14000 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 14504 35000 14504 35000 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 15512 34776 15512 34776 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 30184 30800 30184 30800 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 26040 34832 26040 34832 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
rlabel metal3 24584 36008 24584 36008 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 15176 41832 15176 41832 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 13888 40376 13888 40376 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 13888 17416 13888 17416 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 17080 17864 17080 17864 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 10752 17416 10752 17416 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
rlabel metal3 10304 18424 10304 18424 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 11032 19488 11032 19488 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q
rlabel metal3 11032 20888 11032 20888 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
rlabel metal3 29288 30184 29288 30184 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 10640 2968 10640 2968 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
rlabel metal3 11368 5096 11368 5096 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
rlabel metal3 23856 27832 23856 27832 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 25592 28504 25592 28504 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
rlabel metal3 18424 17640 18424 17640 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q
rlabel metal3 18648 17080 18648 17080 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 31248 10024 31248 10024 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 29064 10192 29064 10192 0 Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 42168 3976 42168 3976 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 43064 5376 43064 5376 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 38864 28840 38864 28840 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q
rlabel metal3 39480 27272 39480 27272 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 36344 25928 36344 25928 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 36008 25144 36008 25144 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 26824 44184 26824 44184 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 26488 43568 26488 43568 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 41272 14784 41272 14784 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 43120 15848 43120 15848 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 37240 29680 37240 29680 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 38360 29120 38360 29120 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 43400 28336 43400 28336 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q
rlabel metal3 28448 26264 28448 26264 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 30408 25984 30408 25984 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 28392 43008 28392 43008 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 29624 42224 29624 42224 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 37912 15680 37912 15680 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 39144 14616 39144 14616 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q
rlabel metal3 30016 28616 30016 28616 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
rlabel metal3 28000 28728 28000 28728 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q
rlabel metal3 28112 19208 28112 19208 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
rlabel metal3 26880 19208 26880 19208 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 44296 28896 44296 28896 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
rlabel metal3 22176 15512 22176 15512 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
rlabel metal3 20160 16072 20160 16072 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 25592 25984 25592 25984 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 28000 27048 28000 27048 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 27720 36344 27720 36344 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 28728 35224 28728 35224 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
rlabel metal3 40376 2968 40376 2968 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 42280 2184 42280 2184 0 Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 28840 13832 28840 13832 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 30520 14224 30520 14224 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 42616 37856 42616 37856 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q
rlabel metal3 42952 35896 42952 35896 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 44128 39032 44128 39032 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 45920 38584 45920 38584 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 24696 18984 24696 18984 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 22456 19208 22456 19208 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q
rlabel metal3 23744 16856 23744 16856 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
rlabel metal3 24976 16856 24976 16856 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q
rlabel metal3 36736 40264 36736 40264 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 35448 40600 35448 40600 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
rlabel metal3 43792 35112 43792 35112 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 36680 37184 36680 37184 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q
rlabel metal3 35168 36456 35168 36456 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q
rlabel metal3 25032 20776 25032 20776 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 22680 20328 22680 20328 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 19992 18144 19992 18144 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
rlabel metal3 20104 19320 20104 19320 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 44408 26656 44408 26656 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 44632 25200 44632 25200 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
rlabel metal3 34440 25480 34440 25480 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 34104 25536 34104 25536 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
rlabel metal3 46648 34776 46648 34776 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
rlabel metal3 28280 22568 28280 22568 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q
rlabel metal3 28896 24584 28896 24584 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
rlabel metal3 45640 32760 45640 32760 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 44128 33320 44128 33320 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 23800 3304 23800 3304 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 23912 2240 23912 2240 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q
rlabel metal3 28112 3752 28112 3752 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 30296 3024 30296 3024 0 Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 32536 39004 32536 39004 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
rlabel metal3 34384 39704 34384 39704 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q
rlabel metal2 32984 38304 32984 38304 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 34104 38360 34104 38360 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 27272 46928 27272 46928 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
rlabel metal3 28056 47544 28056 47544 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 36680 18704 36680 18704 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 38024 18704 38024 18704 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 44520 49952 44520 49952 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
rlabel metal3 41552 50792 41552 50792 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 15736 45360 15736 45360 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 14504 45136 14504 45136 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 25592 45360 25592 45360 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 7784 38472 7784 38472 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 10472 35896 10472 35896 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q
rlabel metal3 18368 47432 18368 47432 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
rlabel metal3 18256 46088 18256 46088 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q
rlabel metal3 10080 26152 10080 26152 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 9184 28616 9184 28616 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 42560 10024 42560 10024 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 43512 10920 43512 10920 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 48328 23408 48328 23408 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 47096 22456 47096 22456 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q
rlabel metal3 28168 44296 28168 44296 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 20776 2576 20776 2576 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
rlabel metal3 20384 2744 20384 2744 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 36680 16968 36680 16968 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 38080 17080 38080 17080 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 28728 50680 28728 50680 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 42280 53032 42280 53032 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 35560 43568 35560 43568 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q
rlabel metal2 39592 43176 39592 43176 0 Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q
rlabel metal3 45584 31528 45584 31528 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q
rlabel metal2 48552 31640 48552 31640 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
rlabel metal2 39088 38584 39088 38584 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q
rlabel metal2 40376 37520 40376 37520 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q
rlabel metal2 40600 40264 40600 40264 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
rlabel metal2 41944 40264 41944 40264 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q
rlabel metal2 21672 44800 21672 44800 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
rlabel metal2 23744 44408 23744 44408 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
rlabel metal2 40376 17360 40376 17360 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
rlabel metal3 42280 17080 42280 17080 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q
rlabel metal2 50680 53592 50680 53592 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q
rlabel metal2 48216 52416 48216 52416 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q
rlabel metal2 40712 33488 40712 33488 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q
rlabel metal2 39144 39368 39144 39368 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q
rlabel metal2 40600 36176 40600 36176 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q
rlabel metal3 39200 40376 39200 40376 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 40824 41048 40824 41048 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 24584 43960 24584 43960 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
rlabel metal3 25032 43400 25032 43400 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
rlabel metal3 42616 19432 42616 19432 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 43288 18928 43288 18928 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 47880 50064 47880 50064 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q
rlabel metal3 47936 49784 47936 49784 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q
rlabel metal2 41776 32536 41776 32536 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q
rlabel metal2 34552 41888 34552 41888 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 40936 43344 40936 43344 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q
rlabel metal2 27104 33320 27104 33320 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
rlabel metal2 28000 33432 28000 33432 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q
rlabel metal2 45080 5488 45080 5488 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
rlabel metal2 45976 9072 45976 9072 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q
rlabel metal3 47824 39704 47824 39704 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
rlabel metal2 46200 39872 46200 39872 0 Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q
rlabel metal2 47544 21224 47544 21224 0 Inst_LUT4AB_switch_matrix.E1BEG0
rlabel metal2 53704 18144 53704 18144 0 Inst_LUT4AB_switch_matrix.E1BEG1
rlabel metal3 43232 22904 43232 22904 0 Inst_LUT4AB_switch_matrix.E1BEG2
rlabel metal2 50008 22064 50008 22064 0 Inst_LUT4AB_switch_matrix.E1BEG3
rlabel metal3 22904 10472 22904 10472 0 Inst_LUT4AB_switch_matrix.E2BEG0
rlabel metal4 41160 19320 41160 19320 0 Inst_LUT4AB_switch_matrix.E2BEG1
rlabel metal3 41272 22456 41272 22456 0 Inst_LUT4AB_switch_matrix.E2BEG2
rlabel metal3 52248 17920 52248 17920 0 Inst_LUT4AB_switch_matrix.E2BEG3
rlabel metal2 55944 25928 55944 25928 0 Inst_LUT4AB_switch_matrix.E2BEG4
rlabel metal3 28392 41104 28392 41104 0 Inst_LUT4AB_switch_matrix.E2BEG5
rlabel metal2 52584 25928 52584 25928 0 Inst_LUT4AB_switch_matrix.E2BEG6
rlabel metal2 55944 19712 55944 19712 0 Inst_LUT4AB_switch_matrix.E2BEG7
rlabel metal2 21672 40936 21672 40936 0 Inst_LUT4AB_switch_matrix.E6BEG0
rlabel metal2 20328 46424 20328 46424 0 Inst_LUT4AB_switch_matrix.E6BEG1
rlabel metal4 49336 38024 49336 38024 0 Inst_LUT4AB_switch_matrix.EE4BEG0
rlabel metal2 31696 42504 31696 42504 0 Inst_LUT4AB_switch_matrix.EE4BEG1
rlabel metal2 54880 48216 54880 48216 0 Inst_LUT4AB_switch_matrix.EE4BEG2
rlabel metal3 44520 39312 44520 39312 0 Inst_LUT4AB_switch_matrix.EE4BEG3
rlabel metal2 11816 22512 11816 22512 0 Inst_LUT4AB_switch_matrix.JN2BEG0
rlabel metal3 40656 27608 40656 27608 0 Inst_LUT4AB_switch_matrix.JN2BEG1
rlabel metal3 40936 23576 40936 23576 0 Inst_LUT4AB_switch_matrix.JN2BEG2
rlabel metal2 44184 22456 44184 22456 0 Inst_LUT4AB_switch_matrix.JN2BEG3
rlabel metal2 17080 44912 17080 44912 0 Inst_LUT4AB_switch_matrix.JN2BEG4
rlabel metal2 41944 36120 41944 36120 0 Inst_LUT4AB_switch_matrix.JN2BEG5
rlabel metal4 17192 45248 17192 45248 0 Inst_LUT4AB_switch_matrix.JN2BEG6
rlabel metal3 20496 40936 20496 40936 0 Inst_LUT4AB_switch_matrix.JN2BEG7
rlabel metal2 2240 2184 2240 2184 0 Inst_LUT4AB_switch_matrix.JS2BEG0
rlabel metal2 25256 5824 25256 5824 0 Inst_LUT4AB_switch_matrix.JS2BEG1
rlabel metal2 24920 2240 24920 2240 0 Inst_LUT4AB_switch_matrix.JS2BEG2
rlabel metal2 26488 3752 26488 3752 0 Inst_LUT4AB_switch_matrix.JS2BEG3
rlabel metal2 24248 2800 24248 2800 0 Inst_LUT4AB_switch_matrix.JS2BEG4
rlabel metal2 18984 28728 18984 28728 0 Inst_LUT4AB_switch_matrix.JS2BEG5
rlabel metal3 26600 2744 26600 2744 0 Inst_LUT4AB_switch_matrix.JS2BEG6
rlabel metal2 5096 5768 5096 5768 0 Inst_LUT4AB_switch_matrix.JS2BEG7
rlabel metal3 4312 37128 4312 37128 0 Inst_LUT4AB_switch_matrix.JW2BEG0
rlabel metal2 30296 2016 30296 2016 0 Inst_LUT4AB_switch_matrix.JW2BEG1
rlabel metal3 23688 22008 23688 22008 0 Inst_LUT4AB_switch_matrix.JW2BEG2
rlabel metal2 15960 6440 15960 6440 0 Inst_LUT4AB_switch_matrix.JW2BEG3
rlabel metal2 25480 11032 25480 11032 0 Inst_LUT4AB_switch_matrix.JW2BEG4
rlabel metal3 2072 1176 2072 1176 0 Inst_LUT4AB_switch_matrix.JW2BEG5
rlabel metal3 1064 16688 1064 16688 0 Inst_LUT4AB_switch_matrix.JW2BEG6
rlabel metal3 6160 22904 6160 22904 0 Inst_LUT4AB_switch_matrix.JW2BEG7
rlabel metal2 19824 42840 19824 42840 0 Inst_LUT4AB_switch_matrix.M_AB
rlabel metal3 19992 48888 19992 48888 0 Inst_LUT4AB_switch_matrix.M_AD
rlabel metal2 20552 42672 20552 42672 0 Inst_LUT4AB_switch_matrix.M_AH
rlabel metal3 17584 23912 17584 23912 0 Inst_LUT4AB_switch_matrix.M_EF
rlabel metal3 1288 31864 1288 31864 0 Inst_LUT4AB_switch_matrix.N1BEG0
rlabel metal2 3080 39480 3080 39480 0 Inst_LUT4AB_switch_matrix.N1BEG1
rlabel metal4 15848 29736 15848 29736 0 Inst_LUT4AB_switch_matrix.N1BEG2
rlabel metal3 5712 40936 5712 40936 0 Inst_LUT4AB_switch_matrix.N1BEG3
rlabel metal2 13832 21560 13832 21560 0 Inst_LUT4AB_switch_matrix.N4BEG0
rlabel metal3 12936 45192 12936 45192 0 Inst_LUT4AB_switch_matrix.N4BEG1
rlabel metal2 14168 30912 14168 30912 0 Inst_LUT4AB_switch_matrix.N4BEG2
rlabel metal3 14168 16408 14168 16408 0 Inst_LUT4AB_switch_matrix.N4BEG3
rlabel metal2 22848 40152 22848 40152 0 Inst_LUT4AB_switch_matrix.NN4BEG0
rlabel metal3 28896 54712 28896 54712 0 Inst_LUT4AB_switch_matrix.NN4BEG1
rlabel metal3 24136 31640 24136 31640 0 Inst_LUT4AB_switch_matrix.NN4BEG2
rlabel metal3 25984 49224 25984 49224 0 Inst_LUT4AB_switch_matrix.NN4BEG3
rlabel metal2 24472 11928 24472 11928 0 Inst_LUT4AB_switch_matrix.S1BEG0
rlabel metal2 23016 7280 23016 7280 0 Inst_LUT4AB_switch_matrix.S1BEG1
rlabel metal2 25704 14560 25704 14560 0 Inst_LUT4AB_switch_matrix.S1BEG2
rlabel metal2 25312 17304 25312 17304 0 Inst_LUT4AB_switch_matrix.S1BEG3
rlabel metal2 37688 2856 37688 2856 0 Inst_LUT4AB_switch_matrix.S4BEG0
rlabel metal3 38360 3304 38360 3304 0 Inst_LUT4AB_switch_matrix.S4BEG1
rlabel metal2 38528 2184 38528 2184 0 Inst_LUT4AB_switch_matrix.S4BEG2
rlabel metal3 39480 2744 39480 2744 0 Inst_LUT4AB_switch_matrix.S4BEG3
rlabel metal3 44576 2744 44576 2744 0 Inst_LUT4AB_switch_matrix.SS4BEG0
rlabel metal4 44296 3696 44296 3696 0 Inst_LUT4AB_switch_matrix.SS4BEG1
rlabel metal2 39816 5936 39816 5936 0 Inst_LUT4AB_switch_matrix.SS4BEG2
rlabel metal3 39032 2856 39032 2856 0 Inst_LUT4AB_switch_matrix.SS4BEG3
rlabel metal2 2968 5096 2968 5096 0 Inst_LUT4AB_switch_matrix.W1BEG0
rlabel metal2 17080 2772 17080 2772 0 Inst_LUT4AB_switch_matrix.W1BEG1
rlabel metal2 12040 3052 12040 3052 0 Inst_LUT4AB_switch_matrix.W1BEG2
rlabel metal3 10248 2744 10248 2744 0 Inst_LUT4AB_switch_matrix.W1BEG3
rlabel metal2 2072 18648 2072 18648 0 Inst_LUT4AB_switch_matrix.W6BEG0
rlabel metal2 2072 20944 2072 20944 0 Inst_LUT4AB_switch_matrix.W6BEG1
rlabel metal3 5936 33320 5936 33320 0 Inst_LUT4AB_switch_matrix.WW4BEG0
rlabel metal3 16240 33768 16240 33768 0 Inst_LUT4AB_switch_matrix.WW4BEG1
rlabel metal2 2184 20608 2184 20608 0 Inst_LUT4AB_switch_matrix.WW4BEG2
rlabel metal2 4984 15568 4984 15568 0 Inst_LUT4AB_switch_matrix.WW4BEG3
rlabel metal2 728 57050 728 57050 0 N1BEG[0]
rlabel metal2 1176 56546 1176 56546 0 N1BEG[1]
rlabel metal2 1624 57218 1624 57218 0 N1BEG[2]
rlabel metal2 2072 55538 2072 55538 0 N1BEG[3]
rlabel metal2 672 2632 672 2632 0 N1END[0]
rlabel metal2 1176 798 1176 798 0 N1END[1]
rlabel metal2 1624 798 1624 798 0 N1END[2]
rlabel metal2 2072 350 2072 350 0 N1END[3]
rlabel metal2 2520 55874 2520 55874 0 N2BEG[0]
rlabel metal2 2968 56714 2968 56714 0 N2BEG[1]
rlabel metal3 2128 49784 2128 49784 0 N2BEG[2]
rlabel metal2 3864 56994 3864 56994 0 N2BEG[3]
rlabel metal3 1064 50568 1064 50568 0 N2BEG[4]
rlabel metal2 2240 49224 2240 49224 0 N2BEG[5]
rlabel metal2 3864 52752 3864 52752 0 N2BEG[6]
rlabel metal2 2240 53928 2240 53928 0 N2BEG[7]
rlabel metal3 2072 33544 2072 33544 0 N2BEGb[0]
rlabel metal2 12824 40712 12824 40712 0 N2BEGb[1]
rlabel metal2 8904 36456 8904 36456 0 N2BEGb[2]
rlabel metal2 3752 52920 3752 52920 0 N2BEGb[3]
rlabel metal2 13160 42896 13160 42896 0 N2BEGb[4]
rlabel metal2 12544 41384 12544 41384 0 N2BEGb[5]
rlabel metal2 8064 36568 8064 36568 0 N2BEGb[6]
rlabel metal2 1512 54992 1512 54992 0 N2BEGb[7]
rlabel metal2 2408 29400 2408 29400 0 N2END[0]
rlabel metal2 6552 2030 6552 2030 0 N2END[1]
rlabel metal2 26824 21224 26824 21224 0 N2END[2]
rlabel metal2 22680 33432 22680 33432 0 N2END[3]
rlabel metal3 17976 15232 17976 15232 0 N2END[4]
rlabel metal2 8344 854 8344 854 0 N2END[5]
rlabel metal3 21000 29400 21000 29400 0 N2END[6]
rlabel metal3 16296 49112 16296 49112 0 N2END[7]
rlabel metal2 2520 350 2520 350 0 N2MID[0]
rlabel metal2 2968 742 2968 742 0 N2MID[1]
rlabel metal4 20104 43288 20104 43288 0 N2MID[2]
rlabel metal2 3864 742 3864 742 0 N2MID[3]
rlabel metal2 26488 2800 26488 2800 0 N2MID[4]
rlabel metal4 16184 30688 16184 30688 0 N2MID[5]
rlabel metal4 1624 48870 1624 48870 0 N2MID[6]
rlabel metal2 25144 27048 25144 27048 0 N2MID[7]
rlabel metal3 7896 36680 7896 36680 0 N4BEG[0]
rlabel metal2 5712 55832 5712 55832 0 N4BEG[10]
rlabel metal2 6328 56000 6328 56000 0 N4BEG[11]
rlabel metal3 9128 55832 9128 55832 0 N4BEG[12]
rlabel metal2 15512 56882 15512 56882 0 N4BEG[13]
rlabel metal2 16184 54432 16184 54432 0 N4BEG[14]
rlabel metal2 16408 56154 16408 56154 0 N4BEG[15]
rlabel metal2 2184 55776 2184 55776 0 N4BEG[1]
rlabel metal2 23352 53704 23352 53704 0 N4BEG[2]
rlabel metal3 17528 54544 17528 54544 0 N4BEG[3]
rlabel metal2 3024 55832 3024 55832 0 N4BEG[4]
rlabel metal2 24920 56392 24920 56392 0 N4BEG[5]
rlabel metal2 2296 56056 2296 56056 0 N4BEG[6]
rlabel metal2 7336 54040 7336 54040 0 N4BEG[7]
rlabel metal2 3696 55944 3696 55944 0 N4BEG[8]
rlabel metal2 4312 55328 4312 55328 0 N4BEG[9]
rlabel metal3 17304 14840 17304 14840 0 N4END[0]
rlabel metal2 14168 518 14168 518 0 N4END[10]
rlabel metal2 14616 854 14616 854 0 N4END[11]
rlabel metal2 15064 854 15064 854 0 N4END[12]
rlabel metal2 15512 406 15512 406 0 N4END[13]
rlabel metal2 15960 854 15960 854 0 N4END[14]
rlabel metal2 16408 854 16408 854 0 N4END[15]
rlabel metal2 19880 15512 19880 15512 0 N4END[1]
rlabel metal2 24696 7616 24696 7616 0 N4END[2]
rlabel metal2 15176 25956 15176 25956 0 N4END[3]
rlabel metal2 11480 854 11480 854 0 N4END[4]
rlabel metal2 11928 406 11928 406 0 N4END[5]
rlabel metal2 12376 854 12376 854 0 N4END[6]
rlabel metal3 8176 55272 8176 55272 0 N4END[7]
rlabel metal2 13272 854 13272 854 0 N4END[8]
rlabel metal2 13720 462 13720 462 0 N4END[9]
rlabel metal2 16856 56882 16856 56882 0 NN4BEG[0]
rlabel metal2 20944 53928 20944 53928 0 NN4BEG[10]
rlabel metal2 19208 55496 19208 55496 0 NN4BEG[11]
rlabel metal2 18872 56336 18872 56336 0 NN4BEG[12]
rlabel metal3 21056 55832 21056 55832 0 NN4BEG[13]
rlabel metal3 22904 55944 22904 55944 0 NN4BEG[14]
rlabel metal2 23352 56336 23352 56336 0 NN4BEG[15]
rlabel metal2 16408 54488 16408 54488 0 NN4BEG[1]
rlabel metal2 17752 56938 17752 56938 0 NN4BEG[2]
rlabel metal2 18200 56994 18200 56994 0 NN4BEG[3]
rlabel metal2 18648 57050 18648 57050 0 NN4BEG[4]
rlabel metal3 17976 55944 17976 55944 0 NN4BEG[5]
rlabel metal2 17864 55328 17864 55328 0 NN4BEG[6]
rlabel metal3 20216 55944 20216 55944 0 NN4BEG[7]
rlabel metal2 18592 55384 18592 55384 0 NN4BEG[8]
rlabel metal2 18200 56000 18200 56000 0 NN4BEG[9]
rlabel metal2 16856 854 16856 854 0 NN4END[0]
rlabel metal2 21336 406 21336 406 0 NN4END[10]
rlabel metal2 21784 854 21784 854 0 NN4END[11]
rlabel metal2 22232 910 22232 910 0 NN4END[12]
rlabel metal2 22680 406 22680 406 0 NN4END[13]
rlabel metal2 23128 518 23128 518 0 NN4END[14]
rlabel metal2 23576 854 23576 854 0 NN4END[15]
rlabel metal2 17304 854 17304 854 0 NN4END[1]
rlabel metal2 17752 910 17752 910 0 NN4END[2]
rlabel metal2 18200 854 18200 854 0 NN4END[3]
rlabel metal2 14504 54208 14504 54208 0 NN4END[4]
rlabel metal2 19096 238 19096 238 0 NN4END[5]
rlabel metal2 19544 742 19544 742 0 NN4END[6]
rlabel metal2 19992 910 19992 910 0 NN4END[7]
rlabel metal2 20440 854 20440 854 0 NN4END[8]
rlabel metal2 20888 798 20888 798 0 NN4END[9]
rlabel metal2 24472 182 24472 182 0 S1BEG[0]
rlabel metal2 24920 294 24920 294 0 S1BEG[1]
rlabel metal2 25368 350 25368 350 0 S1BEG[2]
rlabel metal2 25816 294 25816 294 0 S1BEG[3]
rlabel metal2 16072 42000 16072 42000 0 S1END[0]
rlabel metal2 18200 46536 18200 46536 0 S1END[1]
rlabel metal2 16296 43176 16296 43176 0 S1END[2]
rlabel metal2 19096 43792 19096 43792 0 S1END[3]
rlabel metal2 26264 238 26264 238 0 S2BEG[0]
rlabel metal2 26712 518 26712 518 0 S2BEG[1]
rlabel metal2 27160 294 27160 294 0 S2BEG[2]
rlabel metal2 27608 294 27608 294 0 S2BEG[3]
rlabel metal2 28056 406 28056 406 0 S2BEG[4]
rlabel metal2 28504 182 28504 182 0 S2BEG[5]
rlabel metal2 28952 518 28952 518 0 S2BEG[6]
rlabel metal2 29400 294 29400 294 0 S2BEG[7]
rlabel metal2 29848 1078 29848 1078 0 S2BEGb[0]
rlabel metal2 30296 182 30296 182 0 S2BEGb[1]
rlabel metal2 30744 406 30744 406 0 S2BEGb[2]
rlabel metal2 31192 910 31192 910 0 S2BEGb[3]
rlabel metal2 31640 854 31640 854 0 S2BEGb[4]
rlabel metal2 32088 294 32088 294 0 S2BEGb[5]
rlabel metal2 32536 126 32536 126 0 S2BEGb[6]
rlabel metal2 32984 1078 32984 1078 0 S2BEGb[7]
rlabel metal3 21000 24528 21000 24528 0 S2END[0]
rlabel metal4 17192 16352 17192 16352 0 S2END[1]
rlabel metal4 15624 6216 15624 6216 0 S2END[2]
rlabel metal2 22792 35952 22792 35952 0 S2END[3]
rlabel metal2 22456 16464 22456 16464 0 S2END[4]
rlabel metal2 17304 46760 17304 46760 0 S2END[5]
rlabel metal4 25928 32368 25928 32368 0 S2END[6]
rlabel metal2 15736 53368 15736 53368 0 S2END[7]
rlabel metal2 26264 56434 26264 56434 0 S2MID[0]
rlabel metal3 30632 1176 30632 1176 0 S2MID[1]
rlabel metal2 28728 1232 28728 1232 0 S2MID[2]
rlabel metal2 31360 23016 31360 23016 0 S2MID[3]
rlabel metal3 27888 3080 27888 3080 0 S2MID[4]
rlabel metal2 28448 21224 28448 21224 0 S2MID[5]
rlabel metal3 34272 2744 34272 2744 0 S2MID[6]
rlabel metal3 30352 44184 30352 44184 0 S2MID[7]
rlabel metal2 33432 462 33432 462 0 S4BEG[0]
rlabel metal2 37912 630 37912 630 0 S4BEG[10]
rlabel metal2 38360 406 38360 406 0 S4BEG[11]
rlabel metal2 38808 742 38808 742 0 S4BEG[12]
rlabel metal2 39256 238 39256 238 0 S4BEG[13]
rlabel metal2 39704 1862 39704 1862 0 S4BEG[14]
rlabel metal2 40152 294 40152 294 0 S4BEG[15]
rlabel metal2 33880 966 33880 966 0 S4BEG[1]
rlabel metal2 34328 182 34328 182 0 S4BEG[2]
rlabel metal2 34776 238 34776 238 0 S4BEG[3]
rlabel metal2 35224 1078 35224 1078 0 S4BEG[4]
rlabel metal2 35672 406 35672 406 0 S4BEG[5]
rlabel metal2 36120 1078 36120 1078 0 S4BEG[6]
rlabel metal2 36568 294 36568 294 0 S4BEG[7]
rlabel metal2 37016 406 37016 406 0 S4BEG[8]
rlabel metal2 37464 518 37464 518 0 S4BEG[9]
rlabel metal2 22904 6832 22904 6832 0 S4END[0]
rlabel metal2 37744 56056 37744 56056 0 S4END[10]
rlabel metal2 38472 55496 38472 55496 0 S4END[11]
rlabel metal2 38808 57050 38808 57050 0 S4END[12]
rlabel metal2 39256 56434 39256 56434 0 S4END[13]
rlabel metal2 39480 56336 39480 56336 0 S4END[14]
rlabel metal2 40152 56434 40152 56434 0 S4END[15]
rlabel metal3 20328 39480 20328 39480 0 S4END[1]
rlabel metal2 30520 1680 30520 1680 0 S4END[2]
rlabel metal2 20048 22456 20048 22456 0 S4END[3]
rlabel metal3 34440 55272 34440 55272 0 S4END[4]
rlabel metal2 35448 55440 35448 55440 0 S4END[5]
rlabel metal2 36008 55832 36008 55832 0 S4END[6]
rlabel metal2 35560 56224 35560 56224 0 S4END[7]
rlabel metal3 36736 56056 36736 56056 0 S4END[8]
rlabel metal2 36904 56112 36904 56112 0 S4END[9]
rlabel metal3 44968 2184 44968 2184 0 SS4BEG[0]
rlabel metal2 45080 406 45080 406 0 SS4BEG[10]
rlabel metal2 45528 686 45528 686 0 SS4BEG[11]
rlabel metal2 45976 1246 45976 1246 0 SS4BEG[12]
rlabel metal3 46760 3640 46760 3640 0 SS4BEG[13]
rlabel metal2 46872 518 46872 518 0 SS4BEG[14]
rlabel metal2 47320 574 47320 574 0 SS4BEG[15]
rlabel metal2 46760 728 46760 728 0 SS4BEG[1]
rlabel metal2 41496 574 41496 574 0 SS4BEG[2]
rlabel metal2 47432 1400 47432 1400 0 SS4BEG[3]
rlabel metal3 44296 728 44296 728 0 SS4BEG[4]
rlabel metal2 42840 1246 42840 1246 0 SS4BEG[5]
rlabel metal2 46984 1960 46984 1960 0 SS4BEG[6]
rlabel metal2 43736 182 43736 182 0 SS4BEG[7]
rlabel metal2 44184 238 44184 238 0 SS4BEG[8]
rlabel metal2 44632 350 44632 350 0 SS4BEG[9]
rlabel metal4 22904 33992 22904 33992 0 SS4END[0]
rlabel metal2 44856 3024 44856 3024 0 SS4END[10]
rlabel metal2 46312 1736 46312 1736 0 SS4END[11]
rlabel metal4 45640 20970 45640 20970 0 SS4END[12]
rlabel metal2 46200 3808 46200 3808 0 SS4END[13]
rlabel metal2 46872 3864 46872 3864 0 SS4END[14]
rlabel metal2 48104 1736 48104 1736 0 SS4END[15]
rlabel metal2 18816 15288 18816 15288 0 SS4END[1]
rlabel metal2 41496 56490 41496 56490 0 SS4END[2]
rlabel metal3 40264 30128 40264 30128 0 SS4END[3]
rlabel metal2 42168 2464 42168 2464 0 SS4END[4]
rlabel metal3 43120 2184 43120 2184 0 SS4END[5]
rlabel metal2 42840 3864 42840 3864 0 SS4END[6]
rlabel metal2 44296 2352 44296 2352 0 SS4END[7]
rlabel metal2 44184 56994 44184 56994 0 SS4END[8]
rlabel metal3 44800 3640 44800 3640 0 SS4END[9]
rlabel metal2 47768 406 47768 406 0 UserCLK
rlabel metal2 52248 35616 52248 35616 0 UserCLK_regs
rlabel metal2 47768 56882 47768 56882 0 UserCLKo
rlabel metal2 15288 2240 15288 2240 0 W1BEG[0]
rlabel metal2 15176 840 15176 840 0 W1BEG[1]
rlabel metal3 462 1176 462 1176 0 W1BEG[2]
rlabel metal2 11592 896 11592 896 0 W1BEG[3]
rlabel metal3 53858 280 53858 280 0 W1END[0]
rlabel metal3 50288 2968 50288 2968 0 W1END[1]
rlabel metal3 54068 1064 54068 1064 0 W1END[2]
rlabel metal3 50120 1456 50120 1456 0 W1END[3]
rlabel metal3 1694 2072 1694 2072 0 W2BEG[0]
rlabel metal2 13944 2296 13944 2296 0 W2BEG[1]
rlabel metal2 7784 616 7784 616 0 W2BEG[2]
rlabel metal3 294 3416 294 3416 0 W2BEG[3]
rlabel metal2 7336 3808 7336 3808 0 W2BEG[4]
rlabel metal2 8008 2688 8008 2688 0 W2BEG[5]
rlabel metal2 10920 840 10920 840 0 W2BEG[6]
rlabel metal3 910 5208 910 5208 0 W2BEG[7]
rlabel metal2 11592 4312 11592 4312 0 W2BEGb[0]
rlabel metal2 10920 4760 10920 4760 0 W2BEGb[1]
rlabel metal2 4088 2408 4088 2408 0 W2BEGb[2]
rlabel metal3 406 7000 406 7000 0 W2BEGb[3]
rlabel metal3 1190 7448 1190 7448 0 W2BEGb[4]
rlabel metal3 1722 7896 1722 7896 0 W2BEGb[5]
rlabel metal3 462 8344 462 8344 0 W2BEGb[6]
rlabel metal3 798 8792 798 8792 0 W2BEGb[7]
rlabel metal3 39704 10472 39704 10472 0 W2END[0]
rlabel metal2 8008 16128 8008 16128 0 W2END[1]
rlabel metal2 25704 8064 25704 8064 0 W2END[2]
rlabel metal3 44352 19992 44352 19992 0 W2END[3]
rlabel metal2 20832 16072 20832 16072 0 W2END[4]
rlabel metal2 15736 41160 15736 41160 0 W2END[5]
rlabel metal4 43624 4424 43624 4424 0 W2END[6]
rlabel metal4 44296 19600 44296 19600 0 W2END[7]
rlabel metal3 35224 2408 35224 2408 0 W2MID[0]
rlabel metal3 46144 2968 46144 2968 0 W2MID[1]
rlabel metal3 48944 2632 48944 2632 0 W2MID[2]
rlabel metal3 51688 3304 51688 3304 0 W2MID[3]
rlabel metal3 19208 2520 19208 2520 0 W2MID[4]
rlabel metal2 24024 6608 24024 6608 0 W2MID[5]
rlabel metal3 42840 16744 42840 16744 0 W2MID[6]
rlabel metal3 54096 16632 54096 16632 0 W2MID[7]
rlabel metal3 350 16408 350 16408 0 W6BEG[0]
rlabel metal2 1064 18928 1064 18928 0 W6BEG[10]
rlabel metal3 574 21336 574 21336 0 W6BEG[11]
rlabel metal3 350 16856 350 16856 0 W6BEG[1]
rlabel metal3 1722 17304 1722 17304 0 W6BEG[2]
rlabel metal2 5656 17248 5656 17248 0 W6BEG[3]
rlabel metal3 518 18200 518 18200 0 W6BEG[4]
rlabel metal3 182 18648 182 18648 0 W6BEG[5]
rlabel metal3 462 19096 462 19096 0 W6BEG[6]
rlabel metal3 1722 19544 1722 19544 0 W6BEG[7]
rlabel metal2 3976 19936 3976 19936 0 W6BEG[8]
rlabel metal2 3304 20160 3304 20160 0 W6BEG[9]
rlabel metal3 56266 16408 56266 16408 0 W6END[0]
rlabel metal3 52122 20888 52122 20888 0 W6END[10]
rlabel metal3 56882 21336 56882 21336 0 W6END[11]
rlabel metal2 20440 30072 20440 30072 0 W6END[1]
rlabel metal3 56602 17304 56602 17304 0 W6END[2]
rlabel metal3 57274 17752 57274 17752 0 W6END[3]
rlabel metal3 56434 18200 56434 18200 0 W6END[4]
rlabel metal2 51464 15568 51464 15568 0 W6END[5]
rlabel metal3 57162 19096 57162 19096 0 W6END[6]
rlabel metal2 52808 18648 52808 18648 0 W6END[7]
rlabel metal2 48440 19712 48440 19712 0 W6END[8]
rlabel metal2 46984 18368 46984 18368 0 W6END[9]
rlabel metal2 1624 2464 1624 2464 0 WW4BEG[0]
rlabel metal2 13496 8848 13496 8848 0 WW4BEG[10]
rlabel metal2 9576 14000 9576 14000 0 WW4BEG[11]
rlabel metal3 406 14616 406 14616 0 WW4BEG[12]
rlabel metal2 7952 13160 7952 13160 0 WW4BEG[13]
rlabel metal3 8792 14728 8792 14728 0 WW4BEG[14]
rlabel metal2 9240 15568 9240 15568 0 WW4BEG[15]
rlabel metal2 2128 3752 2128 3752 0 WW4BEG[1]
rlabel metal2 8288 8904 8288 8904 0 WW4BEG[2]
rlabel metal3 1722 10584 1722 10584 0 WW4BEG[3]
rlabel metal3 1120 3752 1120 3752 0 WW4BEG[4]
rlabel metal3 350 11480 350 11480 0 WW4BEG[5]
rlabel metal3 630 11928 630 11928 0 WW4BEG[6]
rlabel metal2 168 6216 168 6216 0 WW4BEG[7]
rlabel metal3 126 12824 126 12824 0 WW4BEG[8]
rlabel metal3 1246 13272 1246 13272 0 WW4BEG[9]
rlabel metal3 19488 25704 19488 25704 0 WW4END[0]
rlabel metal2 49784 12936 49784 12936 0 WW4END[10]
rlabel metal2 56280 2912 56280 2912 0 WW4END[11]
rlabel metal3 57218 14616 57218 14616 0 WW4END[12]
rlabel metal2 49896 14896 49896 14896 0 WW4END[13]
rlabel metal3 56994 15512 56994 15512 0 WW4END[14]
rlabel metal2 50680 15624 50680 15624 0 WW4END[15]
rlabel metal2 23912 33656 23912 33656 0 WW4END[1]
rlabel metal3 43344 23240 43344 23240 0 WW4END[2]
rlabel metal4 26376 22624 26376 22624 0 WW4END[3]
rlabel metal2 51464 7560 51464 7560 0 WW4END[4]
rlabel metal3 55258 11480 55258 11480 0 WW4END[5]
rlabel metal2 56168 2660 56168 2660 0 WW4END[6]
rlabel metal3 56546 12376 56546 12376 0 WW4END[7]
rlabel metal3 53032 9016 53032 9016 0 WW4END[8]
rlabel metal2 54488 4536 54488 4536 0 WW4END[9]
rlabel metal2 45248 49112 45248 49112 0 _0000_
rlabel metal2 49336 16743 49336 16743 0 _0001_
rlabel metal2 52136 24248 52136 24248 0 _0002_
rlabel metal2 46648 26488 46648 26488 0 _0003_
rlabel metal3 46816 37352 46816 37352 0 _0004_
rlabel metal3 49224 51464 49224 51464 0 _0005_
rlabel metal2 49056 48328 49056 48328 0 _0006_
rlabel metal3 44520 52136 44520 52136 0 _0007_
rlabel metal2 20104 6664 20104 6664 0 _0008_
rlabel metal2 20944 3640 20944 3640 0 _0009_
rlabel metal2 21336 5096 21336 5096 0 _0010_
rlabel metal2 21896 6440 21896 6440 0 _0011_
rlabel metal2 20776 4592 20776 4592 0 _0012_
rlabel metal2 20104 4592 20104 4592 0 _0013_
rlabel metal3 20328 4312 20328 4312 0 _0014_
rlabel metal3 21952 2744 21952 2744 0 _0015_
rlabel metal3 21560 2632 21560 2632 0 _0016_
rlabel metal2 22848 2632 22848 2632 0 _0017_
rlabel metal3 33152 2744 33152 2744 0 _0018_
rlabel metal3 27048 2128 27048 2128 0 _0019_
rlabel metal4 3080 20552 3080 20552 0 _0020_
rlabel metal3 37520 4984 37520 4984 0 _0021_
rlabel metal2 38808 4872 38808 4872 0 _0022_
rlabel metal3 47376 10472 47376 10472 0 _0023_
rlabel metal3 46648 4928 46648 4928 0 _0024_
rlabel metal2 54152 5600 54152 5600 0 _0025_
rlabel metal2 53872 6104 53872 6104 0 _0026_
rlabel metal2 7280 6776 7280 6776 0 _0027_
rlabel metal2 9352 7056 9352 7056 0 _0028_
rlabel metal2 7840 5208 7840 5208 0 _0029_
rlabel metal3 8736 5320 8736 5320 0 _0030_
rlabel metal2 4872 6944 4872 6944 0 _0031_
rlabel metal3 8120 5768 8120 5768 0 _0032_
rlabel metal2 7112 6328 7112 6328 0 _0033_
rlabel metal3 6776 6664 6776 6664 0 _0034_
rlabel metal2 44968 13664 44968 13664 0 _0035_
rlabel metal2 26488 22904 26488 22904 0 _0036_
rlabel metal2 14952 6888 14952 6888 0 _0037_
rlabel metal3 15624 6776 15624 6776 0 _0038_
rlabel metal3 16408 3528 16408 3528 0 _0039_
rlabel metal2 16968 4368 16968 4368 0 _0040_
rlabel metal3 15288 5768 15288 5768 0 _0041_
rlabel metal2 17024 5208 17024 5208 0 _0042_
rlabel metal2 16632 5992 16632 5992 0 _0043_
rlabel metal2 15512 6328 15512 6328 0 _0044_
rlabel metal3 45024 15176 45024 15176 0 _0045_
rlabel metal2 43624 13552 43624 13552 0 _0046_
rlabel metal3 45416 16072 45416 16072 0 _0047_
rlabel metal2 48552 10752 48552 10752 0 _0048_
rlabel metal2 50232 11144 50232 11144 0 _0049_
rlabel metal3 52584 8344 52584 8344 0 _0050_
rlabel metal2 52024 9912 52024 9912 0 _0051_
rlabel metal2 51688 10080 51688 10080 0 _0052_
rlabel metal2 51912 13272 51912 13272 0 _0053_
rlabel metal2 52136 12656 52136 12656 0 _0054_
rlabel metal2 52136 13328 52136 13328 0 _0055_
rlabel metal2 52304 10808 52304 10808 0 _0056_
rlabel metal4 49784 10472 49784 10472 0 _0057_
rlabel metal2 50008 9408 50008 9408 0 _0058_
rlabel metal2 52136 6160 52136 6160 0 _0059_
rlabel metal2 50232 9632 50232 9632 0 _0060_
rlabel metal3 48104 10584 48104 10584 0 _0061_
rlabel metal2 48888 10584 48888 10584 0 _0062_
rlabel metal2 48888 16352 48888 16352 0 _0063_
rlabel metal3 47712 15288 47712 15288 0 _0064_
rlabel metal2 46256 16296 46256 16296 0 _0065_
rlabel metal2 50792 16744 50792 16744 0 _0066_
rlabel metal2 43456 15512 43456 15512 0 _0067_
rlabel metal2 45192 14784 45192 14784 0 _0068_
rlabel metal2 47320 16800 47320 16800 0 _0069_
rlabel metal2 52472 17024 52472 17024 0 _0070_
rlabel metal2 52528 18312 52528 18312 0 _0071_
rlabel metal3 53256 21784 53256 21784 0 _0072_
rlabel metal3 54880 18200 54880 18200 0 _0073_
rlabel metal2 53648 17528 53648 17528 0 _0074_
rlabel metal2 53648 17864 53648 17864 0 _0075_
rlabel metal2 51576 16296 51576 16296 0 _0076_
rlabel metal3 53536 22120 53536 22120 0 _0077_
rlabel metal2 47600 15848 47600 15848 0 _0078_
rlabel metal3 53536 20776 53536 20776 0 _0079_
rlabel metal2 49000 14952 49000 14952 0 _0080_
rlabel metal3 54712 16128 54712 16128 0 _0081_
rlabel metal3 52136 18480 52136 18480 0 _0082_
rlabel metal2 48216 11760 48216 11760 0 _0083_
rlabel metal2 47320 12488 47320 12488 0 _0084_
rlabel metal2 47824 12040 47824 12040 0 _0085_
rlabel metal2 48328 12376 48328 12376 0 _0086_
rlabel metal2 48384 12712 48384 12712 0 _0087_
rlabel metal2 48328 9268 48328 9268 0 _0088_
rlabel metal3 50792 13160 50792 13160 0 _0089_
rlabel metal2 55720 13888 55720 13888 0 _0090_
rlabel metal2 55608 14392 55608 14392 0 _0091_
rlabel metal2 52360 17360 52360 17360 0 _0092_
rlabel metal3 51072 18536 51072 18536 0 _0093_
rlabel metal3 54320 21336 54320 21336 0 _0094_
rlabel metal2 52920 20888 52920 20888 0 _0095_
rlabel metal2 54824 17864 54824 17864 0 _0096_
rlabel metal2 56280 18816 56280 18816 0 _0097_
rlabel metal3 53592 20664 53592 20664 0 _0098_
rlabel metal2 52864 20216 52864 20216 0 _0099_
rlabel metal2 54040 24528 54040 24528 0 _0100_
rlabel metal2 10080 48104 10080 48104 0 _0101_
rlabel metal2 10192 46648 10192 46648 0 _0102_
rlabel metal2 8344 48328 8344 48328 0 _0103_
rlabel metal2 9912 46872 9912 46872 0 _0104_
rlabel metal2 13048 40320 13048 40320 0 _0105_
rlabel metal4 10808 41832 10808 41832 0 _0106_
rlabel metal2 12712 46312 12712 46312 0 _0107_
rlabel metal2 12936 45864 12936 45864 0 _0108_
rlabel metal2 44296 32032 44296 32032 0 _0109_
rlabel metal2 7112 20608 7112 20608 0 _0110_
rlabel metal2 21672 25620 21672 25620 0 _0111_
rlabel metal2 25032 25424 25032 25424 0 _0112_
rlabel metal2 21336 24472 21336 24472 0 _0113_
rlabel metal2 21112 25144 21112 25144 0 _0114_
rlabel metal2 21672 27608 21672 27608 0 _0115_
rlabel metal3 21392 26712 21392 26712 0 _0116_
rlabel metal3 22736 25704 22736 25704 0 _0117_
rlabel metal2 24584 25032 24584 25032 0 _0118_
rlabel metal2 40040 21616 40040 21616 0 _0119_
rlabel metal3 15512 17472 15512 17472 0 _0120_
rlabel metal2 25368 32760 25368 32760 0 _0121_
rlabel metal3 44856 32200 44856 32200 0 _0122_
rlabel metal2 43512 35672 43512 35672 0 _0123_
rlabel metal2 16968 30800 16968 30800 0 _0124_
rlabel metal2 19208 29008 19208 29008 0 _0125_
rlabel metal3 19880 29288 19880 29288 0 _0126_
rlabel metal3 19936 28840 19936 28840 0 _0127_
rlabel metal2 20216 30296 20216 30296 0 _0128_
rlabel metal2 19656 28840 19656 28840 0 _0129_
rlabel metal2 20104 28168 20104 28168 0 _0130_
rlabel metal2 19880 28112 19880 28112 0 _0131_
rlabel metal2 27384 32536 27384 32536 0 _0132_
rlabel metal3 19712 17864 19712 17864 0 _0133_
rlabel metal2 16184 50120 16184 50120 0 _0134_
rlabel metal3 18816 46648 18816 46648 0 _0135_
rlabel metal3 20440 46872 20440 46872 0 _0136_
rlabel metal2 16072 49840 16072 49840 0 _0137_
rlabel metal3 15288 43512 15288 43512 0 _0138_
rlabel metal2 16968 44912 16968 44912 0 _0139_
rlabel metal2 16576 44520 16576 44520 0 _0140_
rlabel metal2 15624 45248 15624 45248 0 _0141_
rlabel metal2 30744 2576 30744 2576 0 _0142_
rlabel metal2 28560 33320 28560 33320 0 _0143_
rlabel metal2 43400 36064 43400 36064 0 _0144_
rlabel metal3 51464 43512 51464 43512 0 _0145_
rlabel metal2 53816 34664 53816 34664 0 _0146_
rlabel metal2 53256 29848 53256 29848 0 _0147_
rlabel metal2 43512 31136 43512 31136 0 _0148_
rlabel metal2 51968 33992 51968 33992 0 _0149_
rlabel metal4 44184 30856 44184 30856 0 _0150_
rlabel metal2 51240 35336 51240 35336 0 _0151_
rlabel metal2 50232 30912 50232 30912 0 _0152_
rlabel metal3 54936 24808 54936 24808 0 _0153_
rlabel metal2 49448 26320 49448 26320 0 _0154_
rlabel metal3 50568 35448 50568 35448 0 _0155_
rlabel metal2 50344 32704 50344 32704 0 _0156_
rlabel metal3 40040 35672 40040 35672 0 _0157_
rlabel metal2 38864 35784 38864 35784 0 _0158_
rlabel metal2 2408 40320 2408 40320 0 _0159_
rlabel metal2 2744 39984 2744 39984 0 _0160_
rlabel metal2 2184 39480 2184 39480 0 _0161_
rlabel metal2 4088 38696 4088 38696 0 _0162_
rlabel metal2 3976 40208 3976 40208 0 _0163_
rlabel metal3 4256 49672 4256 49672 0 _0164_
rlabel metal2 5208 41832 5208 41832 0 _0165_
rlabel metal2 4928 40376 4928 40376 0 _0166_
rlabel metal2 42112 36680 42112 36680 0 _0167_
rlabel metal2 39256 28896 39256 28896 0 _0168_
rlabel metal2 39144 27496 39144 27496 0 _0169_
rlabel metal2 39816 28000 39816 28000 0 _0170_
rlabel metal2 39200 25144 39200 25144 0 _0171_
rlabel metal2 39256 24752 39256 24752 0 _0172_
rlabel metal2 23464 21168 23464 21168 0 _0173_
rlabel metal3 47264 26824 47264 26824 0 _0174_
rlabel metal3 52360 28056 52360 28056 0 _0175_
rlabel metal2 52920 44296 52920 44296 0 _0176_
rlabel metal2 33320 13664 33320 13664 0 _0177_
rlabel metal2 39256 39984 39256 39984 0 _0178_
rlabel metal2 8288 39704 8288 39704 0 _0179_
rlabel metal2 3304 38864 3304 38864 0 _0180_
rlabel metal2 9576 38360 9576 38360 0 _0181_
rlabel metal3 8792 38024 8792 38024 0 _0182_
rlabel metal2 9968 41272 9968 41272 0 _0183_
rlabel metal2 9464 36960 9464 36960 0 _0184_
rlabel metal3 8848 38696 8848 38696 0 _0185_
rlabel metal3 9688 38696 9688 38696 0 _0186_
rlabel metal2 43288 39480 43288 39480 0 _0187_
rlabel metal3 36568 28280 36568 28280 0 _0188_
rlabel metal2 35224 23912 35224 23912 0 _0189_
rlabel metal2 35784 23408 35784 23408 0 _0190_
rlabel metal2 35616 23240 35616 23240 0 _0191_
rlabel metal4 39872 20970 39872 20970 0 _0192_
rlabel metal3 48104 39592 48104 39592 0 _0193_
rlabel metal2 25032 44296 25032 44296 0 _0194_
rlabel metal3 16576 41944 16576 41944 0 _0195_
rlabel metal2 8400 31752 8400 31752 0 _0196_
rlabel metal2 9576 30912 9576 30912 0 _0197_
rlabel metal2 10136 31024 10136 31024 0 _0198_
rlabel metal3 10024 30184 10024 30184 0 _0199_
rlabel metal2 9296 29400 9296 29400 0 _0200_
rlabel metal2 7560 32648 7560 32648 0 _0201_
rlabel metal3 8624 30408 8624 30408 0 _0202_
rlabel metal2 9352 29176 9352 29176 0 _0203_
rlabel metal2 20776 47264 20776 47264 0 _0204_
rlabel metal2 26376 44296 26376 44296 0 _0205_
rlabel metal2 50232 47600 50232 47600 0 _0206_
rlabel metal2 51184 48216 51184 48216 0 _0207_
rlabel metal3 54824 48328 54824 48328 0 _0208_
rlabel metal2 43624 47600 43624 47600 0 _0209_
rlabel metal4 50232 40768 50232 40768 0 _0210_
rlabel metal2 52024 43288 52024 43288 0 _0211_
rlabel metal2 49672 43288 49672 43288 0 _0212_
rlabel metal3 50120 41552 50120 41552 0 _0213_
rlabel metal2 41048 17416 41048 17416 0 _0214_
rlabel metal2 40264 16744 40264 16744 0 _0215_
rlabel metal2 40656 16296 40656 16296 0 _0216_
rlabel metal2 3864 34216 3864 34216 0 _0217_
rlabel metal2 2408 34440 2408 34440 0 _0218_
rlabel metal2 2744 34216 2744 34216 0 _0219_
rlabel metal3 3528 34104 3528 34104 0 _0220_
rlabel metal2 3416 35364 3416 35364 0 _0221_
rlabel metal3 6720 35000 6720 35000 0 _0222_
rlabel metal3 5768 34888 5768 34888 0 _0223_
rlabel metal2 5096 34440 5096 34440 0 _0224_
rlabel metal2 43288 17472 43288 17472 0 _0225_
rlabel metal2 42280 17595 42280 17595 0 _0226_
rlabel metal2 41496 20440 41496 20440 0 _0227_
rlabel metal2 41272 17584 41272 17584 0 _0228_
rlabel metal2 53424 46872 53424 46872 0 _0229_
rlabel metal2 54208 42728 54208 42728 0 _0230_
rlabel metal3 53984 42616 53984 42616 0 _0231_
rlabel metal2 51800 44072 51800 44072 0 _0232_
rlabel metal2 52416 45304 52416 45304 0 _0233_
rlabel metal2 52696 47096 52696 47096 0 _0234_
rlabel metal2 55160 45808 55160 45808 0 _0235_
rlabel metal2 53256 45360 53256 45360 0 _0236_
rlabel metal2 51016 44576 51016 44576 0 _0237_
rlabel metal2 49672 50624 49672 50624 0 _0238_
rlabel metal2 2184 48328 2184 48328 0 _0239_
rlabel metal3 6160 47544 6160 47544 0 _0240_
rlabel metal2 7392 39368 7392 39368 0 _0241_
rlabel metal3 3976 47768 3976 47768 0 _0242_
rlabel metal3 16632 48216 16632 48216 0 _0243_
rlabel metal4 15400 55109 15400 55109 0 _0244_
rlabel metal2 3584 49224 3584 49224 0 _0245_
rlabel metal2 3752 46648 3752 46648 0 _0246_
rlabel metal3 46312 34328 46312 34328 0 _0247_
rlabel metal2 46648 34328 46648 34328 0 _0248_
rlabel metal2 46424 34216 46424 34216 0 _0249_
rlabel metal2 47264 33544 47264 33544 0 _0250_
rlabel metal2 47040 30184 47040 30184 0 _0251_
rlabel metal3 42840 28728 42840 28728 0 _0252_
rlabel metal2 47320 30240 47320 30240 0 _0253_
rlabel metal2 19208 35056 19208 35056 0 _0254_
rlabel metal2 19712 34888 19712 34888 0 _0255_
rlabel metal2 20048 35672 20048 35672 0 _0256_
rlabel metal2 19768 35112 19768 35112 0 _0257_
rlabel metal2 20328 33544 20328 33544 0 _0258_
rlabel metal3 21336 34104 21336 34104 0 _0259_
rlabel metal3 20272 34104 20272 34104 0 _0260_
rlabel metal2 19880 33824 19880 33824 0 _0261_
rlabel metal2 44352 30856 44352 30856 0 _0262_
rlabel metal2 30520 31136 30520 31136 0 _0263_
rlabel metal3 29680 30744 29680 30744 0 _0264_
rlabel metal3 28336 30744 28336 30744 0 _0265_
rlabel metal3 44184 30464 44184 30464 0 _0266_
rlabel metal2 46424 29064 46424 29064 0 _0267_
rlabel metal3 47544 29512 47544 29512 0 _0268_
rlabel metal2 49560 29680 49560 29680 0 _0269_
rlabel metal2 49840 26488 49840 26488 0 _0270_
rlabel metal2 52584 29008 52584 29008 0 _0271_
rlabel metal2 52248 26152 52248 26152 0 _0272_
rlabel metal3 56336 30408 56336 30408 0 _0273_
rlabel metal3 54152 34216 54152 34216 0 _0274_
rlabel metal2 55496 34104 55496 34104 0 _0275_
rlabel metal3 54432 29400 54432 29400 0 _0276_
rlabel metal2 53256 32032 53256 32032 0 _0277_
rlabel metal2 52248 30576 52248 30576 0 _0278_
rlabel metal2 52472 30912 52472 30912 0 _0279_
rlabel metal2 35784 28168 35784 28168 0 _0280_
rlabel metal2 35672 29792 35672 29792 0 _0281_
rlabel metal3 33488 28728 33488 28728 0 _0282_
rlabel metal3 33488 27832 33488 27832 0 _0283_
rlabel metal3 36008 23128 36008 23128 0 _0284_
rlabel metal3 33656 29288 33656 29288 0 _0285_
rlabel metal3 32480 30184 32480 30184 0 _0286_
rlabel metal3 33320 29624 33320 29624 0 _0287_
rlabel metal2 36960 23128 36960 23128 0 _0288_
rlabel metal2 41216 6776 41216 6776 0 _0289_
rlabel metal2 33320 9912 33320 9912 0 _0290_
rlabel metal2 44296 7952 44296 7952 0 _0291_
rlabel metal2 3304 42336 3304 42336 0 _0292_
rlabel metal2 3640 42616 3640 42616 0 _0293_
rlabel metal2 4368 42952 4368 42952 0 _0294_
rlabel metal2 3640 43792 3640 43792 0 _0295_
rlabel metal3 4200 44968 4200 44968 0 _0296_
rlabel metal2 5488 44520 5488 44520 0 _0297_
rlabel metal3 2996 45304 2996 45304 0 _0298_
rlabel metal3 4592 43512 4592 43512 0 _0299_
rlabel metal3 29176 3808 29176 3808 0 _0300_
rlabel metal2 42168 22064 42168 22064 0 _0301_
rlabel metal3 42448 8232 42448 8232 0 _0302_
rlabel metal3 43568 8120 43568 8120 0 _0303_
rlabel metal2 43624 9072 43624 9072 0 _0304_
rlabel metal2 42560 24584 42560 24584 0 _0305_
rlabel metal2 44632 28280 44632 28280 0 _0306_
rlabel metal2 52584 30744 52584 30744 0 _0307_
rlabel metal2 56168 27888 56168 27888 0 _0308_
rlabel metal2 55160 24136 55160 24136 0 _0309_
rlabel metal2 56168 26992 56168 26992 0 _0310_
rlabel metal2 54936 28336 54936 28336 0 _0311_
rlabel metal3 54152 27272 54152 27272 0 _0312_
rlabel metal3 53704 26376 53704 26376 0 _0313_
rlabel metal2 54880 27272 54880 27272 0 _0314_
rlabel metal2 51352 32592 51352 32592 0 _0315_
rlabel metal2 49336 28840 49336 28840 0 _0316_
rlabel metal2 39368 44072 39368 44072 0 _0317_
rlabel metal3 40712 35448 40712 35448 0 _0318_
rlabel metal2 45528 42224 45528 42224 0 _0319_
rlabel metal2 25256 42840 25256 42840 0 _0320_
rlabel metal3 42896 47992 42896 47992 0 _0321_
rlabel metal2 39480 43848 39480 43848 0 _0322_
rlabel metal2 39144 43568 39144 43568 0 _0323_
rlabel metal2 42952 47040 42952 47040 0 _0324_
rlabel metal2 39592 46648 39592 46648 0 _0325_
rlabel metal2 42616 46144 42616 46144 0 _0326_
rlabel metal2 42952 43232 42952 43232 0 _0327_
rlabel metal3 43288 45192 43288 45192 0 _0328_
rlabel metal3 43176 45080 43176 45080 0 _0329_
rlabel metal2 43176 45416 43176 45416 0 _0330_
rlabel metal2 43288 42896 43288 42896 0 _0331_
rlabel metal2 43624 42728 43624 42728 0 _0332_
rlabel metal2 43736 18200 43736 18200 0 _0333_
rlabel metal2 42952 17976 42952 17976 0 _0334_
rlabel metal2 43624 18088 43624 18088 0 _0335_
rlabel metal2 43512 18872 43512 18872 0 _0336_
rlabel metal2 48328 43568 48328 43568 0 _0337_
rlabel metal3 45640 41272 45640 41272 0 _0338_
rlabel metal2 48216 42336 48216 42336 0 _0339_
rlabel metal2 47264 49784 47264 49784 0 _0340_
rlabel metal2 46088 42672 46088 42672 0 _0341_
rlabel metal3 46704 42728 46704 42728 0 _0342_
rlabel metal3 48664 43288 48664 43288 0 _0343_
rlabel metal2 43288 41552 43288 41552 0 _0344_
rlabel metal2 46872 42840 46872 42840 0 _0345_
rlabel metal2 46256 41384 46256 41384 0 _0346_
rlabel metal2 46592 42728 46592 42728 0 _0347_
rlabel metal2 47544 48104 47544 48104 0 _0348_
rlabel metal2 44968 50680 44968 50680 0 _0349_
rlabel metal2 48664 46312 48664 46312 0 _0350_
rlabel metal2 39200 46088 39200 46088 0 _0351_
rlabel metal3 11144 50792 11144 50792 0 _0352_
rlabel metal2 9912 53536 9912 53536 0 _0353_
rlabel metal2 12768 52360 12768 52360 0 _0354_
rlabel metal2 13328 54488 13328 54488 0 _0355_
rlabel metal2 13832 51296 13832 51296 0 _0356_
rlabel metal2 13720 53704 13720 53704 0 _0357_
rlabel metal2 21784 54600 21784 54600 0 _0358_
rlabel metal2 12264 54600 12264 54600 0 _0359_
rlabel metal2 36904 40264 36904 40264 0 _0360_
rlabel metal3 35896 40376 35896 40376 0 _0361_
rlabel metal2 36232 39144 36232 39144 0 _0362_
rlabel metal3 38696 26264 38696 26264 0 _0363_
rlabel metal2 39480 39984 39480 39984 0 _0364_
rlabel metal2 34440 41552 34440 41552 0 _0365_
rlabel metal2 15288 39144 15288 39144 0 _0366_
rlabel metal2 16184 39984 16184 39984 0 _0367_
rlabel metal2 39816 40880 39816 40880 0 _0368_
rlabel metal3 39872 42056 39872 42056 0 _0369_
rlabel metal2 40712 42336 40712 42336 0 _0370_
rlabel metal2 41272 43512 41272 43512 0 _0371_
rlabel metal2 41720 44744 41720 44744 0 _0372_
rlabel metal2 39088 45864 39088 45864 0 _0373_
rlabel metal2 33432 34832 33432 34832 0 _0374_
rlabel metal2 25480 36680 25480 36680 0 _0375_
rlabel metal3 19936 52248 19936 52248 0 _0376_
rlabel metal3 18760 51240 18760 51240 0 _0377_
rlabel metal2 21112 51072 21112 51072 0 _0378_
rlabel metal2 21224 51240 21224 51240 0 _0379_
rlabel metal2 16296 52416 16296 52416 0 _0380_
rlabel metal2 18144 49336 18144 49336 0 _0381_
rlabel metal2 20832 48440 20832 48440 0 _0382_
rlabel metal3 18368 51352 18368 51352 0 _0383_
rlabel metal2 35672 37184 35672 37184 0 _0384_
rlabel metal3 1848 24584 1848 24584 0 _0385_
rlabel metal2 38136 46312 38136 46312 0 _0386_
rlabel metal2 32536 54320 32536 54320 0 _0387_
rlabel metal2 27720 43512 27720 43512 0 _0388_
rlabel metal2 22456 42112 22456 42112 0 _0389_
rlabel metal2 25592 51016 25592 51016 0 _0390_
rlabel metal2 24024 51464 24024 51464 0 _0391_
rlabel metal2 25704 51576 25704 51576 0 _0392_
rlabel metal2 26152 53424 26152 53424 0 _0393_
rlabel metal2 24696 50680 24696 50680 0 _0394_
rlabel metal4 25928 54152 25928 54152 0 _0395_
rlabel metal2 25592 53928 25592 53928 0 _0396_
rlabel metal3 25088 53704 25088 53704 0 _0397_
rlabel metal2 18536 20944 18536 20944 0 _0398_
rlabel metal2 28952 42840 28952 42840 0 _0399_
rlabel metal2 39088 48104 39088 48104 0 _0400_
rlabel metal2 35504 51352 35504 51352 0 _0401_
rlabel metal3 33824 53704 33824 53704 0 _0402_
rlabel metal3 32536 49224 32536 49224 0 _0403_
rlabel metal2 39032 53592 39032 53592 0 _0404_
rlabel metal4 1960 20272 1960 20272 0 _0405_
rlabel metal2 13328 13944 13328 13944 0 _0406_
rlabel metal3 16352 17080 16352 17080 0 _0407_
rlabel metal2 16968 16800 16968 16800 0 _0408_
rlabel metal4 19320 15456 19320 15456 0 _0409_
rlabel metal3 36064 18312 36064 18312 0 _0410_
rlabel metal3 4200 51408 4200 51408 0 _0411_
rlabel metal2 4032 51576 4032 51576 0 _0412_
rlabel metal2 6048 51128 6048 51128 0 _0413_
rlabel metal2 5432 51632 5432 51632 0 _0414_
rlabel metal2 7448 38696 7448 38696 0 _0415_
rlabel metal2 5992 45528 5992 45528 0 _0416_
rlabel metal3 6888 51240 6888 51240 0 _0417_
rlabel metal2 6048 51352 6048 51352 0 _0418_
rlabel metal2 39368 18872 39368 18872 0 _0419_
rlabel metal2 38584 16408 38584 16408 0 _0420_
rlabel metal3 37632 17864 37632 17864 0 _0421_
rlabel metal2 32200 53368 32200 53368 0 _0422_
rlabel metal2 34776 54880 34776 54880 0 _0423_
rlabel metal2 35112 54320 35112 54320 0 _0424_
rlabel metal2 37800 54880 37800 54880 0 _0425_
rlabel metal3 36568 50568 36568 50568 0 _0426_
rlabel metal3 36960 47992 36960 47992 0 _0427_
rlabel metal3 36624 50792 36624 50792 0 _0428_
rlabel metal2 41608 54320 41608 54320 0 _0429_
rlabel metal2 38808 44912 38808 44912 0 _0430_
rlabel metal2 37128 41720 37128 41720 0 _0431_
rlabel metal3 37520 43400 37520 43400 0 _0432_
rlabel metal2 35448 44184 35448 44184 0 _0433_
rlabel metal2 39704 43120 39704 43120 0 _0434_
rlabel metal3 38472 48104 38472 48104 0 _0435_
rlabel metal2 36904 47320 36904 47320 0 _0436_
rlabel metal2 38248 44744 38248 44744 0 _0437_
rlabel metal3 30800 44408 30800 44408 0 _0438_
rlabel metal2 30520 43008 30520 43008 0 _0439_
rlabel metal2 34664 52304 34664 52304 0 _0440_
rlabel metal3 34384 44408 34384 44408 0 _0441_
rlabel metal2 35560 48776 35560 48776 0 _0442_
rlabel metal3 31192 47432 31192 47432 0 _0443_
rlabel metal2 35672 48888 35672 48888 0 _0444_
rlabel metal2 30072 49056 30072 49056 0 _0445_
rlabel metal3 30128 47544 30128 47544 0 _0446_
rlabel metal3 32816 47208 32816 47208 0 _0447_
rlabel metal3 37240 18312 37240 18312 0 _0448_
rlabel metal2 38584 47488 38584 47488 0 _0449_
rlabel metal2 38360 48048 38360 48048 0 _0450_
rlabel metal3 37072 47544 37072 47544 0 _0451_
rlabel metal2 33656 47488 33656 47488 0 _0452_
rlabel metal2 31304 44576 31304 44576 0 _0453_
rlabel metal3 31976 46088 31976 46088 0 _0454_
rlabel metal3 34888 46760 34888 46760 0 _0455_
rlabel metal3 36512 44520 36512 44520 0 _0456_
rlabel metal2 35504 47992 35504 47992 0 _0457_
rlabel metal2 35672 45416 35672 45416 0 _0458_
rlabel metal2 36456 46984 36456 46984 0 _0459_
rlabel metal3 41552 48776 41552 48776 0 _0460_
rlabel metal2 42504 48104 42504 48104 0 _0461_
rlabel metal2 18088 48384 18088 48384 0 _0462_
rlabel metal3 18088 49000 18088 49000 0 _0463_
rlabel metal2 16912 47992 16912 47992 0 _0464_
rlabel metal2 11368 44912 11368 44912 0 _0465_
rlabel metal2 11088 45304 11088 45304 0 _0466_
rlabel metal2 48216 31892 48216 31892 0 _0467_
rlabel metal2 48552 30912 48552 30912 0 _0468_
rlabel metal3 46144 30856 46144 30856 0 _0469_
rlabel metal2 48384 30968 48384 30968 0 _0470_
rlabel metal3 48944 31192 48944 31192 0 _0471_
rlabel metal3 55160 35448 55160 35448 0 _0472_
rlabel metal2 52640 38808 52640 38808 0 _0473_
rlabel metal4 53144 46144 53144 46144 0 _0474_
rlabel metal3 51520 38920 51520 38920 0 _0475_
rlabel metal2 53592 39592 53592 39592 0 _0476_
rlabel metal3 54376 36568 54376 36568 0 _0477_
rlabel metal2 52752 35672 52752 35672 0 _0478_
rlabel metal3 55048 39032 55048 39032 0 _0479_
rlabel metal3 55048 38808 55048 38808 0 _0480_
rlabel metal3 55160 38920 55160 38920 0 _0481_
rlabel metal3 53256 35672 53256 35672 0 _0482_
rlabel metal3 45528 4312 45528 4312 0 _0483_
rlabel metal3 45360 10360 45360 10360 0 _0484_
rlabel metal2 44296 6272 44296 6272 0 _0485_
rlabel metal4 50232 19080 50232 19080 0 _0486_
rlabel metal2 50904 34552 50904 34552 0 _0487_
rlabel metal2 52584 37744 52584 37744 0 _0488_
rlabel metal2 55832 35840 55832 35840 0 _0489_
rlabel metal3 55440 35000 55440 35000 0 _0490_
rlabel metal2 51128 38304 51128 38304 0 _0491_
rlabel metal3 55608 34776 55608 34776 0 _0492_
rlabel metal2 54824 37576 54824 37576 0 _0493_
rlabel metal2 51352 40488 51352 40488 0 _0494_
rlabel metal2 47544 36120 47544 36120 0 _0495_
rlabel metal2 10696 42504 10696 42504 0 _0496_
rlabel metal2 10528 42952 10528 42952 0 _0497_
rlabel metal2 9912 45584 9912 45584 0 _0498_
rlabel metal2 8232 43008 8232 43008 0 _0499_
rlabel metal2 4816 25480 4816 25480 0 _0500_
rlabel metal3 4312 27160 4312 27160 0 _0501_
rlabel metal2 3584 26824 3584 26824 0 _0502_
rlabel metal2 4368 25704 4368 25704 0 _0503_
rlabel metal2 3304 27720 3304 27720 0 _0504_
rlabel metal3 3640 28672 3640 28672 0 _0505_
rlabel metal2 3304 28504 3304 28504 0 _0506_
rlabel metal3 4760 26264 4760 26264 0 _0507_
rlabel metal2 7784 21616 7784 21616 0 _0508_
rlabel metal2 5152 24920 5152 24920 0 _0509_
rlabel metal3 5768 24136 5768 24136 0 _0510_
rlabel metal2 5544 25088 5544 25088 0 _0511_
rlabel metal2 6104 24976 6104 24976 0 _0512_
rlabel metal3 9240 23016 9240 23016 0 _0513_
rlabel metal3 8624 23912 8624 23912 0 _0514_
rlabel metal3 7784 24136 7784 24136 0 _0515_
rlabel metal2 6440 24920 6440 24920 0 _0516_
rlabel metal2 4984 31416 4984 31416 0 _0517_
rlabel metal2 3192 33768 3192 33768 0 _0518_
rlabel metal3 3920 32312 3920 32312 0 _0519_
rlabel metal3 4928 31080 4928 31080 0 _0520_
rlabel metal2 3416 30688 3416 30688 0 _0521_
rlabel metal2 3976 32200 3976 32200 0 _0522_
rlabel metal2 4536 29400 4536 29400 0 _0523_
rlabel metal2 4200 30016 4200 30016 0 _0524_
rlabel metal2 13440 27832 13440 27832 0 _0525_
rlabel metal2 12320 25704 12320 25704 0 _0526_
rlabel metal3 12992 26264 12992 26264 0 _0527_
rlabel metal2 13440 26264 13440 26264 0 _0528_
rlabel metal2 14728 28504 14728 28504 0 _0529_
rlabel metal3 13104 27272 13104 27272 0 _0530_
rlabel metal2 13048 26824 13048 26824 0 _0531_
rlabel metal2 12824 26936 12824 26936 0 _0532_
rlabel metal3 9016 26264 9016 26264 0 _0533_
rlabel metal3 9128 26488 9128 26488 0 _0534_
rlabel metal2 7896 27608 7896 27608 0 _0535_
rlabel metal3 9632 27720 9632 27720 0 _0536_
rlabel metal2 9352 28336 9352 28336 0 _0537_
rlabel metal2 9016 28840 9016 28840 0 _0538_
rlabel metal3 10024 43400 10024 43400 0 _0539_
rlabel metal2 11816 43792 11816 43792 0 _0540_
rlabel metal3 11200 43624 11200 43624 0 _0541_
rlabel metal2 7112 45136 7112 45136 0 _0542_
rlabel metal3 5880 42168 5880 42168 0 _0543_
rlabel metal2 5208 43960 5208 43960 0 _0544_
rlabel metal2 9800 43456 9800 43456 0 _0545_
rlabel metal2 9240 42280 9240 42280 0 _0546_
rlabel metal2 8960 42728 8960 42728 0 _0547_
rlabel metal3 2072 14616 2072 14616 0 _0548_
rlabel metal2 1512 14784 1512 14784 0 _0549_
rlabel metal2 4424 13160 4424 13160 0 _0550_
rlabel metal2 4200 15400 4200 15400 0 _0551_
rlabel metal2 5320 13552 5320 13552 0 _0552_
rlabel metal2 4928 13944 4928 13944 0 _0553_
rlabel metal3 4312 14616 4312 14616 0 _0554_
rlabel metal3 2856 14728 2856 14728 0 _0555_
rlabel metal2 7224 9072 7224 9072 0 _0556_
rlabel metal2 5096 7504 5096 7504 0 _0557_
rlabel metal2 4984 9072 4984 9072 0 _0558_
rlabel metal2 7672 9688 7672 9688 0 _0559_
rlabel metal3 8568 13048 8568 13048 0 _0560_
rlabel metal2 6440 11984 6440 11984 0 _0561_
rlabel metal4 4984 12656 4984 12656 0 _0562_
rlabel metal2 5432 11648 5432 11648 0 _0563_
rlabel metal2 5600 11368 5600 11368 0 _0564_
rlabel metal3 8344 12936 8344 12936 0 _0565_
rlabel metal2 11424 9240 11424 9240 0 _0566_
rlabel metal2 11592 9576 11592 9576 0 _0567_
rlabel metal2 11312 10584 11312 10584 0 _0568_
rlabel metal3 10640 10696 10640 10696 0 _0569_
rlabel metal2 12040 10864 12040 10864 0 _0570_
rlabel metal2 12152 10584 12152 10584 0 _0571_
rlabel metal2 9912 11928 9912 11928 0 _0572_
rlabel metal2 9016 11368 9016 11368 0 _0573_
rlabel metal3 10360 18312 10360 18312 0 _0574_
rlabel metal3 12152 19320 12152 19320 0 _0575_
rlabel metal3 12712 19432 12712 19432 0 _0576_
rlabel metal3 11480 19880 11480 19880 0 _0577_
rlabel metal2 11592 20496 11592 20496 0 _0578_
rlabel metal2 8904 16520 8904 16520 0 _0579_
rlabel metal2 9016 16352 9016 16352 0 _0580_
rlabel metal3 10192 17864 10192 17864 0 _0581_
rlabel metal3 9912 16296 9912 16296 0 _0582_
rlabel metal2 9352 20104 9352 20104 0 _0583_
rlabel metal2 16184 24024 16184 24024 0 _0584_
rlabel metal2 16072 24136 16072 24136 0 _0585_
rlabel metal2 16856 22792 16856 22792 0 _0586_
rlabel metal2 15400 24752 15400 24752 0 _0587_
rlabel metal3 18648 23352 18648 23352 0 _0588_
rlabel metal2 19544 24472 19544 24472 0 _0589_
rlabel metal2 17416 22624 17416 22624 0 _0590_
rlabel metal2 17248 22568 17248 22568 0 _0591_
rlabel metal2 6104 18536 6104 18536 0 _0592_
rlabel metal3 4704 17864 4704 17864 0 _0593_
rlabel metal2 6104 19264 6104 19264 0 _0594_
rlabel metal2 5992 19544 5992 19544 0 _0595_
rlabel metal2 17528 20720 17528 20720 0 _0596_
rlabel metal2 16128 18312 16128 18312 0 _0597_
rlabel metal2 3752 22400 3752 22400 0 _0598_
rlabel metal2 1400 22064 1400 22064 0 _0599_
rlabel metal3 17528 40936 17528 40936 0 _0600_
rlabel metal2 17920 43288 17920 43288 0 _0601_
rlabel metal2 7448 34328 7448 34328 0 _0602_
rlabel metal2 8120 33768 8120 33768 0 _0603_
rlabel metal3 30408 20776 30408 20776 0 _0604_
rlabel metal3 29904 22456 29904 22456 0 _0605_
rlabel metal2 38920 9240 38920 9240 0 _0606_
rlabel metal2 38304 8904 38304 8904 0 _0607_
rlabel metal2 33320 2240 33320 2240 0 _0608_
rlabel metal3 32088 4088 32088 4088 0 _0609_
rlabel metal2 31752 17528 31752 17528 0 _0610_
rlabel metal2 33096 16856 33096 16856 0 _0611_
rlabel metal2 31080 19264 31080 19264 0 _0612_
rlabel metal2 32536 16800 32536 16800 0 _0613_
rlabel metal3 33712 16968 33712 16968 0 _0614_
rlabel metal2 32984 17976 32984 17976 0 _0615_
rlabel metal2 43512 2968 43512 2968 0 _0616_
rlabel metal3 20888 46088 20888 46088 0 _0617_
rlabel metal2 19264 46872 19264 46872 0 _0618_
rlabel metal2 19320 46200 19320 46200 0 _0619_
rlabel metal2 21784 49056 21784 49056 0 _0620_
rlabel metal3 23464 47432 23464 47432 0 _0621_
rlabel metal2 20048 45864 20048 45864 0 _0622_
rlabel metal2 23016 40712 23016 40712 0 _0623_
rlabel metal2 22680 41440 22680 41440 0 _0624_
rlabel metal2 21560 40488 21560 40488 0 _0625_
rlabel metal2 20720 41272 20720 41272 0 _0626_
rlabel metal3 30128 38248 30128 38248 0 _0627_
rlabel metal3 29848 38920 29848 38920 0 _0628_
rlabel metal3 35280 31864 35280 31864 0 _0629_
rlabel metal2 38920 32144 38920 32144 0 _0630_
rlabel metal2 35952 30968 35952 30968 0 _0631_
rlabel metal2 38584 32816 38584 32816 0 _0632_
rlabel metal2 38696 31360 38696 31360 0 _0633_
rlabel metal2 38248 30632 38248 30632 0 _0634_
rlabel metal3 52920 29792 52920 29792 0 _0635_
rlabel metal2 31976 41384 31976 41384 0 _0636_
rlabel metal3 31192 41832 31192 41832 0 _0637_
rlabel metal2 15736 38136 15736 38136 0 _0638_
rlabel metal3 15344 37016 15344 37016 0 _0639_
rlabel metal2 27720 48216 27720 48216 0 _0640_
rlabel metal3 26992 49112 26992 49112 0 _0641_
rlabel metal2 25088 31752 25088 31752 0 _0642_
rlabel metal3 25368 30856 25368 30856 0 _0643_
rlabel metal2 30184 51856 30184 51856 0 _0644_
rlabel metal2 29624 52584 29624 52584 0 _0645_
rlabel metal2 25592 36848 25592 36848 0 _0646_
rlabel metal2 25256 37632 25256 37632 0 _0647_
rlabel metal2 35504 50008 35504 50008 0 _0648_
rlabel metal3 40152 18648 40152 18648 0 _0649_
rlabel metal2 42000 20552 42000 20552 0 _0650_
rlabel metal3 41888 20888 41888 20888 0 _0651_
rlabel metal2 42392 20552 42392 20552 0 _0652_
rlabel metal2 40600 21840 40600 21840 0 _0653_
rlabel metal3 41160 21000 41160 21000 0 _0654_
rlabel metal4 39256 21896 39256 21896 0 _0655_
rlabel metal2 41496 22484 41496 22484 0 _0656_
rlabel metal2 41272 21525 41272 21525 0 _0657_
rlabel metal2 48888 21280 48888 21280 0 _0658_
rlabel metal2 44296 51016 44296 51016 0 _0659_
rlabel metal2 41496 25648 41496 25648 0 _0660_
rlabel metal3 42280 25704 42280 25704 0 _0661_
rlabel metal2 40992 27160 40992 27160 0 _0662_
rlabel metal2 43176 26656 43176 26656 0 _0663_
rlabel metal2 43120 26264 43120 26264 0 _0664_
rlabel metal3 40488 25592 40488 25592 0 _0665_
rlabel metal2 41384 25760 41384 25760 0 _0666_
rlabel metal3 42224 24808 42224 24808 0 _0667_
rlabel metal3 42168 25368 42168 25368 0 _0668_
rlabel metal2 41496 26320 41496 26320 0 _0669_
rlabel metal2 42112 26152 42112 26152 0 _0670_
rlabel metal2 51240 21728 51240 21728 0 _0671_
rlabel metal3 46984 51128 46984 51128 0 _0672_
rlabel metal2 44632 50148 44632 50148 0 _0673_
rlabel metal3 45360 51352 45360 51352 0 _0674_
rlabel metal2 49672 20272 49672 20272 0 _0675_
rlabel metal2 49224 16632 49224 16632 0 _0676_
rlabel metal2 50344 17752 50344 17752 0 _0677_
rlabel metal2 49672 16632 49672 16632 0 _0678_
rlabel metal2 52808 22904 52808 22904 0 _0679_
rlabel metal2 51576 22680 51576 22680 0 _0680_
rlabel metal2 53704 24360 53704 24360 0 _0681_
rlabel metal2 47376 25704 47376 25704 0 _0682_
rlabel metal2 52024 28392 52024 28392 0 _0683_
rlabel metal3 46424 26264 46424 26264 0 _0684_
rlabel metal3 48832 27832 48832 27832 0 _0685_
rlabel metal2 47320 27384 47320 27384 0 _0686_
rlabel metal3 47040 38136 47040 38136 0 _0687_
rlabel metal2 47544 37744 47544 37744 0 _0688_
rlabel metal2 48440 40376 48440 40376 0 _0689_
rlabel metal2 47040 36680 47040 36680 0 _0690_
rlabel metal3 47992 37912 47992 37912 0 _0691_
rlabel metal2 23800 54600 23800 54600 0 _0692_
rlabel metal3 44296 45584 44296 45584 0 _0693_
rlabel metal2 48664 53816 48664 53816 0 _0694_
rlabel metal4 50344 51101 50344 51101 0 _0695_
rlabel metal2 50456 51856 50456 51856 0 _0696_
rlabel metal3 47376 49000 47376 49000 0 _0697_
rlabel metal3 47320 46648 47320 46648 0 _0698_
rlabel metal2 49336 51744 49336 51744 0 _0699_
rlabel metal2 48608 49000 48608 49000 0 _0700_
rlabel metal3 49112 49000 49112 49000 0 _0701_
rlabel metal2 43064 54208 43064 54208 0 _0702_
rlabel metal3 36792 51632 36792 51632 0 _0703_
rlabel metal3 32648 51576 32648 51576 0 _0704_
rlabel metal2 44632 51968 44632 51968 0 _0705_
rlabel metal2 43512 51800 43512 51800 0 _0706_
rlabel metal2 35616 39032 35616 39032 0 _0707_
rlabel metal3 44688 33992 44688 33992 0 _0708_
rlabel metal2 16128 11368 16128 11368 0 _0709_
rlabel metal2 17192 10080 17192 10080 0 _0710_
rlabel metal2 35784 26712 35784 26712 0 _0711_
rlabel metal3 37688 25704 37688 25704 0 _0712_
rlabel metal2 12096 8792 12096 8792 0 _0713_
rlabel metal2 13496 2772 13496 2772 0 _0714_
rlabel metal2 19096 12936 19096 12936 0 _0715_
rlabel metal2 35336 25872 35336 25872 0 _0716_
rlabel metal2 27048 4536 27048 4536 0 _0717_
rlabel metal2 20944 2744 20944 2744 0 _0718_
rlabel metal2 20944 5656 20944 5656 0 _0719_
rlabel metal3 20664 3752 20664 3752 0 _0720_
rlabel metal2 36904 5712 36904 5712 0 _0721_
rlabel metal3 36288 10584 36288 10584 0 _0722_
rlabel metal2 32872 5768 32872 5768 0 _0723_
rlabel metal2 34328 5208 34328 5208 0 _0724_
rlabel metal2 36792 4480 36792 4480 0 _0725_
rlabel metal2 14392 3808 14392 3808 0 _0726_
rlabel metal3 16968 2632 16968 2632 0 _0727_
rlabel metal3 9352 7336 9352 7336 0 _0728_
rlabel metal2 8232 5992 8232 5992 0 _0729_
rlabel metal2 52696 11200 52696 11200 0 _0730_
rlabel metal4 9016 53368 9016 53368 0 _0731_
rlabel metal3 12880 51128 12880 51128 0 _0732_
rlabel metal2 41888 25704 41888 25704 0 _0733_
rlabel metal3 49784 15960 49784 15960 0 _0734_
rlabel metal2 48664 13048 48664 13048 0 _0735_
rlabel metal2 46648 14616 46648 14616 0 _0736_
rlabel metal2 4200 49616 4200 49616 0 _0737_
rlabel metal3 6160 49784 6160 49784 0 _0738_
rlabel metal2 29904 30408 29904 30408 0 _0739_
rlabel metal3 19152 34104 19152 34104 0 _0740_
rlabel metal2 19096 34384 19096 34384 0 _0741_
rlabel metal3 10864 48776 10864 48776 0 _0742_
rlabel metal3 8176 47544 8176 47544 0 _0743_
rlabel metal2 20888 24360 20888 24360 0 _0744_
rlabel metal2 25144 24528 25144 24528 0 _0745_
rlabel metal3 16128 48328 16128 48328 0 _0746_
rlabel metal2 16408 43736 16408 43736 0 _0747_
rlabel metal2 16520 29120 16520 29120 0 _0748_
rlabel metal2 20944 28056 20944 28056 0 _0749_
rlabel metal2 5320 45136 5320 45136 0 _0750_
rlabel metal4 3528 49952 3528 49952 0 _0751_
rlabel metal2 34552 28448 34552 28448 0 _0752_
rlabel metal3 3808 41944 3808 41944 0 _0753_
rlabel metal2 4424 38976 4424 38976 0 _0754_
rlabel metal2 51856 34104 51856 34104 0 _0755_
rlabel metal2 50232 43344 50232 43344 0 _0756_
rlabel metal2 54600 42588 54600 42588 0 _0757_
rlabel metal2 8008 39536 8008 39536 0 _0758_
rlabel metal3 8344 38136 8344 38136 0 _0759_
rlabel metal2 7896 29904 7896 29904 0 _0760_
rlabel metal2 10584 30072 10584 30072 0 _0761_
rlabel metal2 5320 33824 5320 33824 0 _0762_
rlabel metal2 6328 29848 6328 29848 0 _0763_
rlabel metal2 13048 17024 13048 17024 0 _0764_
rlabel metal2 54824 46256 54824 46256 0 _0765_
rlabel metal2 42952 40880 42952 40880 0 _0766_
rlabel metal2 42952 42000 42952 42000 0 _0767_
rlabel metal2 39368 45640 39368 45640 0 _0768_
rlabel metal2 20160 53816 20160 53816 0 _0769_
rlabel metal2 20440 53088 20440 53088 0 _0770_
rlabel metal2 24808 53424 24808 53424 0 _0771_
rlabel metal2 27048 53200 27048 53200 0 _0772_
rlabel metal3 7112 36344 7112 36344 0 _0773_
rlabel metal2 31192 52752 31192 52752 0 _0774_
rlabel metal2 39816 44240 39816 44240 0 _0775_
rlabel metal2 42504 47208 42504 47208 0 _0776_
rlabel metal3 3528 32424 3528 32424 0 _0777_
rlabel metal2 5880 30240 5880 30240 0 _0778_
rlabel metal3 12600 27720 12600 27720 0 _0779_
rlabel metal2 12824 28056 12824 28056 0 _0780_
rlabel metal2 4480 25480 4480 25480 0 _0781_
rlabel metal2 4088 25621 4088 25621 0 _0782_
rlabel metal2 11032 42392 11032 42392 0 _0783_
rlabel metal2 1624 14560 1624 14560 0 _0784_
rlabel metal2 11592 11088 11592 11088 0 _0785_
rlabel metal2 17192 20664 17192 20664 0 _0786_
rlabel metal2 20664 12712 20664 12712 0 _0787_
rlabel metal2 20776 12880 20776 12880 0 _0788_
rlabel metal3 20888 12152 20888 12152 0 _0789_
rlabel metal2 19992 12880 19992 12880 0 _0790_
rlabel metal2 23016 13104 23016 13104 0 _0791_
rlabel metal2 23128 13384 23128 13384 0 _0792_
rlabel metal3 19488 11592 19488 11592 0 _0793_
rlabel metal2 19096 13888 19096 13888 0 _0794_
rlabel metal2 48048 19992 48048 19992 0 _0795_
rlabel metal2 32704 24696 32704 24696 0 _0796_
rlabel metal3 33152 25256 33152 25256 0 _0797_
rlabel metal2 33320 25368 33320 25368 0 _0798_
rlabel metal2 32424 22904 32424 22904 0 _0799_
rlabel metal2 23576 39928 23576 39928 0 _0800_
rlabel metal3 27888 6104 27888 6104 0 _0801_
rlabel metal3 27944 5320 27944 5320 0 _0802_
rlabel metal2 26824 4424 26824 4424 0 _0803_
rlabel metal2 26936 4816 26936 4816 0 _0804_
rlabel metal2 25648 6776 25648 6776 0 _0805_
rlabel metal2 26824 5208 26824 5208 0 _0806_
rlabel metal2 26264 5376 26264 5376 0 _0807_
rlabel metal2 26152 4816 26152 4816 0 _0808_
rlabel metal2 45192 19320 45192 19320 0 _0809_
rlabel metal2 44296 19432 44296 19432 0 _0810_
rlabel metal2 47432 10080 47432 10080 0 _0811_
rlabel metal2 16408 12488 16408 12488 0 _0812_
rlabel metal2 15792 10024 15792 10024 0 _0813_
rlabel metal2 16296 9128 16296 9128 0 _0814_
rlabel metal3 15736 10024 15736 10024 0 _0815_
rlabel metal2 17472 9800 17472 9800 0 _0816_
rlabel metal2 14952 8512 14952 8512 0 _0817_
rlabel metal2 16632 8568 16632 8568 0 _0818_
rlabel metal3 16968 9912 16968 9912 0 _0819_
rlabel metal2 49112 11536 49112 11536 0 _0820_
rlabel metal2 44184 25536 44184 25536 0 _0821_
rlabel metal2 12600 5600 12600 5600 0 _0822_
rlabel metal2 11816 6720 11816 6720 0 _0823_
rlabel metal2 11928 6216 11928 6216 0 _0824_
rlabel metal2 12208 5880 12208 5880 0 _0825_
rlabel metal3 12936 6776 12936 6776 0 _0826_
rlabel metal2 11704 6160 11704 6160 0 _0827_
rlabel metal2 10584 7056 10584 7056 0 _0828_
rlabel metal2 11480 6216 11480 6216 0 _0829_
rlabel metal2 46928 9016 46928 9016 0 _0830_
rlabel metal2 46088 13720 46088 13720 0 _0831_
rlabel metal3 46536 13048 46536 13048 0 _0832_
rlabel metal3 47656 8904 47656 8904 0 _0833_
rlabel metal2 54936 4704 54936 4704 0 _0834_
rlabel metal2 56112 4312 56112 4312 0 _0835_
rlabel metal2 36288 10024 36288 10024 0 _0836_
rlabel metal2 37016 6272 37016 6272 0 _0837_
rlabel metal3 34328 6944 34328 6944 0 _0838_
rlabel metal2 33208 5656 33208 5656 0 _0839_
rlabel metal2 33320 6048 33320 6048 0 _0840_
rlabel metal3 35280 6664 35280 6664 0 _0841_
rlabel metal2 34664 7336 34664 7336 0 _0842_
rlabel metal3 33880 6552 33880 6552 0 _0843_
rlabel metal2 33488 5320 33488 5320 0 _0844_
rlabel metal2 33824 6440 33824 6440 0 _0845_
rlabel metal3 36008 5880 36008 5880 0 _0846_
rlabel metal2 36456 9352 36456 9352 0 _0847_
rlabel metal2 36344 6160 36344 6160 0 _0848_
rlabel metal3 36232 11592 36232 11592 0 _0849_
rlabel metal2 39368 5488 39368 5488 0 _0850_
rlabel metal3 20440 16296 20440 16296 0 _0851_
rlabel metal2 36400 3416 36400 3416 0 _0852_
rlabel metal3 37408 3416 37408 3416 0 _0853_
rlabel metal2 38696 4424 38696 4424 0 _0854_
rlabel metal2 39256 5600 39256 5600 0 _0855_
rlabel metal2 17640 2072 17640 2072 0 _0856_
rlabel metal2 21560 2632 21560 2632 0 _0857_
rlabel metal2 20776 5152 20776 5152 0 _0858_
rlabel metal2 48888 54936 48888 54936 0 clknet_0_UserCLK
rlabel metal3 50232 33544 50232 33544 0 clknet_0_UserCLK_regs
rlabel metal2 48104 55496 48104 55496 0 clknet_1_0__leaf_UserCLK
rlabel metal2 48104 23072 48104 23072 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal3 49560 47768 49560 47768 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal3 35056 50008 35056 50008 0 net1
rlabel metal3 56560 23240 56560 23240 0 net10
rlabel metal2 53256 53984 53256 53984 0 net100
rlabel metal3 46256 46760 46256 46760 0 net101
rlabel metal3 19376 40376 19376 40376 0 net102
rlabel metal2 19768 44464 19768 44464 0 net103
rlabel metal3 22176 52920 22176 52920 0 net104
rlabel metal4 19320 42336 19320 42336 0 net105
rlabel metal2 20720 52920 20720 52920 0 net106
rlabel metal3 14168 47096 14168 47096 0 net107
rlabel metal2 5320 39368 5320 39368 0 net108
rlabel metal3 7056 41160 7056 41160 0 net109
rlabel metal3 56448 49560 56448 49560 0 net11
rlabel metal3 1848 49224 1848 49224 0 net110
rlabel metal2 1848 50008 1848 50008 0 net111
rlabel metal2 1512 53200 1512 53200 0 net112
rlabel metal3 18984 52808 18984 52808 0 net113
rlabel metal2 4984 32536 4984 32536 0 net114
rlabel metal2 13160 39396 13160 39396 0 net115
rlabel metal2 16968 40656 16968 40656 0 net116
rlabel metal2 7560 28616 7560 28616 0 net117
rlabel metal2 18760 44240 18760 44240 0 net118
rlabel metal3 16744 41552 16744 41552 0 net119
rlabel metal3 54040 22904 54040 22904 0 net12
rlabel metal3 1512 50736 1512 50736 0 net120
rlabel metal2 1176 54096 1176 54096 0 net121
rlabel metal3 6944 55384 6944 55384 0 net122
rlabel metal2 12488 55216 12488 55216 0 net123
rlabel metal3 11256 51352 11256 51352 0 net124
rlabel metal2 7336 55552 7336 55552 0 net125
rlabel metal2 9688 53704 9688 53704 0 net126
rlabel metal2 15848 53592 15848 53592 0 net127
rlabel metal2 13832 54824 13832 54824 0 net128
rlabel metal3 2604 54264 2604 54264 0 net129
rlabel metal2 56224 21560 56224 21560 0 net13
rlabel metal2 23576 53088 23576 53088 0 net130
rlabel metal2 24808 55216 24808 55216 0 net131
rlabel metal2 2632 55216 2632 55216 0 net132
rlabel metal2 25144 56224 25144 56224 0 net133
rlabel metal2 1960 55272 1960 55272 0 net134
rlabel metal3 8456 54488 8456 54488 0 net135
rlabel metal2 11032 54488 11032 54488 0 net136
rlabel metal2 11088 55384 11088 55384 0 net137
rlabel metal3 12208 55384 12208 55384 0 net138
rlabel metal2 20888 53704 20888 53704 0 net139
rlabel metal2 56168 15288 56168 15288 0 net14
rlabel metal3 20720 54376 20720 54376 0 net140
rlabel metal2 22904 55216 22904 55216 0 net141
rlabel metal2 19320 56112 19320 56112 0 net142
rlabel metal2 22288 55496 22288 55496 0 net143
rlabel metal2 25368 55608 25368 55608 0 net144
rlabel metal2 16072 54544 16072 54544 0 net145
rlabel metal3 15484 55384 15484 55384 0 net146
rlabel metal3 14392 55832 14392 55832 0 net147
rlabel metal2 19320 54040 19320 54040 0 net148
rlabel metal2 19768 54600 19768 54600 0 net149
rlabel metal2 54712 21112 54712 21112 0 net15
rlabel metal3 18536 55384 18536 55384 0 net150
rlabel metal2 20608 55496 20608 55496 0 net151
rlabel metal2 21224 54432 21224 54432 0 net152
rlabel metal3 20328 55384 20328 55384 0 net153
rlabel metal3 22904 4312 22904 4312 0 net154
rlabel metal2 20272 1176 20272 1176 0 net155
rlabel metal2 21168 1176 21168 1176 0 net156
rlabel metal2 21672 1288 21672 1288 0 net157
rlabel metal2 2632 1680 2632 1680 0 net158
rlabel metal2 23128 1568 23128 1568 0 net159
rlabel metal2 55944 21000 55944 21000 0 net16
rlabel metal2 24248 1624 24248 1624 0 net160
rlabel metal3 25592 1176 25592 1176 0 net161
rlabel metal2 25816 1232 25816 1232 0 net162
rlabel metal2 26152 1344 26152 1344 0 net163
rlabel metal2 26936 1848 26936 1848 0 net164
rlabel metal2 28056 1232 28056 1232 0 net165
rlabel metal2 29736 1456 29736 1456 0 net166
rlabel metal3 32256 952 32256 952 0 net167
rlabel metal3 31920 1064 31920 1064 0 net168
rlabel metal3 33600 3640 33600 3640 0 net169
rlabel metal2 56224 23016 56224 23016 0 net17
rlabel metal2 28952 2240 28952 2240 0 net170
rlabel metal3 30772 2072 30772 2072 0 net171
rlabel metal3 35784 1176 35784 1176 0 net172
rlabel metal2 35000 2996 35000 2996 0 net173
rlabel metal3 35112 33992 35112 33992 0 net174
rlabel metal3 38864 2744 38864 2744 0 net175
rlabel metal3 40768 2184 40768 2184 0 net176
rlabel metal2 41496 2352 41496 2352 0 net177
rlabel metal2 43512 1624 43512 1624 0 net178
rlabel metal2 39144 3528 39144 3528 0 net179
rlabel metal3 40936 27664 40936 27664 0 net18
rlabel metal2 45304 1288 45304 1288 0 net180
rlabel metal3 36176 54040 36176 54040 0 net181
rlabel metal2 38248 1512 38248 1512 0 net182
rlabel metal3 36848 2184 36848 2184 0 net183
rlabel metal3 35952 55832 35952 55832 0 net184
rlabel metal3 37240 55832 37240 55832 0 net185
rlabel metal3 38304 2184 38304 2184 0 net186
rlabel metal3 39200 55384 39200 55384 0 net187
rlabel metal3 38080 4312 38080 4312 0 net188
rlabel metal2 40040 1400 40040 1400 0 net189
rlabel metal2 30408 27440 30408 27440 0 net19
rlabel metal2 42504 2240 42504 2240 0 net190
rlabel metal2 47208 2352 47208 2352 0 net191
rlabel metal3 48832 2184 48832 2184 0 net192
rlabel metal3 46872 2520 46872 2520 0 net193
rlabel metal3 48104 3528 48104 3528 0 net194
rlabel metal2 40040 3920 40040 3920 0 net195
rlabel metal3 48216 5096 48216 5096 0 net196
rlabel metal2 43288 1624 43288 1624 0 net197
rlabel metal2 43960 2352 43960 2352 0 net198
rlabel metal2 47656 1400 47656 1400 0 net199
rlabel metal3 46928 21000 46928 21000 0 net2
rlabel metal2 56224 28840 56224 28840 0 net20
rlabel metal2 48664 1344 48664 1344 0 net200
rlabel metal3 43792 2632 43792 2632 0 net201
rlabel metal2 47320 2240 47320 2240 0 net202
rlabel metal2 49224 1568 49224 1568 0 net203
rlabel metal2 49896 1288 49896 1288 0 net204
rlabel metal2 46144 2632 46144 2632 0 net205
rlabel metal3 50008 55832 50008 55832 0 net206
rlabel metal2 15624 2464 15624 2464 0 net207
rlabel metal3 16128 1176 16128 1176 0 net208
rlabel metal3 13608 2184 13608 2184 0 net209
rlabel metal2 56392 29176 56392 29176 0 net21
rlabel metal2 11816 1848 11816 1848 0 net210
rlabel metal2 16520 2296 16520 2296 0 net211
rlabel metal2 13944 3640 13944 3640 0 net212
rlabel metal3 6664 952 6664 952 0 net213
rlabel metal2 13048 2912 13048 2912 0 net214
rlabel metal3 10192 3640 10192 3640 0 net215
rlabel metal2 2072 1512 2072 1512 0 net216
rlabel metal3 6328 1064 6328 1064 0 net217
rlabel metal3 10808 7672 10808 7672 0 net218
rlabel metal2 8344 3920 8344 3920 0 net219
rlabel metal3 53368 49448 53368 49448 0 net22
rlabel metal3 19992 4032 19992 4032 0 net220
rlabel metal2 4424 4088 4424 4088 0 net221
rlabel metal3 23744 5768 23744 5768 0 net222
rlabel metal2 16744 6440 16744 6440 0 net223
rlabel metal3 19432 5376 19432 5376 0 net224
rlabel metal3 7840 4200 7840 4200 0 net225
rlabel metal2 16184 2856 16184 2856 0 net226
rlabel metal3 15736 1008 15736 1008 0 net227
rlabel metal3 1568 18200 1568 18200 0 net228
rlabel metal3 1568 21448 1568 21448 0 net229
rlabel metal4 32872 51184 32872 51184 0 net23
rlabel metal2 16296 21952 16296 21952 0 net230
rlabel metal3 53648 15736 53648 15736 0 net231
rlabel metal2 24584 23912 24584 23912 0 net232
rlabel metal2 1568 13496 1568 13496 0 net233
rlabel metal3 40040 14224 40040 14224 0 net234
rlabel metal3 42616 18760 42616 18760 0 net235
rlabel metal2 46760 18424 46760 18424 0 net236
rlabel metal3 20888 18928 20888 18928 0 net237
rlabel metal2 50456 20776 50456 20776 0 net238
rlabel metal2 1960 1848 1960 1848 0 net239
rlabel metal2 39816 51688 39816 51688 0 net24
rlabel metal3 43624 4592 43624 4592 0 net240
rlabel metal2 50456 15512 50456 15512 0 net241
rlabel metal4 2072 22624 2072 22624 0 net242
rlabel metal2 3864 7280 3864 7280 0 net243
rlabel metal3 8624 15624 8624 15624 0 net244
rlabel metal3 7504 15176 7504 15176 0 net245
rlabel metal2 44072 840 44072 840 0 net246
rlabel metal2 55888 2184 55888 2184 0 net247
rlabel metal3 52304 2632 52304 2632 0 net248
rlabel metal4 1512 5320 1512 5320 0 net249
rlabel metal2 47544 39872 47544 39872 0 net25
rlabel metal3 17864 4592 17864 4592 0 net250
rlabel metal3 21000 12432 21000 12432 0 net251
rlabel metal2 55944 2744 55944 2744 0 net252
rlabel metal3 41832 3304 41832 3304 0 net253
rlabel metal3 13496 11704 13496 11704 0 net254
rlabel metal2 55104 47880 55104 47880 0 net26
rlabel metal2 49112 49924 49112 49924 0 net27
rlabel metal2 50904 44520 50904 44520 0 net28
rlabel metal2 15848 41160 15848 41160 0 net29
rlabel metal2 53424 18200 53424 18200 0 net3
rlabel metal3 15232 38696 15232 38696 0 net30
rlabel metal3 22344 41272 22344 41272 0 net31
rlabel metal2 2744 45864 2744 45864 0 net32
rlabel metal4 18536 48328 18536 48328 0 net33
rlabel metal2 56112 39816 56112 39816 0 net34
rlabel metal3 46480 40712 46480 40712 0 net35
rlabel metal2 54936 38752 54936 38752 0 net36
rlabel metal2 55272 50792 55272 50792 0 net37
rlabel metal2 54936 51296 54936 51296 0 net38
rlabel metal3 55440 48104 55440 48104 0 net39
rlabel metal2 47432 22344 47432 22344 0 net4
rlabel metal2 52360 51800 52360 51800 0 net40
rlabel metal2 56280 40488 56280 40488 0 net41
rlabel metal2 55328 44408 55328 44408 0 net42
rlabel metal3 55496 42952 55496 42952 0 net43
rlabel metal2 56280 41944 56280 41944 0 net44
rlabel metal2 52024 32984 52024 32984 0 net45
rlabel metal2 56280 49224 56280 49224 0 net46
rlabel metal2 55216 47656 55216 47656 0 net47
rlabel metal2 51128 37520 51128 37520 0 net48
rlabel metal3 55720 49224 55720 49224 0 net49
rlabel metal2 48776 20496 48776 20496 0 net5
rlabel metal3 44184 51800 44184 51800 0 net50
rlabel metal3 33152 37576 33152 37576 0 net51
rlabel metal2 44520 37800 44520 37800 0 net52
rlabel metal2 30856 55328 30856 55328 0 net53
rlabel metal2 49896 53368 49896 53368 0 net54
rlabel metal2 29120 55832 29120 55832 0 net55
rlabel metal3 44128 48440 44128 48440 0 net56
rlabel metal3 44352 48328 44352 48328 0 net57
rlabel metal2 52360 52864 52360 52864 0 net58
rlabel metal3 49448 52752 49448 52752 0 net59
rlabel metal2 53704 5824 53704 5824 0 net6
rlabel metal2 47320 53200 47320 53200 0 net60
rlabel metal2 44856 49616 44856 49616 0 net61
rlabel metal2 49112 53760 49112 53760 0 net62
rlabel metal2 46536 52640 46536 52640 0 net63
rlabel metal2 45976 53592 45976 53592 0 net64
rlabel metal2 47208 53760 47208 53760 0 net65
rlabel metal2 46536 53704 46536 53704 0 net66
rlabel metal2 46088 55272 46088 55272 0 net67
rlabel metal3 43680 54376 43680 54376 0 net68
rlabel metal2 45080 55384 45080 55384 0 net69
rlabel metal3 55720 10584 55720 10584 0 net7
rlabel metal3 42840 55384 42840 55384 0 net70
rlabel metal3 43288 54264 43288 54264 0 net71
rlabel metal2 52976 52136 52976 52136 0 net72
rlabel metal2 43848 55328 43848 55328 0 net73
rlabel metal2 41104 54488 41104 54488 0 net74
rlabel metal3 29288 52808 29288 52808 0 net75
rlabel metal3 43176 40880 43176 40880 0 net76
rlabel metal3 52696 48048 52696 48048 0 net77
rlabel metal2 50176 52696 50176 52696 0 net78
rlabel metal2 26152 55720 26152 55720 0 net79
rlabel metal3 46928 24472 46928 24472 0 net8
rlabel metal2 40992 52808 40992 52808 0 net80
rlabel metal3 28448 55944 28448 55944 0 net81
rlabel metal2 46200 43232 46200 43232 0 net82
rlabel metal2 53816 32928 53816 32928 0 net83
rlabel metal2 47656 53312 47656 53312 0 net84
rlabel metal2 45192 56392 45192 56392 0 net85
rlabel metal3 42616 56000 42616 56000 0 net86
rlabel metal2 43848 56168 43848 56168 0 net87
rlabel metal2 46760 55216 46760 55216 0 net88
rlabel metal4 48552 53816 48552 53816 0 net89
rlabel metal2 56000 16632 56000 16632 0 net9
rlabel metal3 40152 49224 40152 49224 0 net90
rlabel metal2 55888 26152 55888 26152 0 net91
rlabel metal3 44464 26600 44464 26600 0 net92
rlabel metal3 51352 55944 51352 55944 0 net93
rlabel metal2 34552 56616 34552 56616 0 net94
rlabel metal2 44296 56224 44296 56224 0 net95
rlabel metal2 26376 54600 26376 54600 0 net96
rlabel metal3 33824 48440 33824 48440 0 net97
rlabel metal4 41384 46144 41384 46144 0 net98
rlabel metal2 50456 49728 50456 49728 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 57456
<< end >>
