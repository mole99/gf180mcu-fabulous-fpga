* NGSPICE file created from RegFile.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VDD VSS W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_3155_ FrameData[19] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2106_ Inst_RegFile_32x4.mem\[26\]\[2\] B_ADR0 _0740_ _0741_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3086_ FrameData[14] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2037_ _1340_ B_ADR0 _0674_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2939_ FrameData[27] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1606_ AD3 BD0 BD2 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ _0263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2724_ Inst_RegFile_32x4.mem\[18\]\[3\] _1198_ _1229_ _0063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2655_ Inst_RegFile_32x4.mem\[27\]\[3\] _1198_ _1208_ _0015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2586_ _1150_ _1152_ _1154_ _0141_ _1155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1537_ N2END[5] E2END[5] SS4END[1] W2END[5] Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q _0197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1468_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0131_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3207_ FrameData[7] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1399_ W6END[0] _1290_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3069_ FrameData[29] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3138_ FrameData[2] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_5_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q _0935_ _1033_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ _1034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2371_ N1END[3] E1END[3] W1END[3] AD2 Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q _0976_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2638_ Inst_RegFile_32x4.mem\[25\]\[0\] _1182_ _1202_ _0004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2569_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0931_ _1137_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ _1138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2707_ _1184_ Inst_RegFile_32x4.mem\[14\]\[1\] _1226_ _0049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput242 net242 WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput220 net220 W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput231 net231 W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput253 net253 WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_559 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1871_ _1265_ _0514_ _1271_ _0515_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1940_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q _0575_ _0578_ _0565_ _0568_ _0581_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_16_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3472_ N2MID[4] net117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2423_ N2END[2] S2END[2] E2END[2] WW4END[2] Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q _1019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_43_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3541_ Inst_RegFile_switch_matrix.S4BEG1 net177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2285_ AD3 BD0 BD1 BD2 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ _0900_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2354_ N2END[0] S2END[0] E2END[0] WW4END[3] Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q _0961_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_529 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2070_ Inst_RegFile_32x4.mem\[0\]\[2\] B_ADR0 _0705_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2972_ FrameData[28] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1785_ _1334_ A_ADR0 _0434_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1854_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _0293_ _0499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1923_ _1287_ Inst_RegFile_switch_matrix.JS2BEG6 _0564_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3386_ Inst_RegFile_switch_matrix.E6BEG0 net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3455_ FrameStrobe[19] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2406_ N1END[0] E1END[0] S1END[0] AD3 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q _1006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3524_ S2MID[4] net169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2268_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0884_ _0883_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q
+ _0885_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2337_ _0468_ _0946_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q _0947_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2199_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0823_ _0824_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_5 FrameStrobe[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3240_ FrameData[8] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1570_ E6END[0] S2END[4] S4END[0] W2END[4] Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q _0229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2122_ _1252_ _0754_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q _0755_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3171_ FrameData[3] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2053_ _0550_ _0684_ _0689_ _0690_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_60_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2955_ FrameData[11] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3507_ Inst_RegFile_switch_matrix.NN4BEG3 net143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1768_ _1321_ A_ADR0 _0419_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1837_ _0478_ _0480_ _0482_ _1260_ _0483_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1906_ _0545_ _0547_ _0548_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2886_ FrameData[6] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3438_ FrameStrobe[2] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3369_ E2MID[1] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1699_ _0348_ _0349_ _0351_ _0180_ _0219_ _0352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput31 net31 E6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput75 net75 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput64 net64 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput53 net53 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput42 net42 EE4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput20 net20 E2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput7 net7 E2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput86 net86 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput97 net97 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1622_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q _0277_ _0278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2740_ _1207_ _1221_ _1233_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2671_ Inst_RegFile_32x4.mem\[30\]\[1\] _1184_ _1214_ _0025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3223_ FrameData[23] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1553_ Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q _0209_ _0211_ _0212_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1484_ A_ADR0 _0147_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3154_ FrameData[18] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2105_ _1323_ B_ADR0 _0740_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3085_ FrameData[13] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2036_ _0670_ _0672_ _0486_ _0673_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2938_ FrameData[26] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_465 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2869_ _0063_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[18\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ Inst_RegFile_32x4.mem\[18\]\[2\] _1186_ _1229_ _0062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1605_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _0261_ _0262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2585_ _1269_ Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ _1153_ _1154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2654_ Inst_RegFile_32x4.mem\[27\]\[2\] _1186_ _1208_ _0014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1536_ N4END[1] W2END[4] SS4END[1] Inst_RegFile_switch_matrix.JS2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q _0196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1398_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _1289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1467_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3137_ FrameData[1] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3206_ FrameData[6] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2019_ _0580_ _0627_ _0638_ _0648_ _0657_ Inst_RegFile_32x4.BD_comb\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3068_ FrameData[28] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2370_ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q _0972_ _0974_ _0975_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_538 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2706_ _1182_ Inst_RegFile_32x4.mem\[14\]\[0\] _1226_ _0048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Left_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1519_ _0162_ _0179_ _0180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2637_ _1135_ _1201_ _1202_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2568_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _1136_ _1137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2499_ BD1 _0468_ Inst_RegFile_switch_matrix.JN2BEG1 _0530_ Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q Inst_RegFile_switch_matrix.E1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput232 net232 W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput210 net210 W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput243 net243 WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput221 net221 W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1870_ NN4END[1] E2END[5] S2END[5] W2END[5] Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q _0514_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3540_ Inst_RegFile_switch_matrix.S4BEG0 net176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2422_ _1018_ _1017_ Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q Inst_RegFile_switch_matrix.NN4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3471_ N2MID[3] net116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2353_ _0960_ _0959_ Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q Inst_RegFile_switch_matrix.WW4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2284_ W1END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ _0899_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1999_ _0631_ _0632_ _0637_ _0517_ _0550_ _0638_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_6_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_70_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_switch_matrix.JW2BEG6
+ _0563_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2971_ FrameData[27] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1853_ _1265_ _0497_ _0498_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1784_ _0424_ _0427_ _0432_ _0218_ _0254_ _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3523_ S2MID[3] net168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3454_ FrameStrobe[18] net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3385_ E6END[11] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2405_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q _1002_ _1004_ _1005_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2336_ N2END[4] E2END[4] SS4END[2] W2END[4] Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q _0946_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2267_ W1END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ _0884_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2198_ W6END[0] AD0 AD2 AD3 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ _0823_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_63_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_6 FrameStrobe[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3170_ FrameData[2] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ AD3 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ _0754_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2052_ _0486_ _0688_ _0686_ _0517_ _0689_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2954_ FrameData[10] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2885_ FrameData[5] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1905_ _1273_ _0546_ _0547_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3506_ Inst_RegFile_switch_matrix.NN4BEG2 net142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1836_ _1261_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ _0481_ _0482_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1767_ Inst_RegFile_32x4.mem\[20\]\[2\] A_ADR0 _0417_ _0418_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1698_ Inst_RegFile_32x4.mem\[4\]\[1\] A_ADR0 _0350_ _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3437_ FrameStrobe[1] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3299_ Inst_RegFile_32x4.BD_comb\[3\] clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.BD_reg\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3368_ E2MID[0] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2319_ _0930_ _0931_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput98 net98 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput65 net65 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput32 net32 E6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput21 net21 E6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput43 net43 EE4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput87 net87 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput54 net54 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput76 net76 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput10 net10 E2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput8 net8 E2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1621_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q _0275_ _0276_ _0277_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1552_ _1267_ Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q
+ _0210_ _0211_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2670_ Inst_RegFile_32x4.mem\[30\]\[0\] _1182_ _1214_ _0024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3222_ FrameData[22] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3153_ FrameData[17] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2104_ Inst_RegFile_32x4.mem\[24\]\[2\] B_ADR0 _0738_ _0739_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1483_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q _0146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2035_ Inst_RegFile_32x4.mem\[26\]\[3\] B_ADR0 _0671_ _0672_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3084_ FrameData[12] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2868_ _0062_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[18\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2937_ FrameData[25] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_20_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1819_ Inst_RegFile_32x4.AD_comb\[3\] Inst_RegFile_32x4.AD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2799_ _1186_ Inst_RegFile_32x4.mem\[11\]\[2\] _1245_ _0122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2722_ Inst_RegFile_32x4.mem\[18\]\[1\] _1184_ _1229_ _0061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1604_ W1END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ _0261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2584_ E2END[3] Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q _1153_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2653_ Inst_RegFile_32x4.mem\[27\]\[1\] _1184_ _1208_ _0013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1535_ Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q _0192_ _0194_ _0195_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3067_ FrameData[27] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1466_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q _0129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1397_ W2END[4] _1288_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3136_ FrameData[0] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3205_ FrameData[5] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2018_ _0550_ _0656_ _0580_ _0657_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2636_ _1142_ _1149_ _1170_ _1201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput200 net200 SS4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2705_ _1203_ _1218_ _1226_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1518_ _0173_ _0176_ _0177_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ _0179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2498_ Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q _1078_ _1076_ Inst_RegFile_switch_matrix.E1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2567_ N2MID[2] W2MID[2] E2MID[2] Inst_RegFile_switch_matrix.E2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q _1136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1449_ Inst_RegFile_32x4.mem\[31\]\[3\] _1340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput211 net211 W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput244 net244 WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput222 net222 W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput233 net233 W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3119_ FrameData[15] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_2_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_14_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_23_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ N2MID[2] net115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2421_ N1END[1] E1END[1] W1END[1] AD0 Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q _1018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_43_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2352_ N1END[2] S1END[2] W1END[2] AD1 Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ _0960_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_29_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q _0896_ _0898_ _0892_ _0894_ Inst_RegFile_switch_matrix.E2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_52_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0486_ _0634_ _0636_ _0637_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2619_ _0921_ _0943_ _0572_ _1185_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q
+ _1186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3599_ WW4END[10] net250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_58_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1921_ _0562_ _0559_ Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q Inst_RegFile_switch_matrix.JN2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1852_ E2MID[4] S2MID[4] W2MID[4] Inst_RegFile_switch_matrix.JS2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q _0497_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_29_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2970_ FrameData[26] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3453_ FrameStrobe[17] net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1783_ _0429_ _0431_ _0181_ _0432_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3522_ S2MID[2] net167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3384_ E6END[10] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2266_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0882_ _0883_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2404_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q _0160_ _1003_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ _1004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2335_ _0945_ _0944_ Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q Inst_RegFile_switch_matrix.WW4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2197_ _0816_ _0818_ _0820_ _0822_ Inst_RegFile_switch_matrix.JN2BEG2 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_7 FrameStrobe[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2120_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0752_ _0753_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2051_ _1327_ B_ADR0 _0687_ _0688_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1835_ N4END[2] Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q _0481_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2953_ FrameData[9] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2884_ FrameData[4] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1904_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q _0546_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3436_ FrameStrobe[0] net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3505_ Inst_RegFile_switch_matrix.NN4BEG1 net141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1766_ _1320_ A_ADR0 _0417_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1697_ _1301_ A_ADR0 _0350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3367_ Inst_RegFile_switch_matrix.E2BEG7 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2249_ W1END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ _0868_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3298_ Inst_RegFile_32x4.BD_comb\[2\] clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.BD_reg\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2318_ N2MID[3] E2MID[3] S2MID[3] W2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q _0930_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_23_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput99 net99 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput55 net55 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput66 net66 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput44 net44 EE4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput88 net88 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput33 net33 EE4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput22 net22 E6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput77 net77 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput9 net9 E2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput11 net11 E2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1352_ Inst_RegFile_switch_matrix.JS2BEG5 _0276_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1551_ Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q Inst_RegFile_switch_matrix.JS2BEG5
+ _0210_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1482_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q _0145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3221_ FrameData[21] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3152_ FrameData[16] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2103_ _1322_ B_ADR0 _0738_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3083_ FrameData[11] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ _1338_ B_ADR0 _0671_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2936_ FrameData[24] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2867_ _0061_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[18\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1818_ _0300_ _0455_ _0466_ _0433_ _0444_ Inst_RegFile_32x4.AD_comb\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2798_ _1184_ Inst_RegFile_32x4.mem\[11\]\[1\] _1245_ _0121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3419_ FrameData[15] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1749_ _1323_ _0147_ _0399_ _0400_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_559 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2721_ Inst_RegFile_32x4.mem\[18\]\[0\] _1182_ _1229_ _0060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2652_ Inst_RegFile_32x4.mem\[27\]\[0\] _1182_ _1208_ _0012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1465_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2583_ _1151_ _1152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1603_ _0183_ _0222_ _0259_ _0218_ _0254_ _0260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1534_ _1288_ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ _0193_ _0194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3204_ FrameData[4] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3066_ FrameData[26] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3135_ FrameData[31] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1396_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _1287_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2017_ _0651_ _0655_ _0517_ _0656_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ FrameData[7] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_56_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2704_ Inst_RegFile_32x4.mem\[23\]\[3\] _1198_ _1225_ _0047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2635_ _1141_ _1199_ _1200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput212 net212 W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput201 net201 SS4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput223 net223 W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput234 net234 W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1517_ _0177_ _0178_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2497_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q BD2 _1077_ _1078_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2566_ _1122_ _1134_ _1135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput245 net245 WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1448_ Inst_RegFile_32x4.mem\[29\]\[3\] _1339_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1379_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q _1270_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3049_ FrameData[9] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3118_ FrameData[14] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_2_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_529 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ BD0 _0213_ _0497_ _1016_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ _1017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2351_ BD1 _0930_ _0936_ _0514_ Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q
+ _0959_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2282_ _0135_ _0897_ _0898_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1997_ Inst_RegFile_32x4.mem\[29\]\[1\] B_ADR0 _0486_ _0635_ _0636_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_15_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3598_ WW4END[9] net249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2549_ _0144_ _1058_ _1118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2618_ N4END[1] W6END[1] E6END[1] Inst_RegFile_switch_matrix.JS2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q _1185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_58_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_28_Left_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1851_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q _0494_ _0496_ _0490_ _0492_ Inst_RegFile_switch_matrix.JS2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1920_ _0560_ _0561_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q _0562_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_12_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3383_ E6END[9] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3452_ FrameStrobe[16] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2403_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q BD3 _1003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1782_ _1340_ _0147_ _0430_ _0431_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3521_ S2MID[1] net166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2265_ _0881_ _0882_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2196_ _0128_ _0821_ _0129_ _0822_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2334_ N1END[1] S1END[1] W1END[1] AD0 Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ _0945_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_8 FrameStrobe[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ Inst_RegFile_32x4.mem\[4\]\[3\] B_ADR0 _0687_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_2_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_2_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2952_ FrameData[8] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2883_ FrameData[3] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1834_ _0479_ _0480_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1765_ _0180_ _0415_ _0413_ _0218_ _0416_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1903_ Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q _0542_ _0544_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q
+ _0545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3504_ Inst_RegFile_switch_matrix.NN4BEG0 net140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3435_ FrameData[31] net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3366_ Inst_RegFile_switch_matrix.E2BEG6 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1696_ Inst_RegFile_32x4.mem\[7\]\[1\] A_ADR0 _0162_ _0179_ _0349_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2248_ AD3 BD0 BD1 BD2 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ _0867_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_68_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ Inst_RegFile_32x4.BD_comb\[1\] clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.BD_reg\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2179_ _0806_ _0803_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q Inst_RegFile_switch_matrix.JS2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2317_ AD0 AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ _0929_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput34 net34 EE4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput23 net23 E6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput12 net12 E2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput89 net89 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput67 net67 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput56 net56 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput78 net78 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput45 net45 EE4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3220_ FrameData[20] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1550_ N2MID[4] S2MID[4] Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q _0209_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q _0144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3151_ FrameData[15] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2102_ _0550_ _0731_ _0736_ _0737_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3082_ FrameData[10] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2033_ Inst_RegFile_32x4.mem\[24\]\[3\] B_ADR0 _0669_ _0670_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2935_ FrameData[23] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2866_ _0060_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[18\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1748_ Inst_RegFile_32x4.mem\[26\]\[2\] _0147_ _0399_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_15_Left_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1817_ _0253_ _0460_ _0465_ _0466_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2797_ _1182_ Inst_RegFile_32x4.mem\[11\]\[0\] _1245_ _0120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3418_ FrameData[14] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3349_ _0121_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[11\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1679_ Inst_RegFile_32x4.AD_comb\[0\] Inst_RegFile_32x4.AD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2582_ WW4END[2] Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ _1151_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2720_ _1204_ _1221_ _1229_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1602_ _0256_ _0258_ _0181_ _0259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2651_ _1135_ _1207_ _1208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1464_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _1355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1533_ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q Inst_RegFile_switch_matrix.JS2BEG3
+ _0193_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1395_ Inst_RegFile_32x4.mem\[15\]\[0\] _1286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3203_ FrameData[3] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_70_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3065_ FrameData[25] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3134_ FrameData[30] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2016_ _0654_ _0652_ _0486_ _0655_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2918_ FrameData[6] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2849_ _0043_ clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.mem\[22\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_519 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1516_ N2END[3] E2END[3] S2END[3] WW4END[1] Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q _0177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2703_ Inst_RegFile_32x4.mem\[23\]\[2\] _1186_ _1225_ _0046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2634_ _1149_ _1170_ _1199_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2565_ _1132_ _1131_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _1134_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput213 net213 W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput246 net246 WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput224 net224 W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput202 net202 SS4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput235 net235 W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1378_ SS4END[3] _1269_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2496_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q _0573_ _1077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3117_ FrameData[13] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1447_ Inst_RegFile_32x4.mem\[27\]\[3\] _1338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3048_ FrameData[8] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_2_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_69_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2281_ E2END[1] S2END[1] E6END[1] W2END[1] Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q _0897_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2350_ _0958_ _0957_ Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q Inst_RegFile_switch_matrix.WW4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1996_ _1309_ B_ADR0 _0635_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_15_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2617_ Inst_RegFile_32x4.mem\[24\]\[1\] _1184_ _1174_ _0001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3597_ WW4END[8] net248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2548_ _0144_ _1114_ _1117_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_58_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q BD3 _1063_ _0139_ _1064_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_66_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkload0 clknet_4_0_0_UserCLK_regs clkload0/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_11_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_10_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_3_Left_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_541 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _1266_ _0495_ _0496_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3520_ S2MID[0] net165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1781_ Inst_RegFile_32x4.mem\[30\]\[3\] _0147_ _0430_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3451_ FrameStrobe[15] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3382_ E6END[8] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2402_ _0468_ _1001_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q _1002_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2333_ BD0 _0213_ _0497_ _0943_ Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ _0944_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2264_ AD3 BD0 BD1 BD2 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ _0881_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2195_ E6END[1] S2END[3] W2END[3] WW4END[2] Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q _0821_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1979_ _1304_ B_ADR0 _0618_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_9 N2MID[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2951_ FrameData[7] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1902_ _1274_ Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q
+ _0543_ _0544_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_15_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q W2END[2] Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ _0479_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1764_ Inst_RegFile_32x4.mem\[16\]\[2\] A_ADR0 _0414_ _0415_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2882_ FrameData[2] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3503_ NN4END[15] net139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3434_ FrameData[30] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3296_ Inst_RegFile_32x4.BD_comb\[0\] clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.BD_reg\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2316_ NN4END[1] E1END[3] SS4END[1] W1END[3] Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0928_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3365_ Inst_RegFile_switch_matrix.E2BEG5 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1695_ Inst_RegFile_32x4.mem\[6\]\[1\] _0147_ _0348_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2178_ _0805_ _0804_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0806_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2247_ _0866_ _0863_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q Inst_RegFile_switch_matrix.JW2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_23_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput35 net35 EE4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput57 net57 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput46 net46 EE4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput24 net24 E6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput13 net13 E2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput68 net68 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput79 net79 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3150_ FrameData[14] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q _0143_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2101_ _0486_ _0735_ _0733_ _0517_ _0736_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3081_ FrameData[9] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2032_ _1337_ B_ADR0 _0669_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2934_ FrameData[22] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2865_ _0059_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[16\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1678_ _0300_ _0321_ _0332_ _0311_ _0260_ Inst_RegFile_32x4.AD_comb\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1816_ _0461_ _0462_ _0464_ _0180_ _0219_ _0465_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2796_ _1206_ _1216_ _1245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1747_ _0390_ _0393_ _0397_ _0218_ _0253_ _0398_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3417_ FrameData[13] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3279_ FrameData[15] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3348_ _0120_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[11\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_503 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_521 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_539 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2581_ _0816_ _0818_ _0820_ _0822_ Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q _1150_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1601_ _1299_ _0147_ _0257_ _0258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2650_ _1141_ _1149_ _1170_ _1207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1532_ N4END[1] SS4END[1] Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q _0192_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_517 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q _1354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3133_ FrameData[29] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1394_ Inst_RegFile_32x4.mem\[13\]\[0\] _1285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3202_ FrameData[2] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3064_ FrameData[24] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_33_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2015_ _1303_ B_ADR0 _0653_ _0654_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2848_ _0042_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[22\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2917_ FrameData[5] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2779_ _1186_ Inst_RegFile_32x4.mem\[7\]\[2\] _1241_ _0106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2702_ Inst_RegFile_32x4.mem\[23\]\[1\] _1184_ _1225_ _0045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1515_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _0175_ _0176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2495_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q Inst_RegFile_switch_matrix.JN2BEG2
+ _1075_ Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q _1076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2633_ Inst_RegFile_32x4.mem\[24\]\[3\] _1198_ _1174_ _0003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput236 net236 W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2564_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _1131_ _1125_ _1133_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput225 net225 W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput214 net214 W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput203 net203 SS4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput247 net247 WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3116_ FrameData[12] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1377_ WW4END[3] _1268_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1446_ Inst_RegFile_32x4.mem\[25\]\[3\] _1337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3047_ FrameData[7] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_11_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_528 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2280_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0895_ _0896_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2616_ _0570_ _0936_ _1016_ _1183_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q
+ _1184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1995_ Inst_RegFile_32x4.mem\[30\]\[1\] B_ADR0 _0633_ _0634_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1429_ Inst_RegFile_32x4.mem\[21\]\[2\] _1320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2478_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q _0573_ _1063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3596_ WW4END[7] net247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2547_ _1109_ _1111_ _1113_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q _1116_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_66_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkload1 clknet_4_1_0_UserCLK_regs clkload1/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ _1339_ _0147_ _0428_ _0429_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3450_ FrameStrobe[14] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3381_ E6END[7] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2401_ NN4END[3] E2END[6] S2END[6] W2END[6] Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q _1001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2332_ N2END[4] S2END[4] EE4END[0] W2END[4] Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q _0943_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2194_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0819_ _0820_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2263_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q _0878_ _0880_ _0874_ _0876_ Inst_RegFile_switch_matrix.JS2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_63_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1978_ Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q _0616_ _0617_ BD0 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3579_ W2MID[6] net224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1832_ _0471_ _0473_ _0475_ _0477_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q _0478_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2881_ _0075_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[21\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ FrameData[6] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1901_ N2MID[0] Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q _0543_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3433_ FrameData[29] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1763_ _1318_ A_ADR0 _0414_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3502_ NN4END[14] net138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1694_ _0345_ _0346_ _0180_ _0347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2315_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q _0912_ _0914_ _0925_ _0927_ Inst_RegFile_switch_matrix.W6BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3364_ Inst_RegFile_switch_matrix.E2BEG4 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3295_ FrameData[31] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2246_ _0864_ _0865_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0866_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2177_ N2END[3] E2END[3] E1END[1] EE4END[2] Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput69 net69 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput58 net58 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput25 net25 E6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput47 net47 EE4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput36 net36 EE4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput14 net14 E2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ _1320_ B_ADR0 _0734_ _0735_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3080_ FrameData[8] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2031_ _0550_ _0662_ _0667_ _0668_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ FrameData[21] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2864_ _0058_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[16\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1815_ Inst_RegFile_32x4.mem\[4\]\[3\] A_ADR0 _0463_ _0464_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2795_ _1198_ Inst_RegFile_32x4.mem\[10\]\[3\] _1244_ _0119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3416_ FrameData[12] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1677_ _0323_ _0326_ _0331_ _0218_ _0254_ _0332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1746_ _0394_ _0396_ _0181_ _0397_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2229_ EE4END[1] E6END[0] S2END[2] W2END[2] Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q _0851_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3347_ _0119_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[10\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3278_ FrameData[14] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1462_ S2END[0] _1353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1531_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q _0189_ _0191_ _0185_ _0187_ Inst_RegFile_switch_matrix.JS2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2580_ _1148_ _1147_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q _1149_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ Inst_RegFile_32x4.mem\[30\]\[0\] _0147_ _0257_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3132_ FrameData[28] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3063_ FrameData[23] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3201_ FrameData[1] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1393_ Inst_RegFile_32x4.mem\[11\]\[0\] _1284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2014_ Inst_RegFile_32x4.mem\[12\]\[1\] B_ADR0 _0653_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2847_ _0041_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[22\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2916_ FrameData[4] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2778_ _1184_ Inst_RegFile_32x4.mem\[7\]\[1\] _1241_ _0105_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1729_ _0162_ _0179_ _0378_ _0379_ _0380_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_46_529 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2701_ Inst_RegFile_32x4.mem\[23\]\[0\] _1182_ _1225_ _0044_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2632_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q _1195_ _1197_ _1190_ _1191_ _1198_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1514_ NN4END[2] Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q _0174_ _0175_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1445_ Inst_RegFile_32x4.mem\[22\]\[3\] _1336_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q _1041_ _1075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2563_ _0142_ _0922_ _1124_ _1132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput215 net215 W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput248 net248 WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput204 net204 SS4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput237 net237 W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput226 net226 W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3115_ FrameData[11] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1376_ W2MID[4] _1267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3046_ FrameData[6] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1994_ _1310_ B_ADR0 _0633_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2615_ EE4END[2] W2END[7] S4END[2] Inst_RegFile_switch_matrix.E2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q _1183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3595_ WW4END[6] net246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1428_ Inst_RegFile_32x4.mem\[18\]\[2\] _1319_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2546_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q _1113_ _1115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2477_ E6END[1] S4END[1] S2END[2] AD0 Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q Inst_RegFile_switch_matrix.S4BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_66_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1359_ WW4END[0] _1250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3029_ FrameData[21] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkload2 clknet_4_2_0_UserCLK_regs clkload2/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_42_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2400_ _1000_ _0999_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q Inst_RegFile_switch_matrix.EE4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ E6END[6] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2331_ _0928_ _0929_ _0942_ _0941_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q
+ Inst_RegFile_switch_matrix.W6BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2262_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0879_ _0880_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2193_ N2END[3] E1END[1] N4END[3] E2END[3] Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q _0819_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1977_ Inst_RegFile_32x4.BD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q _0617_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2529_ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q Inst_RegFile_switch_matrix.JW2BEG3
+ _1098_ Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q _1099_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3578_ W2MID[5] net223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0471_ _0473_ _0475_ _0477_ Inst_RegFile_switch_matrix.E2BEG4 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2880_ _0074_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[21\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1900_ W2MID[0] Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q
+ _0542_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3432_ FrameData[28] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1762_ Inst_RegFile_32x4.mem\[19\]\[2\] A_ADR0 _0162_ _0179_ _0412_ _0413_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3363_ Inst_RegFile_switch_matrix.E2BEG3 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3501_ NN4END[13] net152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1693_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] A_ADR0 _0346_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_69_Left_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2176_ E6END[1] S2END[3] S4END[3] W2END[3] Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q _0804_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2314_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q _0926_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q
+ _0927_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3294_ FrameData[30] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2245_ S2END[1] S4END[1] SS4END[0] W2END[1] Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q _0865_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput37 net37 EE4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput59 net59 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput26 net26 E6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput48 net48 EE4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput15 net15 E2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ _0486_ _0666_ _0664_ _0517_ _0667_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2932_ FrameData[20] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2863_ _0057_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[16\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1745_ _1313_ A_ADR0 _0395_ _0396_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1814_ _1327_ A_ADR0 _0463_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2794_ _1186_ Inst_RegFile_32x4.mem\[10\]\[2\] _1244_ _0118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3415_ FrameData[11] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _0328_ _0330_ _0181_ _0331_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3346_ _0118_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[10\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2228_ N2END[2] E1END[0] N4END[2] E2END[2] Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q _0850_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2159_ Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q _0788_ _0787_ _0789_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3277_ FrameData[13] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_505 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1461_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _1352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1530_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _0190_ _0191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1392_ Inst_RegFile_32x4.mem\[9\]\[0\] _1283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3200_ FrameData[0] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3131_ FrameData[27] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3062_ FrameData[22] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2013_ Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] B_ADR0 _0652_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2915_ FrameData[3] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2846_ _0040_ clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.mem\[22\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1728_ Inst_RegFile_32x4.mem\[8\]\[2\] _0147_ _0379_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2777_ _1182_ Inst_RegFile_32x4.mem\[7\]\[0\] _1241_ _0104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3329_ _0101_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[6\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1659_ _1253_ A_ADR0 _0314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput205 net205 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2700_ _1207_ _1223_ _1225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2562_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q _0946_ _1130_ _1131_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2631_ _0138_ _1196_ _1197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput216 net216 W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1513_ _1344_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q
+ _0174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1375_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _1266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1444_ Inst_RegFile_32x4.mem\[21\]\[3\] _1335_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput227 net227 W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput249 net249 WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput238 net238 WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2493_ _1072_ _1074_ Inst_RegFile_switch_matrix.S1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3114_ FrameData[10] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3045_ FrameData[5] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0023_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[2\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Left_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_60_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1993_ _0517_ _0629_ _0632_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_15_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2614_ Inst_RegFile_32x4.mem\[24\]\[0\] _1182_ _1174_ _0000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3594_ WW4END[5] net245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2545_ N2MID[0] W2MID[0] S2MID[0] Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q _1114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_7_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1427_ Inst_RegFile_32x4.mem\[17\]\[2\] _1318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1358_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q _1249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2476_ E6END[0] S2END[3] S4END[2] AD1 Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q Inst_RegFile_switch_matrix.S4BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ FrameData[20] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkload3 clknet_4_3_0_UserCLK_regs clkload3/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ _0128_ _0817_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q _0818_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2330_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ _0942_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2261_ N2END[1] E2END[1] E1END[3] E6END[1] Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q _0879_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_63_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1976_ _0616_ Inst_RegFile_32x4.BD_comb\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_536 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q _1053_ _1098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3577_ W2MID[4] net222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2459_ _1047_ _1049_ Inst_RegFile_switch_matrix.W1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _1319_ A_ADR0 _0412_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1830_ _1262_ _0476_ _1263_ _0477_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ NN4END[12] net151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3431_ FrameData[27] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2313_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ _0926_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1692_ _1300_ A_ADR0 _0344_ _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3362_ Inst_RegFile_switch_matrix.E2BEG2 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2175_ _0802_ _0801_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q _0803_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3293_ FrameData[29] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2244_ N1END[3] N2END[1] E2END[1] E6END[1] Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q _0864_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_23_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1959_ _1272_ B_ADR0 _0486_ _0599_ _0600_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput27 net27 E6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput49 net49 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput38 net38 EE4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput16 net16 E2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2931_ FrameData[19] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2862_ _0056_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[16\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1744_ Inst_RegFile_32x4.mem\[7\]\[2\] A_ADR0 _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1813_ Inst_RegFile_32x4.mem\[7\]\[3\] A_ADR0 _0162_ _0179_ _0462_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2793_ _1184_ Inst_RegFile_32x4.mem\[10\]\[1\] _1244_ _0117_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3414_ FrameData[10] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_517 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3276_ FrameData[12] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1675_ _1286_ _0147_ _0329_ _0330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3345_ _0117_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[10\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2227_ _0847_ _0848_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0849_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2158_ N2MID[7] E2MID[7] Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q _0788_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _0723_ _0721_ _0486_ _0724_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_509 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ FrameData[26] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1460_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _1351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1391_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q _1282_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3061_ FrameData[21] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2012_ _0650_ _0649_ _0486_ _0651_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2845_ _0039_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[17\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ FrameData[2] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1658_ _1264_ A_ADR0 _0181_ _0312_ _0313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2776_ _1206_ _1237_ _1241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1727_ Inst_RegFile_32x4.mem\[9\]\[2\] A_ADR0 _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1589_ _1348_ _0244_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q _0247_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3259_ FrameData[27] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3328_ _0100_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[6\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1512_ Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q _0171_ _0172_ _0173_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2561_ _1126_ _1127_ _1129_ Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q
+ _1130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput206 net206 W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2630_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q _1196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput217 net217 W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput239 net239 WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput228 net228 W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2492_ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q Inst_RegFile_switch_matrix.E2BEG3
+ _1073_ Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q _1074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1443_ Inst_RegFile_32x4.mem\[18\]\[3\] _1334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3113_ FrameData[9] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1374_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _1265_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ FrameData[4] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_18_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2828_ _0022_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[2\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ _1198_ Inst_RegFile_32x4.mem\[3\]\[3\] _1236_ _0091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkload10 clknet_4_12_0_UserCLK_regs clkload10/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_1992_ _1308_ B_ADR0 _0486_ _0630_ _0631_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2613_ _1176_ _1181_ _1182_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2475_ S2END[0] W6END[1] S4END[3] AD2 Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q Inst_RegFile_switch_matrix.S4BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3593_ WW4END[4] net238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2544_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q _0272_ _1113_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1357_ S2MID[7] _1248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1426_ Inst_RegFile_32x4.mem\[15\]\[2\] _1317_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3027_ FrameData[19] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkload4 clknet_4_4_0_UserCLK_regs clkload4/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_57_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2191_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ _0817_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _0134_ _0877_ _0878_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_23_Left_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1975_ _0556_ _0593_ _0603_ _0615_ _0616_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2527_ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q AD2 _1096_ _1097_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3576_ W2MID[3] net221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2458_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q Inst_RegFile_switch_matrix.JS2BEG0
+ _1048_ Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q _1049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1409_ Inst_RegFile_32x4.mem\[2\]\[1\] _1300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2389_ AD0 AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ _0991_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1760_ _0253_ _0404_ _0410_ _0411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ Inst_RegFile_32x4.mem\[3\]\[1\] A_ADR0 _0344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3430_ FrameData[26] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2312_ _0916_ _0924_ _0136_ _0925_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3292_ FrameData[28] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3361_ Inst_RegFile_switch_matrix.E2BEG1 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2174_ W6END[1] AD0 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2243_ _0861_ _0862_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q _0863_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput39 net39 EE4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput28 net28 E6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput17 net17 E2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1889_ _0530_ _0531_ _1273_ _0532_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1958_ Inst_RegFile_32x4.mem\[7\]\[0\] B_ADR0 _0599_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_9_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_9_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3559_ Inst_RegFile_switch_matrix.SS4BEG3 net195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ FrameData[18] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2861_ _0055_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[15\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3413_ FrameData[9] net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1743_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] A_ADR0 _0394_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1674_ Inst_RegFile_32x4.mem\[14\]\[0\] _0147_ _0329_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1812_ Inst_RegFile_32x4.mem\[6\]\[3\] _0147_ _0461_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2792_ _1182_ Inst_RegFile_32x4.mem\[10\]\[0\] _1244_ _0116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2226_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ _0848_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3275_ FrameData[11] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3344_ _0116_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[10\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2157_ _1248_ Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ _0786_ _0787_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_36_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2088_ Inst_RegFile_32x4.mem\[12\]\[2\] B_ADR0 _0722_ _0723_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_10_Left_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1390_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _1281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3060_ FrameData[20] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2011_ Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] B_ADR0 _0650_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2844_ _0038_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[17\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2913_ FrameData[1] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1588_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0245_ _0246_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2775_ _1198_ Inst_RegFile_32x4.mem\[6\]\[3\] _1240_ _0103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1657_ Inst_RegFile_32x4.mem\[3\]\[0\] A_ADR0 _0312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1726_ _1315_ _0147_ _0376_ _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3189_ FrameData[21] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3258_ FrameData[26] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3327_ _0099_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[5\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2209_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ _0833_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_47_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1511_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q S4END[2] _0172_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1442_ Inst_RegFile_32x4.mem\[17\]\[3\] _1333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2560_ NN4END[1] Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q _1128_ _1129_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2491_ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q _1053_ _1073_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput218 net218 W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput229 net229 W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput207 net207 W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3112_ FrameData[8] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3043_ FrameData[3] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_4_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1373_ Inst_RegFile_32x4.mem\[2\]\[0\] _1264_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_546 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2827_ _0021_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[2\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2758_ _1186_ Inst_RegFile_32x4.mem\[3\]\[2\] _1236_ _0090_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2689_ _1201_ _1221_ _1222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1709_ _1310_ _0147_ _0361_ _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_44_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkload11 clknet_4_13_0_UserCLK_regs clkload11/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_2612_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _1177_ _1180_ _1181_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1991_ Inst_RegFile_32x4.mem\[27\]\[1\] B_ADR0 _0630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3592_ Inst_RegFile_switch_matrix.W6BEG1 net228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2474_ S2END[1] W6END[0] S4END[0] AD3 Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q Inst_RegFile_switch_matrix.S4BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1425_ Inst_RegFile_32x4.mem\[13\]\[2\] _1316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2543_ _1109_ _1111_ _1112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3026_ FrameData[18] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1356_ E2MID[6] _1247_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkload5 clknet_4_7_0_UserCLK_regs clkload5/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_11_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_557 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2190_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0815_ _0816_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _0549_ _0614_ _0581_ _0615_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_538 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3575_ W2MID[2] net220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2388_ NN4END[0] SS4END[0] E1END[3] W1END[3] Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q _0990_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2526_ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q _1058_ Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q
+ _1096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1408_ Inst_RegFile_32x4.mem\[31\]\[0\] _1299_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2457_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q _0195_ _1048_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3009_ FrameData[1] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ _0219_ _0337_ _0342_ _0254_ _0343_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3291_ FrameData[27] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2311_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0920_ _0923_ _0924_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_29_Left_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3360_ Inst_RegFile_switch_matrix.E2BEG0 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2242_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ _0862_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2173_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ _0801_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_18_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0486_ _0595_ _0597_ _0518_ _0598_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput29 net29 E6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput18 net18 E2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2509_ _1084_ _1086_ Inst_RegFile_switch_matrix.E1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3558_ Inst_RegFile_switch_matrix.SS4BEG2 net194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1888_ N2END[1] S2END[1] EE4END[3] W2END[1] Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q _0531_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3489_ Inst_RegFile_switch_matrix.N4BEG1 net125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2860_ _0054_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[15\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1811_ _0180_ _0457_ _0458_ _0459_ _0218_ _0460_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2791_ _1203_ _1216_ _1244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3412_ FrameData[8] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1673_ _1285_ _0147_ _0327_ _0328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1742_ _0180_ _0392_ _0218_ _0393_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2225_ W6END[0] AD0 AD2 AD3 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ _0847_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3274_ FrameData[10] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3343_ _0115_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[0\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2156_ W2MID[7] Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q _0786_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ _1316_ B_ADR0 _0722_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2989_ FrameData[13] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_42_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ Inst_RegFile_32x4.mem\[10\]\[1\] Inst_RegFile_32x4.mem\[11\]\[1\] B_ADR0 _0649_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_544 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2912_ FrameData[0] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_41_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2843_ _0037_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[17\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2774_ _1186_ Inst_RegFile_32x4.mem\[6\]\[2\] _1240_ _0102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1725_ Inst_RegFile_32x4.mem\[10\]\[2\] _0147_ _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1587_ S1END[0] S2END[6] S1END[2] W1END[2] Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q _0245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1656_ _0253_ _0305_ _0310_ _0300_ _0311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3326_ _0098_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[5\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3188_ FrameData[20] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3257_ FrameData[25] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2139_ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q _0768_ _0770_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ _0771_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2208_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0831_ _0832_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1510_ _0164_ _0166_ _0168_ _0170_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q _0171_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_4_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput219 net219 W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1441_ Inst_RegFile_32x4.mem\[15\]\[3\] _1332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput208 net208 W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2490_ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q BD0 _1071_ _1072_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1372_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q _1263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3111_ FrameData[7] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3042_ FrameData[2] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1708_ Inst_RegFile_32x4.mem\[30\]\[1\] _0147_ _0361_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2688_ _1134_ _1220_ _1221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2757_ _1184_ Inst_RegFile_32x4.mem\[3\]\[1\] _1236_ _0089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2826_ _0020_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[2\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1639_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _0293_ _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3309_ _0081_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[29\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ Inst_RegFile_32x4.mem\[25\]\[1\] B_ADR0 _0486_ _0628_ _0629_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_15_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkload12 clknet_4_14_0_UserCLK_regs clkload12/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2611_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _1179_ Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ _1180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3591_ Inst_RegFile_switch_matrix.W6BEG0 net227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2542_ Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q _1110_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q
+ _1111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2473_ _1060_ _1062_ Inst_RegFile_switch_matrix.W1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1424_ Inst_RegFile_32x4.mem\[11\]\[2\] _1315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3025_ FrameData[17] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkload6 clknet_4_8_0_UserCLK_regs clkload6/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_2809_ _0003_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[24\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _0608_ _0613_ _0517_ _0614_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2525_ _1091_ _1093_ _1095_ Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q Inst_RegFile_switch_matrix.N1BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3574_ W2MID[1] net219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2387_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q _0980_ _0982_ _0987_ _0989_ Inst_RegFile_switch_matrix.E6BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1407_ Inst_RegFile_32x4.mem\[29\]\[0\] _1298_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2456_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q BD2 _1046_ _1047_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ FrameData[0] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3290_ FrameData[26] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2172_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q _0798_ _0800_ _0794_ _0796_ Inst_RegFile_switch_matrix.JW2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2310_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0922_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ _0923_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2241_ W6END[1] AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ _0861_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1887_ NN4END[0] E6END[0] W2END[0] Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q _0530_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1956_ _1264_ B_ADR0 _0486_ _0596_ _0597_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3488_ Inst_RegFile_switch_matrix.N4BEG0 net124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput19 net19 E2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2508_ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q Inst_RegFile_switch_matrix.JN2BEG3
+ _1085_ Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q _1086_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3557_ Inst_RegFile_switch_matrix.SS4BEG1 net193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2439_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q BD1 _1033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1810_ Inst_RegFile_32x4.mem\[3\]\[3\] A_ADR0 _0162_ _0179_ _0459_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2790_ _1198_ Inst_RegFile_32x4.mem\[0\]\[3\] _1243_ _0115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1741_ Inst_RegFile_32x4.mem\[0\]\[2\] A_ADR0 _0391_ _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3411_ FrameData[7] net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1672_ Inst_RegFile_32x4.mem\[12\]\[0\] _0147_ _0327_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3342_ _0114_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[0\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3273_ FrameData[9] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2155_ N2MID[6] E2MID[6] W2MID[6] Inst_RegFile_switch_matrix.JN2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q _0785_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2224_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q _0844_ _0846_ _0840_ _0842_ Inst_RegFile_switch_matrix.E2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_36_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2086_ Inst_RegFile_32x4.mem\[14\]\[2\] B_ADR0 _0720_ _0721_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2988_ FrameData[12] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1939_ _0576_ _0579_ _0569_ _0580_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_48_Left_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Left_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_5_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_5_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Left_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2911_ FrameData[31] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2842_ _0036_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[17\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_41_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1724_ Inst_RegFile_32x4.AD_comb\[1\] Inst_RegFile_32x4.AD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2773_ _1184_ Inst_RegFile_32x4.mem\[6\]\[1\] _1240_ _0101_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1586_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q _0244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3256_ FrameData[24] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1655_ _0180_ _0307_ _0309_ _0219_ _0310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3325_ _0097_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[5\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2069_ Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q _0703_ _0704_ BD3 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3187_ FrameData[19] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2138_ _1247_ Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q
+ _0769_ _0770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2207_ W6END[0] AD0 AD2 AD3 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ _0831_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_47_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1371_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _1262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3110_ FrameData[6] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput209 net209 W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1440_ Inst_RegFile_32x4.mem\[13\]\[3\] _1331_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3041_ FrameData[1] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2825_ _0019_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[28\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1707_ _1309_ A_ADR0 _0359_ _0360_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1638_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q _0293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2687_ _1107_ _1120_ _1220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2756_ _1182_ Inst_RegFile_32x4.mem\[3\]\[0\] _1236_ _0088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3308_ _0080_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[29\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1569_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _0227_ _0228_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3239_ FrameData[7] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkload13 clknet_4_15_0_UserCLK_regs clkload13/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2610_ _1178_ _1179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2472_ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q Inst_RegFile_switch_matrix.JS2BEG3
+ _1061_ Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q _1062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3590_ W6END[11] net237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2541_ N4END[0] SS4END[0] Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q _1110_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1423_ Inst_RegFile_32x4.mem\[9\]\[2\] _1314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ FrameData[16] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkload7 clknet_4_9_0_UserCLK_regs clkload7/Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2808_ _0002_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[24\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2739_ Inst_RegFile_32x4.mem\[21\]\[3\] _1198_ _1232_ _0075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_6_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ _0612_ _0610_ _0486_ _0613_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3573_ W2MID[0] net218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2455_ Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q _0789_ Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q
+ _1046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2524_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q AD3 _1094_ _1095_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2386_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0988_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ _0989_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1406_ Inst_RegFile_32x4.mem\[27\]\[0\] _1297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3007_ FrameData[31] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2171_ _1354_ _0799_ _0800_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2240_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q _0858_ _0860_ _0854_ _0856_ Inst_RegFile_switch_matrix.JW2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XPHY_EDGE_ROW_27_Left_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q _0527_ _0529_ _0523_ _0525_ Inst_RegFile_switch_matrix.JW2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_31_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1955_ Inst_RegFile_32x4.mem\[3\]\[0\] B_ADR0 _0596_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2438_ _0930_ _0484_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q _1032_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2507_ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q _1053_ _1085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3487_ N4END[15] net123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3556_ Inst_RegFile_switch_matrix.SS4BEG0 net192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q _0922_ _0973_ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ _0974_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_4_13_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_13_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_22_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1671_ _0180_ _0325_ _0218_ _0326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1740_ _1311_ A_ADR0 _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3410_ FrameData[6] net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3272_ FrameData[8] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3341_ _0113_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[0\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2154_ _0783_ _0784_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ _1317_ B_ADR0 _0720_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2223_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q _0845_ _0846_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ FrameData[11] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1869_ _0510_ _0512_ _0513_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1938_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q _0578_ _0579_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3608_ Inst_RegFile_switch_matrix.WW4BEG3 net244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3539_ S4END[15] net175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_70_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_546 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2910_ FrameData[30] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2841_ _0035_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[13\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1654_ Inst_RegFile_32x4.mem\[23\]\[0\] A_ADR0 _0162_ _0179_ _0308_ _0309_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_41_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1723_ _0300_ _0343_ _0353_ _0364_ _0375_ Inst_RegFile_32x4.AD_comb\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2772_ _1182_ Inst_RegFile_32x4.mem\[6\]\[0\] _1240_ _0100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3255_ FrameData[23] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1585_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0242_ _1349_ _0243_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3324_ _0096_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[5\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2206_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q _0828_ _0830_ _0824_ _0826_ Inst_RegFile_switch_matrix.JW2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2068_ Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q Inst_RegFile_32x4.BD_reg\[3\] _0704_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3186_ FrameData[18] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2137_ N2MID[6] Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q _0769_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_502 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1370_ SS4END[2] _1261_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3040_ FrameData[0] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2824_ _0018_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[28\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1637_ _0287_ _0289_ _0291_ _0292_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1706_ Inst_RegFile_32x4.mem\[29\]\[1\] A_ADR0 _0359_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2686_ _1198_ Inst_RegFile_32x4.mem\[13\]\[3\] _1219_ _0035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2755_ _1206_ _1212_ _1236_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1499_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _0160_ Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ _0161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3307_ _0079_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[19\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1568_ N1END[2] N2END[4] NN4END[3] E2END[4] Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q _0227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3169_ FrameData[1] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3238_ FrameData[6] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2471_ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q _1053_ _1061_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1422_ Inst_RegFile_32x4.mem\[6\]\[2\] _1313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_switch_matrix.JW2BEG2
+ _1108_ _1109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3023_ FrameData[15] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkload8 clknet_4_10_0_UserCLK_regs clkload8/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2738_ Inst_RegFile_32x4.mem\[21\]\[2\] _1186_ _1232_ _0074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2807_ _0001_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[24\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2669_ _1204_ _1209_ _1214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_390 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ Inst_RegFile_32x4.mem\[12\]\[0\] B_ADR0 _0611_ _0612_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3572_ Inst_RegFile_switch_matrix.JW2BEG7 net217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2385_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ _0988_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1405_ Inst_RegFile_32x4.mem\[25\]\[0\] _1296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2454_ BD3 _0468_ Inst_RegFile_switch_matrix.JS2BEG1 _0530_ Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q Inst_RegFile_switch_matrix.W1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2523_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q _0789_ _1094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3006_ FrameData[30] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_62_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Left_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ E6END[1] S2END[3] S4END[3] W2END[3] Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0799_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1954_ _1253_ B_ADR0 _0594_ _0595_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3555_ SS4END[15] net191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1885_ _1281_ _0528_ _0529_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2437_ _1031_ _1030_ Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q Inst_RegFile_switch_matrix.NN4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2506_ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q AD3 _1083_ _1084_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3486_ N4END[14] net122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2368_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q _0238_ _0973_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2299_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q _0911_ _0912_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput190 net190 SS4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1670_ Inst_RegFile_32x4.mem\[8\]\[0\] A_ADR0 _0324_ _0325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3271_ FrameData[7] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2222_ N1END[0] N2END[2] N4END[2] NN4END[1] Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q _0845_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3340_ _0112_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[0\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2153_ N2END[7] S2END[7] EE4END[2] W2END[7] Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2084_ _0716_ _0718_ _0486_ _0719_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2986_ FrameData[10] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1937_ N2END[2] _1287_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _0577_ _0578_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3538_ S4END[14] net174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1868_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q _0511_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ _0512_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3607_ Inst_RegFile_switch_matrix.WW4BEG2 net243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1799_ _1329_ _0147_ _0180_ _0447_ _0448_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3469_ N2MID[1] net114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_70_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_503 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2840_ _0034_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[13\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2771_ _1203_ _1237_ _1240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1584_ AD3 BD0 BD2 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ _0242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1653_ _1295_ A_ADR0 _0308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1722_ _0253_ _0369_ _0374_ _0300_ _0375_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_7_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3254_ FrameData[22] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3185_ FrameData[17] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3323_ _0095_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[4\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2205_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0829_ _0830_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2067_ _0703_ Inst_RegFile_32x4.BD_comb\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2136_ S2MID[6] Inst_RegFile_switch_matrix.JN2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q
+ _0768_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2969_ FrameData[25] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_1_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_46_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2823_ _0017_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[28\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1705_ _0180_ _0357_ _0218_ _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2754_ Inst_RegFile_32x4.mem\[31\]\[3\] _1198_ _1235_ _0087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1636_ _1254_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q
+ _0290_ _0291_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3306_ _0078_ clknet_4_10_0_UserCLK_regs Inst_RegFile_32x4.mem\[19\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1567_ _1351_ _0225_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q _0226_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2685_ _1186_ Inst_RegFile_32x4.mem\[13\]\[2\] _1219_ _0034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2119_ W1END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ _0752_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1498_ Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q _0157_ _0159_ _0160_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3168_ FrameData[0] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3237_ FrameData[5] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_52_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3099_ FrameData[27] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ Inst_RegFile_32x4.mem\[2\]\[2\] _1312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2470_ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q BD1 _1059_ _1060_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3022_ FrameData[14] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkload9 clknet_4_11_0_UserCLK_regs clkload9/ZN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_2737_ Inst_RegFile_32x4.mem\[21\]\[1\] _1184_ _1232_ _0073_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2806_ _0000_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[24\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2668_ _1198_ Inst_RegFile_32x4.mem\[2\]\[3\] _1213_ _0023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1619_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q Inst_RegFile_switch_matrix.JW2BEG5
+ _0275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2599_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q _1167_ _1168_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _1285_ B_ADR0 _0611_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3571_ Inst_RegFile_switch_matrix.JW2BEG6 net216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2522_ Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q _1092_ _1093_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1404_ Inst_RegFile_32x4.mem\[22\]\[0\] _1295_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2384_ _0984_ _0986_ _0137_ _0987_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2453_ Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q _1045_ _1043_ Inst_RegFile_switch_matrix.W1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3005_ FrameData[29] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_36_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1884_ S1END[1] S2END[5] S1END[3] W1END[1] Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q _0528_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1953_ Inst_RegFile_32x4.mem\[0\]\[0\] B_ADR0 _0594_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ SS4END[14] net190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2505_ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q _1058_ Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q
+ _1083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3485_ N4END[13] net136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2436_ N1END[3] E1END[3] W1END[3] AD2 Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q _1031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2298_ NN4END[2] E1END[2] SS4END[2] W1END[2] Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q _0911_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2367_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q BD2 _0971_ _0972_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput180 net180 S4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput191 net191 SS4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2152_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _0781_ _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3270_ FrameData[6] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2221_ _0132_ _0843_ _0844_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2083_ Inst_RegFile_32x4.mem\[10\]\[2\] B_ADR0 _0717_ _0718_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1867_ E6END[1] S4END[1] Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q _0511_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2985_ FrameData[9] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1936_ S2END[2] Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _0577_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3537_ S4END[13] net188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3468_ N2MID[0] net113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3606_ Inst_RegFile_switch_matrix.WW4BEG1 net242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1798_ Inst_RegFile_32x4.mem\[8\]\[3\] _0147_ _0447_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3399_ EE4END[15] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2419_ NN4END[0] S2END[2] E2END[2] W2END[2] Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q _1016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_29_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_541 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1721_ _0180_ _0371_ _0373_ _0219_ _0374_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_41_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2770_ _1198_ Inst_RegFile_32x4.mem\[5\]\[3\] _1239_ _0099_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ _1348_ _0240_ _0241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1652_ Inst_RegFile_32x4.mem\[20\]\[0\] A_ADR0 _0306_ _0307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_44_Left_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3322_ _0094_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[4\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3253_ FrameData[21] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3184_ FrameData[16] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_53_Left_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2135_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q _0766_ _0765_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q
+ _0767_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2204_ N1END[0] E2END[2] N2END[2] E6END[0] Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q _0829_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2066_ _0668_ _0680_ _0690_ _0702_ _0703_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1919_ E2END[7] S1END[3] S2END[7] W1END[1] Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0561_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_62_Left_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2899_ FrameData[19] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2968_ FrameData[24] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ Inst_RegFile_32x4.mem\[25\]\[1\] A_ADR0 _0356_ _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2822_ _0016_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[28\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2753_ Inst_RegFile_32x4.mem\[31\]\[2\] _1186_ _1235_ _0086_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2684_ _1184_ Inst_RegFile_32x4.mem\[13\]\[1\] _1219_ _0033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1635_ N2MID[2] Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q _0290_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3305_ _0077_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[19\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1497_ _1259_ Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ _0158_ _0159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1566_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ _0225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3167_ FrameData[31] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2118_ Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q _0750_ _0751_ BD2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3098_ FrameData[26] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3236_ FrameData[4] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2049_ _1328_ B_ADR0 _0486_ _0685_ _0686_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_52_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_515 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ Inst_RegFile_32x4.mem\[1\]\[2\] _1311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3021_ FrameData[13] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_36_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ _1198_ Inst_RegFile_32x4.mem\[12\]\[3\] _1246_ _0127_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2736_ Inst_RegFile_32x4.mem\[21\]\[0\] _1182_ _1232_ _0072_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1618_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q Inst_RegFile_switch_matrix.JN2BEG5
+ _0273_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q _0274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2667_ _1186_ Inst_RegFile_32x4.mem\[2\]\[2\] _1213_ _0022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_470 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3219_ FrameData[19] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1549_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q _0206_ _0208_ _0202_ _0204_ Inst_RegFile_switch_matrix.JS2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2598_ _0141_ _1166_ _1167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q _0195_ _1092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3570_ Inst_RegFile_switch_matrix.JW2BEG5 net215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1403_ Inst_RegFile_32x4.mem\[21\]\[0\] _1294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2383_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0920_ _0985_ _0986_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2452_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q AD0 _1044_ _1045_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3004_ FrameData[28] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ Inst_RegFile_32x4.mem\[16\]\[3\] _1198_ _1228_ _0059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1883_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _0526_ _0527_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1952_ _0549_ _0592_ _0580_ _0593_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3553_ SS4END[13] net204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2435_ _1027_ _1029_ _1030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3484_ N4END[12] net135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2504_ _1080_ _1082_ Inst_RegFile_switch_matrix.E1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_554 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2297_ _0910_ _0907_ Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q Inst_RegFile_switch_matrix.JN2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2366_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q _0920_ _0971_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput170 net170 S2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput181 net181 S4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput192 net192 SS4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2151_ _0780_ _0781_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2220_ E2END[2] S2END[2] E6END[0] W2END[2] Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q _0843_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2082_ _1315_ B_ADR0 _0717_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2984_ FrameData[8] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q Inst_RegFile_switch_matrix.JS2BEG4
+ _0509_ _0510_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1935_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _0571_ _0574_ _0576_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3605_ Inst_RegFile_switch_matrix.WW4BEG0 net241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1797_ Inst_RegFile_32x4.mem\[10\]\[3\] A_ADR0 _0445_ _0446_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3536_ S4END[12] net187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3467_ Inst_RegFile_switch_matrix.JN2BEG7 net112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3398_ EE4END[14] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2418_ _1015_ _1014_ Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q Inst_RegFile_switch_matrix.EE4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2349_ N1END[3] S1END[3] W1END[3] AD2 Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ _0958_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_70_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_502 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1651_ _1294_ A_ADR0 _0306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1720_ Inst_RegFile_32x4.mem\[22\]\[1\] _0147_ _0162_ _0179_ _0372_ _0373_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3252_ FrameData[20] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1582_ WW4END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3321_ _0093_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[4\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3183_ FrameData[15] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2134_ N2END[7] E2END[7] S2END[7] WW4END[0] Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q _0766_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2203_ _0130_ _0827_ _0828_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2065_ _0549_ _0701_ _0581_ _0702_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ FrameData[23] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1849_ S1END[3] S2END[7] SS4END[1] W1END[1] Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q _0495_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1918_ N1END[3] N2END[7] NN4END[1] E1END[3] Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q _0560_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2898_ FrameData[18] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3519_ Inst_RegFile_switch_matrix.JS2BEG7 net164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_4_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2821_ _0015_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[27\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1634_ _1258_ _0288_ _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1703_ _1307_ A_ADR0 _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ Inst_RegFile_32x4.mem\[31\]\[1\] _1184_ _1235_ _0085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2683_ _1182_ Inst_RegFile_32x4.mem\[13\]\[0\] _1219_ _0032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3304_ _0076_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[19\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1496_ W2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q _0158_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1565_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q _0223_ _0224_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3235_ FrameData[3] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_18_Left_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3166_ FrameData[30] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2117_ Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q Inst_RegFile_32x4.BD_reg\[2\] _0751_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3097_ FrameData[25] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2048_ Inst_RegFile_32x4.mem\[7\]\[3\] B_ADR0 _0685_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ FrameData[12] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_48_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _1186_ Inst_RegFile_32x4.mem\[12\]\[2\] _1246_ _0126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1617_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _0272_ _0273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2735_ _1201_ _1223_ _1232_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2597_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q _1166_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2666_ _1184_ Inst_RegFile_32x4.mem\[2\]\[1\] _1213_ _0021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3218_ FrameData[18] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_57_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1548_ _1346_ _0207_ _0208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3149_ FrameData[13] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1479_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q _0142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_65_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_28_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1402_ Inst_RegFile_32x4.mem\[18\]\[0\] _1293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2451_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q _0573_ _1044_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2520_ Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q Inst_RegFile_switch_matrix.JW2BEG0
+ _1091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0922_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ _0985_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3003_ FrameData[27] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_62_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ Inst_RegFile_32x4.mem\[16\]\[2\] _1186_ _1228_ _0058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2649_ _1142_ _1199_ _1206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3552_ SS4END[12] net203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1882_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q _0526_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1951_ _0586_ _0591_ _0517_ _0592_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_544 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q _0922_ _1028_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ _1029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3483_ N4END[11] net134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2365_ _0970_ Inst_RegFile_switch_matrix.SS4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2503_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q Inst_RegFile_switch_matrix.JN2BEG0
+ _1081_ Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q _1082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_39_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2296_ _0909_ _0908_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0910_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_20 W6END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput182 net182 S4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput171 net171 S2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput160 net160 S2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput193 net193 SS4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ N4END[3] E2END[3] W2END[3] Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ Inst_RegFile_32x4.mem\[8\]\[2\] B_ADR0 _0715_ _0716_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ FrameData[7] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1934_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _0571_ _0574_ _0575_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3535_ S4END[11] net186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1865_ Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q _1268_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q
+ _0509_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3604_ WW4END[15] net240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1796_ _1330_ A_ADR0 _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3397_ EE4END[13] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3466_ Inst_RegFile_switch_matrix.JN2BEG6 net111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2417_ N1END[2] E1END[2] S1END[2] AD1 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q _1015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2348_ Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q _0954_ _0956_ _0957_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ N1END[3] N2END[1] N4END[1] NN4END[0] Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q _0895_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_543 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ _0180_ _0304_ _0302_ _0218_ _0305_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1581_ _0232_ _0234_ _0238_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q
+ _0239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3182_ FrameData[14] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3251_ FrameData[19] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3320_ _0092_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[4\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2202_ S2END[2] S4END[2] SS4END[1] W2END[2] Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q _0827_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_49_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2133_ Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q _0764_ _0762_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ _0765_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ _0695_ _0700_ _0517_ _0701_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1917_ _0557_ _0558_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q _0559_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2897_ FrameData[17] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2966_ FrameData[22] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1848_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0493_ _0494_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1779_ Inst_RegFile_32x4.mem\[28\]\[3\] _0147_ _0428_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3518_ Inst_RegFile_switch_matrix.JS2BEG6 net163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3449_ FrameStrobe[13] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_4_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2820_ _0014_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[27\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ Inst_RegFile_32x4.mem\[31\]\[0\] _1182_ _1235_ _0084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_9_Left_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1633_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q W2MID[2] _0288_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1564_ W6END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ _0223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1702_ _1308_ A_ADR0 _0181_ _0354_ _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2682_ _1200_ _1218_ _1219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3165_ FrameData[29] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1495_ N2MID[3] E2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q _0157_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3303_ Inst_RegFile_32x4.AD_comb\[3\] clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.AD_reg\[3\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3234_ FrameData[2] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2116_ _0750_ Inst_RegFile_32x4.BD_comb\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3096_ FrameData[24] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_1_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2047_ _0486_ _0681_ _0683_ _0518_ _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_13_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ FrameData[5] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_476 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ Inst_RegFile_32x4.mem\[20\]\[3\] _1198_ _1231_ _0071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2803_ _1184_ Inst_RegFile_32x4.mem\[12\]\[1\] _1246_ _0125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1547_ S1END[2] S2END[6] SS4END[2] W1END[0] Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q _0207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2596_ _1158_ _1159_ _1163_ _1165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1616_ Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q _0271_ _0270_ _0272_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2665_ _1182_ Inst_RegFile_32x4.mem\[2\]\[0\] _1213_ _0020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3217_ FrameData[17] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3148_ FrameData[12] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_57_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1478_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q _0141_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ FrameData[7] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1401_ Inst_RegFile_32x4.mem\[17\]\[0\] _1292_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2381_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0212_ _0983_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ _0984_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2450_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q Inst_RegFile_switch_matrix.JS2BEG2
+ _1042_ Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q _1043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_5_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3002_ FrameData[26] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_36_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_523 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ Inst_RegFile_32x4.mem\[16\]\[1\] _1184_ _1228_ _0057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2648_ Inst_RegFile_32x4.mem\[26\]\[3\] _1198_ _1205_ _0011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2579_ N2END[3] S2END[3] _1136_ _1123_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q
+ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q _1148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1950_ _0590_ _0588_ _0486_ _0591_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3551_ SS4END[11] net202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1881_ _1281_ _0524_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q _0525_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2502_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q _0195_ _1081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2433_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q _0178_ _1028_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2364_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q _0969_ _0968_ _0970_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_22_Left_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3482_ N4END[10] net133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2295_ N2END[1] N4END[1] E1END[3] E2END[1] Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q _0909_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_10 W6END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_21 WW4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput150 net150 NN4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput161 net161 S2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput172 net172 S2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput183 net183 S4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput194 net194 SS4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ _1314_ B_ADR0 _0715_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2982_ FrameData[6] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1933_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _0572_ _0574_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3534_ S4END[10] net185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1864_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q _0506_ _0508_ _0502_ _0504_ Inst_RegFile_switch_matrix.JS2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3465_ Inst_RegFile_switch_matrix.JN2BEG5 net110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1795_ _0253_ _0438_ _0443_ _0300_ _0444_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3603_ WW4END[14] net239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3396_ EE4END[12] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2416_ BD1 _0930_ _0936_ _0766_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q
+ _1014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2278_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0893_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q
+ _0894_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2347_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q _0922_ _0955_ Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ _0956_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_70_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q _0235_ _0237_ _0238_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3181_ FrameData[13] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3250_ FrameData[18] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2132_ N4END[3] Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q _0763_ _0764_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2201_ _0130_ _0825_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q _0826_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2063_ _0699_ _0697_ _0486_ _0700_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1916_ AD3 BD0 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ _0558_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1847_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q _0493_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2896_ FrameData[16] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2965_ FrameData[21] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3448_ FrameStrobe[12] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_31_Left_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1778_ _0180_ _0426_ _0218_ _0427_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3517_ Inst_RegFile_switch_matrix.JS2BEG5 net162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3379_ E6END[5] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_40_Left_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1701_ Inst_RegFile_32x4.mem\[27\]\[1\] A_ADR0 _0354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2750_ _1207_ _1209_ _1235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2681_ _1134_ _1215_ _1218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1632_ _0280_ _0282_ _0284_ _0286_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q _0287_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1494_ N2MID[2] S2MID[2] E2MID[2] Inst_RegFile_switch_matrix.E2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q _0156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1563_ _0180_ _0221_ _0218_ _0222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3302_ Inst_RegFile_32x4.AD_comb\[2\] clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.AD_reg\[2\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3164_ FrameData[28] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2115_ _0714_ _0726_ _0737_ _0749_ _0750_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3095_ FrameData[23] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3233_ FrameData[1] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2046_ _1326_ B_ADR0 _0486_ _0682_ _0683_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_17_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2879_ _0073_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[21\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ FrameData[4] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_9_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2733_ Inst_RegFile_32x4.mem\[20\]\[2\] _1186_ _1231_ _0070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2802_ _1182_ Inst_RegFile_32x4.mem\[12\]\[0\] _1246_ _0124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_14_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2664_ _1203_ _1212_ _1213_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1546_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _0205_ _0206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2595_ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _1160_ _1162_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q
+ _1164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1477_ Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q _0140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1615_ S2END[0] W2END[0] Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q _0271_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3216_ FrameData[16] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_57_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3147_ FrameData[11] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3078_ FrameData[6] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2029_ _1335_ B_ADR0 _0665_ _0666_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1400_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q _1291_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2380_ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0497_ _0983_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ FrameData[25] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2716_ Inst_RegFile_32x4.mem\[16\]\[0\] _1182_ _1228_ _0056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2647_ Inst_RegFile_32x4.mem\[26\]\[2\] _1186_ _1205_ _0010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1529_ N2END[4] E2END[4] E1END[2] EE4END[3] Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q _0190_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2578_ _1143_ _1144_ _1145_ _1146_ _1147_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1880_ AD3 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ _0524_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3550_ SS4END[10] net201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3481_ N4END[9] net132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2501_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q BD0 _1079_ _1080_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2432_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q BD2 _1026_ _1027_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2363_ N1END[0] E1END[0] W1END[0] AD3 Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q _0969_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ EE4END[0] E6END[1] S2END[1] W2END[1] Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q _0908_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_22 WW4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_11 W6END[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput140 net140 NN4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput151 net151 NN4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput184 net184 S4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput162 net162 S2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput173 net173 S4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput195 net195 SS4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1863_ _1270_ _0507_ _0508_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1932_ _0572_ _0573_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3602_ WW4END[13] net253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2981_ FrameData[5] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3533_ S4END[9] net184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ Inst_RegFile_switch_matrix.JN2BEG4 net109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1794_ _0180_ _0440_ _0442_ _0219_ _0443_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2415_ _1013_ _1012_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q Inst_RegFile_switch_matrix.EE4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3395_ EE4END[11] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2277_ W6END[1] AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ _0893_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2346_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q _0198_ _0955_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3180_ FrameData[12] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_49_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2131_ _1251_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q _0763_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2062_ Inst_RegFile_32x4.mem\[12\]\[3\] B_ADR0 _0698_ _0699_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2200_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ _0825_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2964_ FrameData[20] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1846_ _1266_ _0491_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q _0492_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1915_ W1END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ _0557_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2895_ FrameData[15] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1777_ Inst_RegFile_32x4.mem\[24\]\[3\] A_ADR0 _0425_ _0426_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3378_ E6END[4] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3447_ FrameStrobe[11] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3516_ Inst_RegFile_switch_matrix.JS2BEG4 net161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2329_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0940_ _0938_ _0941_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _0280_ _0282_ _0284_ _0286_ Inst_RegFile_switch_matrix.E2BEG6 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _1198_ Inst_RegFile_32x4.mem\[9\]\[3\] _1217_ _0031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1700_ _0219_ _0347_ _0352_ _0253_ _0353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1493_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q _0153_ _0155_ _0149_ _0151_ Inst_RegFile_switch_matrix.E2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1562_ Inst_RegFile_32x4.mem\[24\]\[0\] A_ADR0 _0220_ _0221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3301_ Inst_RegFile_32x4.AD_comb\[1\] clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.AD_reg\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3232_ FrameData[0] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3163_ FrameData[27] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2114_ _0549_ _0748_ _0580_ _0749_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3094_ FrameData[22] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2045_ Inst_RegFile_32x4.mem\[3\]\[3\] B_ADR0 _0682_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2947_ FrameData[3] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1829_ EE4END[3] S1END[1] S1END[3] S2END[5] Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q _0476_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2878_ _0072_ clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.mem\[21\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_8_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_8_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_68_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _1172_ _1218_ _1246_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ Inst_RegFile_32x4.mem\[20\]\[1\] _1184_ _1231_ _0069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2594_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q _1162_ _1163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1614_ _1255_ Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q
+ _0269_ _0270_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2663_ _1133_ _1211_ _1212_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1545_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q _0205_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_57_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1476_ Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q _0139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3215_ FrameData[15] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_65_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ Inst_RegFile_32x4.mem\[20\]\[3\] B_ADR0 _0665_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3146_ FrameData[10] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3077_ FrameData[5] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_24_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3000_ FrameData[24] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2646_ Inst_RegFile_32x4.mem\[26\]\[1\] _1184_ _1205_ _0009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2715_ _1173_ _1221_ _1228_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2577_ _0145_ _0531_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q _1146_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1528_ _1347_ _0188_ _0189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1459_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _1350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3129_ FrameData[25] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_529 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2431_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q _0920_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ _1026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3480_ N4END[8] net131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2500_ Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q _0789_ Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q
+ _1079_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2362_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q _0967_ _0965_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q
+ _0968_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2293_ _0905_ _0906_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q _0907_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_23 E6END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_12 W6END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput141 net141 NN4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput152 net152 NN4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput130 net130 N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2629_ Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q _1192_ _1194_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ _1195_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput185 net185 S4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput163 net163 S2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput196 net196 SS4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput174 net174 S4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ FrameData[4] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1862_ S1END[1] S2END[5] SS4END[3] W1END[1] Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q _0507_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1793_ Inst_RegFile_32x4.mem\[23\]\[3\] A_ADR0 _0162_ _0179_ _0441_ _0442_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3601_ WW4END[12] net252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1931_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q _0572_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3532_ S4END[8] net183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3394_ EE4END[10] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3463_ Inst_RegFile_switch_matrix.JN2BEG3 net108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2414_ N1END[3] E1END[3] S1END[3] AD2 Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q _1013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2276_ _0135_ _0891_ _0892_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2345_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q BD2 _0953_ _0954_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_491 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2130_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q S4END[3] Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ _0761_ _0762_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2061_ _1331_ B_ADR0 _0698_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1914_ _0521_ _0550_ _0555_ _0556_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2963_ FrameData[19] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1845_ AD3 BD0 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ _0491_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2894_ FrameData[14] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1776_ _1337_ A_ADR0 _0425_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3515_ Inst_RegFile_switch_matrix.JS2BEG3 net160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3377_ E6END[3] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3446_ FrameStrobe[10] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2328_ Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q _0468_ _0939_ _0940_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2259_ S2END[1] W2END[1] S4END[1] WW4END[0] Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q _0877_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1630_ _1256_ _0285_ _1257_ _0286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3231_ FrameData[31] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1492_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q _0154_ _0155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3162_ FrameData[26] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1561_ _1296_ A_ADR0 _0220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3300_ Inst_RegFile_32x4.AD_comb\[0\] clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.AD_reg\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2113_ _0742_ _0747_ _0517_ _0748_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3093_ FrameData[21] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2044_ Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] B_ADR0 _0681_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2877_ _0071_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[20\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2946_ FrameData[2] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _0474_ _0475_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1759_ _0180_ _0409_ _0407_ _0218_ _0410_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_9_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3429_ FrameData[25] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2731_ Inst_RegFile_32x4.mem\[20\]\[0\] _1182_ _1231_ _0068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2800_ _1198_ Inst_RegFile_32x4.mem\[11\]\[3\] _1245_ _0123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1544_ _1346_ _0203_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q _0204_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2593_ _1247_ _0140_ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _1161_ _1162_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1613_ N2END[0] Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q _0269_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _1107_ _1121_ _1211_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3145_ FrameData[9] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3214_ FrameData[14] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q _0138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_65_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2027_ _1336_ B_ADR0 _0486_ _0663_ _0664_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3076_ FrameData[4] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2929_ FrameData[17] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2714_ _1198_ Inst_RegFile_32x4.mem\[15\]\[3\] _1227_ _0055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1527_ E6END[0] S2END[4] S4END[0] W2END[4] Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q _0188_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2645_ Inst_RegFile_32x4.mem\[26\]\[0\] _1182_ _1205_ _0008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2576_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q Inst_RegFile_switch_matrix.JN2BEG0
+ _1145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1458_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q _1349_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3128_ FrameData[24] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1389_ E6END[0] _1280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3059_ FrameData[19] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2430_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q _1023_ _1025_ Inst_RegFile_switch_matrix.NN4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2361_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q BD3 _0966_ _0967_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2292_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ _0906_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_22_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_13 W6END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_24 E6END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput142 net142 NN4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput131 net131 N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput120 net120 N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2559_ _1255_ Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q _1128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput153 net153 S1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2628_ _1274_ Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q
+ _1193_ _1194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput164 net164 S2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput186 net186 S4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput175 net175 S4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput197 net197 SS4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _1287_ _0570_ _0571_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3531_ S4END[7] net182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1792_ _1336_ A_ADR0 _0441_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1861_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q _0505_ _0506_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_26_Left_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3600_ WW4END[11] net251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3462_ Inst_RegFile_switch_matrix.JN2BEG2 net107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3393_ EE4END[9] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2413_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q _1009_ _1011_ _1012_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2344_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q _0920_ _0953_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2275_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ _0891_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2060_ Inst_RegFile_32x4.mem\[14\]\[3\] B_ADR0 _0696_ _0697_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1913_ _0486_ _0554_ _0552_ _0517_ _0555_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2962_ FrameData[18] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2893_ FrameData[13] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1844_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0489_ _0490_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3445_ FrameStrobe[9] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1775_ _1338_ _0147_ _0181_ _0423_ _0424_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3514_ Inst_RegFile_switch_matrix.JS2BEG2 net159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3376_ E6END[2] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2327_ Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q _0160_ _0939_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2258_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0875_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q
+ _0876_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2189_ W6END[1] AD0 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ _0815_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1560_ _0200_ _0217_ _0219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3230_ FrameData[30] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1491_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q _0154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3161_ FrameData[25] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2112_ _0746_ _0744_ _0486_ _0747_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3092_ FrameData[20] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2043_ _0549_ _0679_ _0580_ _0680_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1827_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q _0474_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2876_ _0070_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[20\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2945_ FrameData[1] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3428_ FrameData[24] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1758_ _1325_ _0147_ _0408_ _0409_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1689_ _0338_ _0339_ _0341_ _0180_ _0219_ _0342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_68_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3359_ Inst_RegFile_switch_matrix.E1BEG3 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_13_Left_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _1173_ _1223_ _1231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2661_ Inst_RegFile_32x4.mem\[28\]\[3\] _1198_ _1210_ _0019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_14_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1612_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q _0266_ _0268_ _0262_ _0264_ Inst_RegFile_switch_matrix.JN2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1543_ AD3 BD0 BD2 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ _0203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1474_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2592_ S2MID[6] _0140_ _1161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3144_ FrameData[8] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3075_ FrameData[3] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3213_ FrameData[13] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_65_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ Inst_RegFile_32x4.mem\[23\]\[3\] B_ADR0 _0663_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2928_ FrameData[16] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2859_ _0053_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[15\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_4_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_4_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_14_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ _1135_ _1204_ _1205_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2713_ _1186_ Inst_RegFile_32x4.mem\[15\]\[2\] _1227_ _0054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1457_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _1348_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1526_ _1347_ _0186_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q _0187_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2575_ _0145_ Inst_RegFile_switch_matrix.JS2BEG0 _0146_ _1144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3058_ FrameData[18] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1388_ S2END[1] _1279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3127_ FrameData[23] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ _0550_ _0642_ _0647_ _0648_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_2_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Left_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _0160_ _0966_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_47_Left_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2291_ W6END[1] AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ _0905_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_56_Left_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_25 EE4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_14 W6END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput143 net143 NN4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput132 net132 N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_65_Left_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput121 net121 N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput110 net110 N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2627_ N2MID[0] Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q _1193_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1509_ _0164_ _0166_ _0168_ _0170_ Inst_RegFile_switch_matrix.E2BEG3 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2558_ S4END[1] Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q
+ _1127_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput187 net187 S4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput154 net154 S1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput165 net165 S2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput176 net176 S4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput198 net198 SS4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2489_ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q _1058_ Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ _1071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1860_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q _0505_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_1_Left_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3530_ S4END[6] net181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3461_ Inst_RegFile_switch_matrix.JN2BEG1 net106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1791_ Inst_RegFile_32x4.mem\[20\]\[3\] A_ADR0 _0439_ _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2274_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q _0890_ _0885_ Inst_RegFile_switch_matrix.E2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3392_ EE4END[8] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2412_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q _0922_ _1010_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ _1011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2343_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q _0950_ _0952_ Inst_RegFile_switch_matrix.WW4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1989_ _1307_ B_ADR0 _0628_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1843_ W1END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ _0489_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1912_ _1294_ B_ADR0 _0553_ _0554_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2892_ FrameData[12] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2961_ FrameData[17] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3444_ FrameStrobe[8] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3513_ Inst_RegFile_switch_matrix.JS2BEG1 net158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1774_ Inst_RegFile_32x4.mem\[26\]\[3\] _0147_ _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3375_ E2MID[7] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2326_ Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q _0930_ _0937_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ _0938_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2257_ W6END[1] AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ _0875_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2188_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q _0812_ _0814_ _0808_ _0810_ Inst_RegFile_switch_matrix.E2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_40_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1490_ _1343_ _0152_ _0153_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3160_ FrameData[24] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3091_ FrameData[19] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ Inst_RegFile_32x4.mem\[28\]\[2\] B_ADR0 _0745_ _0746_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2042_ _0673_ _0678_ _0517_ _0679_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1826_ _1262_ _0472_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q _0473_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2875_ _0069_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[20\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2944_ FrameData[0] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3427_ FrameData[23] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ Inst_RegFile_32x4.mem\[30\]\[2\] _0147_ _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1688_ Inst_RegFile_32x4.mem\[12\]\[1\] A_ADR0 _0340_ _0341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3358_ Inst_RegFile_switch_matrix.E1BEG2 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3289_ FrameData[25] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2309_ N2MID[4] S2MID[4] E2MID[4] Inst_RegFile_switch_matrix.JS2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q _0922_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_12_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_12_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_8_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _0267_ _0268_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2660_ Inst_RegFile_32x4.mem\[28\]\[2\] _1186_ _1210_ _0018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1542_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _0201_ _0202_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2591_ W2MID[6] Inst_RegFile_switch_matrix.JN2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q
+ _1160_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1473_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q _0136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3212_ FrameData[12] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2025_ _0486_ _0659_ _0661_ _0518_ _0662_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3143_ FrameData[7] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3074_ FrameData[2] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2927_ FrameData[15] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ _0052_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[15\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1809_ Inst_RegFile_32x4.mem\[2\]\[3\] _0147_ _0458_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2789_ _1186_ Inst_RegFile_32x4.mem\[0\]\[2\] _1243_ _0114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2643_ _1141_ _1149_ _1169_ _1204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2712_ _1184_ Inst_RegFile_32x4.mem\[15\]\[1\] _1227_ _0053_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2574_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q Inst_RegFile_switch_matrix.JW2BEG0
+ _1143_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1525_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ _0186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1456_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _1347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1387_ S2MID[1] _1278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3057_ FrameData[17] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3126_ FrameData[22] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2008_ _0486_ _0646_ _0644_ _0517_ _0647_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _0904_ _0901_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q Inst_RegFile_switch_matrix.JN2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_15 WW4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput100 net100 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput144 net144 NN4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput122 net122 N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput133 net133 N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput111 net111 N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2557_ _0143_ Inst_RegFile_switch_matrix.JS2BEG2 _1126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2626_ S2MID[0] Inst_RegFile_switch_matrix.JW2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q
+ _1192_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput155 net155 S1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput166 net166 S2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput177 net177 S4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1508_ _1289_ _0169_ _1291_ _0170_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput188 net188 S4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1439_ Inst_RegFile_32x4.mem\[11\]\[3\] _1330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput199 net199 SS4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2488_ Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q _1070_ _1068_ Inst_RegFile_switch_matrix.S1BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3109_ FrameData[5] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1790_ _1335_ A_ADR0 _0439_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3460_ Inst_RegFile_switch_matrix.JN2BEG0 net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3391_ EE4END[7] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2411_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q _0784_ _1010_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2273_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0889_ _0888_ _0890_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2342_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q _0951_ _0952_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1988_ _0621_ _0622_ _0626_ _0517_ _0549_ _0627_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2609_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q _1178_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3589_ W6END[10] net236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2960_ FrameData[16] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1911_ Inst_RegFile_32x4.mem\[20\]\[0\] B_ADR0 _0553_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1842_ _1293_ B_ADR0 _0486_ _0487_ _0488_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2891_ FrameData[11] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_40_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1773_ Inst_RegFile_32x4.AD_comb\[2\] Inst_RegFile_32x4.AD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ AD2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3443_ FrameStrobe[7] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3374_ E2MID[6] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3512_ Inst_RegFile_switch_matrix.JS2BEG0 net157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2187_ _1355_ _0813_ _0814_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2325_ Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q _0935_ _0937_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2256_ _0134_ _0873_ _0874_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3090_ FrameData[18] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2110_ _1324_ B_ADR0 _0745_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2041_ _0677_ _0675_ _0486_ _0678_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2943_ FrameData[31] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1825_ AD3 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ _0472_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2874_ _0068_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[20\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1756_ _0162_ _0179_ _0405_ _0406_ _0407_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3426_ FrameData[22] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2308_ _0920_ _0921_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1687_ _1303_ A_ADR0 _0340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3357_ Inst_RegFile_switch_matrix.E1BEG1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3288_ FrameData[24] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2239_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0859_ _0860_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ N1END[2] NN4END[2] N2END[6] E1END[2] Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q _0267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2590_ W2MID[6] Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q
+ _1159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_14_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1541_ W1END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ _0201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3211_ FrameData[11] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3142_ FrameData[6] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1472_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2024_ _1334_ B_ADR0 _0486_ _0660_ _0661_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3073_ FrameData[1] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ FrameData[14] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2857_ _0051_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[14\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2788_ _1184_ Inst_RegFile_32x4.mem\[0\]\[1\] _1243_ _0113_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1739_ _1312_ A_ADR0 _0181_ _0389_ _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1808_ Inst_RegFile_32x4.mem\[1\]\[3\] _0147_ _0456_ _0457_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3409_ FrameData[5] net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2711_ _1182_ Inst_RegFile_32x4.mem\[15\]\[0\] _1227_ _0052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1524_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q _0184_ _0185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2573_ _1138_ _1140_ _1142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2642_ _1142_ _1171_ _1203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1455_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _1346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1386_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q _1277_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3125_ FrameData[21] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3056_ FrameData[16] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ _1301_ B_ADR0 _0645_ _0646_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2909_ FrameData[29] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_0_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_17_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_16 WW4END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput145 net145 NN4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput134 net134 N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput123 net123 N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1507_ E6END[0] S2END[4] SS4END[3] W2END[4] Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q _0169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput101 net101 N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput112 net112 N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2556_ _0142_ _0922_ _1124_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _1125_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2625_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q _0961_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q
+ _1191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput156 net156 S1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput167 net167 S2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput178 net178 S4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2487_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q BD1 _1069_ _1070_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput189 net189 SS4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1369_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _1260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3108_ FrameData[4] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1438_ Inst_RegFile_32x4.mem\[9\]\[3\] _1329_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3039_ FrameData[31] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_21_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3390_ EE4END[6] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2410_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q BD2 _1008_ _1009_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2341_ N1END[0] S1END[0] W1END[0] AD3 Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ _0951_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_6_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2272_ N1END[0] E1END[0] N2END[0] E2END[0] Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q _0889_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_35_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1987_ _0625_ _0623_ _0486_ _0626_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2608_ N2MID[6] S2MID[6] W2MID[6] Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q _1177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3588_ W6END[9] net235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2539_ _1290_ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ _1108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1910_ _1295_ B_ADR0 _0486_ _0551_ _0552_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2890_ FrameData[10] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1841_ Inst_RegFile_32x4.mem\[19\]\[0\] B_ADR0 _0487_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1772_ _0300_ _0388_ _0398_ _0411_ _0422_ Inst_RegFile_32x4.AD_comb\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3511_ Inst_RegFile_switch_matrix.S1BEG3 net156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2324_ _0935_ _0936_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3442_ FrameStrobe[6] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3373_ E2MID[5] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2186_ E6END[1] S2END[3] SS4END[2] W2END[3] Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q _0813_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2255_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ _0873_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ Inst_RegFile_32x4.mem\[28\]\[3\] B_ADR0 _0676_ _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2942_ FrameData[30] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2873_ _0067_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[1\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1824_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _0470_ _0471_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1755_ Inst_RegFile_32x4.mem\[28\]\[2\] _0147_ _0406_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1686_ Inst_RegFile_32x4.mem\[15\]\[1\] A_ADR0 _0162_ _0179_ _0339_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3425_ FrameData[21] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2238_ N1END[0] E1END[0] N2END[0] E2END[0] Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q _0859_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2307_ Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q _0917_ _0919_ _0920_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3287_ FrameData[23] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3356_ Inst_RegFile_switch_matrix.E1BEG0 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2169_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q _0797_ _0798_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1540_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q _0196_ _0199_ _0200_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3210_ FrameData[10] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3141_ FrameData[5] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1471_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q _0134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2023_ Inst_RegFile_32x4.mem\[19\]\[3\] B_ADR0 _0660_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3072_ FrameData[0] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2925_ FrameData[13] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2856_ _0050_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[14\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_17_Left_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1807_ Inst_RegFile_32x4.mem\[0\]\[3\] A_ADR0 _0456_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3408_ FrameData[4] net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2787_ _1182_ Inst_RegFile_32x4.mem\[0\]\[0\] _1243_ _0112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1738_ Inst_RegFile_32x4.mem\[3\]\[2\] A_ADR0 _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1669_ _1283_ A_ADR0 _0324_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _0111_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[8\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2710_ _1206_ _1218_ _1227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1523_ W6END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ _0184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2641_ Inst_RegFile_32x4.mem\[25\]\[3\] _1198_ _1202_ _0007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2572_ _1138_ _1140_ _1141_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1454_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q _1345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3124_ FrameData[20] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3055_ FrameData[15] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1385_ WW4END[1] _1276_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_471 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ Inst_RegFile_32x4.mem\[4\]\[1\] B_ADR0 _0645_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2908_ FrameData[28] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2839_ _0033_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[13\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q _1187_ _1189_ _0138_ _1190_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_17 WW4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput135 net135 N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput124 net124 N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput146 net146 NN4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1506_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _0167_ _0168_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput113 net113 N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput102 net102 N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_34_Left_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2555_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q _1123_ _1124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput168 net168 S2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput157 net157 S2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1437_ Inst_RegFile_32x4.mem\[6\]\[3\] _1328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput179 net179 S4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2486_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q _0789_ _1069_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3107_ FrameData[3] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_38_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1368_ S2MID[3] _1259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3038_ FrameData[30] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_43_Left_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Left_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_70_Left_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2271_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0887_ _0888_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q _0947_ _0949_ _0950_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1986_ _1306_ B_ADR0 _0624_ _0625_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2607_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _0998_ _1175_ Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ _1176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3587_ W6END[8] net234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2538_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q _1101_ _1103_ _1106_ _1107_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2469_ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q _1058_ Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ _1059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_547 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1840_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q _0467_ _0469_ _0483_ _0485_ _0486_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_32_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3441_ FrameStrobe[5] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1771_ _0253_ _0416_ _0421_ _0300_ _0422_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_40_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3510_ Inst_RegFile_switch_matrix.S1BEG2 net155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2254_ _0872_ _0869_ Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q Inst_RegFile_switch_matrix.JS2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3372_ E2MID[4] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2323_ Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q _0932_ _0934_ _0935_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2185_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0811_ _0812_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ Inst_RegFile_32x4.mem\[14\]\[0\] B_ADR0 _0609_ _0610_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1823_ W1END[1] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ _0470_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_539 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2872_ _0066_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[1\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2941_ FrameData[29] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3424_ FrameData[20] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1754_ Inst_RegFile_32x4.mem\[29\]\[2\] A_ADR0 _0405_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1685_ Inst_RegFile_32x4.mem\[14\]\[1\] _0147_ _0338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2237_ _0133_ _0857_ _0858_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2306_ _1267_ Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q
+ _0918_ _0919_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_503 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3286_ FrameData[22] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3355_ _0127_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[12\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2099_ Inst_RegFile_32x4.mem\[20\]\[2\] B_ADR0 _0734_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2168_ N1END[1] N2END[3] NN4END[2] E2END[3] Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q _0797_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1470_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3140_ FrameData[4] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3071_ FrameData[31] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2022_ _1333_ B_ADR0 _0658_ _0659_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2924_ FrameData[12] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2855_ _0049_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[14\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1806_ _0448_ _0449_ _0454_ _0254_ _0455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2786_ _1172_ _1212_ _1243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3407_ FrameData[3] net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1599_ _1298_ _0147_ _0255_ _0256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1668_ _1284_ _0147_ _0181_ _0322_ _0323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1737_ _0253_ _0381_ _0387_ _0388_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3338_ _0110_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[8\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3269_ FrameData[5] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2640_ Inst_RegFile_32x4.mem\[25\]\[2\] _1186_ _1202_ _0006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1453_ E2END[2] _1344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1522_ _1297_ _0147_ _0181_ _0182_ _0183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2571_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _1053_ _1139_ _1140_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3123_ FrameData[19] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1384_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _1275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3054_ FrameData[14] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2005_ _1302_ B_ADR0 _0486_ _0643_ _0644_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2907_ FrameData[27] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_61_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2838_ _0032_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[13\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2769_ _1186_ Inst_RegFile_32x4.mem\[5\]\[2\] _1239_ _0098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_18 EE4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput125 net125 N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput114 net114 N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput103 net103 N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2554_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q _1123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2623_ _1280_ Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q
+ _1188_ _1189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput147 net147 NN4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1367_ Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q _1258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput136 net136 N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1505_ N1END[2] N2END[4] N4END[0] E2END[4] Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q _0167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1436_ Inst_RegFile_32x4.mem\[5\]\[3\] _1327_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput169 net169 S2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput158 net158 S2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2485_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q Inst_RegFile_switch_matrix.E2BEG0
+ _1067_ Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q _1068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3106_ FrameData[2] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_55_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3037_ FrameData[29] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0886_ _0887_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1985_ Inst_RegFile_32x4.mem\[20\]\[1\] B_ADR0 _0624_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2606_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q _1041_ _1175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2537_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q _1105_ _1106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3586_ W6END[7] net233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_21_Left_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2399_ N1END[1] E1END[1] S1END[1] AD0 Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q _1000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1419_ Inst_RegFile_32x4.mem\[31\]\[1\] _1310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2468_ _1054_ _1056_ _1057_ Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q _1058_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_43_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_545 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0180_ _0418_ _0420_ _0219_ _0421_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_32_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3440_ FrameStrobe[4] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_40_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3371_ E2MID[3] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2253_ _0871_ _0870_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q _0872_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2184_ N1END[1] N2END[3] N4END[3] E2END[3] Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q _0811_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2322_ _1259_ Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ _0933_ _0934_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1899_ _0536_ _0537_ _0540_ _0541_ Inst_RegFile_switch_matrix.JW2BEG6 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1968_ _1286_ B_ADR0 _0609_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3569_ Inst_RegFile_switch_matrix.JW2BEG4 net214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2940_ FrameData[28] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1822_ _1260_ _0468_ _0469_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1753_ _0180_ _0400_ _0403_ _0219_ _0404_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2871_ _0065_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[1\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3423_ FrameData[19] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3354_ _0126_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[12\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1684_ _0180_ _0334_ _0335_ _0336_ _0337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2167_ _1354_ _0795_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q _0796_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2236_ S1END[0] S2END[0] S1END[2] W1END[0] Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q _0857_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2305_ Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q Inst_RegFile_switch_matrix.JS2BEG3
+ _0918_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3285_ FrameData[21] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2098_ _1321_ B_ADR0 _0486_ _0732_ _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_0_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ Inst_RegFile_32x4.mem\[16\]\[3\] B_ADR0 _0658_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3070_ FrameData[30] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2923_ FrameData[11] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2854_ _0048_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[14\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1805_ _0450_ _0451_ _0453_ _0180_ _0219_ _0454_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2785_ _1198_ Inst_RegFile_32x4.mem\[8\]\[3\] _1242_ _0111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1736_ _0180_ _0383_ _0386_ _0218_ _0387_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3406_ FrameData[2] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1598_ Inst_RegFile_32x4.mem\[28\]\[0\] _0147_ _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1667_ Inst_RegFile_32x4.mem\[10\]\[0\] _0147_ _0322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3337_ _0109_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[8\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3199_ FrameData[31] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3268_ FrameData[4] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2219_ _0132_ _0841_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q _0842_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2570_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _1019_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ _1139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1452_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q _1343_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3122_ FrameData[18] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1383_ E2MID[0] _1274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1521_ Inst_RegFile_32x4.mem\[26\]\[0\] _0147_ _0182_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3053_ FrameData[13] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_23_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2004_ Inst_RegFile_32x4.mem\[7\]\[1\] B_ADR0 _0643_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2906_ FrameData[26] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2699_ Inst_RegFile_32x4.mem\[22\]\[3\] _1198_ _1224_ _0043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1719_ Inst_RegFile_32x4.mem\[23\]\[1\] A_ADR0 _0372_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2768_ _1184_ Inst_RegFile_32x4.mem\[5\]\[1\] _1239_ _0097_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2837_ _0031_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[9\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_19 FrameStrobe[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput126 net126 N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput148 net148 NN4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput137 net137 NN4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1504_ _1289_ _0165_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q _0166_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput115 net115 N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput104 net104 N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2553_ _1107_ _1121_ _1122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2622_ N4END[0] Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q _1188_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput159 net159 S2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1366_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q _1257_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3105_ FrameData[1] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_28_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q _0195_ _1067_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1435_ Inst_RegFile_32x4.mem\[2\]\[3\] _1326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_38_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3036_ FrameData[28] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_21_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ Inst_RegFile_32x4.mem\[22\]\[1\] Inst_RegFile_32x4.mem\[23\]\[1\] B_ADR0 _0623_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2536_ _1353_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ _1104_ _1105_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2605_ _1135_ _1173_ _1174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_509 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2467_ N2MID[1] E2MID[1] Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q _1057_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3585_ W6END[6] net232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2398_ BD0 _0213_ _0497_ _0998_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ _0999_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1418_ Inst_RegFile_32x4.mem\[28\]\[1\] _1309_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3019_ FrameData[11] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_59_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3370_ E2MID[2] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2321_ W2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q _0933_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2252_ N1END[0] E1END[0] N2END[0] E2END[0] Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q _0871_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2183_ _1355_ _0809_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q _0810_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_48_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1898_ _1275_ _0538_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q _0541_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1967_ _0605_ _0607_ _0486_ _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2519_ BD0 _0468_ Inst_RegFile_switch_matrix.JW2BEG1 _0530_ Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q Inst_RegFile_switch_matrix.N1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3568_ Inst_RegFile_switch_matrix.JW2BEG3 net213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3499_ NN4END[11] net150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_516 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Left_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2870_ _0064_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[1\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1821_ N2MID[3] E2MID[3] S2MID[3] W2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q _0468_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1752_ _0162_ _0179_ _0401_ _0402_ _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1683_ Inst_RegFile_32x4.mem\[11\]\[1\] A_ADR0 _0162_ _0179_ _0336_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3422_ FrameData[18] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2304_ N2MID[4] E2MID[4] Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q _0917_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3284_ FrameData[20] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3353_ _0125_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[12\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2097_ Inst_RegFile_32x4.mem\[23\]\[2\] B_ADR0 _0732_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2166_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ _0795_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2235_ _0133_ _0855_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q _0856_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2999_ FrameData[23] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2020_ Inst_RegFile_32x4.BD_comb\[1\] Inst_RegFile_32x4.BD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ BD1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2853_ _0047_ clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.mem\[23\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2922_ FrameData[10] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ Inst_RegFile_32x4.mem\[12\]\[3\] A_ADR0 _0452_ _0453_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1735_ _0162_ _0179_ _0384_ _0385_ _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1666_ _0313_ _0316_ _0320_ _0218_ _0253_ _0321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2784_ _1186_ Inst_RegFile_32x4.mem\[8\]\[2\] _1242_ _0110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3405_ FrameData[1] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3267_ FrameData[3] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1597_ _0239_ _0252_ _0254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3336_ _0108_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[8\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3198_ FrameData[30] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2149_ _0779_ _0776_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q Inst_RegFile_switch_matrix.JN2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ _0841_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1520_ _0162_ _0179_ _0181_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3121_ FrameData[17] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1451_ W2END[7] _1342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1382_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q _1273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3052_ FrameData[12] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2003_ _0486_ _0639_ _0641_ _0518_ _0642_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_61_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2905_ FrameData[25] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2836_ _0030_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[9\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2698_ Inst_RegFile_32x4.mem\[22\]\[2\] _1186_ _1224_ _0042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1649_ Inst_RegFile_32x4.mem\[16\]\[0\] A_ADR0 _0303_ _0304_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1718_ Inst_RegFile_32x4.mem\[20\]\[1\] A_ADR0 _0370_ _0371_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2767_ _1182_ Inst_RegFile_32x4.mem\[5\]\[0\] _1239_ _0096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3319_ _0091_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[3\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput138 net138 NN4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput149 net149 NN4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput127 net127 N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1503_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ _0165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput116 net116 N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput105 net105 N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2621_ S4END[0] Inst_RegFile_switch_matrix.JW2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q
+ _1187_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2483_ BD2 _0468_ Inst_RegFile_switch_matrix.E2BEG1 _0530_ Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q Inst_RegFile_switch_matrix.S1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2552_ _1112_ _1115_ _1119_ _1121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_533 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1365_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _1256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3104_ FrameData[0] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1434_ Inst_RegFile_32x4.mem\[31\]\[2\] _1325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3035_ FrameData[27] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ _0013_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[27\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_547 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1983_ _0517_ _0619_ _0622_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2604_ _1142_ _1149_ _1169_ _1173_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1417_ Inst_RegFile_32x4.mem\[26\]\[1\] _1308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2535_ N2END[0] Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _1104_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2466_ Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q _1055_ _1056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3584_ W6END[5] net231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2397_ N2END[6] E2END[6] SS4END[3] W2END[6] Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q _0998_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3018_ FrameData[10] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_43_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_536 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_514 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_539 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ S1END[0] S2END[0] SS4END[0] W1END[0] Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q _0870_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2320_ N2MID[3] E2MID[3] Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q _0932_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2182_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ _0809_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1966_ Inst_RegFile_32x4.mem\[10\]\[0\] B_ADR0 _0606_ _0607_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1897_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0539_ _0540_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3567_ Inst_RegFile_switch_matrix.JW2BEG2 net212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2518_ Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q _1090_ _1088_ Inst_RegFile_switch_matrix.N1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2449_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q _1041_ _1042_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3498_ NN4END[10] net149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1820_ _0287_ _0289_ _0291_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0467_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_45_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ FrameData[17] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1751_ Inst_RegFile_32x4.mem\[24\]\[2\] _0147_ _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1682_ Inst_RegFile_32x4.mem\[10\]\[1\] _0147_ _0335_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3283_ FrameData[19] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2234_ AD3 BD0 BD1 BD2 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ _0855_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2303_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0212_ _0915_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ _0916_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3352_ _0124_ clknet_4_5_0_UserCLK_regs Inst_RegFile_32x4.mem\[12\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2165_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q _0793_ _0794_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2096_ _0486_ _0728_ _0730_ _0518_ _0731_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2998_ FrameData[22] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1949_ Inst_RegFile_32x4.mem\[28\]\[0\] B_ADR0 _0589_ _0590_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_16_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_528 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2852_ _0046_ clknet_4_14_0_UserCLK_regs Inst_RegFile_32x4.mem\[23\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2921_ FrameData[9] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2783_ _1184_ Inst_RegFile_32x4.mem\[8\]\[1\] _1242_ _0109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1803_ _1331_ A_ADR0 _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_68_Left_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3404_ FrameData[0] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1665_ _0317_ _0319_ _0181_ _0320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1596_ _0239_ _0252_ _0253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1734_ Inst_RegFile_32x4.mem\[12\]\[2\] _0147_ _0385_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3197_ FrameData[29] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3266_ FrameData[2] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3335_ _0107_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[7\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2217_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q _0839_ _0840_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2148_ _0777_ _0778_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q _0779_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2079_ _0550_ _0709_ _0713_ _0714_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1450_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q _1341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_10_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3120_ FrameData[16] FrameStrobe[5] Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3051_ FrameData[11] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1381_ Inst_RegFile_32x4.mem\[6\]\[0\] _1272_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_61_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2002_ _1300_ B_ADR0 _0486_ _0640_ _0641_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2904_ FrameData[24] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2766_ _1200_ _1237_ _1239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2835_ _0029_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[9\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1648_ _1292_ A_ADR0 _0303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1717_ _1306_ A_ADR0 _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2697_ Inst_RegFile_32x4.mem\[22\]\[1\] _1184_ _1224_ _0041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1579_ _1279_ Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ _0236_ _0237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3318_ _0090_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.mem\[3\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3249_ FrameData[17] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ Inst_RegFile_32x4.mem\[24\]\[2\] _1186_ _1174_ _0002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput139 net139 NN4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput128 net128 N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput117 net117 N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1502_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _0163_ _0164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput106 net106 N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1433_ Inst_RegFile_32x4.mem\[29\]\[2\] _1324_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2482_ _1064_ _1066_ Inst_RegFile_switch_matrix.S1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2551_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q _1117_ _1118_ _1116_ _1120_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3034_ FrameData[26] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1364_ EE4END[1] _1255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3103_ FrameData[31] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2818_ _0012_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[27\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2749_ Inst_RegFile_32x4.mem\[29\]\[3\] _1198_ _1234_ _0083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_7_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_7_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_52_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1982_ _1305_ B_ADR0 _0486_ _0620_ _0621_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_43_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2534_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _0156_ _1102_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ _1103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2603_ _1141_ _1171_ _1172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3583_ W6END[4] net230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2396_ _0990_ _0991_ _0997_ _0996_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q
+ Inst_RegFile_switch_matrix.E6BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1416_ Inst_RegFile_32x4.mem\[24\]\[1\] _1307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2465_ W2MID[1] Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q _1055_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3017_ FrameData[9] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_6_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2250_ _0868_ _0867_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q _0869_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2181_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q _0807_ _0808_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Left_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1965_ _1284_ B_ADR0 _0606_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1896_ S1END[1] S2END[7] S1END[3] W1END[3] Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q _0539_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2517_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q BD1 _1089_ _1090_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3566_ Inst_RegFile_switch_matrix.JW2BEG1 net211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3497_ NN4END[9] net148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2379_ _0137_ _0981_ _0982_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2448_ Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q _1038_ _1040_ _1041_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1750_ Inst_RegFile_32x4.mem\[25\]\[2\] A_ADR0 _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3420_ FrameData[16] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ _0123_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[11\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1681_ Inst_RegFile_32x4.mem\[9\]\[1\] _0147_ _0333_ _0334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3282_ FrameData[18] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2164_ W6END[1] AD0 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ _0793_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2302_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0497_ _0915_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2233_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q _0853_ _0854_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2095_ _1319_ B_ADR0 _0486_ _0729_ _0730_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1879_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q _0522_ _0523_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2997_ FrameData[21] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1948_ _1298_ B_ADR0 _0589_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3549_ SS4END[9] net200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2920_ FrameData[8] FrameStrobe[11] Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2851_ _0045_ clknet_4_11_0_UserCLK_regs Inst_RegFile_32x4.mem\[23\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2782_ _1182_ Inst_RegFile_32x4.mem\[8\]\[0\] _1242_ _0108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1733_ Inst_RegFile_32x4.mem\[13\]\[2\] A_ADR0 _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1802_ Inst_RegFile_32x4.mem\[15\]\[3\] A_ADR0 _0162_ _0179_ _0451_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3403_ Inst_RegFile_switch_matrix.EE4BEG3 net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1664_ _1272_ A_ADR0 _0318_ _0319_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3334_ _0106_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[7\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1595_ _0250_ _0251_ _0252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3196_ FrameData[28] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2147_ E6END[0] S2END[4] W2END[4] WW4END[3] Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q _0778_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3265_ FrameData[1] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2216_ W6END[0] AD0 AD2 AD3 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ _0839_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_64_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2078_ _0486_ _0712_ _0711_ _0517_ _0713_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1380_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q _1271_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3050_ FrameData[10] FrameStrobe[7] Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2001_ Inst_RegFile_32x4.mem\[3\]\[1\] B_ADR0 _0640_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2903_ FrameData[23] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2696_ Inst_RegFile_32x4.mem\[22\]\[0\] _1182_ _1224_ _0040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1716_ _0180_ _0368_ _0366_ _0218_ _0369_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2765_ _1198_ Inst_RegFile_32x4.mem\[4\]\[3\] _1238_ _0095_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2834_ _0028_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[9\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1647_ Inst_RegFile_32x4.mem\[19\]\[0\] A_ADR0 _0162_ _0179_ _0301_ _0302_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3317_ _0089_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[3\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1578_ W2END[1] Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q _0236_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3248_ FrameData[16] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3179_ FrameData[11] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_15_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_26_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput107 net107 N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2550_ _0144_ _1114_ _1118_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q _1119_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput129 net129 N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput118 net118 N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1363_ S2MID[2] _1254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1501_ W6END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ _0163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1432_ Inst_RegFile_32x4.mem\[27\]\[2\] _1323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2481_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q Inst_RegFile_switch_matrix.E2BEG2
+ _1065_ Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q _1066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3033_ FrameData[25] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3102_ FrameData[30] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2748_ Inst_RegFile_32x4.mem\[29\]\[2\] _1186_ _1234_ _0082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2817_ _0011_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[26\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2679_ _1186_ Inst_RegFile_32x4.mem\[9\]\[2\] _1217_ _0030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_549 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ Inst_RegFile_32x4.mem\[19\]\[1\] B_ADR0 _0620_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2533_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q _0215_ _1102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2602_ _1149_ _1169_ _1171_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3582_ W6END[3] net229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2395_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ _0997_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1415_ Inst_RegFile_32x4.mem\[21\]\[1\] _1306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2464_ _1278_ Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q _1054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3016_ FrameData[8] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2180_ W6END[1] AD0 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ _0807_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_0_Left_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_65_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1895_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q _0538_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1964_ Inst_RegFile_32x4.mem\[8\]\[0\] B_ADR0 _0604_ _0605_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2516_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q _0573_ _1089_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2447_ _1250_ Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q
+ _1039_ _1040_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3565_ Inst_RegFile_switch_matrix.JW2BEG0 net210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3496_ NN4END[8] net147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2378_ AD0 AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ _0981_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_47_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2301_ _0136_ _0913_ _0914_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1680_ Inst_RegFile_32x4.mem\[8\]\[1\] A_ADR0 _0333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3350_ _0122_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[11\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2163_ _0791_ _0792_ A_ADR0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2232_ WW4END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ _0853_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3281_ FrameData[17] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2094_ Inst_RegFile_32x4.mem\[19\]\[2\] B_ADR0 _0729_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1878_ WW4END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ _0522_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2996_ FrameData[20] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1947_ Inst_RegFile_32x4.mem\[30\]\[0\] B_ADR0 _0587_ _0588_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3548_ SS4END[8] net199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_59_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3479_ N4END[7] net130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2850_ _0044_ clknet_4_15_0_UserCLK_regs Inst_RegFile_32x4.mem\[23\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1663_ Inst_RegFile_32x4.mem\[7\]\[0\] A_ADR0 _0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1732_ _1317_ _0147_ _0382_ _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1801_ Inst_RegFile_32x4.mem\[14\]\[3\] _0147_ _0450_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2781_ _1172_ _1216_ _1242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3402_ Inst_RegFile_switch_matrix.EE4BEG2 net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3264_ FrameData[0] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3333_ _0105_ clknet_4_4_0_UserCLK_regs Inst_RegFile_32x4.mem\[7\]\[1\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1594_ _1350_ _0248_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q _0251_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3195_ FrameData[27] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2146_ N2END[4] N4END[0] E1END[2] E2END[4] Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q _0777_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] B_ADR0 _0712_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2215_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q _0836_ _0838_ _0832_ _0834_ Inst_RegFile_switch_matrix.JS2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_64_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2979_ FrameData[3] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2000_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] B_ADR0 _0639_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2902_ FrameData[22] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_61_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2833_ _0027_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[30\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1646_ _1293_ A_ADR0 _0301_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2695_ _1204_ _1223_ _1224_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1715_ Inst_RegFile_32x4.mem\[17\]\[1\] A_ADR0 _0367_ _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2764_ _1186_ Inst_RegFile_32x4.mem\[4\]\[2\] _1238_ _0094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3247_ FrameData[15] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1577_ NN4END[2] E2END[1] Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q _0235_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3316_ _0088_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[3\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3178_ FrameData[10] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2129_ Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q _0760_ _0761_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput119 net119 N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1500_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _0156_ _0161_ _0162_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput108 net108 N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2480_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q _1041_ _1065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput90 net90 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1431_ Inst_RegFile_32x4.mem\[25\]\[2\] _1322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3101_ FrameData[29] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1362_ Inst_RegFile_32x4.mem\[1\]\[0\] _1253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3032_ FrameData[24] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2816_ _0010_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[26\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1629_ EE4END[1] S1END[1] S1END[3] S2END[7] Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q _0285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2747_ Inst_RegFile_32x4.mem\[29\]\[1\] _1184_ _1234_ _0081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2678_ _1184_ Inst_RegFile_32x4.mem\[9\]\[1\] _1217_ _0029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ Inst_RegFile_32x4.mem\[17\]\[1\] B_ADR0 _0486_ _0618_ _0619_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q _1164_ _1167_ _1155_ _1156_ _1170_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2532_ _1100_ _1101_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2463_ Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q _1050_ _1051_ _1052_ _1053_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3581_ W6END[2] net226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2394_ _0993_ _0995_ _0996_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1414_ Inst_RegFile_32x4.mem\[18\]\[1\] _1305_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3015_ FrameData[7] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_3_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1894_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0534_ _1277_ _0537_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1963_ _1283_ B_ADR0 _0604_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2515_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q Inst_RegFile_switch_matrix.JW2BEG2
+ _1087_ Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q _1088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2446_ Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q Inst_RegFile_switch_matrix.JN2BEG1
+ _1039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3495_ NN4END[7] net146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3564_ Inst_RegFile_switch_matrix.W1BEG3 net209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2377_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0979_ _0980_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2231_ _0852_ _0849_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q Inst_RegFile_switch_matrix.JN2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3280_ FrameData[16] FrameStrobe[0] Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2300_ AD0 AD2 AD1 AD3 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ _0913_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2093_ _1318_ B_ADR0 _0727_ _0728_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2162_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _0783_ _0782_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ _0792_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2995_ FrameData[19] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_16_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3547_ SS4END[7] net198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1877_ _0486_ _0520_ _0518_ _0488_ _0521_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_8_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1946_ _1299_ B_ADR0 _0587_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2429_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q _1024_ _1025_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_59_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3478_ N4END[6] net129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0181_ _0446_ _0218_ _0449_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3401_ Inst_RegFile_switch_matrix.EE4BEG1 net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2780_ _1198_ Inst_RegFile_32x4.mem\[7\]\[3\] _1241_ _0107_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1662_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] A_ADR0 _0317_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1731_ Inst_RegFile_32x4.mem\[14\]\[2\] _0147_ _0382_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3194_ FrameData[26] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_37_Left_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3263_ FrameData[31] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3332_ _0104_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[7\]\[0\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1593_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _0249_ _0250_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2214_ _0131_ _0837_ _0838_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2145_ _0774_ _0775_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q _0776_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2076_ _1313_ B_ADR0 _0486_ _0710_ _0711_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_46_Left_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2978_ FrameData[2] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1929_ E2MID[2] W2MID[2] S2MID[2] Inst_RegFile_switch_matrix.E2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q _0570_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_523 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Left_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2901_ FrameData[21] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2832_ _0026_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[30\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2763_ _1184_ Inst_RegFile_32x4.mem\[4\]\[1\] _1238_ _0093_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1645_ _0274_ _0278_ _0299_ _0300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1714_ _1304_ A_ADR0 _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2694_ _1133_ _1220_ _1223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1576_ Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q _0233_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ _0234_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3177_ FrameData[9] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3246_ FrameData[14] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3315_ _0087_ clknet_4_7_0_UserCLK_regs Inst_RegFile_32x4.mem\[31\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2128_ Inst_RegFile_switch_matrix.JN2BEG4 _0760_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_24_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ _1332_ B_ADR0 _0696_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1430_ Inst_RegFile_32x4.mem\[22\]\[2\] _1321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput109 net109 N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput1 net1 E1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput91 net91 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3031_ FrameData[23] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput80 net80 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1361_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _1252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3100_ FrameData[28] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2815_ _0009_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[26\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2746_ Inst_RegFile_32x4.mem\[29\]\[0\] _1182_ _1234_ _0080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_21_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1628_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0283_ _0284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1559_ _0200_ _0217_ _0218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2677_ _1182_ Inst_RegFile_32x4.mem\[9\]\[0\] _1217_ _0028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3229_ FrameData[29] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_11_0_UserCLK_regs clknet_0_UserCLK_regs clknet_4_11_0_UserCLK_regs VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2600_ _1165_ _1168_ _1157_ _1169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3580_ W2MID[7] net225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2393_ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q _0468_ _0994_ _0995_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1413_ Inst_RegFile_32x4.mem\[16\]\[1\] _1304_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2531_ _0961_ Inst_RegFile_switch_matrix.JN2BEG7 Inst_RegFile_switch_matrix.JS2BEG7
+ Inst_RegFile_switch_matrix.JW2BEG7 Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ _1100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2462_ _1342_ Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q
+ _1052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3014_ FrameData[6] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2729_ _1198_ Inst_RegFile_32x4.mem\[1\]\[3\] _1230_ _0067_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_554 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0550_ _0598_ _0602_ _0603_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_18_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _1275_ _0535_ _0536_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3563_ Inst_RegFile_switch_matrix.W1BEG2 net208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2376_ NN4END[3] SS4END[3] E1END[2] W1END[2] Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q _0979_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2514_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q _1041_ _1087_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2445_ NN4END[3] S4END[3] Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q _1038_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3494_ NN4END[6] net145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _0850_ _0851_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0852_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2092_ Inst_RegFile_32x4.mem\[16\]\[2\] B_ADR0 _0727_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2161_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _0785_ _0790_ _0791_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2994_ FrameData[18] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1945_ _0583_ _0585_ _0486_ _0586_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_16_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3546_ SS4END[6] net197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1876_ _1292_ B_ADR0 _0519_ _0520_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_8_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2428_ N1END[0] E1END[0] W1END[0] AD3 Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q _1024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2359_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _0468_ _0964_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ _0965_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ N4END[5] net128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3400_ Inst_RegFile_switch_matrix.EE4BEG0 net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1592_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q _0249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3331_ _0103_ clknet_4_1_0_UserCLK_regs Inst_RegFile_32x4.mem\[6\]\[3\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ _0180_ _0315_ _0218_ _0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1730_ _0180_ _0377_ _0380_ _0219_ _0381_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3193_ FrameData[25] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2144_ BD0 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ _0775_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3262_ FrameData[30] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2213_ S2END[2] S4END[2] W2END[2] WW4END[1] Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q _0837_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_64_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2075_ Inst_RegFile_32x4.mem\[7\]\[2\] B_ADR0 _0710_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1859_ _1270_ _0503_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q _0504_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2977_ FrameData[1] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1928_ _0565_ _0568_ _0569_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3529_ S4END[5] net180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ FrameData[20] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1713_ Inst_RegFile_32x4.mem\[19\]\[1\] A_ADR0 _0162_ _0179_ _0365_ _0366_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2831_ _0025_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[30\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2762_ _1182_ Inst_RegFile_32x4.mem\[4\]\[0\] _1238_ _0092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1644_ _0294_ _0295_ _0298_ _0299_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2693_ Inst_RegFile_32x4.mem\[17\]\[3\] _1198_ _1222_ _0039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3314_ _0086_ clknet_4_6_0_UserCLK_regs Inst_RegFile_32x4.mem\[31\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1575_ EE4END[3] S4END[0] Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q _0233_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3176_ FrameData[8] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2127_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q _0757_ _0759_ _0753_ _0755_ Inst_RegFile_switch_matrix.JN2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3245_ FrameData[13] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_16_Left_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2058_ _0692_ _0694_ _0486_ _0695_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput70 net70 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1360_ EE4END[0] _1251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput2 net2 E1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput92 net92 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput81 net81 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3030_ FrameData[22] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_31_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _0008_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[26\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2745_ _1201_ _1209_ _1234_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2676_ _1200_ _1216_ _1217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1489_ EE4END[2] S1END[0] S1END[2] S2END[6] Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q _0152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1627_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q _0283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1558_ _1345_ _0213_ _0216_ Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q _0217_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3228_ FrameData[28] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3159_ FrameData[23] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2530_ _1097_ _1099_ Inst_RegFile_switch_matrix.N1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q _0160_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ _0994_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2461_ Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q Inst_RegFile_switch_matrix.E2BEG2
+ _1051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1412_ Inst_RegFile_32x4.mem\[13\]\[1\] _1303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_552 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3013_ FrameData[5] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2659_ Inst_RegFile_32x4.mem\[28\]\[1\] _1184_ _1210_ _0017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2728_ _1186_ Inst_RegFile_32x4.mem\[1\]\[2\] _1230_ _0066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_19_Left_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ WW4END[1] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ _0535_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ _0486_ _0601_ _0600_ _0517_ _0602_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ N2END[2] N4END[1] E6END[1] BD0 Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q Inst_RegFile_switch_matrix.N4BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3493_ NN4END[5] net144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3562_ Inst_RegFile_switch_matrix.W1BEG1 net207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2444_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q _1035_ _1037_ Inst_RegFile_switch_matrix.NN4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2375_ _0978_ _0977_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q Inst_RegFile_switch_matrix.SS4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2160_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q _0789_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ _0790_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ _0549_ _0725_ _0581_ _0726_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1875_ Inst_RegFile_32x4.mem\[16\]\[0\] B_ADR0 _0519_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2993_ FrameData[17] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1944_ Inst_RegFile_32x4.mem\[26\]\[0\] B_ADR0 _0584_ _0585_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_16_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3545_ SS4END[5] net196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2427_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q _1020_ _1022_ _1023_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3476_ N4END[4] net121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2289_ _0903_ _0902_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q _0904_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2358_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _0272_ _0964_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ _0102_ clknet_4_0_0_UserCLK_regs Inst_RegFile_32x4.mem\[6\]\[2\] VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1591_ E2MID[0] W2MID[0] S2MID[0] Inst_RegFile_switch_matrix.JW2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q _0248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1660_ Inst_RegFile_32x4.mem\[0\]\[0\] A_ADR0 _0314_ _0315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3192_ FrameData[24] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2143_ W6END[0] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ _0774_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3261_ FrameData[29] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2212_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0835_ _0836_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2074_ _0486_ _0706_ _0708_ _0518_ _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1858_ AD3 BD2 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ _0503_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2976_ FrameData[0] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1927_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _0566_ _0567_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q
+ _0568_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3528_ S4END[4] net173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3459_ Inst_RegFile_switch_matrix.N1BEG3 net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1789_ _0180_ _0437_ _0435_ _0218_ _0438_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_57_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_469 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2830_ _0024_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[30\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_1 E6END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1643_ _0296_ _0297_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q _0298_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1712_ _1305_ A_ADR0 _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2692_ Inst_RegFile_32x4.mem\[17\]\[2\] _1186_ _1222_ _0038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2761_ _1172_ _1237_ _1238_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3244_ FrameData[12] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3313_ _0085_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.mem\[31\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1574_ Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q Inst_RegFile_switch_matrix.JW2BEG3
+ _0231_ _0232_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2126_ _1252_ _0758_ _0759_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2057_ Inst_RegFile_32x4.mem\[10\]\[3\] B_ADR0 _0693_ _0694_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3175_ FrameData[7] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2959_ FrameData[15] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput93 net93 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput82 net82 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput60 net60 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput71 net71 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput3 net3 E1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ _0007_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[25\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1626_ _1256_ _0281_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q _0282_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2744_ Inst_RegFile_32x4.mem\[19\]\[3\] _1198_ _1233_ _0079_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2675_ _1133_ _1215_ _1216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1488_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q _0150_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q
+ _0151_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3227_ FrameData[27] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1557_ _1345_ _0215_ _0216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3158_ FrameData[22] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3089_ FrameData[17] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2109_ Inst_RegFile_32x4.mem\[30\]\[2\] B_ADR0 _0743_ _0744_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ N4END[2] E2END[2] Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q _1050_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2391_ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q _0930_ _0992_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ _0993_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1411_ Inst_RegFile_32x4.mem\[6\]\[1\] _1302_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3012_ FrameData[4] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2589_ _0140_ Inst_RegFile_switch_matrix.JN2BEG4 _1158_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1609_ _1341_ _0265_ _0266_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2658_ Inst_RegFile_32x4.mem\[28\]\[0\] _1182_ _1210_ _0016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2727_ _1184_ Inst_RegFile_32x4.mem\[1\]\[1\] _1230_ _0065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_509 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1891_ AD3 BD0 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ _0534_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] B_ADR0 _0601_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2443_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q _1036_ _1037_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2512_ N2END[3] N4END[2] E6END[0] BD1 Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q Inst_RegFile_switch_matrix.N4BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3492_ NN4END[4] net137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3561_ Inst_RegFile_switch_matrix.W1BEG0 net206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2374_ N1END[2] E1END[2] W1END[2] AD1 Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q _0978_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_523 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput250 net250 WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _0719_ _0724_ _0517_ _0725_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2992_ FrameData[16] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q _0498_ _0499_ _0516_ _0518_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1943_ _1297_ B_ADR0 _0584_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3544_ SS4END[4] net189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3475_ N2MID[7] net120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2426_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q _0160_ _1021_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ _1022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2288_ N1END[0] N2END[0] NN4END[0] E1END[0] Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q _0903_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_67_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2357_ _0963_ _0962_ Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q Inst_RegFile_switch_matrix.SS4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_50_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ _0241_ _0243_ _0246_ _0247_ Inst_RegFile_switch_matrix.JW2BEG5 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3260_ FrameData[28] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3191_ FrameData[23] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2142_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q _0771_ _0773_ _0767_ B_ADR0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_22_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2073_ _1312_ B_ADR0 _0486_ _0707_ _0708_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2211_ N2END[2] E2END[2] E1END[0] E6END[0] Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q _0835_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_64_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2975_ FrameData[31] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1857_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q _0501_ _0502_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1788_ Inst_RegFile_32x4.mem\[16\]\[3\] A_ADR0 _0436_ _0437_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3527_ S2MID[7] net172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1926_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_switch_matrix.JN2BEG6
+ _0567_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3389_ EE4END[5] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3458_ Inst_RegFile_switch_matrix.N1BEG2 net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2409_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q _0920_ _1008_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Left_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_2 FrameStrobe[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1642_ S2END[1] Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ _0297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2691_ Inst_RegFile_32x4.mem\[17\]\[1\] _1184_ _1222_ _0037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1711_ _0355_ _0358_ _0363_ _0218_ _0254_ _0364_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2760_ _1134_ _1211_ _1237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_60_Left_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3243_ FrameData[11] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3312_ _0084_ clknet_4_12_0_UserCLK_regs Inst_RegFile_32x4.mem\[31\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1573_ _1276_ Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q
+ _0231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2125_ E2END[5] S1END[1] S2END[5] W1END[1] Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q _0758_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3174_ FrameData[6] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2056_ _1330_ B_ADR0 _0693_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1909_ Inst_RegFile_32x4.mem\[23\]\[0\] B_ADR0 _0551_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2958_ FrameData[14] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2889_ FrameData[9] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput94 net94 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput61 net61 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput50 net50 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput72 net72 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput83 net83 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput4 net4 E1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2743_ Inst_RegFile_32x4.mem\[19\]\[2\] _1186_ _1233_ _0078_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2812_ _0006_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[25\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1625_ AD3 BD0 BD1 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ _0281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1556_ _0214_ _0215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2674_ _1107_ _1120_ _1215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_67_551 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1487_ W1END[2] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ _0150_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3226_ FrameData[26] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3157_ FrameData[21] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3088_ FrameData[16] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2108_ _1325_ B_ADR0 _0743_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2039_ _1339_ B_ADR0 _0676_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1410_ Inst_RegFile_32x4.mem\[5\]\[1\] _1301_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2390_ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q _0935_ _0992_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3011_ FrameData[3] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_64_543 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2726_ _1182_ Inst_RegFile_32x4.mem\[1\]\[0\] _1230_ _0064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1608_ E2END[6] S1END[2] S2END[6] W1END[0] Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q _0265_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2588_ _1155_ _1156_ _1157_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2657_ _1173_ _1209_ _1210_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1539_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q _0198_ Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q
+ _0199_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3209_ FrameData[9] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_47_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_535 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3560_ clknet_1_0__leaf_UserCLK net205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _1282_ _0532_ _0533_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3491_ Inst_RegFile_switch_matrix.N4BEG3 net127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2442_ N1END[2] E1END[2] W1END[2] AD1 Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q _1036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2511_ N2END[0] W6END[1] N4END[3] BD2 Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q Inst_RegFile_switch_matrix.N4BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2373_ BD1 _0930_ _0936_ _0531_ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ _0977_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2709_ _1198_ Inst_RegFile_32x4.mem\[14\]\[3\] _1226_ _0051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput251 net251 WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput240 net240 WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_557 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ FrameData[15] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ Inst_RegFile_32x4.mem\[24\]\[0\] B_ADR0 _0582_ _0583_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ _1271_ _0500_ _0513_ _0515_ _0517_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3543_ Inst_RegFile_switch_matrix.S4BEG3 net179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2425_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q BD3 _1021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3474_ N2MID[6] net119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2356_ N1END[1] E1END[1] W1END[1] AD0 Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q _0963_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_67_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2287_ E2END[0] S2END[0] S1END[0] W1END[0] Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q _0902_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_50_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_516 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3190_ FrameData[22] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2210_ _0131_ _0833_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q _0834_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _1249_ _0772_ _0773_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2072_ Inst_RegFile_32x4.mem\[3\]\[2\] B_ADR0 _0707_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2974_ FrameData[30] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1925_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q _0238_ _0566_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1856_ W1END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ _0501_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1787_ _1333_ A_ADR0 _0436_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3526_ S2MID[6] net171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3388_ EE4END[4] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3457_ Inst_RegFile_switch_matrix.N1BEG1 net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2408_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q _1005_ _1007_ Inst_RegFile_switch_matrix.EE4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2339_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q _0160_ _0948_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ _0949_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_3 FrameStrobe[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1641_ N2END[1] _1352_ _0296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2690_ Inst_RegFile_32x4.mem\[17\]\[0\] _1182_ _1222_ _0036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1572_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q _0228_ _0230_ _0224_ _0226_ Inst_RegFile_switch_matrix.JW2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1710_ _0360_ _0362_ _0181_ _0363_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3311_ _0083_ clknet_4_13_0_UserCLK_regs Inst_RegFile_32x4.mem\[29\]\[3\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2124_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0756_ _0757_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3242_ FrameData[10] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3173_ FrameData[5] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2055_ Inst_RegFile_32x4.mem\[8\]\[3\] B_ADR0 _0691_ _0692_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1839_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0484_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q
+ _0485_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2957_ FrameData[13] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1908_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q _0548_ _0533_ _0550_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2888_ FrameData[8] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3509_ Inst_RegFile_switch_matrix.S1BEG1 net154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput5 net5 E2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput95 net95 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput84 net84 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput62 net62 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput73 net73 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput51 net51 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput40 net40 EE4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2742_ Inst_RegFile_32x4.mem\[19\]\[1\] _1184_ _1233_ _0077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2811_ _0005_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.mem\[25\]\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1624_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0279_ _0280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1555_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q _0214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2673_ Inst_RegFile_32x4.mem\[30\]\[3\] _1198_ _1214_ _0027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1486_ _1343_ _0148_ _0149_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3225_ FrameData[25] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3156_ FrameData[20] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2107_ _0739_ _0741_ _0486_ _0742_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3087_ FrameData[15] FrameStrobe[6] Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2038_ Inst_RegFile_32x4.mem\[30\]\[3\] B_ADR0 _0674_ _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3010_ FrameData[2] FrameStrobe[8] Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2656_ _1122_ _1133_ _1209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2725_ _1200_ _1212_ _1230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1607_ _1341_ _0263_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q _0264_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2587_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q _1001_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ _1156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1538_ _0197_ _0198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1469_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q _0132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3208_ FrameData[8] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3139_ FrameData[3] FrameStrobe[4] Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3490_ Inst_RegFile_switch_matrix.N4BEG2 net126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2510_ N2END[1] N4END[0] W6END[0] BD3 Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q Inst_RegFile_switch_matrix.N4BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2441_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q _1032_ _1034_ _1035_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2372_ _0976_ _0975_ Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q Inst_RegFile_switch_matrix.SS4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2639_ Inst_RegFile_32x4.mem\[25\]\[1\] _1184_ _1202_ _0005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput241 net241 WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput252 net252 WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput230 net230 W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2708_ _1186_ Inst_RegFile_32x4.mem\[14\]\[2\] _1226_ _0050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2990_ FrameData[14] FrameStrobe[9] Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1872_ _0510_ _0512_ _0515_ _0516_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1941_ _1296_ B_ADR0 _0582_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3473_ N2MID[5] net118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3542_ Inst_RegFile_switch_matrix.S4BEG2 net178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2286_ _0899_ _0900_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q _0901_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2424_ _0468_ _1019_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q _1020_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2355_ BD0 _0213_ _0497_ _0961_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ _0962_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_67_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_28_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_539 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2140_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q _0772_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2071_ _1311_ B_ADR0 _0705_ _0706_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1855_ _1265_ _0497_ _0499_ _0500_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1924_ Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q _0563_ _0564_ _0565_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2973_ FrameData[29] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1786_ Inst_RegFile_32x4.mem\[19\]\[3\] A_ADR0 _0162_ _0179_ _0434_ _0435_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3456_ Inst_RegFile_switch_matrix.N1BEG0 net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3525_ S2MID[5] net170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2269_ EE4END[0] S1END[2] S1END[0] S2END[0] Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q _0886_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3387_ Inst_RegFile_switch_matrix.E6BEG1 net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2407_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q _1006_ _1007_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2338_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q BD3 _0948_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_4 FrameStrobe[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1640_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _0292_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ _0295_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1571_ _1351_ _0229_ _0230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3310_ _0082_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[29\]\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2123_ N1END[1] N2END[5] NN4END[3] E1END[1] Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q _0756_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3241_ FrameData[9] FrameStrobe[1] Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3172_ FrameData[4] FrameStrobe[3] Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2054_ _1329_ B_ADR0 _0691_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1838_ N2END[3] E2END[3] SS4END[0] W2END[3] Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q
+ Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q _0484_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2956_ FrameData[12] FrameStrobe[10] Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1907_ _0532_ _0548_ _1282_ _0549_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2887_ FrameData[7] FrameStrobe[12] Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_3439_ FrameStrobe[3] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1769_ Inst_RegFile_32x4.mem\[23\]\[2\] A_ADR0 _0162_ _0179_ _0419_ _0420_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3508_ Inst_RegFile_switch_matrix.S1BEG0 net153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 E6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput52 net52 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput41 net41 EE4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput6 net6 E2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput96 net96 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput85 net85 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput63 net63 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput74 net74 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ Inst_RegFile_32x4.mem\[19\]\[0\] _1182_ _1233_ _0076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2810_ _0004_ clknet_4_3_0_UserCLK_regs Inst_RegFile_32x4.mem\[25\]\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2672_ Inst_RegFile_32x4.mem\[30\]\[2\] _1186_ _1214_ _0026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1485_ AD3 BD0 BD2 BD3 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ _0148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3224_ FrameData[24] FrameStrobe[2] Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1623_ W1END[3] AD0 AD1 AD2 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ _0279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1554_ N2MID[4] W2MID[4] S2MID[4] Inst_RegFile_switch_matrix.JS2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q _0213_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
.ends

