* NGSPICE file created from LUT4AB.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VDD VSS W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_2106_ FrameData[3] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2037_ FrameData[30] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1270_ E2MID[6] S2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q _0247_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0985_ _0824_ _0825_ _0827_ _0829_ Inst_LUT4AB_switch_matrix.JN2BEG1 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2655_ W2MID[7] net226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1606_ S2END[1] W2END[1] S4END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0562_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1468_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0432_ _0434_ _0775_ _0435_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1399_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0365_ _0370_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1537_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0500_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2586_ Inst_LUT4AB_switch_matrix.S1BEG3 net157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ Inst_LUT4AB_switch_matrix.E2BEG5 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2371_ FrameData[12] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1253_ _0231_ _0213_ _0176_ _0232_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1322_ S1END[1] S2END[5] S1END[3] W1END[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q _0297_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1184_ _0160_ _0162_ _0165_ _0166_ Inst_LUT4AB_switch_matrix.JN2BEG5 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0968_ F G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q _0814_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2569_ NN4END[6] net146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0899_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q _0747_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput220 net220 W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2638_ Inst_LUT4AB_switch_matrix.W1BEG2 net209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput253 net253 WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput242 net242 WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput231 net231 W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ FrameData[29] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1871_ FrameData[24] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_16_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0000_ clknet_1_1__leaf_UserCLK_regs Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_24_Left_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_69_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1305_ F G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0281_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2285_ FrameData[22] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2354_ FrameData[27] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1236_ _0215_ _0216_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1167_ _0142_ _0143_ _0133_ _0132_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q
+ _0150_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1098_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q _0083_ _0735_ _0086_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ FrameData[31] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1021_ N2END[4] E1END[2] E2END[4] E6END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _0013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1923_ FrameData[12] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1785_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q _0671_ _0689_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1854_ FrameData[7] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2406_ FrameData[15] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_65_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_470 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2337_ FrameData[10] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2268_ FrameData[5] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1219_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_29_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2199_ FrameData[0] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_5 N4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1570_ N1END[0] N2END[0] E1END[0] E2END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q _0530_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2122_ FrameData[19] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2053_ FrameData[14] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1004_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q
+ _0847_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1906_ FrameData[27] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1837_ FrameData[22] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1768_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q _0671_ _0675_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _0637_ _0636_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q Inst_LUT4AB_switch_matrix.EE4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_11_Left_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput75 net75 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput64 net64 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput42 net42 EE4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput20 net20 E2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput31 net31 E6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput7 net7 E2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput86 net86 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput97 net97 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2671_ WW4END[7] net248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1622_ _0575_ _0576_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1484_ _0449_ _0450_ _0451_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1553_ _0513_ _0514_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0515_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2105_ FrameData[2] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2036_ FrameData[29] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0984_ _0713_ _0828_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q _0829_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1536_ _0498_ _0499_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q Inst_LUT4AB_switch_matrix.M_AD
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2654_ W2MID[6] net225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2585_ Inst_LUT4AB_switch_matrix.S1BEG2 net156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1605_ NN4END[1] E2END[1] E1END[3] E6END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0561_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1398_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0363_ _0368_ _0369_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1467_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0367_ _0433_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q
+ _0434_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2019_ FrameData[12] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ FrameData[11] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1321_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q _0296_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1252_ _0757_ _0208_ _0229_ _0206_ _0230_ _0231_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1183_ _0753_ _0163_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q _0166_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0967_ _0709_ _0812_ _0813_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2568_ NN4END[5] net145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2499_ FrameData[20] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0898_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0746_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_58_Left_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput221 net221 W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput210 net210 W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2637_ Inst_LUT4AB_switch_matrix.W1BEG1 net208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1519_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q _0291_ _0483_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q
+ _0484_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput254 net254 WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput243 net243 WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput232 net232 W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Left_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1870_ FrameData[23] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2353_ FrameData[26] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2422_ FrameData[31] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2284_ FrameData[21] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1166_ _0148_ _0149_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1304_ A B D E Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0280_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1235_ NN4END[2] E2END[1] S2END[1] W2END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q _0215_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_50_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1097_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q _0830_ _0084_ _0085_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1999_ FrameData[24] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_7_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1020_ _0719_ _0011_ _0012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1922_ FrameData[11] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1784_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop _0687_ _0688_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1853_ FrameData[6] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2336_ FrameData[9] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2405_ FrameData[14] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2267_ FrameData[4] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1218_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0198_ _0761_ _0199_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2198_ FrameData[31] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1149_ N2END[4] E2END[4] SS4END[2] W2END[4] Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q _0133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_35_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_6 N4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ FrameData[18] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2052_ FrameData[13] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1003_ _0840_ _0841_ _0843_ _0845_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q _0846_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_485 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1905_ FrameData[26] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1767_ _0776_ _0659_ _0673_ _0674_ _0000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1698_ N1END[3] E1END[3] S1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0637_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1836_ FrameData[21] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2319_ FrameData[24] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput87 net87 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput98 net98 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput76 net76 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput54 net54 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput65 net65 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput43 net43 EE4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput21 net21 E2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput32 net32 E6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput8 net8 E2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput10 net10 E2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ S1END[0] S1END[2] S2END[0] W1END[0] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q _0514_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2670_ WW4END[6] net247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1621_ F G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0575_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1483_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0442_ _0445_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0450_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2104_ FrameData[1] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2035_ FrameData[28] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1819_ FrameData[4] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0983_ N2END[2] E1END[0] N4END[2] E2END[2] Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q _0828_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1535_ Inst_LUT4AB_switch_matrix.M_AB _0498_ _0496_ _0499_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2584_ Inst_LUT4AB_switch_matrix.S1BEG1 net155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2653_ W2MID[5] net224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1604_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0556_ _0559_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ _0560_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1466_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0365_ _0433_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1397_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0364_ _0368_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2018_ FrameData[11] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1320_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q _0294_ _0751_ _0295_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1182_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0164_ _0165_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1251_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0209_ _0211_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0230_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_62_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0897_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q _0745_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2636_ Inst_LUT4AB_switch_matrix.W1BEG0 net207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput200 net200 SS4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0966_ A B C E Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ _0812_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2498_ FrameData[19] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2567_ NN4END[4] net138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1449_ _0773_ _0417_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0418_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1518_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q _0289_ _0483_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput222 net222 W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput211 net211 W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput233 net233 W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput244 net244 WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ FrameData[20] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1303_ _0277_ _0278_ _0271_ _0279_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2352_ FrameData[25] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2421_ FrameData[30] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1165_ _0109_ _0110_ _0121_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q
+ _0148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1096_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q _0832_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q
+ _0084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1234_ EE4END[3] WW4END[1] S4END[0] Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q _0214_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_50_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1998_ FrameData[23] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0949_ N2MID[3] E2MID[3] Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q _0796_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2619_ SS4END[4] net190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1921_ FrameData[10] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1852_ FrameData[5] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1783_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q _0658_ _0687_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2266_ FrameData[3] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2335_ FrameData[8] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2404_ FrameData[13] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1148_ NN4END[1] EE4END[1] S4END[1] Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q _0132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1217_ E G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2197_ FrameData[30] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1079_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q _0035_ _0067_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_7 N4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ FrameData[17] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2051_ FrameData[12] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1002_ _0840_ _0841_ _0843_ _0845_ Inst_LUT4AB_switch_matrix.JS2BEG1 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_19_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ FrameData[25] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ FrameData[20] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1766_ Inst_LH_LUT4c_frame_config_dffesr.c_reset_value _0672_ _0659_ _0674_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1697_ H _0018_ _0142_ _0158_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0636_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2249_ FrameData[18] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2318_ FrameData[23] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_23_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput88 net88 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput55 net55 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput66 net66 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput99 net99 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput33 net33 E6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput77 net77 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput44 net44 EE4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput22 net22 E6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput9 net9 E2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput11 net11 E2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1482_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0441_ _0444_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0449_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1551_ N1END[0] NN4END[0] E1END[0] E2END[0] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q _0513_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1620_ B D C E Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ _0574_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2103_ FrameData[0] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ FrameData[27] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1818_ FrameData[3] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1749_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0656_ _0657_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0826_ _0827_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2652_ W2MID[4] net223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1534_ C D _0497_ _0498_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1465_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0363_ _0431_ _0432_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2583_ Inst_LUT4AB_switch_matrix.S1BEG0 net154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0558_ _0559_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1396_ _0366_ _0367_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2017_ FrameData[10] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1250_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0193_ _0229_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1181_ S1END[2] W1END[0] S2END[6] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q _0164_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2635_ clknet_1_0__leaf_UserCLK net206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0896_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q _0744_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput223 net223 W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput201 net201 SS4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput212 net212 W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput234 net234 W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0965_ _0795_ _0800_ _0810_ _0809_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q
+ _0811_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2566_ Inst_LUT4AB_switch_matrix.N4BEG3 net128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2497_ FrameData[18] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1448_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0417_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _0481_ _0482_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput245 net245 WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1379_ _0317_ _0323_ _0325_ _0351_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_53_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ FrameData[29] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2282_ FrameData[19] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1233_ _0756_ _0208_ _0210_ _0212_ _0213_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_49_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1302_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0153_ _0272_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0278_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2351_ FrameData[24] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1164_ _0122_ _0144_ _0147_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1095_ _0820_ _0821_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q _0083_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_50_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1997_ FrameData[22] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0948_ E2MID[2] S2MID[2] W2MID[2] Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q _0795_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2549_ N2MID[6] net120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2618_ Inst_LUT4AB_switch_matrix.S4BEG3 net180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0879_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0727_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1920_ FrameData[9] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1851_ FrameData[4] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1782_ _0682_ _0685_ _0686_ _0683_ _0003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2403_ FrameData[12] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2265_ FrameData[2] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1216_ _0760_ _0196_ _0197_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2196_ FrameData[29] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2334_ FrameData[7] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_35_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1147_ _0125_ _0127_ _0129_ _0131_ Inst_LUT4AB_switch_matrix.JS2BEG2 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1078_ _0736_ _0047_ _0065_ _0066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_8 N4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ FrameData[11] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1001_ _0723_ _0844_ _0724_ _0845_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1765_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q _0671_ _0460_ _0673_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1903_ FrameData[24] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1834_ FrameData[19] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1696_ _0635_ Inst_LUT4AB_switch_matrix.EE4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2179_ FrameData[12] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2317_ FrameData[22] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2248_ FrameData[17] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput23 net23 E6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput34 net34 EE4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 E2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput89 net89 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput67 net67 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput78 net78 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput56 net56 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput45 net45 EE4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1550_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0509_ _0511_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ _0512_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1481_ _0419_ _0420_ _0410_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q
+ _0448_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2102_ FrameData[31] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2033_ FrameData[26] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1817_ FrameData[2] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_15_Left_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1748_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q Inst_LUT4AB_switch_matrix.JS2BEG2
+ _0655_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q _0656_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1679_ _0620_ _0621_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q _0622_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0981_ E6END[0] S2END[2] W2END[2] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q _0826_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2582_ Inst_LUT4AB_switch_matrix.NN4BEG3 net144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2651_ W2MID[3] net222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1602_ _0557_ _0558_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1533_ _0465_ _0496_ _0783_ _0497_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1464_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0364_ _0431_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1395_ N2END[7] E2END[7] S2END[7] WW4END[0] Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q _0366_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ FrameData[9] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1180_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0163_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0964_ NN4END[0] S2END[2] E2END[2] W2END[2] Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q _0810_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2565_ Inst_LUT4AB_switch_matrix.N4BEG2 net127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0895_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0743_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1516_ _0479_ _0480_ _0472_ _0481_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2634_ Inst_LUT4AB_switch_matrix.SS4BEG3 net196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput246 net246 WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput202 net202 SS4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput213 net213 W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput224 net224 W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput235 net235 W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2496_ FrameData[17] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1378_ Inst_LF_LUT4c_frame_config_dffesr.c_out_mux _0349_ _0350_ F VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1447_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0415_ _0416_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_48_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2281_ FrameData[18] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_63_Left_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1232_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0209_ _0211_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0212_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1301_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0151_ _0274_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ _0277_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2350_ FrameData[23] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1163_ _0122_ _0144_ _0146_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1094_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0076_ _0080_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0071_ _0082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1996_ FrameData[21] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_15_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0947_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q _0792_ _0794_ _0788_ _0790_ Inst_LUT4AB_switch_matrix.E2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2548_ N2MID[5] net119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2617_ Inst_LUT4AB_switch_matrix.S4BEG2 net179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0878_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0726_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2479_ FrameData[0] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1781_ Inst_LC_LUT4c_frame_config_dffesr.c_reset_value _0684_ _0686_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1850_ FrameData[3] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2402_ FrameData[11] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ FrameData[6] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1215_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2195_ FrameData[28] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1146_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0130_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
+ _0131_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2264_ FrameData[1] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_35_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1077_ _0736_ _0045_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q _0065_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ FrameData[4] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_26_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_9 N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1000_ S4END[2] SS4END[2] W2END[2] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _0844_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1902_ FrameData[23] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_42_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q _0671_ _0672_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1833_ FrameData[18] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2316_ FrameData[21] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1695_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q _0634_ _0633_ _0635_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_48_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2178_ FrameData[11] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1129_ N1END[1] N4END[3] N2END[3] E2END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q _0115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2247_ FrameData[16] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_23_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput57 net57 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput24 net24 E6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput35 net35 EE4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput46 net46 EE4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput13 net13 E2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput79 net79 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput68 net68 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1480_ _0443_ _0446_ _0447_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2101_ FrameData[30] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2032_ FrameData[25] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1678_ _0018_ _0142_ _0204_ _0398_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0621_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1747_ _0284_ _0288_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0655_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1816_ FrameData[1] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_469 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0980_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0822_ _0714_ _0825_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2581_ Inst_LUT4AB_switch_matrix.NN4BEG2 net143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1532_ Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_switch_matrix.JS2BEG5
+ Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q
+ _0496_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2650_ W2MID[2] net221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1601_ F G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q _0557_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1463_ _0317_ _0323_ _0386_ _0400_ _0325_ _0430_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1394_ N4END[3] EE4END[0] S4END[3] Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q _0365_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2015_ FrameData[8] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_56_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0894_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0742_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0963_ EE4END[2] S4END[2] W2END[7] Inst_LUT4AB_switch_matrix.E2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q _0809_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2495_ FrameData[16] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2564_ Inst_LUT4AB_switch_matrix.N4BEG1 net126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1515_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0147_ _0473_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0480_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2633_ Inst_LUT4AB_switch_matrix.SS4BEG2 net195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput225 net225 W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput214 net214 W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput203 net203 SS4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput247 net247 WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput236 net236 W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1446_ S1END[1] S1END[3] S2END[7] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0415_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1377_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ _0350_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2280_ FrameData[17] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1162_ _0122_ _0144_ _0145_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1231_ _0193_ _0206_ _0211_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1300_ _0273_ _0275_ _0276_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1093_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0077_ _0079_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1995_ FrameData[20] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0877_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q _0725_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2616_ Inst_LUT4AB_switch_matrix.S4BEG1 net178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0946_ _0715_ _0793_ _0794_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2478_ Inst_LUT4AB_switch_matrix.EE4BEG3 net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2547_ N2MID[4] net118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1429_ E2MID[4] W2MID[4] S2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q _0398_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q _0671_ _0316_ _0685_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2401_ FrameData[10] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2332_ FrameData[5] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_65_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1214_ N2END[5] E2END[5] SS4END[1] W2END[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q _0195_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1145_ S2END[3] W2END[3] S4END[3] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q _0130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2194_ FrameData[27] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2263_ FrameData[0] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1076_ Inst_LA_LUT4c_frame_config_dffesr.c_out_mux _0063_ _0064_ A VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1978_ FrameData[3] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0929_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0777_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1901_ FrameData[22] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1832_ FrameData[17] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1694_ N1END[0] S1END[0] E1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ _0634_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1763_ _0661_ _0664_ _0670_ _0671_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2315_ FrameData[20] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2246_ FrameData[15] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2177_ FrameData[10] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1128_ _0744_ _0113_ _0745_ _0114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1059_ _0045_ _0046_ _0036_ _0035_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q
+ _0048_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_31_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput69 net69 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput58 net58 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput25 net25 E6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput47 net47 EE4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput36 net36 EE4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput14 net14 E2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2100_ FrameData[29] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2031_ FrameData[24] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1815_ FrameData[0] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1677_ G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q _0620_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1746_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0119_ _0653_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ _0654_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2229_ FrameData[30] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2580_ Inst_LUT4AB_switch_matrix.NN4BEG1 net142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1462_ _0429_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ G VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1531_ _0495_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ D VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1600_ B D C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ _0556_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1393_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q _0364_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2014_ FrameData[7] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ E _0173_ Inst_LUT4AB_switch_matrix.JN2BEG0 _0194_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q Inst_LUT4AB_switch_matrix.E1BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_56_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0893_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q _0741_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2632_ Inst_LUT4AB_switch_matrix.SS4BEG1 net194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0962_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q _0806_ _0808_ _0802_ _0804_ Inst_LUT4AB_switch_matrix.E2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_9_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2494_ FrameData[15] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2563_ Inst_LUT4AB_switch_matrix.N4BEG0 net125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1445_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0413_ _0412_ _0414_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1514_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0146_ _0475_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ _0479_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput215 net215 W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput226 net226 W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput204 net204 SS4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput248 net248 WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput237 net237 W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1376_ _0340_ _0348_ _0349_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_61_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1230_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0193_ _0207_ _0210_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1161_ _0142_ _0143_ _0133_ _0132_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q
+ _0144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1092_ _0072_ _0074_ _0080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1994_ FrameData[19] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2615_ Inst_LUT4AB_switch_matrix.S4BEG0 net177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0876_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q _0724_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0945_ E6END[0] S2END[4] W2END[4] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _0793_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1428_ _0391_ _0393_ _0396_ _0397_ Inst_LUT4AB_switch_matrix.JS2BEG6 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2477_ Inst_LUT4AB_switch_matrix.EE4BEG2 net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2546_ N2MID[3] net117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1359_ _0319_ _0331_ _0332_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ FrameData[9] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2331_ FrameData[4] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2262_ FrameData[31] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1213_ N4END[1] SS4END[1] W2END[4] Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q _0194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1144_ _0748_ _0128_ _0129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2193_ FrameData[26] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1075_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ _0064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1977_ FrameData[2] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0928_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop _0776_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0859_ S2MID[6] _0707_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2529_ FrameStrobe[18] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ FrameData[21] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1831_ FrameData[16] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1693_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q _0632_ _0630_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ _0633_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1762_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q _0666_ _0669_ _0670_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_69_Left_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2314_ FrameData[19] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2245_ FrameData[14] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2176_ FrameData[9] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1127_ A B D E Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ _0113_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1058_ _0046_ _0047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput59 net59 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput37 net37 EE4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput26 net26 E6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput48 net48 EE4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 E2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ FrameData[23] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q Inst_LUT4AB_switch_matrix.JN2BEG2
+ _0653_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1814_ FrameData[31] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1676_ _0617_ _0618_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q _0619_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2159_ FrameData[24] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2228_ FrameData[29] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1461_ _0428_ _0425_ _0421_ _0429_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1392_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q _0360_ _0362_ _0363_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1530_ _0478_ _0482_ _0486_ _0494_ _0495_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2013_ FrameData[6] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1728_ F Inst_LUT4AB_switch_matrix.JN2BEG1 _0385_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q Inst_LUT4AB_switch_matrix.E1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1659_ _0605_ _0604_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q Inst_LUT4AB_switch_matrix.SS4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0961_ _0717_ _0807_ _0808_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ N4END[15] net124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0892_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0740_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput205 net205 SS4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2631_ Inst_LUT4AB_switch_matrix.SS4BEG0 net193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput216 net216 W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2493_ FrameData[14] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1444_ E H F Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q _0413_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1375_ _0336_ _0342_ _0345_ _0347_ _0348_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1513_ _0472_ _0477_ _0478_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput227 net227 W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput249 net249 WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput238 net238 W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1160_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q _0143_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Left_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1091_ _0073_ _0075_ _0079_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_41_Left_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1993_ FrameData[18] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0944_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _0791_ _0792_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2614_ S4END[15] net176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2545_ N2MID[2] net116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0875_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _0723_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1427_ _0771_ _0394_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q _0397_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2476_ Inst_LUT4AB_switch_matrix.EE4BEG1 net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1358_ _0326_ _0330_ _0331_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_50_Left_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1289_ NN4END[3] E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q _0265_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_21_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1212_ _0187_ _0192_ _0178_ _0177_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q
+ _0193_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2330_ FrameData[3] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2261_ FrameData[30] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2192_ FrameData[25] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1143_ NN4END[3] E1END[1] E2END[3] E6END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1074_ _0048_ _0052_ _0057_ _0062_ _0063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0927_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0775_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1976_ FrameData[1] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2528_ FrameStrobe[17] net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2459_ E6END[10] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q Inst_LUT4AB_switch_matrix.JN2BEG1
+ _0668_ _0669_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1830_ FrameData[15] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2313_ FrameData[18] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1692_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q C _0631_ _0632_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2244_ FrameData[13] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1126_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q _0111_ _0112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2175_ FrameData[8] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1057_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q _0046_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1959_ FrameData[16] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput38 net38 EE4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput49 net49 EE4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput27 net27 E6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput16 net16 E2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1813_ FrameData[30] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1744_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0227_ _0651_ _0652_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1675_ C D E F Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0618_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ FrameData[23] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2089_ FrameData[18] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2227_ FrameData[28] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1109_ _0096_ _0097_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1460_ _0427_ _0426_ _0373_ _0428_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1391_ _0707_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
+ _0361_ _0362_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2012_ FrameData[5] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ G _0020_ Inst_LUT4AB_switch_matrix.JN2BEG2 _0830_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q Inst_LUT4AB_switch_matrix.E1BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1658_ N1END[1] E1END[1] W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0605_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1589_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0546_ _0547_ _0545_ Inst_LUT4AB_switch_matrix.M_AH
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_26_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0960_ E6END[0] S2END[2] W2END[2] WW4END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _0807_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput206 net206 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2561_ N4END[14] net123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2492_ FrameData[13] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1512_ _0474_ _0476_ _0477_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0891_ S2END[6] _0739_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2630_ SS4END[15] net192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput239 net239 WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput217 net217 W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput228 net228 W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1443_ _0773_ _0411_ _0412_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1374_ _0329_ _0343_ _0346_ _0323_ _0347_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1090_ _0072_ _0074_ _0078_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1992_ FrameData[17] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0874_ E6END[1] _0722_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0943_ N1END[2] N2END[4] N4END[0] E2END[4] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _0791_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2613_ S4END[14] net175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2475_ Inst_LUT4AB_switch_matrix.EE4BEG0 net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2544_ N2MID[1] net115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1426_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0395_ _0396_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1357_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0327_ _0329_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0330_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1288_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q _0739_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q
+ _0263_ _0264_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1211_ _0191_ _0192_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1142_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0126_ _0749_ _0127_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2191_ FrameData[24] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2260_ FrameData[29] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1073_ _0048_ _0061_ _0062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_23_Left_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0926_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0774_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1975_ FrameData[0] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2527_ FrameStrobe[16] net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1409_ S1END[1] S1END[3] S2END[7] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0380_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2458_ E6END[9] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2389_ FrameData[30] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1691_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0191_ _0631_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1760_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0667_ _0668_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2312_ FrameData[17] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2243_ FrameData[12] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1125_ F G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2174_ FrameData[7] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1056_ N2MID[0] E2MID[0] S2MID[0] Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q _0045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput39 net39 EE4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1958_ FrameData[15] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput28 net28 E6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0909_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0757_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1889_ FrameData[10] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput17 net17 E2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1674_ E1END[2] W1END[2] A B Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0617_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1812_ FrameData[29] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1743_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0301_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ _0651_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2226_ FrameData[27] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2157_ FrameData[22] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1039_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0029_ _0729_ _0030_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2088_ FrameData[17] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1108_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0076_ _0077_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0079_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0096_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai222_1
XPHY_EDGE_ROW_10_Left_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q Inst_LUT4AB_switch_matrix.JN2BEG6
+ _0361_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2011_ FrameData[4] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_462 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1588_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0542_ _0547_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1657_ E _0204_ _0398_ _0036_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0604_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1726_ E Inst_LUT4AB_switch_matrix.E2BEG3 _0301_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q Inst_LUT4AB_switch_matrix.S1BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2209_ FrameData[10] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0890_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0738_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2491_ FrameData[12] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2560_ N4END[13] net137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1442_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0411_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1511_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0147_ _0475_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0476_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput207 net207 W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput218 net218 W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput229 net229 W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1373_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0319_ _0346_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1709_ H _0018_ _0142_ _0178_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0644_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2612_ S4END[13] net189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1991_ FrameData[16] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0873_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q _0721_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0942_ _0715_ _0789_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q _0790_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1425_ S1END[3] W1END[1] S2END[7] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0395_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2474_ EE4END[15] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2543_ N2MID[0] net114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1356_ _0328_ _0329_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1287_ W2END[6] Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q _0263_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1141_ F G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1210_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q _0190_ _0189_ _0191_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1072_ _0023_ _0060_ _0061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2190_ FrameData[23] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ FrameData[31] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0925_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0773_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2526_ FrameStrobe[15] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1408_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q _0376_ _0770_ _0379_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2457_ E6END[8] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2388_ FrameData[29] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1339_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0151_ _0272_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0313_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0385_ _0629_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ _0630_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2311_ FrameData[16] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2242_ FrameData[11] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_29_Left_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1124_ N2MID[3] E2MID[3] S2MID[3] W2MID[3] Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q _0110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2173_ FrameData[6] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1055_ _0038_ _0040_ _0043_ _0044_ Inst_LUT4AB_switch_matrix.JW2BEG3 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1957_ FrameData[14] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput29 net29 E6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2509_ FrameData[30] net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1888_ FrameData[9] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0908_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0756_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput18 net18 E2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1811_ FrameData[28] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1673_ _0616_ Inst_LUT4AB_switch_matrix.SS4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1742_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0047_ _0649_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ _0650_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2225_ FrameData[26] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2156_ FrameData[21] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1038_ F G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q _0029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2087_ FrameData[16] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1107_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0079_ _0080_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0071_ _0095_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ FrameData[3] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1725_ F _0173_ Inst_LUT4AB_switch_matrix.E2BEG0 _0194_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q Inst_LUT4AB_switch_matrix.S1BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1587_ _0783_ _0543_ _0546_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1656_ _0603_ _0602_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q Inst_LUT4AB_switch_matrix.WW4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2208_ FrameData[9] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2139_ FrameData[4] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2490_ FrameData[11] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1510_ _0123_ _0144_ _0475_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput219 net219 W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput208 net208 W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1441_ _0409_ _0410_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1372_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0319_ _0327_ _0344_
+ _0345_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1708_ _0643_ _0642_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q Inst_LUT4AB_switch_matrix.NN4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1639_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q _0585_ _0587_ _0589_ _0591_ Inst_LUT4AB_switch_matrix.W6BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_64_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1990_ FrameData[15] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_15_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0941_ F G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _0789_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2611_ S4END[12] net188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2542_ Inst_LUT4AB_switch_matrix.JN2BEG7 net113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0872_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q _0720_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1424_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q _0394_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1355_ _0321_ _0322_ _0328_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2473_ EE4END[14] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1286_ E2END[3] WW4END[2] SS4END[3] Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q _0262_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1140_ _0748_ _0124_ _0125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1071_ _0059_ _0058_ _0811_ _0060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0924_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q _0772_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1973_ FrameData[30] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2525_ FrameStrobe[14] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1407_ _0769_ _0377_ _0378_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2456_ E6END[7] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1338_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0153_ _0274_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ _0312_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ FrameData[28] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1269_ _0241_ _0242_ _0244_ _0246_ Inst_LUT4AB_switch_matrix.JN2BEG4 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2310_ FrameData[15] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2172_ FrameData[5] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2241_ FrameData[10] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1123_ N2MID[2] W2MID[2] E2MID[2] Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q _0109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1054_ _0726_ _0041_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0044_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1956_ FrameData[13] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0907_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux _0755_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1887_ FrameData[8] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_21_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2508_ FrameData[29] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput19 net19 E2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2439_ Inst_LUT4AB_switch_matrix.E2BEG4 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1810_ FrameData[27] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1741_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0419_ _0649_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1672_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q _0615_ _0614_ _0616_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2155_ FrameData[20] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1106_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0076_ _0077_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2224_ FrameData[25] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2086_ FrameData[15] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1037_ _0728_ _0027_ _0028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1939_ FrameData[28] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_48_Left_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Left_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_66_Left_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1724_ G Inst_LUT4AB_switch_matrix.E2BEG1 _0385_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q Inst_LUT4AB_switch_matrix.S1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1586_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0544_ _0545_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1655_ N1END[2] S1END[2] W1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0603_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2138_ FrameData[3] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2069_ FrameData[30] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2207_ FrameData[8] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1371_ _0766_ _0319_ _0344_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput209 net209 W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1440_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q _0406_ _0408_ _0409_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_390 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1707_ N1END[0] W1END[0] E1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ _0643_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1638_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0590_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ _0591_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1569_ S1END[0] S1END[2] SS4END[0] WW4END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q _0529_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0940_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _0787_ _0788_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_15_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2610_ S4END[11] net187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2541_ Inst_LUT4AB_switch_matrix.JN2BEG6 net112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2472_ EE4END[13] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0871_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _0719_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1423_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0392_ _0772_ _0393_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1354_ _0321_ _0322_ _0327_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1285_ _0255_ _0257_ _0260_ _0261_ Inst_LUT4AB_switch_matrix.JN2BEG2 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_66_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_485 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1070_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0834_ _0059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0923_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0771_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1972_ FrameData[29] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2524_ FrameStrobe[13] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2455_ E6END[6] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1406_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0377_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1268_ _0737_ _0245_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0246_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1337_ _0271_ _0310_ _0311_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2386_ FrameData[27] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_64_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1199_ _0758_ _0180_ _0181_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1122_ _0102_ _0104_ _0106_ _0108_ Inst_LUT4AB_switch_matrix.E2BEG4 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2171_ FrameData[4] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_27_Left_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2240_ FrameData[9] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1053_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0042_ _0043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1955_ FrameData[12] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1886_ FrameData[7] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0906_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q _0754_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2507_ FrameData[28] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2438_ Inst_LUT4AB_switch_matrix.E2BEG3 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2369_ FrameData[10] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1740_ _0444_ _0648_ net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ N1END[2] W1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ _0615_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2154_ FrameData[19] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ FrameData[24] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1105_ _0081_ _0082_ _0092_ _0093_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2085_ FrameData[14] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1036_ A D C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ _0027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1938_ FrameData[27] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1869_ FrameData[22] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1654_ G _0800_ _0110_ _0389_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0602_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1723_ H _0020_ Inst_LUT4AB_switch_matrix.E2BEG2 _0830_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q Inst_LUT4AB_switch_matrix.S1BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1585_ _0499_ _0543_ _0538_ _0544_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2206_ FrameData[7] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2137_ FrameData[2] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1019_ S2END[4] W2END[4] S4END[0] WW4END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _0011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2068_ FrameData[29] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_14_Left_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0319_ _0343_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1706_ C _0192_ _0385_ _0121_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ _0642_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1637_ G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q _0590_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_69_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
+ _0465_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1568_ _0779_ _0525_ _0780_ _0528_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0870_ E2MID[4] _0718_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1422_ E H F Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0392_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2471_ EE4END[12] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2540_ Inst_LUT4AB_switch_matrix.JN2BEG5 net111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1353_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0323_ _0324_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0326_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1284_ _0740_ _0258_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q _0261_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0999_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _0842_ _0843_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2669_ WW4END[5] net246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0922_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q _0770_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1971_ FrameData[28] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2523_ FrameStrobe[12] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2454_ E6END[5] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1405_ E H F Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q _0376_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2385_ FrameData[26] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_68_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1267_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0245_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1198_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1336_ _0308_ _0309_ _0310_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1121_ _0742_ _0107_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0108_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2170_ FrameData[3] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1052_ S2END[4] W2END[4] S4END[0] WW4END[2] Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1954_ FrameData[11] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0905_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0753_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1885_ FrameData[6] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2506_ FrameData[27] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2437_ Inst_LUT4AB_switch_matrix.E2BEG2 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2368_ FrameData[9] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1319_ F G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q _0294_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_39_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2299_ FrameData[4] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_50 N4END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput190 net190 SS4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_45_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q _0613_ _0611_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
+ _0614_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2222_ FrameData[23] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2153_ FrameData[18] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1035_ _0835_ _0025_ _0811_ _0026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2084_ FrameData[13] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1104_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0079_ _0091_ _0070_
+ _0092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1937_ FrameData[26] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1799_ Inst_LF_LUT4c_frame_config_dffesr.c_reset_value _0699_ _0701_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1868_ FrameData[21] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1584_ Inst_LUT4AB_switch_matrix.M_EF _0542_ _0539_ _0543_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1653_ _0601_ _0600_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q Inst_LUT4AB_switch_matrix.WW4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1722_ E6END[1] S4END[1] S2END[2] A Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ Inst_LUT4AB_switch_matrix.S4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2205_ FrameData[6] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_64_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2136_ FrameData[1] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1018_ _0719_ _0858_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q _0010_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2067_ FrameData[28] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1705_ _0641_ _0640_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q Inst_LUT4AB_switch_matrix.NN4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_61_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1567_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0526_ _0527_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1636_ _0786_ _0588_ _0589_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _0462_ _0463_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q _0464_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2119_ FrameData[16] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1421_ _0771_ _0390_ _0391_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2470_ EE4END[11] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_462 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1352_ _0324_ _0325_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1283_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0259_ _0260_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2668_ WW4END[4] net239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0998_ NN4END[2] EE4END[2] E1END[0] E6END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _0842_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2599_ S2MID[4] net170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1619_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q _0571_ _0573_ _0567_ _0569_ Inst_LUT4AB_switch_matrix.E2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_67_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0921_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q _0769_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ FrameData[27] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2522_ FrameStrobe[11] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ E6END[4] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1404_ N2END[3] SS4END[0] E2END[3] W2END[3] Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q _0375_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2384_ FrameData[25] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1335_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0153_ _0272_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0309_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1266_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q _0243_ _0244_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1197_ E G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1120_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0107_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_48_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1051_ N1END[2] E2END[4] N2END[4] E6END[0] Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1953_ FrameData[10] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1884_ FrameData[5] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0904_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q _0752_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_31_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2505_ FrameData[26] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1318_ _0750_ _0292_ _0293_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2298_ FrameData[3] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2367_ FrameData[8] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2436_ Inst_LUT4AB_switch_matrix.E2BEG1 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1249_ _0225_ _0226_ _0215_ _0214_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q
+ _0228_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_51 NN4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_40 SS4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput191 net191 SS4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput180 net180 S4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2152_ FrameData[17] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2221_ FrameData[22] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1034_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0834_ _0025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2083_ FrameData[12] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1103_ _0090_ _0091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1936_ FrameData[25] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1867_ FrameData[20] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1798_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q _0671_ _0348_ _0340_ _0700_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2419_ FrameData[28] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_4_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Left_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1721_ E6END[0] S4END[2] S2END[3] B Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ Inst_LUT4AB_switch_matrix.S4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1583_ H G _0541_ _0542_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1652_ N1END[3] S1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0601_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_44_Left_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Left_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2135_ FrameData[0] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2204_ FrameData[5] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_64_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1017_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _0008_ _0009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2066_ FrameData[27] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_62_Left_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1919_ FrameData[8] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1704_ N1END[1] E1END[1] W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ _0641_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_69_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ _0463_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1566_ E G F Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q _0526_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1635_ _0018_ _0142_ _0204_ _0398_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0588_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2118_ FrameData[15] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2049_ FrameData[10] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_1_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0390_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1351_ _0320_ _0322_ _0324_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1282_ E6END[1] S2END[3] W2END[3] WW4END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0259_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0997_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _0838_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q
+ _0841_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1618_ _0785_ _0572_ _0573_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2667_ Inst_LUT4AB_switch_matrix.W6BEG1 net229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1549_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0510_ _0511_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2598_ S2MID[3] net169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0920_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux _0768_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2521_ FrameStrobe[10] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1265_ S1END[1] S2END[5] W1END[1] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0243_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2452_ E6END[3] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1403_ N4END[2] W2END[2] SS4END[2] Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q _0374_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1334_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0151_ _0274_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0308_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2383_ FrameData[24] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ N2END[3] S2END[3] E2END[3] WW4END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q _0178_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1050_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0039_ _0727_ _0040_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0903_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q _0751_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1952_ FrameData[9] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1883_ FrameData[4] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2504_ FrameData[25] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2435_ Inst_LUT4AB_switch_matrix.E2BEG0 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1317_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0292_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_39_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2297_ FrameData[2] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2366_ FrameData[7] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_2_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1248_ _0226_ _0227_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1179_ _0753_ _0161_ _0754_ _0162_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_30 SS4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_52 net239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_41 W2MID[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput192 net192 SS4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput181 net181 S4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput170 net170 S2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2151_ FrameData[16] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2220_ FrameData[21] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1102_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0076_ _0077_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0080_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0090_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_2082_ FrameData[11] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1033_ _0850_ _0854_ _0019_ _0021_ _0024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1797_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q _0671_ _0699_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1935_ FrameData[24] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1866_ FrameData[19] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2418_ FrameData[27] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_37_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2349_ FrameData[22] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ H _0018_ _0142_ _0195_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0600_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_41_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1720_ S2END[0] W6END[1] S4END[3] C Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ Inst_LUT4AB_switch_matrix.S4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1582_ _0783_ _0539_ _0540_ _0541_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2134_ FrameData[31] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2203_ FrameData[4] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2065_ FrameData[26] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_21_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1016_ A B C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ _0008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1918_ FrameData[7] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_out_mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1849_ FrameData[2] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1703_ E _0204_ _0398_ _0810_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ _0640_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1634_ _0786_ _0586_ _0587_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2683_ Inst_LUT4AB_switch_matrix.WW4BEG3 net245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1496_ Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ _0462_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1565_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0525_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_18_Left_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2117_ FrameData[14] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_52_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ FrameData[9] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_1_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1350_ _0320_ _0322_ _0323_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1281_ N2END[3] N4END[3] E1END[1] E2END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0258_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_66_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0996_ _0723_ _0839_ _0840_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2597_ S2MID[2] net168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1617_ E6END[1] W2END[1] S2END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0572_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2666_ Inst_LUT4AB_switch_matrix.W6BEG0 net228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1479_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0444_ _0445_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0446_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1548_ E G F Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q _0510_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2520_ FrameStrobe[9] net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2451_ E6END[2] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1402_ _0768_ _0351_ _0372_ _0373_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1264_ _0737_ _0239_ _0738_ _0242_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1333_ _0271_ _0276_ _0279_ _0306_ _0307_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2382_ FrameData[23] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1195_ NN4END[2] S4END[2] E2END[2] Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q _0177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_34_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0979_ _0713_ _0823_ _0824_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2649_ W2MID[1] net220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0902_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q _0750_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1951_ FrameData[8] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1882_ FrameData[3] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2503_ FrameData[24] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2434_ Inst_LUT4AB_switch_matrix.E1BEG3 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2365_ FrameData[6] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1178_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0161_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_39_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2296_ FrameData[1] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1316_ _0290_ _0291_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1247_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q _0226_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_20 NN4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_31 SS4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_42 W2MID[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_53 net250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput193 net193 SS4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput182 net182 S4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput160 net160 S2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput171 net171 S2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_6_Left_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2081_ FrameData[10] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1032_ _0855_ _0022_ _0023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1101_ _0735_ _0087_ _0088_ _0085_ _0086_ _0089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2150_ FrameData[15] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1934_ FrameData[23] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1796_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop _0697_ _0698_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1865_ FrameData[18] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2348_ FrameData[21] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2417_ FrameData[26] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2279_ FrameData[16] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1581_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0466_ _0540_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1650_ _0599_ _0598_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q Inst_LUT4AB_switch_matrix.WW4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2202_ FrameData[3] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2133_ FrameData[30] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1015_ F G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _0858_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ FrameData[25] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1917_ FrameData[6] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1848_ FrameData[1] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1779_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q _0671_ _0684_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1702_ _0639_ _0638_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q Inst_LUT4AB_switch_matrix.EE4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1564_ _0519_ _0520_ _0522_ _0524_ Inst_LUT4AB_switch_matrix.JN2BEG7 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1633_ C D E F Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0586_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2682_ Inst_LUT4AB_switch_matrix.WW4BEG2 net244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1495_ _0776_ Inst_LH_LUT4c_frame_config_dffesr.c_out_mux _0461_ H VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_52_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2116_ FrameData[13] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2047_ FrameData[8] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_1_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1280_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0256_ _0741_ _0257_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0995_ F G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _0839_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1547_ _0508_ _0509_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2665_ W6END[11] net238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2596_ S2MID[1] net167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1616_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q _0570_ _0571_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1478_ _0437_ _0439_ _0445_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_59_Left_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1401_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q _0369_ _0371_ _0768_ _0372_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2450_ E2MID[7] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2381_ FrameData[22] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1194_ _0755_ _0145_ _0156_ _0175_ _0176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1263_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q _0240_ _0241_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1332_ _0305_ _0306_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0978_ A D C E Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ _0823_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2579_ Inst_LUT4AB_switch_matrix.NN4BEG0 net141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2648_ W2MID[0] net219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1950_ FrameData[7] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2502_ FrameData[23] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1881_ FrameData[2] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0901_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q _0749_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2364_ FrameData[5] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2433_ Inst_LUT4AB_switch_matrix.E1BEG2 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1315_ N2END[0] S2END[0] EE4END[1] W2END[0] Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q _0290_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_22_Left_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1177_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0159_ _0160_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_464 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ FrameData[0] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1246_ E2MID[0] S2MID[0] W2MID[0] Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q _0225_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_21 NN4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_10 N4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_32 SS4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_43 net232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput150 net150 NN4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput161 net161 S2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput194 net194 SS4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput183 net183 S4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput172 net172 S2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1031_ _0019_ _0021_ _0022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1100_ _0811_ _0024_ Ci _0088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2080_ FrameData[9] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1933_ FrameData[22] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1795_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q _0658_ _0697_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1864_ FrameData[17] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2347_ FrameData[20] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2278_ FrameData[15] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2416_ FrameData[25] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1229_ _0193_ _0207_ _0209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0538_ _0496_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0539_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2132_ FrameData[29] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2201_ FrameData[2] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1014_ _0718_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
+ _0856_ _0857_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_19_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2063_ FrameData[24] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1916_ FrameData[5] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1847_ FrameData[0] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_30_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop _0682_ _0683_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_31_Left_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_40_Left_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1701_ N1END[2] S1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ _0639_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2681_ Inst_LUT4AB_switch_matrix.WW4BEG1 net243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1494_ Inst_LH_LUT4c_frame_config_dffesr.c_out_mux _0460_ _0461_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1563_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0523_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ _0524_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1632_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0584_ _0585_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2115_ FrameData[12] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2046_ FrameData[7] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0994_ A D C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ _0838_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_14_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2664_ W6END[10] net237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1477_ _0438_ _0440_ _0444_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2595_ S2MID[0] net166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1615_ N1END[3] N2END[1] N4END[1] EE4END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0570_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1546_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0508_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2029_ FrameData[22] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_11_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2380_ FrameData[21] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1400_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0367_ _0370_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q
+ _0371_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1331_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q _0304_ _0303_ _0305_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1262_ F G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0240_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1193_ _0755_ _0174_ _0175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2647_ Inst_LUT4AB_switch_matrix.JW2BEG7 net218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0977_ F G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q _0822_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2578_ NN4END[15] net140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1529_ _0486_ _0489_ _0493_ _0494_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ FrameData[1] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_out_mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0900_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0748_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ FrameData[22] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2363_ FrameData[4] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1314_ N4END[0] W6END[0] SS4END[0] Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q _0289_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2294_ FrameData[31] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2432_ Inst_LUT4AB_switch_matrix.E1BEG1 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1176_ E G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0159_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1245_ _0219_ _0220_ _0223_ _0224_ Inst_LUT4AB_switch_matrix.JW2BEG5 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_11 N4END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_22 NN4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_33 SS4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_44 net233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput151 net151 NN4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput140 net140 NN4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput184 net184 S4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput173 net173 S2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput162 net162 S2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput195 net195 SS4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1030_ _0721_ _0020_ _0725_ _0021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1932_ FrameData[21] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1863_ FrameData[16] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1794_ _0692_ _0695_ _0696_ _0693_ _0005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2415_ FrameData[24] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2346_ FrameData[19] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1228_ _0193_ _0206_ _0208_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2277_ FrameData[14] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1159_ N2MID[4] E2MID[4] S2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q _0142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2131_ FrameData[28] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2200_ FrameData[1] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2062_ FrameData[23] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1013_ N2MID[4] Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q _0856_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1915_ FrameData[4] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1846_ FrameData[31] FrameStrobe[18] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1777_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q _0658_ _0682_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ FrameData[2] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1700_ G _0800_ _0110_ _0366_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ _0638_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2680_ Inst_LUT4AB_switch_matrix.WW4BEG0 net242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1631_ E1END[2] W1END[2] A B Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0584_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1493_ _0459_ _0452_ _0448_ _0460_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1562_ S1END[0] W1END[0] S2END[0] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q _0523_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ FrameData[11] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2045_ FrameData[6] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_60_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1829_ FrameData[14] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0993_ _0722_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q
+ _0836_ _0837_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_14_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2594_ Inst_LUT4AB_switch_matrix.JS2BEG7 net165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1614_ _0785_ _0568_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q _0569_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2663_ W6END[9] net236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1476_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0441_ _0442_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0443_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1545_ _0502_ _0503_ _0506_ _0507_ Inst_LUT4AB_switch_matrix.JS2BEG7 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2028_ FrameData[21] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1261_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0239_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1330_ _0300_ _0301_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0304_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1192_ _0167_ _0173_ _0158_ _0157_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q
+ _0174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0976_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q _0821_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2577_ NN4END[14] net139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2646_ Inst_LUT4AB_switch_matrix.JW2BEG6 net217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1459_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0386_ _0400_ _0427_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1528_ _0472_ _0492_ _0493_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ FrameData[21] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2431_ Inst_LUT4AB_switch_matrix.E1BEG0 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1244_ _0762_ _0221_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q _0224_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2362_ FrameData[3] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1313_ _0284_ _0288_ Inst_LUT4AB_switch_matrix.JW2BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2293_ FrameData[30] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_64_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1175_ N2END[7] S2END[7] EE4END[2] W2END[7] Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q _0158_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_23 NN4END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_12 N4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_34 SS4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0959_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _0805_ _0806_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_45 net248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput141 net141 NN4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput152 net152 NN4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput130 net130 N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2629_ SS4END[14] net191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput185 net185 S4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput196 net196 SS4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput163 net163 S2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput174 net174 S4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1793_ Inst_LE_LUT4c_frame_config_dffesr.c_reset_value _0694_ _0696_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1931_ FrameData[20] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1862_ FrameData[15] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2414_ FrameData[23] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2276_ FrameData[13] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2345_ FrameData[18] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1227_ _0206_ _0207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1158_ _0136_ _0137_ _0140_ _0141_ Inst_LUT4AB_switch_matrix.JS2BEG4 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1089_ _0072_ _0075_ _0077_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1012_ _0850_ _0854_ _0855_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2061_ FrameData[22] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2130_ FrameData[27] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1914_ FrameData[3] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ FrameData[30] FrameStrobe[18] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1776_ _0681_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop _0679_ _0002_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2328_ FrameData[1] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_55_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2259_ FrameData[28] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1630_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q _0583_ _0578_ Inst_LUT4AB_switch_matrix.JN2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1492_ _0458_ _0455_ _0436_ _0459_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1561_ _0777_ _0521_ _0522_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2113_ FrameData[10] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2044_ FrameData[5] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1759_ _0733_ Inst_LUT4AB_switch_matrix.E2BEG1 _0667_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_9_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1828_ FrameData[13] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0992_ N4END[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q _0836_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_14_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1544_ _0781_ _0504_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q _0507_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2593_ Inst_LUT4AB_switch_matrix.JS2BEG6 net164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1613_ F G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0568_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2662_ W6END[8] net235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1475_ _0438_ _0439_ _0442_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2027_ FrameData[20] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_20_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1260_ _0238_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ E VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1191_ _0169_ _0171_ _0173_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0975_ N2MID[6] S2MID[6] W2MID[6] Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q _0820_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2576_ NN4END[13] net153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1527_ _0490_ _0491_ _0492_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2645_ Inst_LUT4AB_switch_matrix.JW2BEG5 net216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1458_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0386_ _0400_ _0426_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1389_ N2MID[6] E2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q _0360_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2430_ _0007_ clknet_1_1__leaf_UserCLK_regs Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2361_ FrameData[2] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1243_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0222_ _0223_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1174_ N4END[3] W2END[3] E2END[3] Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q _0157_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1312_ _0752_ _0285_ _0287_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0288_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_2_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ FrameData[29] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_13 N4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_24 NN4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_46 EE4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0889_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q _0737_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_30_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_35 SS4END[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0958_ N1END[0] N2END[2] N4END[2] E2END[2] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _0805_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput142 net142 NN4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput153 net153 NN4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput131 net131 N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2559_ N4END[12] net136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput120 net120 N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2628_ SS4END[13] net205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput175 net175 S4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput197 net197 SS4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput186 net186 S4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput164 net164 S2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1930_ FrameData[19] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1792_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q _0671_ _0238_ _0695_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1861_ FrameData[14] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_26_Left_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2413_ FrameData[22] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2344_ FrameData[17] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2275_ FrameData[12] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1226_ _0204_ _0205_ _0195_ _0194_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
+ _0206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1157_ _0746_ _0138_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q _0141_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1088_ _0073_ _0074_ _0076_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1011_ _0853_ _0854_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2060_ FrameData[21] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1913_ FrameData[2] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1775_ Inst_LB_LUT4c_frame_config_dffesr.c_reset_value _0100_ _0680_ _0681_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1844_ FrameData[29] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2327_ FrameData[0] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2258_ FrameData[27] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_55_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1209_ N2MID[3] E2MID[3] Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q _0190_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2189_ FrameData[22] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1560_ N1END[0] N2END[0] E1END[0] EE4END[0] Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q _0521_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1491_ _0456_ _0457_ _0458_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2112_ FrameData[9] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2043_ FrameData[4] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_60_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1827_ FrameData[12] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1689_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0266_ _0629_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1758_ _0733_ Inst_LUT4AB_switch_matrix.JW2BEG1 _0665_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ _0666_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_68_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_13_Left_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0991_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0834_ _0835_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2661_ W6END[7] net234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1474_ _0437_ _0440_ _0441_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1543_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q _0505_ _0506_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2592_ Inst_LUT4AB_switch_matrix.JS2BEG5 net163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1612_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q _0566_ _0567_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ FrameData[19] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1190_ _0169_ _0171_ _0172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2644_ Inst_LUT4AB_switch_matrix.JW2BEG4 net215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0974_ _0813_ _0815_ _0818_ _0819_ Inst_LUT4AB_switch_matrix.JN2BEG3 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1457_ _0424_ _0404_ _0373_ _0425_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2575_ NN4END[12] net152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1526_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0473_ _0475_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0491_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1388_ _0353_ _0355_ _0358_ _0359_ Inst_LUT4AB_switch_matrix.JN2BEG6 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2009_ FrameData[2] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_33_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_47_Left_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1311_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q _0286_ _0287_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2360_ FrameData[1] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2291_ FrameData[28] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_56_Left_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1242_ S1END[0] S1END[2] S2END[6] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0222_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1173_ _0122_ _0144_ _0151_ _0154_ _0152_ _0156_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_2_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_14 N4END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_25 NN4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_36 SS4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_47 net231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput143 net143 NN4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput132 net132 N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput121 net121 N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_65_Left_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput110 net110 N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0957_ _0717_ _0803_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q _0804_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2627_ SS4END[12] net204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0888_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q _0736_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2558_ N4END[11] net135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2489_ FrameData[10] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1509_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0146_ _0473_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0474_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput154 net154 S1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput198 net198 SS4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput176 net176 S4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput187 net187 S4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput165 net165 S2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ FrameData[13] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_1_Left_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1791_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q _0671_ _0694_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2274_ FrameData[11] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2412_ FrameData[21] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2343_ FrameData[16] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1156_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0139_ _0140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1225_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q _0205_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_35_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1087_ _0074_ _0075_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ FrameData[14] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_58_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1010_ _0725_ _0852_ _0853_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_6_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1912_ FrameData[1] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1843_ FrameData[28] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1774_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q _0671_ _0680_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1208_ _0716_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ _0188_ _0189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2326_ FrameData[31] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2257_ FrameData[26] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2188_ FrameData[21] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1139_ A B D E Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ _0124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0442_ _0445_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0457_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2111_ FrameData[8] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2042_ FrameData[3] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ FrameData[11] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1688_ _0628_ _0627_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q Inst_LUT4AB_switch_matrix.EE4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q Inst_LUT4AB_switch_matrix.JS2BEG1
+ _0665_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_68_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ FrameData[14] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_48_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2660_ W6END[6] net233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0990_ _0833_ Ci Inst_LA_LUT4c_frame_config_dffesr.c_I0mux _0834_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1611_ B D C E Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ _0566_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1473_ _0439_ _0440_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1542_ S1END[0] W1END[0] S2END[0] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0505_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2591_ Inst_LUT4AB_switch_matrix.JS2BEG4 net162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2025_ FrameData[18] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1809_ FrameData[26] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_28_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2574_ NN4END[11] net151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2643_ Inst_LUT4AB_switch_matrix.JW2BEG3 net214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0973_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0816_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
+ _0819_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1456_ _0774_ _0401_ _0422_ _0423_ _0424_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1387_ _0731_ _0356_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0359_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1525_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0146_ _0147_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0490_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2008_ FrameData[1] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_25_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1241_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0221_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1310_ S4END[3] W2END[3] SS4END[3] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q _0286_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2290_ FrameData[27] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1172_ _0151_ _0154_ _0152_ _0155_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_48 EE4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_26 NN4END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_15 N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_37 SS4END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0956_ F G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _0803_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_22_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput133 net133 N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput144 net144 NN4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput100 net100 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2557_ N4END[10] net134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput111 net111 N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput122 net122 N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput166 net166 S2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2626_ SS4END[11] net203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput177 net177 S4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput155 net155 S1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0887_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0735_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2488_ FrameData[9] net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1508_ _0123_ _0144_ _0473_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput188 net188 S4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput199 net199 SS4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1439_ _0764_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q
+ _0407_ _0408_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1790_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop _0692_ _0693_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2411_ FrameData[20] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ FrameData[10] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2342_ FrameData[15] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_28_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1224_ N2MID[4] W2MID[4] S2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q _0204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1155_ S1END[1] S2END[5] W1END[1] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1086_ _0795_ _0800_ _0810_ _0809_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q
+ _0074_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1988_ FrameData[13] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0939_ A B C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ _0787_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2609_ S4END[10] net186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_58_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1911_ FrameData[0] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1842_ FrameData[27] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1773_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q _0658_ _0679_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2187_ FrameData[20] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1207_ W2MID[3] Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q _0188_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2325_ FrameData[30] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2256_ FrameData[25] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1138_ _0122_ _0123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1069_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0834_ _0058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2110_ FrameData[7] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2041_ FrameData[2] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_22_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1756_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q _0663_ _0664_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ FrameData[10] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_reset_value
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2308_ FrameData[13] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1687_ N1END[1] E1END[1] S1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0628_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ FrameData[8] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2590_ Inst_LUT4AB_switch_matrix.JS2BEG3 net161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1610_ _0560_ _0565_ Inst_LUT4AB_switch_matrix.JS2BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1472_ _0384_ _0385_ _0375_ _0374_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q
+ _0439_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1541_ N1END[0] N2END[0] E1END[0] E2END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q _0504_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2024_ FrameData[17] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1739_ _0401_ _0430_ _0445_ _0648_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1808_ FrameData[25] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0972_ _0709_ _0817_ _0818_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2573_ NN4END[10] net150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1524_ _0487_ _0488_ _0472_ _0489_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2642_ Inst_LUT4AB_switch_matrix.JW2BEG2 net213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1455_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0402_ _0403_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0423_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1386_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q _0357_ _0358_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2007_ FrameData[0] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_25_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1240_ _0762_ _0217_ _0763_ _0220_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1171_ _0078_ _0087_ _0088_ _0080_ _0154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_16 N4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_27 NN4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_49 Inst_LUT4AB_switch_matrix.E2BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_38 SS4END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0955_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _0801_ _0802_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0886_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop _0734_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput101 net101 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput123 net123 N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput134 net134 N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2556_ N4END[9] net133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput145 net145 NN4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2487_ FrameData[8] net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput112 net112 N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1507_ _0471_ _0155_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux _0472_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2625_ SS4END[10] net202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput178 net178 S4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput189 net189 S4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput156 net156 S1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput167 net167 S2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1369_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0319_ _0324_ _0341_
+ _0342_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_38_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1438_ W2END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q _0407_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_495 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ FrameData[19] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2341_ FrameData[14] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1154_ N1END[1] N2END[5] E1END[1] E2END[5] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1223_ _0197_ _0199_ _0202_ _0203_ Inst_LUT4AB_switch_matrix.JS2BEG5 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2272_ FrameData[9] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1085_ _0072_ _0073_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1987_ FrameData[12] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0869_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _0717_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0938_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0786_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2608_ S4END[9] net185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2539_ Inst_LUT4AB_switch_matrix.JN2BEG4 net110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_41_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ FrameData[31] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1772_ _0734_ _0676_ _0678_ _0001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1841_ FrameData[26] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2324_ FrameData[29] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2186_ FrameData[19] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1206_ N2MID[2] S2MID[2] E2MID[2] Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q _0187_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1137_ _0109_ _0110_ _0121_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q
+ _0122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2255_ FrameData[24] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_63_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1068_ _0023_ _0056_ _0057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ FrameData[1] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1686_ E _0204_ _0398_ _0831_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0627_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1755_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0172_ _0662_ _0663_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1824_ FrameData[9] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_I0mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2307_ FrameData[12] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2238_ FrameData[7] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ FrameData[2] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1540_ _0781_ _0500_ _0782_ _0503_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ _0437_ _0438_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ FrameData[16] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1807_ FrameData[24] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_17_Left_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1738_ C Inst_LUT4AB_switch_matrix.JW2BEG3 _0301_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q Inst_LUT4AB_switch_matrix.N1BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1669_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q G _0612_ _0613_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0971_ N2END[4] E1END[2] N4END[0] E2END[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _0817_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2572_ NN4END[9] net149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1454_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0387_ _0400_ _0422_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1523_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0473_ _0475_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ _0488_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2641_ Inst_LUT4AB_switch_matrix.JW2BEG1 net212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1385_ S1END[3] W1END[1] S2END[7] W1END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q _0357_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2006_ FrameData[31] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1170_ _0152_ _0153_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_17 NN4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_28 NN4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0885_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0733_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2624_ SS4END[9] net201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_39 SS4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0954_ A D C E Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ _0801_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput146 net146 NN4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput124 net124 N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput102 net102 N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2555_ N4END[8] net132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput135 net135 N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2486_ FrameData[7] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput113 net113 N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1506_ _0468_ _0470_ _0471_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Left_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput179 net179 S4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput157 net157 S1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput168 net168 S2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1437_ N2END[1] EE4END[3] Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q _0406_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1368_ _0767_ _0319_ _0341_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1299_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0153_ _0274_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0275_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_43_Left_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Left_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2340_ FrameData[13] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2271_ FrameData[8] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1153_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0134_ _0747_ _0137_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1222_ _0760_ _0200_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q _0203_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1084_ _0018_ _0020_ _0851_ _0849_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q
+ _0072_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1986_ FrameData[11] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ S4END[8] net184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0868_ S2MID[3] _0716_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0937_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q _0785_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2538_ Inst_LUT4AB_switch_matrix.JN2BEG3 net109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2469_ EE4END[10] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ FrameData[25] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1771_ Inst_LA_LUT4c_frame_config_dffesr.c_reset_value _0675_ _0676_ _0677_ _0678_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2254_ FrameData[23] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2323_ FrameData[28] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2185_ FrameData[18] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1205_ _0181_ _0182_ _0184_ _0186_ Inst_LUT4AB_switch_matrix.E2BEG5 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1136_ N2END[2] E2END[2] S2END[2] WW4END[2] Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q _0121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1067_ _0811_ _0054_ _0055_ _0053_ _0056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1969_ FrameData[26] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_3_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1823_ FrameData[8] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_out_mux VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1685_ _0623_ _0624_ _0626_ _0625_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ Inst_LUT4AB_switch_matrix.E6BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1754_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0252_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ _0662_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2306_ FrameData[11] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2237_ FrameData[6] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1119_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0105_ _0106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2099_ FrameData[28] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_13_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ FrameData[1] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1470_ _0398_ _0399_ _0389_ _0388_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q
+ _0437_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ FrameData[15] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1806_ _0702_ _0705_ _0706_ _0703_ _0007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1737_ D _0173_ Inst_LUT4AB_switch_matrix.JW2BEG0 _0194_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q Inst_LUT4AB_switch_matrix.N1BEG1 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1599_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q _0553_ _0555_ _0549_ _0551_ Inst_LUT4AB_switch_matrix.JW2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1668_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0799_ _0612_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2640_ Inst_LUT4AB_switch_matrix.JW2BEG0 net211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0970_ E6END[0] S2END[4] W2END[4] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q _0816_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2571_ NN4END[8] net148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1522_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0146_ _0147_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0487_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1453_ _0419_ _0420_ _0410_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q
+ _0421_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1384_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0356_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2005_ FrameData[30] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_18 NN4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_29 SS4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput125 net125 N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2554_ N4END[7] net131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput103 net103 N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0884_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0732_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput114 net114 N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0953_ _0799_ _0800_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2623_ SS4END[8] net200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput147 net147 NN4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput136 net136 N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2485_ FrameData[6] net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1367_ _0332_ _0336_ _0339_ _0340_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1505_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0266_ _0469_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ _0470_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput158 net158 S2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput169 net169 S2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1436_ NN4END[0] W2END[0] E6END[0] Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q _0405_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1298_ _0149_ _0150_ _0274_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_21_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1221_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0201_ _0202_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2270_ FrameData[7] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1152_ _0746_ _0135_ _0136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1083_ _0066_ _0069_ _0071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1985_ FrameData[10] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0936_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0784_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2606_ S4END[7] net183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2537_ Inst_LUT4AB_switch_matrix.JN2BEG2 net108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0867_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _0715_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_21_Left_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2468_ EE4END[9] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1419_ NN4END[1] S2END[5] E2END[5] W2END[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q _0389_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2399_ FrameData[8] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0063_ _0675_ _0677_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2253_ FrameData[22] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1204_ _0758_ _0185_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q _0186_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2322_ FrameData[27] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2184_ FrameData[17] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1135_ N4END[2] E2END[2] W2END[7] Inst_LUT4AB_switch_matrix.E2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q _0120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1066_ _0730_ _0834_ _0811_ _0055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1899_ FrameData[20] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0919_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0767_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1968_ FrameData[25] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1753_ _0733_ _0821_ _0660_ _0661_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1822_ FrameData[7] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1684_ G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0626_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2305_ FrameData[10] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2236_ FrameData[5] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2167_ FrameData[0] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1118_ S1END[1] S2END[5] S1END[3] W1END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q _0105_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2098_ FrameData[27] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1049_ F G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q _0039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ FrameData[14] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1805_ Inst_LG_LUT4c_frame_config_dffesr.c_reset_value _0704_ _0706_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1736_ E Inst_LUT4AB_switch_matrix.JW2BEG1 _0385_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q Inst_LUT4AB_switch_matrix.N1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1598_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0554_ _0555_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1667_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0110_ _0610_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ _0611_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2219_ FrameData[20] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_11_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2570_ NN4END[7] net147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1383_ _0731_ _0354_ _0732_ _0355_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1521_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q _0485_ _0484_ _0486_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1452_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q _0420_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2004_ FrameData[29] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1719_ S2END[1] S4END[0] W6END[0] D Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ Inst_LUT4AB_switch_matrix.S4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_19 NN4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0952_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q _0796_ _0798_ _0799_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput148 net148 NN4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput126 net126 N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput137 net137 N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2553_ N4END[6] net130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput104 net104 N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0883_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q _0731_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput115 net115 N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1504_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0262_ _0469_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2622_ SS4END[7] net199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput159 net159 S2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1435_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0386_ _0400_ _0404_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2484_ FrameData[5] net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1366_ _0337_ _0338_ _0319_ _0339_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1297_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0151_ _0272_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0273_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1151_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ _0135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1220_ S1END[2] W1END[0] S2END[6] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _0201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1082_ _0066_ _0069_ _0070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0935_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0783_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1984_ FrameData[9] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_33_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0866_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q _0714_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2605_ S4END[6] net182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2536_ Inst_LUT4AB_switch_matrix.JN2BEG1 net107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2467_ EE4END[8] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1349_ _0187_ _0192_ _0178_ _0177_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q
+ _0322_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1418_ E6END[1] S4END[1] WW4END[3] Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q _0388_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2398_ FrameData[7] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2321_ FrameData[26] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1203_ N1END[2] N2END[6] E1END[2] E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0185_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2252_ FrameData[21] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1134_ Inst_LUT4AB_switch_matrix.E2BEG2 _0119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2183_ FrameData[16] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_33_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1065_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0834_ _0054_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1898_ FrameData[19] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0918_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0766_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1967_ FrameData[24] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2519_ FrameStrobe[8] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Left_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1683_ _0800_ _0110_ _0192_ _0385_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0625_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1752_ _0733_ _0363_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0660_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1821_ FrameData[6] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2304_ FrameData[9] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1117_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0103_ _0743_ _0104_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2097_ FrameData[26] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2235_ FrameData[4] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2166_ FrameData[31] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1048_ _0726_ _0037_ _0038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2020_ FrameData[13] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1804_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q _0671_ _0429_ _0705_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1735_ F _0020_ Inst_LUT4AB_switch_matrix.JW2BEG2 _0830_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q Inst_LUT4AB_switch_matrix.N1BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1666_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0409_ _0610_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1597_ N1END[3] E2END[1] N2END[1] E6END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _0554_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ FrameData[19] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2149_ FrameData[14] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1520_ _0300_ _0301_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q _0485_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1382_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0354_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1451_ N2MID[0] E2MID[0] W2MID[0] Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q _0419_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2003_ FrameData[28] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_35_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1718_ F Inst_LUT4AB_switch_matrix.JS2BEG3 _0301_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q Inst_LUT4AB_switch_matrix.W1BEG0 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1649_ N1END[0] W1END[0] S1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ _0599_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0951_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q _0716_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ _0797_ _0798_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0882_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0730_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2483_ FrameData[4] net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput149 net149 NN4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput138 net138 NN4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput105 net105 N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2552_ N4END[5] net129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput127 net127 N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput116 net116 N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1503_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0250_ _0467_ _0468_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2621_ SS4END[6] net198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1434_ _0386_ _0400_ _0403_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1365_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0327_ _0329_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0338_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1296_ _0149_ _0150_ _0272_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1150_ F G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_45_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1081_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q _0067_ _0068_ _0069_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2604_ S4END[5] net181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1983_ FrameData[8] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0934_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q _0782_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0865_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0713_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1417_ _0386_ _0387_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2535_ Inst_LUT4AB_switch_matrix.JN2BEG0 net106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2466_ EE4END[7] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1348_ _0320_ _0321_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1279_ F G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0256_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2397_ FrameData[6] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_28_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2251_ FrameData[20] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2320_ FrameData[25] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1202_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0183_ _0184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1133_ _0112_ _0114_ _0117_ _0118_ Inst_LUT4AB_switch_matrix.E2BEG2 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1064_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0834_ _0053_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2182_ FrameData[15] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_18_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1966_ FrameData[23] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0917_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0765_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1897_ FrameData[18] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2518_ FrameStrobe[7] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2449_ E2MID[6] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1820_ FrameData[5] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1751_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q _0658_ _0659_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1682_ C D E F Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0624_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_68_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ FrameData[3] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_31_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2303_ FrameData[8] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1116_ F G H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2096_ FrameData[25] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2165_ FrameData[30] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1047_ A B C E Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1949_ FrameData[6] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q _0671_ _0704_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_68_Left_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1665_ _0609_ _0608_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q Inst_LUT4AB_switch_matrix.SS4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1596_ _0784_ _0552_ _0553_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1734_ N2END[2] N4END[1] E6END[1] E Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ Inst_LUT4AB_switch_matrix.N4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2217_ FrameData[18] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2148_ FrameData[13] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2079_ FrameData[8] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0414_ _0416_ _0418_ Inst_LUT4AB_switch_matrix.JW2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1381_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q _0352_ _0353_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2002_ FrameData[27] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0535_ _0537_ _0538_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1648_ C _0192_ _0385_ _0133_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ _0598_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1717_ G _0173_ Inst_LUT4AB_switch_matrix.JS2BEG0 _0194_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q Inst_LUT4AB_switch_matrix.W1BEG1 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0950_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q W2MID[3] _0797_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2620_ SS4END[5] net197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0881_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0729_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput128 net128 N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2551_ N4END[4] net122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1433_ _0387_ _0400_ _0402_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2482_ FrameData[3] net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput106 net106 N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput139 net139 NN4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput117 net117 N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1502_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0252_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ _0467_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1364_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0323_ _0324_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0337_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_38_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1295_ _0269_ _0270_ _0271_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1080_ _0736_ _0036_ _0068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1982_ FrameData[7] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_43_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2603_ S4END[4] net174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2534_ Inst_LUT4AB_switch_matrix.N1BEG3 net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0933_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q _0781_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0864_ S2MID[7] _0712_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2465_ EE4END[6] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1347_ _0204_ _0205_ _0195_ _0194_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
+ _0320_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1416_ _0384_ _0385_ _0375_ _0374_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q
+ _0386_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2396_ FrameData[5] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1278_ _0740_ _0254_ _0255_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1201_ S1END[0] S1END[2] S2END[6] W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2250_ FrameData[19] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1132_ _0744_ _0115_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q _0118_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1063_ _0026_ _0051_ _0023_ _0052_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2181_ FrameData[14] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_25_Left_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1965_ FrameData[22] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0916_ S2END[1] _0764_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1896_ FrameData[17] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2517_ FrameStrobe[6] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2379_ FrameData[20] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2448_ E2MID[5] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1750_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0650_ _0652_ _0654_ _0657_ _0658_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1681_ E1END[3] W1END[3] A B Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0623_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2233_ FrameData[2] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2164_ FrameData[29] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2302_ FrameData[7] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1115_ _0742_ _0101_ _0102_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2095_ FrameData[24] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1046_ N2END[0] S2END[0] E2END[0] WW4END[3] Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q _0036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_0_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1948_ FrameData[5] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1879_ FrameData[0] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1802_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop _0702_ _0703_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1733_ N2END[3] N4END[2] E6END[0] F Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ Inst_LUT4AB_switch_matrix.N4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_13_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1664_ N1END[3] E1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ _0609_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1595_ S2END[1] W2END[1] S4END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _0552_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2147_ FrameData[12] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2216_ FrameData[17] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1029_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q _0020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2078_ FrameData[7] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_12_Left_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1380_ E H F Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q _0352_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ FrameData[26] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_63_476 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1716_ H Inst_LUT4AB_switch_matrix.JS2BEG1 _0385_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q Inst_LUT4AB_switch_matrix.W1BEG2 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1578_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q Inst_LUT4AB_switch_matrix.JS2BEG7
+ _0536_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0537_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1647_ _0597_ _0596_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q Inst_LUT4AB_switch_matrix.WW4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ N2MID[7] net121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput107 net107 N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0880_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0728_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput129 net129 N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2481_ FrameData[2] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1432_ _0386_ _0400_ _0401_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1501_ E F _0466_ Inst_LUT4AB_switch_matrix.M_EF VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput118 net118 N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1363_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0335_ _0334_ _0336_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1294_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux _0154_ _0270_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_46_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2679_ WW4END[15] net241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ FrameData[6] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_43_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0932_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q _0780_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2533_ Inst_LUT4AB_switch_matrix.N1BEG2 net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0863_ N2MID[7] _0711_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2602_ S2MID[7] net173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1346_ _0318_ _0317_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux _0319_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2464_ EE4END[5] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1415_ N2MID[3] E2MID[3] S2MID[3] W2MID[3] Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q _0385_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2395_ FrameData[4] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1277_ A B D E Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ _0254_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2180_ FrameData[13] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1200_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0179_ _0759_ _0182_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_0_Left_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1131_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q _0116_ _0117_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1062_ _0049_ _0050_ _0811_ _0051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1895_ FrameData[16] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1964_ FrameData[21] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0915_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q _0763_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2516_ FrameStrobe[5] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2447_ E2MID[4] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2378_ FrameData[19] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1329_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0291_ _0302_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
+ _0303_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1680_ _0619_ _0622_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q Inst_LUT4AB_switch_matrix.E6BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2301_ FrameData[6] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1114_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0101_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ FrameData[28] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2232_ FrameData[1] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2094_ FrameData[23] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1045_ N4END[0] E6END[0] S4END[0] Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q _0035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1947_ FrameData[4] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1878_ FrameData[31] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q _0658_ _0702_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1732_ N2END[0] N4END[3] W6END[1] G Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ Inst_LUT4AB_switch_matrix.N4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1663_ H _0018_ _0142_ _0215_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ _0608_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_13_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1594_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0550_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ _0551_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ FrameData[11] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ FrameData[6] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2215_ FrameData[16] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1028_ _0015_ _0017_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q _0857_ _0019_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_70_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2000_ FrameData[25] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_31_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1715_ A _0020_ Inst_LUT4AB_switch_matrix.JS2BEG2 _0830_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q Inst_LUT4AB_switch_matrix.W1BEG3 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1646_ N1END[1] S1END[1] W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ _0597_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1577_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q _0516_ _0536_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2129_ FrameData[26] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ FrameData[1] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1500_ _0464_ _0465_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0466_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput119 net119 N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput108 net108 N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput90 net90 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1431_ _0398_ _0399_ _0389_ _0388_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q
+ _0400_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1293_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux _0253_ _0268_ _0269_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1362_ _0225_ _0226_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0335_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2678_ WW4END[14] net240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1629_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0582_ _0581_ _0583_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ FrameData[5] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0931_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0779_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0862_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q _0710_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2532_ Inst_LUT4AB_switch_matrix.N1BEG1 net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2463_ EE4END[4] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2601_ S2MID[6] net172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1345_ _0167_ _0173_ _0158_ _0157_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q
+ _0318_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1414_ N2MID[2] W2MID[2] S2MID[2] Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q _0384_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2394_ FrameData[3] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1276_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0252_ _0251_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ _0253_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1130_ E6END[1] S2END[3] W2END[3] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1061_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0834_ _0050_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1894_ FrameData[15] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1963_ FrameData[20] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0914_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0762_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2515_ FrameStrobe[4] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2446_ E2MID[3] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2377_ FrameData[18] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1259_ _0232_ _0237_ _0228_ _0238_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1328_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0289_ _0302_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2231_ FrameData[0] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2300_ FrameData[5] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_7_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2093_ FrameData[22] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1113_ _0100_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1044_ _0028_ _0030_ _0033_ _0034_ Inst_LUT4AB_switch_matrix.JW2BEG1 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2162_ FrameData[27] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1946_ FrameData[3] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1877_ FrameData[30] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2429_ _0006_ clknet_1_1__leaf_UserCLK_regs Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1800_ _0697_ _0700_ _0701_ _0698_ _0006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_13_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1662_ _0607_ _0606_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q Inst_LUT4AB_switch_matrix.SS4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1731_ N2END[1] W6END[0] N4END[0] H Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ Inst_LUT4AB_switch_matrix.N4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2214_ FrameData[15] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_37_Left_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1593_ B D C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ _0550_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2145_ FrameData[10] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_26_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1027_ N2MID[4] E2MID[4] W2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q _0018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2076_ FrameData[5] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1929_ FrameData[18] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_46_Left_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_55_Left_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Left_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _0647_ _0646_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q Inst_LUT4AB_switch_matrix.NN4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1576_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q Inst_LUT4AB_switch_matrix.JN2BEG7
+ _0534_ _0535_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1645_ E _0204_ _0398_ _0851_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ _0596_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2128_ FrameData[25] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_49_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ FrameData[20] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput1 net1 Co VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1430_ N2MID[5] E2MID[5] S2MID[5] W2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q _0399_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput109 net109 N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput80 net80 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput91 net91 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1292_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0262_ _0267_ _0268_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1361_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0216_ _0333_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q
+ _0334_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_46_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1559_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0517_ _0778_ _0520_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2677_ WW4END[13] net254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1628_ N2END[1] E1END[3] N4END[1] E2END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _0582_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0930_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q _0778_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2600_ S2MID[5] net171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0861_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0709_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2462_ Inst_LUT4AB_switch_matrix.E6BEG1 net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1413_ _0378_ _0379_ _0382_ _0383_ Inst_LUT4AB_switch_matrix.E2BEG6 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2531_ Inst_LUT4AB_switch_matrix.N1BEG0 net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2393_ FrameData[2] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1344_ _0145_ _0156_ _0208_ _0211_ _0317_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1275_ N2MID[7] E2MID[7] S2MID[7] W2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q _0252_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1060_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0834_ _0049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1962_ FrameData[19] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_18_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ FrameData[14] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0913_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q _0761_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2514_ FrameStrobe[3] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2376_ FrameData[17] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2445_ E2MID[2] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1258_ _0236_ _0233_ _0176_ _0237_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_54_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1189_ _0711_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q _0170_ _0171_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1327_ N2MID[1] E2MID[1] S2MID[1] W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q _0301_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2230_ FrameData[31] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2092_ FrameData[21] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1043_ _0728_ _0031_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0034_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2161_ FrameData[26] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1112_ _0093_ _0099_ _0089_ _0100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1945_ FrameData[2] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1876_ FrameData[29] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2428_ _0005_ clknet_1_1__leaf_UserCLK_regs Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2359_ FrameData[0] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1730_ D Inst_LUT4AB_switch_matrix.JN2BEG3 _0301_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q Inst_LUT4AB_switch_matrix.E1BEG0 VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1661_ N1END[0] W1END[0] E1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ _0607_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1592_ _0784_ _0548_ _0549_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2213_ FrameData[14] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2144_ FrameData[9] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_64_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1026_ _0016_ _0017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2075_ FrameData[4] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1928_ FrameData[17] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1859_ FrameData[12] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1713_ N1END[2] W1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ _0647_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1575_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q _0533_ _0534_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1644_ _0592_ _0593_ _0595_ _0594_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ Inst_LUT4AB_switch_matrix.W6BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2127_ FrameData[24] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_49_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2058_ FrameData[19] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1009_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q _0851_ _0852_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput2 net2 E1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1360_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0214_ _0333_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput81 net81 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput92 net92 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1291_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0266_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ _0267_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_46_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2676_ WW4END[12] net253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1489_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0441_ _0444_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0456_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1558_ _0777_ _0518_ _0519_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1627_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0580_ _0581_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0860_ W2MID[6] _0708_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2530_ FrameStrobe[19] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2461_ Inst_LUT4AB_switch_matrix.E6BEG0 net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1412_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q _0380_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q
+ _0383_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1343_ _0316_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ C VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2392_ FrameData[1] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1274_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0250_ _0251_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0989_ _0820_ _0821_ _0831_ _0830_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q
+ _0833_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2659_ W6END[5] net232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_19_Left_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1892_ FrameData[13] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0912_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0760_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1961_ FrameData[18] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2513_ FrameStrobe[2] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2375_ FrameData[16] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2444_ E2MID[1] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1326_ N2MID[0] S2MID[0] W2MID[0] Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q _0300_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1257_ _0765_ _0208_ _0235_ _0236_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1188_ E2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ _0170_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2160_ FrameData[25] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_51_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ FrameData[20] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1111_ _0094_ _0095_ _0098_ _0099_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1042_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0032_ _0033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1944_ FrameData[1] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1875_ FrameData[28] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_16_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2427_ _0004_ clknet_1_0__leaf_UserCLK_regs Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1309_ N1END[1] N2END[3] EE4END[3] E6END[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0285_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2358_ FrameData[31] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2289_ FrameData[26] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_8_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_470 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1660_ C _0192_ _0385_ _0290_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ _0606_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1591_ F G H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q _0548_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2143_ FrameData[8] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2212_ FrameData[13] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1025_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q W2MID[4] Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
+ _0016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2074_ FrameData[3] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1927_ FrameData[16] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1858_ FrameData[11] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1789_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q _0658_ _0692_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_1 net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1712_ G _0800_ _0110_ _0375_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ _0646_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_6_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1643_ G H Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0595_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1574_ Inst_LUT4AB_switch_matrix.E2BEG7 _0533_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2057_ FrameData[18] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2126_ FrameData[23] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_49_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1008_ N2END[4] S2END[4] EE4END[0] W2END[4] Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q _0851_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_24_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput93 net93 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput82 net82 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput71 net71 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput60 net60 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput3 net3 E1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1290_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q _0265_ _0264_ _0266_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_46_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ WW4END[11] net252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1626_ _0579_ _0580_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1488_ _0453_ _0454_ _0455_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1557_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0518_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2109_ FrameData[6] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2460_ E6END[11] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1411_ _0769_ _0381_ _0382_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1273_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q _0247_ _0249_ _0250_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1342_ _0311_ _0315_ _0307_ _0316_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2391_ FrameData[0] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0988_ _0831_ _0832_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2589_ Inst_LUT4AB_switch_matrix.JS2BEG2 net160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2658_ W6END[4] net231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1609_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0561_ _0564_ _0565_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1891_ FrameData[12] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1960_ FrameData[17] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0911_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q _0759_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ FrameStrobe[1] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2443_ E2MID[0] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1256_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0209_ _0211_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0234_ _0235_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_56_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1325_ _0293_ _0295_ _0298_ _0299_ Inst_LUT4AB_switch_matrix.JW2BEG4 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2374_ FrameData[15] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_62_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1187_ _0712_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ _0168_ _0169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput250 net250 WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ FrameData[19] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1110_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0080_ _0097_ _0070_
+ _0098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1041_ S2END[2] W2END[2] S4END[2] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q _0032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_16_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1943_ FrameData[0] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1874_ FrameData[27] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2426_ _0003_ clknet_1_0__leaf_UserCLK_regs Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1239_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0218_ _0219_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2288_ FrameData[25] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1308_ _0752_ _0280_ _0283_ _0284_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2357_ FrameData[30] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_70_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1590_ A B _0465_ Inst_LUT4AB_switch_matrix.M_AB VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2142_ FrameData[7] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2211_ FrameData[12] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1024_ _0009_ _0010_ _0012_ _0014_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q _0015_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2073_ FrameData[2] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1926_ FrameData[15] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1788_ _0687_ _0690_ _0691_ _0688_ _0004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1857_ FrameData[10] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2409_ FrameData[18] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_70_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Left_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Left_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1711_ _0645_ _0644_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q Inst_LUT4AB_switch_matrix.NN4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_2 E6END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1642_ _0800_ _0110_ _0192_ _0385_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0594_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_60_Left_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1573_ _0527_ _0528_ _0531_ _0532_ Inst_LUT4AB_switch_matrix.E2BEG7 VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2056_ FrameData[17] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2125_ FrameData[22] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_49_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1007_ _0846_ _0848_ _0721_ _0837_ _0850_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1909_ FrameData[30] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput83 net83 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput94 net94 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput61 net61 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput50 net50 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput72 net72 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput4 net4 E1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_46_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1556_ E G F Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q _0517_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2674_ WW4END[10] net251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1625_ E6END[1] SS4END[1] W2END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0579_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1487_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0442_ _0444_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0454_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2108_ FrameData[5] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2039_ FrameData[0] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ N1END[3] N2END[7] E1END[3] E2END[7] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0381_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_5_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1272_ _0708_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
+ _0248_ _0249_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1341_ _0269_ _0270_ _0314_ _0305_ _0315_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2390_ FrameData[31] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0987_ N2END[6] SS4END[3] E2END[6] W2END[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q _0831_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1539_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q _0501_ _0502_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2588_ Inst_LUT4AB_switch_matrix.JS2BEG1 net159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2657_ W6END[3] net230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1608_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0563_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ _0564_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ FrameData[11] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0910_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0758_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2511_ FrameStrobe[0] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2373_ FrameData[14] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2442_ Inst_LUT4AB_switch_matrix.E2BEG7 net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1255_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0193_ _0207_ _0234_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1324_ _0750_ _0296_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q _0299_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1186_ W2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q _0168_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput251 net251 WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput240 net240 WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1040_ N1END[0] E2END[2] N2END[2] E6END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q _0031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1942_ FrameData[31] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_46_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ FrameData[26] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2425_ _0002_ clknet_1_0__leaf_UserCLK_regs Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2356_ FrameData[29] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1238_ E G H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0218_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1169_ _0148_ _0150_ _0152_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2287_ FrameData[24] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_37_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1307_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0282_ _0283_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ FrameData[11] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2141_ FrameData[6] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_64_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1023_ _0009_ _0010_ _0012_ _0014_ Inst_LUT4AB_switch_matrix.JS2BEG3 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2072_ FrameData[1] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1925_ FrameData[14] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ Inst_LD_LUT4c_frame_config_dffesr.c_reset_value _0689_ _0691_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1856_ FrameData[9] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2339_ FrameData[12] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2408_ FrameData[17] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_70_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1710_ N1END[3] E1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0645_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_3 EE4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1572_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0529_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ _0532_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1641_ C D E F Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0593_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2124_ FrameData[21] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2055_ FrameData[16] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1006_ N4END[1] E6END[1] W6END[1] Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q _0849_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1908_ FrameData[29] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1839_ FrameData[24] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput5 net5 E1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput84 net84 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput73 net73 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput95 net95 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput40 net40 EE4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput51 net51 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput62 net62 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1555_ _0516_ Inst_LUT4AB_switch_matrix.JW2BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2673_ WW4END[9] net250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1624_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0574_ _0577_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
+ _0578_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1486_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0441_ _0445_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0453_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2107_ FrameData[4] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_37_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2038_ FrameData[31] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1340_ _0312_ _0313_ _0314_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1271_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q Inst_LUT4AB_switch_matrix.JN2BEG4
+ _0248_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0986_ NN4END[3] WW4END[0] S4END[3] Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q _0830_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2656_ W6END[2] net227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1469_ _0775_ _0401_ _0430_ _0435_ _0436_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1538_ E G F Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0501_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2587_ Inst_LUT4AB_switch_matrix.JS2BEG0 net158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1607_ _0562_ _0563_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ FrameData[31] net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1323_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q _0297_ _0298_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2372_ FrameData[13] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2441_ Inst_LUT4AB_switch_matrix.E2BEG6 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1254_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0193_ _0206_ _0233_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1185_ N2MID[6] W2MID[6] E2MID[6] Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_62_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput230 net230 W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput252 net252 WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2639_ Inst_LUT4AB_switch_matrix.W1BEG3 net210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0969_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0814_ _0710_ _0815_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput241 net241 WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1941_ FrameData[30] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1872_ FrameData[25] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2286_ FrameData[23] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1306_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q _0281_ _0282_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2355_ FrameData[28] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2424_ _0001_ clknet_1_0__leaf_UserCLK_regs Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1237_ A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0217_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1168_ _0148_ _0150_ _0151_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1099_ _0811_ _0024_ _0087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_2140_ FrameData[5] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1022_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _0013_ _0720_ _0014_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2071_ FrameData[0] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1924_ FrameData[13] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1855_ FrameData[8] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1786_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q _0671_ _0495_ _0690_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2338_ FrameData[11] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2269_ FrameData[6] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_2407_ FrameData[16] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_4 EE4END[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_1571_ _0779_ _0530_ _0531_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1640_ E1END[3] W1END[3] A B Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0592_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ FrameData[20] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_469 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ FrameData[15] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1005_ _0847_ _0848_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1907_ FrameData[28] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1838_ FrameData[23] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1769_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q _0658_ _0676_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput41 net41 EE4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput52 net52 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput30 net30 E6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput6 net6 E2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput85 net85 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput96 net96 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput74 net74 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput63 net63 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ WW4END[8] net249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1485_ _0451_ _0447_ _0436_ _0452_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1554_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q _0515_ _0512_ _0516_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1623_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0576_ _0577_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

