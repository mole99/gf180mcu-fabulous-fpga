* NGSPICE file created from GF_SRAM.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

.subckt GF_SRAM A_SRAM0 A_SRAM1 A_SRAM2 A_SRAM3 A_SRAM4 A_SRAM5 A_SRAM6 A_SRAM7 A_SRAM8
+ CEN_SRAM CLK_SRAM CONFIGURED_top D_SRAM0 D_SRAM1 D_SRAM2 D_SRAM3 D_SRAM4 D_SRAM5
+ D_SRAM6 D_SRAM7 GWEN_SRAM Q_SRAM0 Q_SRAM1 Q_SRAM2 Q_SRAM3 Q_SRAM4 Q_SRAM5 Q_SRAM6
+ Q_SRAM7 Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3] Tile_X0Y0_E2END[4]
+ Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0] Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5] Tile_X0Y0_E2MID[6]
+ Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0] Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1]
+ Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3] Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6]
+ Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10]
+ Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14]
+ Tile_X0Y0_EE4END[15] Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7]
+ Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10]
+ Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14]
+ Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18]
+ Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21]
+ Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25]
+ Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29]
+ Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3]
+ Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7]
+ Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10]
+ Tile_X0Y0_FrameData_O[11] Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14]
+ Tile_X0Y0_FrameData_O[15] Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18]
+ Tile_X0Y0_FrameData_O[19] Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21]
+ Tile_X0Y0_FrameData_O[22] Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25]
+ Tile_X0Y0_FrameData_O[26] Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29]
+ Tile_X0Y0_FrameData_O[2] Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3]
+ Tile_X0Y0_FrameData_O[4] Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7]
+ Tile_X0Y0_FrameData_O[8] Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3]
+ Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0]
+ Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5]
+ Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11]
+ Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5]
+ Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo
+ Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2] Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0]
+ Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5]
+ Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2]
+ Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6]
+ Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10] Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1]
+ Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4] Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6]
+ Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10]
+ Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14]
+ Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3]
+ Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7]
+ Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9] Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11]
+ Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5]
+ Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11] Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15] Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6]
+ Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8] Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0]
+ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13]
+ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17]
+ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20]
+ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24]
+ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28]
+ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31]
+ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6]
+ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0]
+ Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11] Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13]
+ Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15] Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17]
+ Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19] Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20]
+ Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22] Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24]
+ Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26] Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28]
+ Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2] Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31]
+ Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4] Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6]
+ Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8] Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0]
+ Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13]
+ Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15] Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17]
+ Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2]
+ Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6]
+ Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2] Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1]
+ Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3] Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6]
+ Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0] Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3]
+ Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5] Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0]
+ Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11] Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13]
+ Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15] Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3]
+ Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5] Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8]
+ Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3]
+ Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4]
+ Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1]
+ Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3] Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5]
+ Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7] Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11]
+ Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13] Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15]
+ Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3] Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5]
+ Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8] Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK
+ Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2] Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0]
+ Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5]
+ Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2]
+ Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6]
+ Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10] Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1]
+ Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4] Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6]
+ Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10]
+ Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14]
+ Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3]
+ Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7]
+ Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9] VDD VSS WEN_SRAM0 WEN_SRAM1 WEN_SRAM2 WEN_SRAM3
+ WEN_SRAM4 WEN_SRAM5 WEN_SRAM6 WEN_SRAM7
X_0298_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 Tile_X0Y0_S2MID[1]
+ Tile_X0Y1_N2MID[1] Tile_X0Y0_S2END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0367_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Left_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1270_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11 net132 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0221_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q _0150_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_74_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0985_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0419_ _0152_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 _0035_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_97_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1399_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12 net261 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0770_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1253_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2 net124 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1322_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3 net193 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1184_ Tile_X0Y1_FrameStrobe[2] net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_121_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0968_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput242 net242 Tile_X0Y1_W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput220 net220 Tile_X0Y1_S4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0899_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput264 net264 Tile_X0Y1_WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput231 net231 Tile_X0Y1_W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput275 net275 WEN_SRAM1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput253 net253 Tile_X0Y1_W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_104_Right_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0822_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_80_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0684_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0753_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_54_Left_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1236_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2 net98 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1305_ Tile_X0Y1_FrameData[18] net167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1167_ Tile_X0Y0_FrameData[17] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1098_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_118_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1021_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_46_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0805_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_62_Left_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0736_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0667_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_71_Left_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0598_ _0139_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0118_ _0119_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1219_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 net90 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_119_Left_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_128_Left_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0452_ _0057_ _0056_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
+ net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_5 Tile_X0Y0_S2MID[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0521_ Tile_X0Y1_N1END[2] Tile_X0Y1_N4END[2] _0194_ Tile_X0Y0_S4END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_137_Left_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0383_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_49_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1004_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0719_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput53 net53 Tile_X0Y0_FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput64 net64 Tile_X0Y0_FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput75 net75 Tile_X0Y0_N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput42 net42 Tile_X0Y0_FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput31 net31 Tile_X0Y0_FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput20 net20 GWEN_SRAM VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput7 net7 A_SRAM6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput97 net97 Tile_X0Y0_N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput86 net86 Tile_X0Y0_N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0435_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0022_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q _0046_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0504_ Q_SRAM1 _0001_ Q_SRAM2 _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_136_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0366_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0297_ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[6] _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0220_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q _0149_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_74_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0984_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0418_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q _0034_
+ _0033_ _0032_ net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_97_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0349_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 Q_SRAM5 Tile_X0Y0_S1END[3]
+ Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1398_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11 net260 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_118_Right_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1252_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1 net123 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1321_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2 net192 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1183_ Tile_X0Y1_FrameStrobe[1] net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0967_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_101_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput243 net243 Tile_X0Y1_W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput265 net265 Tile_X0Y1_WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput221 net221 Tile_X0Y1_S4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput210 net210 Tile_X0Y1_S4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput232 net232 Tile_X0Y1_W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput276 net276 WEN_SRAM2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput254 net254 Tile_X0Y1_W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0898_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Right_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_100_Left_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0821_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0752_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_127_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0683_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1235_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1 net97 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1166_ Tile_X0Y0_FrameData[16] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1304_ Tile_X0Y1_FrameData[17] net166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1097_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_109_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1020_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_61_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0735_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0804_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_115_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0666_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0597_ Tile_X0Y1_N2END[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ _0118_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1218_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 net89 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1149_ clknet_1_0__leaf_Tile_X0Y1_UserCLK net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_6 Tile_X0Y0_S2MID[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0451_ Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[12]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ _0057_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0382_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0520_ Q_SRAM0 Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1003_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0718_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0649_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_82_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput87 net87 Tile_X0Y0_N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput98 net98 Tile_X0Y0_N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput54 net54 Tile_X0Y0_FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput65 net65 Tile_X0Y0_FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput76 net76 Tile_X0Y0_N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput43 net43 Tile_X0Y0_FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput32 net32 Tile_X0Y0_FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput21 net21 Tile_X0Y0_FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput10 net10 CEN_SRAM VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput8 net8 A_SRAM7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_54_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0434_ _0045_ _0044_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0365_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_68_Right_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0503_ Q_SRAM0 Q_SRAM3 _0002_ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_136_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0296_ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1
+ Tile_X0Y0_S2MID[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q _0000_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_77_Right_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_86_Right_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_95_Right_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0983_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_66_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0417_ Tile_X0Y0_E2END[2] _0151_ _0034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0348_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 Q_SRAM4 Tile_X0Y0_S1END[2]
+ Q_SRAM6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1397_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10 net259 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0279_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1320_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1 net191 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1182_ Tile_X0Y1_FrameStrobe[0] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1251_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0 net122 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0966_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput200 net200 Tile_X0Y1_S2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0897_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_59_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput244 net244 Tile_X0Y1_W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput211 net211 Tile_X0Y1_S4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput266 net266 Tile_X0Y1_WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput222 net222 Tile_X0Y1_S4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput233 net233 Tile_X0Y1_W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput277 net277 WEN_SRAM3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput255 net255 Tile_X0Y1_W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0820_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0751_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0682_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1303_ Tile_X0Y1_FrameData[16] net165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1234_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0 net96 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1165_ Tile_X0Y0_FrameData[15] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1096_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0949_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0665_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0734_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0803_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_84_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0596_ Tile_X0Y1_E2MID[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0108_ _0116_ _0117_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1217_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 net88 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1079_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1148_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_37_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_7 Tile_X0Y0_S2MID[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0381_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0450_ Tile_X0Y0_E6END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_E6END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
+ _0056_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1002_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_17_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0648_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0717_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_122_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0579_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 _0185_ _0074_
+ _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ _0103_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput55 net55 Tile_X0Y0_FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput66 net66 Tile_X0Y0_FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput99 net99 Tile_X0Y0_N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput44 net44 Tile_X0Y0_FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput77 net77 Tile_X0Y0_N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput88 net88 Tile_X0Y0_N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput33 net33 Tile_X0Y0_FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput22 net22 Tile_X0Y0_FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput9 net9 A_SRAM8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput11 net11 CLK_SRAM VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0502_ Q_SRAM0 Q_SRAM3 _0002_ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0433_ Tile_X0Y0_E1END[2] Tile_X0Y0_E6END[10] Tile_X0Y0_EE4END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ _0045_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0295_ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[9] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0364_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_77_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_68_Left_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_77_Left_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_Right_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_101_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0982_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_42_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0416_ Tile_X0Y0_E2MID[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q _0033_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0347_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 Q_SRAM5 Tile_X0Y0_S1END[1]
+ Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_65_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0278_ Tile_X0Y1_E1END[2] _0195_ Tile_X0Y1_E6END[6] _0199_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1396_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9 net273 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1181_ Tile_X0Y0_FrameData[31] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1250_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7 net121 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0896_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0965_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput234 net234 Tile_X0Y1_W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput223 net223 Tile_X0Y1_S4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput201 net201 Tile_X0Y1_S2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput212 net212 Tile_X0Y1_S4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput245 net245 Tile_X0Y1_W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput267 net267 Tile_X0Y1_WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput278 net278 WEN_SRAM4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput256 net256 Tile_X0Y1_W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1379_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4 net252 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Left_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0681_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0750_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_96_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1302_ Tile_X0Y1_FrameData[15] net164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1233_ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_23_Left_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1164_ Tile_X0Y0_FrameData[14] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_32_Left_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1095_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_118_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0948_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0879_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_133_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_41_Left_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_50_Left_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_141_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0802_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_91_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0664_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0733_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1216_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 net87 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0595_ _0140_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0116_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1078_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1147_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_8 Tile_X0Y1_FrameStrobe[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0380_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1001_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_89_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0647_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0716_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_103_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0578_ Tile_X0Y1_E1END[1] Tile_X0Y1_EE4END[13] Tile_X0Y1_E6END[5] _0078_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q _0102_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_139_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput34 net34 Tile_X0Y0_FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput23 net23 Tile_X0Y0_FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput12 net12 D_SRAM0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput56 net56 Tile_X0Y0_FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput67 net67 Tile_X0Y0_FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput89 net89 Tile_X0Y0_N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput45 net45 Tile_X0Y0_FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput78 net78 Tile_X0Y0_N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Right_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0432_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0023_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q _0044_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0501_ Q_SRAM1 _0001_ Q_SRAM2 _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0294_ Tile_X0Y0_E2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_77_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0363_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0981_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_42_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0415_ _0151_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 _0032_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1395_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8 net272 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0346_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 Q_SRAM4 Tile_X0Y0_S1END[0]
+ Q_SRAM6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0277_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q _0198_
+ _0197_ _0196_ _0199_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1180_ Tile_X0Y0_FrameData[30] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0964_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0895_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput268 net268 Tile_X0Y1_WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput202 net202 Tile_X0Y1_S2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput224 net224 Tile_X0Y1_S4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput213 net213 Tile_X0Y1_S4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput235 net235 Tile_X0Y1_W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput246 net246 Tile_X0Y1_W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput257 net257 Tile_X0Y1_W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0329_ Tile_X0Y0_E2MID[0] Tile_X0Y0_E2END[0] Tile_X0Y0_E6END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1378_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3 net251 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput279 net279 WEN_SRAM5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0680_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1232_ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1301_ Tile_X0Y1_FrameData[14] net163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1163_ Tile_X0Y0_FrameData[13] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1094_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_118_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0947_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0878_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_18_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0801_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0663_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_123_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0732_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0594_ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ _0115_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1215_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1 net86 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_127_Right_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1146_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1077_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_9 Tile_X0Y1_FrameStrobe[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1000_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0715_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_143_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0646_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0577_ _0101_ _0100_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_139_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1129_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_0_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput57 net57 Tile_X0Y0_FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput35 net35 Tile_X0Y0_FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput24 net24 Tile_X0Y0_FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput46 net46 Tile_X0Y0_FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput13 net13 D_SRAM1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput68 net68 Tile_X0Y0_FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput79 net79 Tile_X0Y0_N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0431_ _0043_ _0042_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0362_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_28_Right_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0500_ Q_SRAM1 _0000_ Q_SRAM2 _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0293_ Tile_X0Y0_E1END[3] Tile_X0Y0_E6END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0203_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_62_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Right_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Right_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0629_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_55_Right_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_125_Left_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Right_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_134_Left_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_Right_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_143_Left_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_141_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0980_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_94_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_91_Right_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0414_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q _0031_
+ _0030_ _0029_ net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1394_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7 net271 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0345_ _0018_ _0019_ _0021_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0276_ _0158_ _0194_ _0198_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0894_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0963_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_99_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput258 net258 Tile_X0Y1_WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput225 net225 Tile_X0Y1_S4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput214 net214 Tile_X0Y1_S4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput203 net203 Tile_X0Y1_S2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput269 net269 Tile_X0Y1_WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput236 net236 Tile_X0Y1_W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput247 net247 Tile_X0Y1_W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0328_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 Tile_X0Y0_S2MID[7]
+ Tile_X0Y1_N2MID[7] Tile_X0Y0_S2END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1377_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2 net250 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0259_ Tile_X0Y0_E1END[1] Tile_X0Y0_E6END[9] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0183_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
+ _0184_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_120_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Right_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1231_ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A net108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1162_ Tile_X0Y0_FrameData[12] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1300_ Tile_X0Y1_FrameData[13] net162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1093_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0877_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0946_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_7_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0800_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0731_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0662_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_27_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0593_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q _0110_
+ _0113_ _0114_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1214_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 net85 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1145_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1076_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_136_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0929_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0645_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_128_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0714_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_57_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0576_ Tile_X0Y1_E1END[0] Tile_X0Y1_EE4END[12] Tile_X0Y1_E6END[4] _0079_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q _0101_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_122_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1128_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1059_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_38_Left_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput69 net69 Tile_X0Y0_FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput58 net58 Tile_X0Y0_FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput36 net36 Tile_X0Y0_FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput25 net25 Tile_X0Y0_FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput47 net47 Tile_X0Y0_FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput14 net14 D_SRAM2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_47_Left_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0430_ Tile_X0Y0_E1END[1] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ _0043_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0361_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_104_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0292_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0628_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_68_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0559_ _0163_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ _0002_ _0089_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0413_ Tile_X0Y0_E2END[1] _0150_ _0031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0275_ Tile_X0Y1_N1END[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q _0197_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1393_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6 net270 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0344_ Tile_X0Y1_E1END[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ _0020_ _0021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_132_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0893_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0962_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_99_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput259 net259 Tile_X0Y1_WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput204 net204 Tile_X0Y1_S2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput215 net215 Tile_X0Y1_S4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput237 net237 Tile_X0Y1_W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput226 net226 Tile_X0Y1_W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput248 net248 Tile_X0Y1_W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0258_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q _0181_
+ _0182_ _0180_ _0183_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1376_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1 net249 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0327_ Tile_X0Y1_E2MID[0] Tile_X0Y1_E2END[0] Tile_X0Y1_E6END[0] _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_120_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1230_ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A net107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1161_ Tile_X0Y0_FrameData[11] net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1092_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_49_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0876_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0945_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_10_Left_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1359_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0 net230 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_141_Right_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0661_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0730_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_6_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1213_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7 net84 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0592_ Tile_X0Y1_E2END[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q _0112_ _0113_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1144_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1075_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_37_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0859_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0928_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0644_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0713_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0575_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 _0012_ _0075_
+ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ _0100_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_107_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1058_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1127_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput59 net59 Tile_X0Y0_FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput37 net37 Tile_X0Y0_FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput26 net26 Tile_X0Y0_FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput48 net48 Tile_X0Y0_FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 D_SRAM3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0360_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0291_ Tile_X0Y1_E1END[3] _0205_ Tile_X0Y1_E6END[7] _0209_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0627_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0558_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q _0087_
+ _0088_ _0086_ net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_97_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0489_ Tile_X0Y1_N1END[2] Q_SRAM0 _0194_ Q_SRAM2 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_2_Left_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0412_ Tile_X0Y0_E2MID[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q _0030_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1392_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5 net269 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0274_ Tile_X0Y1_E6END[2] _0158_ _0196_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0343_ _0154_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ _0020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0961_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_65_Left_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput216 net216 Tile_X0Y1_S4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput205 net205 Tile_X0Y1_S2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0892_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_101_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Left_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1375_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0 net246 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput238 net238 Tile_X0Y1_W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput227 net227 Tile_X0Y1_W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput249 net249 Tile_X0Y1_W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0257_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 _0182_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0326_ Tile_X0Y1_N2MID[7] Tile_X0Y1_N2END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q _0006_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_120_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_122_Right_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_104_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_92_Left_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1160_ Tile_X0Y0_FrameData[10] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1091_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0944_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0875_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_95_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1358_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3 net229 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0309_ Tile_X0Y0_E2MID[4] Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1289_ Tile_X0Y1_FrameData[2] net180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0660_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0591_ _0142_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ _0111_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0112_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1212_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6 net83 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1143_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1074_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0927_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0858_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0789_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_75_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0643_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0712_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0574_ _0099_ _0098_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1126_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_48_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1057_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput38 net38 Tile_X0Y0_FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput27 net27 Tile_X0Y0_FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput49 net49 Tile_X0Y0_FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput16 net16 D_SRAM4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0290_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q _0207_
+ _0208_ _0206_ _0209_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_39_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0557_ Tile_X0Y1_E2END[2] _0162_ _0088_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0626_ _0138_ _0137_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1109_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0488_ Tile_X0Y1_N1END[1] Q_SRAM1 _0184_ Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_24_Right_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Right_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_67_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_103_Left_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Right_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_112_Left_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0411_ _0150_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 _0029_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1391_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4 net268 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0342_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q _0012_
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q _0019_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_121_Left_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_60_Right_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0273_ Tile_X0Y1_N1END[2] Tile_X0Y1_N4END[2] _0194_ Tile_X0Y0_S4END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q _0195_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_130_Left_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_103_Right_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_85_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0609_ Tile_X0Y1_E6END[2] _0077_ Tile_X0Y1_E6END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
+ _0127_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_123_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0960_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput239 net239 Tile_X0Y1_W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput217 net217 Tile_X0Y1_S4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput206 net206 Tile_X0Y1_S2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput228 net228 Tile_X0Y1_W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0891_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0325_ Tile_X0Y0_E1END[3] Tile_X0Y0_E2MID[0] Tile_X0Y0_E2END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1374_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7 net245 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0256_ _0145_ Tile_X0Y0_S1END[1] _0181_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1090_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0874_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0943_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_62_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0308_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3 Tile_X0Y1_N2MID[3]
+ Tile_X0Y0_S2MID[3] Tile_X0Y0_S2END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1288_ Tile_X0Y1_FrameData[1] net169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1357_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2 net228 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0239_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0 Tile_X0Y0_S2MID[0]
+ Tile_X0Y1_N2MID[0] Tile_X0Y0_S2END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_1__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_1__leaf_Tile_X0Y1_UserCLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0590_ Tile_X0Y1_E2END[5] _0164_ _0111_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1211_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5 net82 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1142_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1073_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0857_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0926_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_89_Right_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0788_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_98_Right_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0711_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0642_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0573_ Tile_X0Y1_E1END[3] Tile_X0Y1_E6END[11] Tile_X0Y1_EE4END[3] _0076_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q _0099_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1125_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1056_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_33_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput39 net39 Tile_X0Y0_FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput28 net28 Tile_X0Y0_FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0909_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput17 net17 D_SRAM5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_16_Left_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_117_Right_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_112_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0625_ Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[11] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0138_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0487_ Tile_X0Y1_N1END[0] Q_SRAM0 _0011_ Q_SRAM2 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0556_ Tile_X0Y1_E2MID[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
+ _0087_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_135_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1039_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_13_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1108_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_83_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0410_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q _0028_
+ _0027_ _0026_ net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1390_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3 net267 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0341_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q _0013_
+ _0016_ _0018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_132_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0272_ Tile_X0Y0_E1END[2] Tile_X0Y0_E6END[10] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0193_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ _0194_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_100_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0608_ _0126_ _0125_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ net275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0539_ Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 _0072_
+ _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0890_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput207 net207 Tile_X0Y1_S2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput218 net218 Tile_X0Y1_S4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput229 net229 Tile_X0Y1_W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0255_ Tile_X0Y0_E6END[1] _0145_ _0180_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0324_ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2END[1] Tile_X0Y0_E6END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1373_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6 net244 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Left_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0873_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0942_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_55_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1356_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1 net227 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0238_ Tile_X0Y1_E2MID[7] Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[7] _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0307_ Tile_X0Y1_E2MID[4] Tile_X0Y1_E6END[4] Tile_X0Y1_E2END[4] _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1287_ Tile_X0Y1_FrameData[0] net158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1210_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4 net81 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1141_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1072_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0856_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0787_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0925_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_28_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1339_ Tile_X0Y0_S4END[8] net210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_Left_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_98_Left_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_86_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0710_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_128_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0641_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0572_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 _0205_ _0072_
+ _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ _0098_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1055_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1124_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput29 net29 Tile_X0Y0_FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0839_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_102_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0908_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput18 net18 D_SRAM6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0624_ Tile_X0Y1_E6END[3] _0076_ Tile_X0Y1_E6END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0137_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_5_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0555_ _0162_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ _0001_ _0086_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0486_ Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0] Tile_X0Y1_E2MID[0] _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_135_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1107_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1038_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_122_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0271_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q _0191_
+ _0192_ _0190_ _0193_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_79_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0340_ _0013_ _0016_ _0017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_35_Left_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_100_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0538_ Tile_X0Y1_N4END[3] Tile_X0Y0_S4END[7] _0075_ _0012_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0607_ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[9] Tile_X0Y1_EE4END[13]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
+ _0126_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_44_Left_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0469_ Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[14]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ _0069_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_53_Left_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput219 net219 Tile_X0Y1_S4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput208 net208 Tile_X0Y1_S2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0323_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 Tile_X0Y0_S2MID[6]
+ Tile_X0Y1_N2MID[6] Tile_X0Y0_S2END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1372_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5 net243 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0254_ _0143_ _0172_ _0174_ _0179_ _0144_ net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_135_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Left_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0941_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0872_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_118_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Left_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_87_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1355_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0 net226 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1286_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15 net148 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0306_ Tile_X0Y1_N2MID[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3
+ Tile_X0Y1_N2END[3] Tile_X0Y0_S2MID[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q _0002_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0237_ Tile_X0Y1_N2MID[0] Tile_X0Y1_N2END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0
+ Tile_X0Y0_S2MID[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q _0165_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_127_Left_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_136_Left_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_119_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1071_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1140_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0924_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_28_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0855_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0786_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1338_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7 net209 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1269_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10 net131 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0640_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0571_ _0097_ _0096_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1054_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_16_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1123_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0907_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0838_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_131_Right_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0769_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput19 net19 D_SRAM7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_138_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_70 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0554_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q _0084_
+ _0085_ _0083_ net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_0623_ _0136_ _0135_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_135_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0485_ Tile_X0Y1_E1END[2] Tile_X0Y1_E2MID[1] Tile_X0Y1_E2END[1] _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1106_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_103_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1037_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_130_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_113_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Right_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0270_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 _0192_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0537_ Tile_X0Y1_N4END[2] Tile_X0Y0_S4END[6] _0074_ _0185_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0606_ Tile_X0Y1_E6END[1] _0078_ Tile_X0Y1_E6END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ _0125_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0468_ Tile_X0Y0_E6END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_E6END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
+ _0068_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0399_ Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 _0022_
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0322_ Tile_X0Y1_E2MID[1] Tile_X0Y1_E6END[1] Tile_X0Y1_E2END[1] _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1371_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4 net242 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput209 net209 Tile_X0Y1_S2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0253_ _0176_ _0178_ _0143_ _0179_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0940_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0871_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_126_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0305_ Tile_X0Y0_E2MID[4] Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[11] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1285_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14 net147 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1354_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 net216 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0236_ Tile_X0Y0_E2MID[7] Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1070_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0854_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_112_Right_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0923_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0785_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Right_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_114_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1268_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9 net141 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_58_Right_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1337_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 net208 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1199_ Tile_X0Y1_FrameStrobe[17] net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0219_ Tile_X0Y0_E2END[4] _0148_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_67_Right_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_76_Right_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0570_ Tile_X0Y1_E1END[2] Tile_X0Y1_E6END[10] Tile_X0Y1_EE4END[2] _0077_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q _0097_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_94_Right_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_65_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1122_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_115_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1053_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0837_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0906_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0699_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0768_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_8_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_60 Tile_X0Y1_N4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0622_ Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[14]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0136_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0553_ Tile_X0Y1_E2END[1] _0161_ _0085_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0484_ Tile_X0Y1_E1END[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2END[2] _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_76_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1105_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_103_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1036_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_123_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_126_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0467_ _0067_ _0066_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ net279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0536_ Tile_X0Y1_N4END[1] Tile_X0Y0_S4END[5] _0073_ _0195_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0605_ _0124_ _0123_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
+ net274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0398_ Tile_X0Y1_N4END[7] Tile_X0Y0_S4END[3] _0025_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1019_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_118_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0321_ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q _0005_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1370_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3 net241 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0252_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q _0175_
+ _0177_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q _0178_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_31_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0519_ Tile_X0Y1_N1END[3] Tile_X0Y1_N4END[3] _0204_ Tile_X0Y0_S4END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_126_Right_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_120_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0870_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_70_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0304_ Tile_X0Y0_E2MID[5] Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1284_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13 net146 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1353_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2 net215 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0235_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q _0164_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_117_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0853_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0922_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0784_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1198_ Tile_X0Y1_FrameStrobe[16] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1267_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8 net140 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0218_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q _0147_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1336_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 net207 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_58_Left_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_67_Left_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_76_Left_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_111_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1121_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1052_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_115_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0836_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0767_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0905_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0698_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_138_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1319_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0 net190 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_61 Tile_X0Y1_N4END[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_50 Q_SRAM5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput190 net190 Tile_X0Y1_S1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0621_ Tile_X0Y1_E6END[2] _0077_ Tile_X0Y1_E6END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0135_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0552_ Tile_X0Y1_E2MID[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
+ _0084_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0483_ Tile_X0Y1_E1END[0] Tile_X0Y1_E2END[3] Tile_X0Y1_E2MID[3] _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1035_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_16_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1104_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_103_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0819_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_115_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0604_ Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[8] Tile_X0Y1_EE4END[12]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ _0124_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0397_ Tile_X0Y1_N4END[6] Tile_X0Y0_S4END[2] _0024_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0466_ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[9] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
+ _0067_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Right_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0535_ Tile_X0Y1_N4END[0] Tile_X0Y0_S4END[4] _0072_ _0205_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_13_Left_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1018_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_22_Left_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Left_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0320_ Tile_X0Y0_E1END[2] Tile_X0Y0_E2MID[1] Tile_X0Y0_E2END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0251_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y1_E2END[3] _0177_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0518_ Q_SRAM0 Q_SRAM3 _0075_ _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0449_ _0055_ _0054_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0303_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2 Tile_X0Y1_N2MID[2]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1283_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12 net145 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1352_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1 net214 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0234_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q _0163_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0998_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_86_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0921_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_65_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0852_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0783_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1335_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 net206 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1197_ Tile_X0Y1_FrameStrobe[15] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0217_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q _0146_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1266_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7 net139 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_120_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1120_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1051_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_115_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0904_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_142_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0697_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0835_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0766_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_138_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1318_ Tile_X0Y1_FrameData[31] net182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1249_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6 net120 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_40 Tile_X0Y1_N4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_51 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_62 net212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput180 net180 Tile_X0Y1_FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput191 net191 Tile_X0Y1_S1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0551_ _0161_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ _0000_ _0083_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0620_ _0134_ _0133_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0482_ Tile_X0Y1_E2MID[4] Tile_X0Y1_E6END[11] Tile_X0Y1_E2END[4] _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1034_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1103_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0818_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_107_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0749_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_95_Left_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0534_ Q_SRAM0 Q_SRAM3 _0079_ _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0603_ Tile_X0Y1_E6END[0] _0079_ Tile_X0Y1_E6END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
+ _0123_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0465_ Tile_X0Y0_E6END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_E6END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ _0066_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0396_ Tile_X0Y1_N4END[5] Tile_X0Y0_S4END[1] _0023_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_131_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1017_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0250_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q _0142_
+ _0176_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_140_Right_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0517_ Tile_X0Y1_N1END[0] Tile_X0Y1_N4END[0] _0011_ Tile_X0Y0_S4END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q _0075_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0448_ Tile_X0Y0_E1END[3] Tile_X0Y0_E6END[7] Tile_X0Y0_EE4END[15] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ _0055_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0379_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0302_ Tile_X0Y1_E2MID[5] Tile_X0Y1_E6END[5] Tile_X0Y1_E2END[5] _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1351_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0 net213 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1282_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11 net144 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0233_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q _0162_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0997_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_39_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0920_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0851_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0782_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1265_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6 net138 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1334_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3 net205 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_18_Right_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_28_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1196_ Tile_X0Y1_FrameStrobe[14] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0216_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q _0145_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_27_Right_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_36_Right_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_113_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Right_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Right_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_115_Left_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_111_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_124_Left_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1050_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0834_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0903_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_133_Left_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0696_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0765_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_72_Right_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_142_Left_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1317_ Tile_X0Y1_FrameData[30] net181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_81_Right_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1248_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5 net119 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1179_ Tile_X0Y0_FrameData[29] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_41 Tile_X0Y1_N4END[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_52 Tile_X0Y1_FrameStrobe[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_30 Tile_X0Y1_N4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_90_Right_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_63 net225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput181 net181 Tile_X0Y1_FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput170 net170 Tile_X0Y1_FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput192 net192 Tile_X0Y1_S1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0550_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q _0081_
+ _0082_ _0080_ net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1102_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0481_ Tile_X0Y1_E2MID[5] Tile_X0Y1_E6END[10] Tile_X0Y1_E2END[5] _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_143_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1033_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0817_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_107_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0679_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0748_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_121_Right_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0464_ _0065_ _0064_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
+ net278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0533_ Tile_X0Y1_N1END[0] Tile_X0Y1_N4END[0] _0011_ Tile_X0Y0_S4END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q _0079_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0602_ _0122_ net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0395_ Tile_X0Y1_N4END[4] Tile_X0Y0_S4END[0] _0022_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_131_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1016_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0447_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0022_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q _0054_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0516_ Q_SRAM1 _0074_ Q_SRAM2 _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0378_ Q_SRAM4 Q_SRAM7 _0025_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1350_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3 net212 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1281_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10 net143 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0301_ Tile_X0Y1_N2MID[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2
+ Tile_X0Y1_N2END[2] Tile_X0Y0_S2MID[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q _0001_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0232_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q _0161_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0996_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_132_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_19_Left_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Left_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_37_Left_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0850_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Left_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0781_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1402_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15 net264 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1264_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5 net137 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1333_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 net204 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0215_ CONFIGURED_top _0144_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1195_ Tile_X0Y1_FrameStrobe[13] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0979_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_105_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0833_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0902_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_142_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_135_Right_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0695_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0764_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_51_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1178_ Tile_X0Y0_FrameData[28] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1316_ Tile_X0Y1_FrameData[29] net179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1247_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4 net118 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_31 Tile_X0Y1_N4END[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_20 Tile_X0Y1_N2MID[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_53 Tile_X0Y1_FrameStrobe[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_42 Tile_X0Y1_N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_64 net225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Right_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput182 net182 Tile_X0Y1_FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput171 net171 Tile_X0Y1_FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput160 net160 Tile_X0Y1_FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput193 net193 Tile_X0Y1_S1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0480_ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[9] _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1101_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_53_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1032_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0816_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0747_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0678_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_123_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0601_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q _0121_
+ _0114_ _0122_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0463_ Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[12]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ _0065_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0394_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0532_ Q_SRAM1 _0078_ Q_SRAM2 _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1015_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0446_ _0053_ _0052_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0377_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q _0025_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0515_ Tile_X0Y1_N1END[1] Tile_X0Y1_N4END[1] _0184_ Tile_X0Y0_S4END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q _0074_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0300_ Tile_X0Y0_E2MID[5] Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[10] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1280_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9 net157 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0231_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q _0160_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0995_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_117_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0429_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0024_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q _0042_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0780_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_116_Right_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1401_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14 net263 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1194_ Tile_X0Y1_FrameStrobe[12] net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1263_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4 net136 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1332_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1 net203 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0214_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q _0143_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0978_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_109_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0832_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0763_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0901_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0694_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1315_ Tile_X0Y1_FrameData[28] net178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1177_ Tile_X0Y0_FrameData[27] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1246_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3 net117 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_10 Tile_X0Y1_FrameStrobe[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_54 Tile_X0Y1_FrameStrobe[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_32 Tile_X0Y1_N4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_21 Tile_X0Y1_N2MID[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_43 Tile_X0Y1_N4END[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_65 net278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput150 net150 Tile_X0Y0_WW4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput161 net161 Tile_X0Y1_FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput172 net172 Tile_X0Y1_FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput183 net183 Tile_X0Y1_FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput194 net194 Tile_X0Y1_S2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1031_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1100_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_143_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0746_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0815_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0677_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_130_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1229_ Tile_X0Y1_N4END[15] net106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_134_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Left_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_73_Left_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Left_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_91_Left_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0531_ Tile_X0Y1_N1END[1] Tile_X0Y1_N4END[1] _0184_ Tile_X0Y0_S4END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q _0078_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0600_ _0117_ _0120_ _0121_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0462_ Tile_X0Y0_E6END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_E6END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
+ _0064_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0393_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_96_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1014_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_139_Left_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0729_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_134_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0514_ Q_SRAM1 _0073_ Q_SRAM2 _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0445_ Tile_X0Y0_E1END[2] Tile_X0Y0_E6END[6] Tile_X0Y0_EE4END[14] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
+ _0053_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0376_ Q_SRAM5 _0024_ Q_SRAM6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0230_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q _0159_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0994_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_140_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0428_ _0041_ _0040_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0359_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1331_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 net202 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1400_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13 net262 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1193_ Tile_X0Y1_FrameStrobe[11] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1262_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3 net135 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0213_ Tile_X0Y0_S2MID[2] _0142_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0977_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_142_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_23_Right_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_132_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0900_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_32_Right_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0693_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0831_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0762_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_102_Left_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ Tile_X0Y1_FrameData[27] net177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_41_Right_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1176_ Tile_X0Y0_FrameData[26] net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1245_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2 net116 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_50_Right_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_33 Tile_X0Y1_N4END[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_11 Tile_X0Y1_FrameStrobe[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_55 Tile_X0Y1_FrameStrobe[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_44 Tile_X0Y1_N4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Left_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_66 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_22 Tile_X0Y1_N2MID[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_120_Left_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput140 net140 Tile_X0Y0_W6BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput151 net151 Tile_X0Y0_WW4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput173 net173 Tile_X0Y1_FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput162 net162 Tile_X0Y1_FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput184 net184 Tile_X0Y1_FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput195 net195 Tile_X0Y1_S2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1030_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_36_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0814_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_115_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0745_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0676_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1228_ Tile_X0Y1_N4END[14] net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1159_ Tile_X0Y0_FrameData[9] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0530_ Q_SRAM1 _0077_ Q_SRAM2 _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0461_ _0063_ _0062_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0392_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1013_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_19_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0728_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0659_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_122_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0444_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0023_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q _0052_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0513_ Tile_X0Y1_N1END[2] Tile_X0Y1_N4END[2] _0194_ Tile_X0Y0_S4END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q _0073_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0375_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q _0024_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_79_Right_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_57_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_88_Right_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_141_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Right_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0993_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_117_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0427_ Tile_X0Y0_E1END[0] Tile_X0Y0_EE4END[0] Tile_X0Y0_E6END[8] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ _0041_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0358_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0289_ Tile_X0Y1_N1END[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q _0208_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_130_Right_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1261_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2 net134 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1330_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7 net201 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1192_ Tile_X0Y1_FrameStrobe[10] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0212_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q _0141_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0976_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_67_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0830_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_92_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0761_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0692_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_41_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1313_ Tile_X0Y1_FrameData[26] net176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1244_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1 net115 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1175_ Tile_X0Y0_FrameData[25] net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_114_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_34 Tile_X0Y1_N4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_56 Tile_X0Y1_FrameStrobe[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_45 Tile_X0Y1_N4END[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_12 Tile_X0Y1_FrameStrobe[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_23 Tile_X0Y1_N2MID[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_67 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0959_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput141 net141 Tile_X0Y0_W6BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput130 net130 Tile_X0Y0_W6BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput152 net152 Tile_X0Y0_WW4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput174 net174 Tile_X0Y1_FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput163 net163 Tile_X0Y1_FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput185 net185 Tile_X0Y1_FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput196 net196 Tile_X0Y1_S2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0813_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0744_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0675_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1227_ Tile_X0Y1_N4END[13] net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1158_ Tile_X0Y0_FrameData[8] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1089_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0460_ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
+ _0063_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0391_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_96_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1012_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0727_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_7_Left_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0658_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_84_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0589_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 _0108_ _0109_
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ _0110_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_84_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0443_ _0051_ _0050_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0374_ Q_SRAM4 Q_SRAM6 _0023_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0512_ Q_SRAM0 Q_SRAM3 _0072_ _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Left_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Left_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0992_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_97_Left_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0426_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ _0025_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q _0040_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0357_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0288_ _0159_ _0204_ _0207_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1191_ Tile_X0Y1_FrameStrobe[9] net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1260_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1 net133 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0211_ Tile_X0Y1_N2END[3] _0140_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0975_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_59_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0409_ Tile_X0Y0_E2END[0] _0149_ _0028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1389_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2 net266 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0760_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_127_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0691_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1174_ Tile_X0Y0_FrameData[24] net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1312_ Tile_X0Y1_FrameData[25] net175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1243_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0 net114 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_13 Tile_X0Y1_FrameStrobe[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_35 Tile_X0Y1_N4END[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_46 Tile_X0Y1_FrameStrobe[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_57 Tile_X0Y1_FrameStrobe[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_68 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0889_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_24 Tile_X0Y1_N2MID[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0958_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_25_Left_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput131 net131 Tile_X0Y0_W6BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput142 net142 Tile_X0Y0_WW4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput153 net153 Tile_X0Y0_WW4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput175 net175 Tile_X0Y1_FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput120 net120 Tile_X0Y0_W2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput164 net164 Tile_X0Y1_FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput186 net186 Tile_X0Y1_FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput197 net197 Tile_X0Y1_S2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_34_Left_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Left_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0743_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0812_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0674_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_99_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1226_ Tile_X0Y1_N4END[12] net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1157_ Tile_X0Y0_FrameData[7] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_102_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1088_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_125_Right_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0390_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_60_Left_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1011_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0726_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_108_Left_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0657_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0588_ Tile_X0Y1_E2END[4] Tile_X0Y0_S2MID[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ _0109_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1209_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3 net80 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_117_Left_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_126_Left_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0511_ Tile_X0Y1_N1END[3] Tile_X0Y1_N4END[3] _0204_ Tile_X0Y0_S4END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q _0072_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0373_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q _0023_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0442_ Tile_X0Y0_E1END[1] Tile_X0Y0_E6END[5] Tile_X0Y0_EE4END[13] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ _0051_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0709_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0991_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_5_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0425_ _0148_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q _0038_ _0039_
+ net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_0356_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0287_ Tile_X0Y1_E6END[3] _0159_ _0206_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1190_ Tile_X0Y1_FrameStrobe[8] net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0210_ Tile_X0Y1_N2MID[6] _0139_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0974_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_113_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0408_ Tile_X0Y0_E2MID[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q _0027_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1388_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1 net265 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0339_ Tile_X0Y1_E6END[0] _0156_ _0015_ _0016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0690_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1311_ Tile_X0Y1_FrameData[24] net174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_139_Right_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1173_ Tile_X0Y0_FrameData[23] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1242_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3 net113 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_47 Tile_X0Y1_FrameStrobe[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_36 Tile_X0Y1_N4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_14 Tile_X0Y1_FrameStrobe[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_25 Tile_X0Y1_N2MID[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_58 Tile_X0Y1_FrameStrobe[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput132 net132 Tile_X0Y0_W6BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput143 net143 Tile_X0Y0_WW4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput121 net121 Tile_X0Y0_W2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput110 net110 Tile_X0Y0_W1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_69 Tile_X0Y0_S4END[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0888_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0957_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_30_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput154 net154 Tile_X0Y0_WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput176 net176 Tile_X0Y1_FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput165 net165 Tile_X0Y1_FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput187 net187 Tile_X0Y1_FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput198 net198 Tile_X0Y1_S2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_137_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Right_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0673_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0742_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0811_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_99_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1225_ Tile_X0Y1_N4END[11] net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1156_ Tile_X0Y0_FrameData[6] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1087_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_102_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1010_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_32_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0656_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0725_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1208_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2 net79 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0587_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q _0164_
+ _0108_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1139_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0510_ Q_SRAM0 Q_SRAM3 _0012_ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0441_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0024_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q _0050_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0372_ Q_SRAM4 Q_SRAM7 _0022_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0639_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0708_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_97_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_39_Right_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Right_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0990_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0424_ Tile_X0Y0_E2MID[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q _0039_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Right_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_Right_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0355_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0286_ Tile_X0Y1_N1END[3] Tile_X0Y1_N4END[3] _0204_ Tile_X0Y0_S4END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q _0205_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Right_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0973_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0407_ _0149_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0 _0026_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1387_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0 net258 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0269_ _0146_ Tile_X0Y0_S1END[2] _0191_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0338_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q _0014_
+ _0015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1310_ Tile_X0Y1_FrameData[23] net173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1241_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2 net112 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1172_ Tile_X0Y0_FrameData[22] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_15 Tile_X0Y1_FrameStrobe[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_37 Tile_X0Y1_N4END[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_59 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_48 Tile_X0Y1_N2MID[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0956_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XANTENNA_26 Tile_X0Y1_N2MID[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput100 net100 Tile_X0Y0_N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput133 net133 Tile_X0Y0_W6BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput144 net144 Tile_X0Y0_WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput155 net155 Tile_X0Y0_WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput177 net177 Tile_X0Y1_FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput122 net122 Tile_X0Y0_W2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput166 net166 Tile_X0Y1_FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput111 net111 Tile_X0Y0_W1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0887_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_7_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput188 net188 Tile_X0Y1_FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput199 net199 Tile_X0Y1_S2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0810_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0672_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0741_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1224_ Tile_X0Y1_N4END[10] net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1155_ Tile_X0Y0_FrameData[5] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1086_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_37_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0939_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0655_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0724_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_69_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0586_ _0107_ _0106_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1207_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1 net78 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1138_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1069_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_40_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Left_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0440_ _0049_ _0048_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_92_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0371_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q _0022_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0707_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0638_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0569_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 _0195_ _0073_
+ _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ _0096_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Left_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0423_ _0153_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 _0038_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_66_Left_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0354_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0285_ Tile_X0Y0_E1END[3] Tile_X0Y0_E6END[11] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0203_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ _0204_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0972_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_58_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0406_ Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1386_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11 net248 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0337_ Tile_X0Y1_N1END[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ _0014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0268_ Tile_X0Y0_E6END[2] _0146_ _0190_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1171_ Tile_X0Y0_FrameData[21] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_79_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1240_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1 net111 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_38 Tile_X0Y1_N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_16 Tile_X0Y1_FrameStrobe[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_27 Tile_X0Y1_N2MID[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Right_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_49 Tile_X0Y1_N2MID[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0955_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0886_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_32_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput101 net101 Tile_X0Y0_N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput134 net134 Tile_X0Y0_W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput156 net156 Tile_X0Y0_WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput145 net145 Tile_X0Y0_WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput178 net178 Tile_X0Y1_FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput123 net123 Tile_X0Y0_W2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput167 net167 Tile_X0Y1_FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput112 net112 Tile_X0Y0_W1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput189 net189 Tile_X0Y1_FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1369_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2 net240 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_105_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_12_Left_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Left_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0740_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_14_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_30_Left_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0671_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1223_ Tile_X0Y1_N4END[9] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1154_ Tile_X0Y0_FrameData[4] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1085_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0869_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0938_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_121_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0723_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0654_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_103_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0585_ Tile_X0Y1_E1END[3] Tile_X0Y1_EE4END[15] Tile_X0Y1_E6END[7] _0076_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q _0107_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1206_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0 net77 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1137_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1068_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_124_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0370_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_92_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0706_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0637_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0568_ _0095_ _0094_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0499_ Q_SRAM0 Q_SRAM3 _0165_ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0422_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q _0037_
+ _0036_ _0035_ net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_0353_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_79_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0284_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q _0201_
+ _0202_ _0200_ _0203_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_134_Right_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_101_Right_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0971_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_113_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0267_ Tile_X0Y0_E1END[1] Tile_X0Y0_E6END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0183_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0405_ Q_SRAM6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1385_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10 net247 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0336_ _0156_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0011_ _0013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1170_ Tile_X0Y0_FrameData[20] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_79_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_39 Tile_X0Y1_N4END[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_17 Tile_X0Y1_N2END[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_28 Tile_X0Y1_N2MID[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0885_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_30_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0954_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput102 net102 Tile_X0Y0_N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput135 net135 Tile_X0Y0_W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput146 net146 Tile_X0Y0_WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput157 net157 Tile_X0Y0_WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput179 net179 Tile_X0Y1_FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput124 net124 Tile_X0Y0_W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput168 net168 Tile_X0Y1_FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput113 net113 Tile_X0Y0_W1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0319_ Tile_X0Y0_E2MID[2] Tile_X0Y0_E2END[2] Tile_X0Y0_E6END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1299_ Tile_X0Y1_FrameData[12] net161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1368_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1 net239 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0670_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_12_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1222_ Tile_X0Y1_N4END[8] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_119_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1153_ Tile_X0Y0_FrameData[3] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1084_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_142_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0799_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0868_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0937_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_87_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_81_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0653_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0722_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_6_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0584_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 _0205_ _0072_
+ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ _0106_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1205_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3 net76 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1067_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1136_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_138_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_92_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0636_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0705_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_115_Right_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0567_ Tile_X0Y1_E1END[1] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[1] _0078_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q _0095_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0498_ Q_SRAM0 Q_SRAM3 _0165_ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1119_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_17_Right_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_119_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Right_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_105_Left_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0352_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0421_ Tile_X0Y0_E2END[3] _0152_ _0037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0283_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 _0202_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_79_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Right_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Right_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_114_Left_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_123_Left_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_62_Right_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0619_ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[9] Tile_X0Y1_EE4END[13]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0134_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_132_Left_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Right_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_141_Left_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_80_Right_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0970_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0404_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0266_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1 Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0335_ Tile_X0Y1_N1END[0] Tile_X0Y1_N4END[0] _0011_ Tile_X0Y0_S4END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q _0012_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1384_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9 net257 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_29 Tile_X0Y1_N2MID[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_18 Tile_X0Y1_N2END[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput103 net103 Tile_X0Y0_N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0884_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput125 net125 Tile_X0Y0_W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput114 net114 Tile_X0Y0_W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0953_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput136 net136 Tile_X0Y0_W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput147 net147 Tile_X0Y0_WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput169 net169 Tile_X0Y1_FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput158 net158 Tile_X0Y1_FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1367_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0 net238 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0318_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5 Tile_X0Y0_S2MID[5]
+ Tile_X0Y1_N2MID[5] Tile_X0Y0_S2END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1298_ Tile_X0Y1_FrameData[11] net160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0249_ _0141_ Tile_X0Y1_E2END[5] _0175_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1221_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7 net92 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1152_ Tile_X0Y0_FrameData[2] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1083_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_142_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0936_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0867_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0798_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_3_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_129_Right_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0721_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0652_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0583_ _0105_ _0104_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1204_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2 net75 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1066_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1135_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0919_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_140_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Left_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0635_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0704_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0566_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 _0185_ _0074_
+ _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ _0094_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_36_Left_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_57_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0497_ Q_SRAM1 _0000_ Q_SRAM2 _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1049_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1118_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_135_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0420_ Tile_X0Y0_E2MID[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q _0036_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0351_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0282_ _0147_ Tile_X0Y0_S1END[3] _0201_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0549_ Tile_X0Y1_E2END[0] _0160_ _0082_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0618_ Tile_X0Y1_E6END[1] _0078_ Tile_X0Y1_E6END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ _0133_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0403_ Q_SRAM4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1383_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8 net256 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0334_ Tile_X0Y0_E1END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_E6END[8] _0010_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q _0011_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0265_ Tile_X0Y1_E1END[1] _0185_ Tile_X0Y1_E6END[5] _0189_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_19 Tile_X0Y1_N2END[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0952_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput104 net104 Tile_X0Y0_N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0883_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput137 net137 Tile_X0Y0_W6BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput148 net148 Tile_X0Y0_WW4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput126 net126 Tile_X0Y0_W2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput115 net115 Tile_X0Y0_W2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput159 net159 Tile_X0Y1_FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1366_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7 net237 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0317_ Tile_X0Y1_E2MID[2] Tile_X0Y1_E6END[2] Tile_X0Y1_E2END[2] _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1297_ Tile_X0Y1_FrameData[10] net159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0248_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0 _0168_ _0173_
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ _0174_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_38_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1220_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6 net91 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1151_ Tile_X0Y0_FrameData[1] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1082_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_35_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0866_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0935_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0797_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1349_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2 net211 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0720_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_111_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0651_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0582_ Tile_X0Y1_E1END[2] Tile_X0Y1_EE4END[14] Tile_X0Y1_E6END[6] _0077_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q _0105_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_6_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1203_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1 net74 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_95_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1134_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_122_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1065_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_33_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0849_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0918_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_75_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0703_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0634_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0496_ Q_SRAM1 _0001_ Q_SRAM2 _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0565_ _0093_ _0092_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1117_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_110_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1048_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0350_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0281_ Tile_X0Y0_E6END[3] _0147_ _0200_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0617_ _0132_ _0131_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0548_ Tile_X0Y1_E2MID[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
+ _0081_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0479_ Tile_X0Y1_E2MID[7] Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[8] _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_55_Left_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0333_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q _0008_
+ _0009_ _0007_ _0010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_0402_ Q_SRAM4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 _0025_
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1382_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7 net255 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0264_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q _0187_
+ _0188_ _0186_ _0189_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_63_Left_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Left_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0882_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_15_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0951_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput105 net105 Tile_X0Y0_N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput138 net138 Tile_X0Y0_W6BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput149 net149 Tile_X0Y0_WW4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput127 net127 Tile_X0Y0_W2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_81_Left_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput116 net116 Tile_X0Y0_W2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1296_ Tile_X0Y1_FrameData[9] net189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1365_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6 net236 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0316_ Tile_X0Y1_N2MID[5] Tile_X0Y1_N2END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q _0004_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_38_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0247_ Tile_X0Y1_E2END[4] Tile_X0Y0_S2MID[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ _0173_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_129_Left_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_84_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_Left_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1150_ Tile_X0Y0_FrameData[0] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1081_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_60_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0865_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0934_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_20_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_143_Right_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_114_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0796_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1348_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1 net225 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1279_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8 net156 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_110_Right_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0650_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0581_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 _0195_ _0073_
+ _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ _0104_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1202_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0 net73 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1064_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1133_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_122_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0848_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_108_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0779_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0917_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_24_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0633_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0702_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_97_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0495_ Q_SRAM0 Q_SRAM3 _0002_ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0564_ Tile_X0Y1_E1END[0] Tile_X0Y1_E6END[8] Tile_X0Y1_EE4END[0] _0079_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q _0093_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1116_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1047_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0280_ Tile_X0Y0_E1END[2] Tile_X0Y0_E6END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0193_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_79_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_22_Right_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_116_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0616_ Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[8] Tile_X0Y1_EE4END[12]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0132_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0478_ Tile_X0Y1_E1END[3] Tile_X0Y1_E6END[11] _0205_ _0209_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0547_ _0160_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ _0165_ _0080_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_31_Right_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_101_Left_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_110_Left_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0332_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 _0009_ VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0401_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 _0024_
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0263_ Tile_X0Y1_N1END[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q _0188_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1381_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6 net254 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0881_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_124_Right_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0950_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_141_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput106 net106 Tile_X0Y0_N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput139 net139 Tile_X0Y0_W6BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput128 net128 Tile_X0Y0_W2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput117 net117 Tile_X0Y0_W2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0315_ Tile_X0Y0_E1END[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1295_ Tile_X0Y1_FrameData[8] net188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1364_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5 net235 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0246_ _0141_ _0166_ _0168_ _0169_ _0171_ _0172_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_38_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0864_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0795_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0933_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1347_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0 net224 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_98_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1278_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7 net155 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0229_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q _0158_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_Right_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1201_ Tile_X0Y1_FrameStrobe[19] net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_69_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0580_ _0102_ _0103_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_87_Right_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1063_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_25_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1132_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0916_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0847_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_96_Right_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0778_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_124_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0632_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_128_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0701_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0563_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 _0012_ _0075_
+ _0165_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ _0092_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0494_ Q_SRAM0 Q_SRAM3 _0002_ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1115_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1046_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_21_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0546_ Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 _0079_
+ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0615_ Tile_X0Y1_E6END[0] _0079_ Tile_X0Y1_E6END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0131_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0477_ Tile_X0Y1_E1END[2] Tile_X0Y1_E6END[10] _0195_ _0199_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_138_Right_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1029_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_105_Right_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0400_ Q_SRAM6 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6 _0023_
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1380_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5 net253 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0331_ Tile_X0Y0_S1END[0] _0155_ _0008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0262_ _0157_ _0184_ _0187_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0529_ Tile_X0Y1_N1END[2] Tile_X0Y1_N4END[2] _0194_ Tile_X0Y0_S4END[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q _0077_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_87_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0880_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xoutput107 net107 Tile_X0Y0_N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput129 net129 Tile_X0Y0_W2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput118 net118 Tile_X0Y0_W2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1363_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4 net234 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0314_ Tile_X0Y0_E2MID[3] Tile_X0Y0_E2END[3] Tile_X0Y0_E6END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1294_ Tile_X0Y1_FrameData[7] net187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0245_ _0139_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ _0170_ _0171_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0932_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0863_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0794_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_54_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1346_ Tile_X0Y0_S4END[15] net223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1277_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6 net154 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0228_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q _0157_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1200_ Tile_X0Y1_FrameStrobe[18] net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_69_Left_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1062_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_18_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1131_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_78_Left_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0915_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0846_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0777_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_124_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_83_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1329_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6 net200 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_96_Left_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_83_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0700_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0631_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0562_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q _0090_
+ _0091_ _0089_ net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_119_Right_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1114_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_17_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0493_ Q_SRAM1 _0001_ Q_SRAM2 _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1045_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_134_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0829_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0476_ Tile_X0Y1_E1END[1] Tile_X0Y1_E6END[9] _0185_ _0189_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0545_ Q_SRAM2 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 _0078_
+ _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0614_ _0130_ _0129_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ net277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1028_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_15_Left_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_91_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_24_Left_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0330_ Tile_X0Y0_E6END[0] _0155_ _0007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0261_ Tile_X0Y1_E6END[1] _0157_ _0186_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_84_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0459_ Tile_X0Y0_E6END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_E6END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ _0062_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0528_ Q_SRAM0 Q_SRAM3 _0076_ _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput108 net108 Tile_X0Y0_N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput119 net119 Tile_X0Y0_W2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput90 net90 Tile_X0Y0_N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0313_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4 Tile_X0Y0_S2MID[4]
+ Tile_X0Y1_N2MID[4] Tile_X0Y0_S2END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1293_ Tile_X0Y1_FrameData[6] net186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1362_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3 net233 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0244_ Tile_X0Y1_N2END[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ _0170_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_31_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Left_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_116_Left_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0862_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_102_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0931_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_43_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0793_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_47_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1345_ Tile_X0Y0_S4END[14] net222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_98_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1276_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5 net153 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0227_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q _0156_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1130_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1061_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_31_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0845_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0914_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0776_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1259_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0 net130 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1328_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5 net199 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput280 net280 WEN_SRAM6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0630_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0492_ Q_SRAM1 _0000_ Q_SRAM2 _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0561_ Tile_X0Y1_E2END[3] _0163_ _0091_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_91_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1113_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1044_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0759_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0828_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_88_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0613_ Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[11] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
+ _0130_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0475_ Tile_X0Y1_E1END[0] Tile_X0Y1_E6END[8] _0012_ _0017_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0544_ Q_SRAM1 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 _0077_
+ _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1027_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_38_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0260_ Tile_X0Y1_N1END[1] Tile_X0Y1_N4END[1] _0184_ Tile_X0Y0_S4END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q _0185_ VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0389_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2 Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0458_ _0061_ _0060_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
+ net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0527_ Tile_X0Y1_N1END[3] Tile_X0Y1_N4END[3] _0204_ Tile_X0Y0_S4END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q _0076_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput109 net109 Tile_X0Y0_UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput1 net1 A_SRAM0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput80 net80 Tile_X0Y0_N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput91 net91 Tile_X0Y0_N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1292_ Tile_X0Y1_FrameData[5] net185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1361_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2 net232 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0243_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q _0140_
+ _0167_ _0169_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0312_ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2END[3] Tile_X0Y1_E6END[3] _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0861_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0792_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0930_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_13_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1344_ Tile_X0Y0_S4END[13] net221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0226_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q _0155_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1275_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4 net152 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_29_Right_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_47_Right_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_Right_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0844_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0775_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0913_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_124_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Right_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1189_ Tile_X0Y1_FrameStrobe[7] net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1258_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7 net129 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1327_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4 net198 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_135_Left_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_74_Right_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput270 net270 Tile_X0Y1_WW4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput281 net281 WEN_SRAM7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_133_Right_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_92_Right_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0491_ Q_SRAM0 Q_SRAM3 _0165_ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0560_ Tile_X0Y1_E2MID[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
+ _0090_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_91_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1043_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1112_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_100_Right_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0827_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0758_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0689_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_56_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0612_ Tile_X0Y1_E6END[3] _0076_ Tile_X0Y1_E6END[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ _0129_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0474_ Tile_X0Y0_E1END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_E6END[4] _0010_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0543_ Q_SRAM0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7 _0076_
+ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1026_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_139_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0526_ Q_SRAM0 Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ _0003_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0457_ Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[14]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ _0061_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0388_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1009_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_135_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput70 net70 Tile_X0Y0_FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1360_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1 net231 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput2 net2 A_SRAM1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput92 net92 Tile_X0Y0_N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput81 net81 Tile_X0Y0_N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1291_ Tile_X0Y1_FrameData[4] net184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0311_ Tile_X0Y1_N2MID[4] Tile_X0Y1_N2END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q _0003_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0242_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q _0141_
+ _0168_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0509_ Q_SRAM1 _0185_ Q_SRAM2 _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0791_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0860_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_11_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1343_ Tile_X0Y0_S4END[12] net220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_39_Left_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1274_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3 net151 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0225_ Tile_X0Y1_E6END[4] _0154_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_48_Left_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0989_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_114_Right_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0912_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0843_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0774_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_52_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1326_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3 net197 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1188_ Tile_X0Y1_FrameStrobe[6] net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1257_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6 net128 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_56_Left_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput271 net271 Tile_X0Y1_WW4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput260 net260 Tile_X0Y1_WW4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0490_ Tile_X0Y1_N1END[3] Q_SRAM1 _0204_ Q_SRAM3 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_91_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1042_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1111_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_142_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0688_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0757_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0826_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1309_ Tile_X0Y1_FrameData[22] net172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0611_ _0128_ _0127_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
+ net276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0542_ Q_SRAM0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4 _0075_
+ _0002_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0473_ _0071_ _0070_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ net281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1025_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0809_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_29_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_1 Tile_X0Y0_S2END[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0456_ Tile_X0Y0_E6END[2] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_E6END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
+ _0060_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0525_ Tile_X0Y1_N1END[0] Tile_X0Y1_N4END[0] _0011_ Tile_X0Y0_S4END[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_20_Left_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0387_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3 Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1008_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_106_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net93 Tile_X0Y0_N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput71 net71 Tile_X0Y0_FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput60 net60 Tile_X0Y0_FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput82 net82 Tile_X0Y0_N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_128_Right_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0310_ Tile_X0Y0_E1END[0] Tile_X0Y0_E2END[3] Tile_X0Y0_E2MID[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput3 net3 A_SRAM2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1290_ Tile_X0Y1_FrameData[3] net183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0241_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_E2MID[0]
+ _0167_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0439_ Tile_X0Y0_E1END[0] Tile_X0Y0_EE4END[12] Tile_X0Y0_E6END[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ _0049_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0508_ Q_SRAM1 _0195_ Q_SRAM2 _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_142_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0790_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_11_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1342_ Tile_X0Y0_S4END[11] net219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1273_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2 net150 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0224_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q _0153_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0988_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_113_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0842_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_71_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0911_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0773_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_45_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1256_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5 net127 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1325_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2 net196 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_3_Left_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_1187_ Tile_X0Y1_FrameStrobe[5] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput261 net261 Tile_X0Y1_WW4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput272 net272 Tile_X0Y1_WW4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput250 net250 Tile_X0Y1_W6BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1110_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_80_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1041_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_119_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0825_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0687_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0756_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1308_ Tile_X0Y1_FrameData[21] net171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1239_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0 net110 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0472_ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
+ _0071_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_109_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_Left_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0610_ Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[14]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ _0128_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0541_ Q_SRAM1 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 _0074_
+ _0001_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1024_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_93_Left_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0808_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_130_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0739_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_76_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Right_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_2 Tile_X0Y0_S2MID[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0455_ _0059_ _0058_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0524_ Q_SRAM1 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5 Q_SRAM2
+ _0004_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_108_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0386_ Q_SRAM4 Q_SRAM7 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1007_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_9_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput72 net72 Tile_X0Y0_FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput94 net94 Tile_X0Y0_N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput61 net61 Tile_X0Y0_FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput83 net83 Tile_X0Y0_N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput50 net50 Tile_X0Y0_FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput4 net4 A_SRAM3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0240_ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2]
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ _0166_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0438_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ _0025_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q _0048_ VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0369_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_69_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0507_ Q_SRAM0 Q_SRAM3 _0205_ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_37_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_142_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1341_ Tile_X0Y0_S4END[10] net218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0223_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q _0152_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1272_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1 net149 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0987_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_120_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_80_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_130_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0841_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0772_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0910_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_25_Right_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1186_ Tile_X0Y1_FrameStrobe[4] net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_94_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1255_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4 net126 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1324_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1 net195 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_34_Right_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_121_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_104_Left_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_Right_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput262 net262 Tile_X0Y1_WW4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput240 net240 Tile_X0Y1_W2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput273 net273 Tile_X0Y1_WW4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput251 net251 Tile_X0Y1_W6BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_113_Left_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_122_Left_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Right_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_131_Left_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_65_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1040_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_0_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_140_Left_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0824_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0755_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0686_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1238_ clknet_1_1__leaf_Tile_X0Y1_UserCLK net109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1169_ Tile_X0Y0_FrameData[19] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1307_ Tile_X0Y1_FrameData[20] net170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0471_ Tile_X0Y0_E6END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_E6END[7] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ _0070_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0540_ Q_SRAM2 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 _0073_
+ _0000_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1023_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0738_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0807_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0669_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_84_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_3 Tile_X0Y0_S2MID[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0454_ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[9] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
+ _0059_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0385_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0 Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0523_ Tile_X0Y1_N1END[1] Tile_X0Y1_N4END[1] _0184_ Tile_X0Y0_S4END[5] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1006_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_34_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_142_Right_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput5 net5 A_SRAM4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput95 net95 Tile_X0Y0_N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput62 net62 Tile_X0Y0_FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput73 net73 Tile_X0Y0_N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput40 net40 Tile_X0Y0_FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput84 net84 Tile_X0Y0_N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput51 net51 Tile_X0Y0_FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_46_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_Right_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_68_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0506_ Q_SRAM0 Q_SRAM3 _0165_ _0006_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0437_ _0047_ _0046_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0368_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_0299_ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1340_ Tile_X0Y0_S4END[9] net217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0222_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q _0151_
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1271_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0 net142 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_133_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_74_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Left_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0986_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_113_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0840_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0771_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_1323_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0 net194 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1185_ Tile_X0Y1_FrameStrobe[3] net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_94_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1254_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3 net125 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput241 net241 Tile_X0Y1_W2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput230 net230 Tile_X0Y1_W2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput252 net252 Tile_X0Y1_W6BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0969_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_114_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput263 net263 Tile_X0Y1_WW4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput274 net274 WEN_SRAM0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0823_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0685_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0754_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_50_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1306_ Tile_X0Y1_FrameData[19] net168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1237_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3 net99 VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1168_ Tile_X0Y0_FrameData[18] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1099_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_109_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0470_ _0069_ _0068_ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
+ net280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1022_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XPHY_EDGE_ROW_123_Right_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_0737_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0668_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0806_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_0599_ _0164_ _0115_ _0119_ _0120_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_9_Left_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_4 Tile_X0Y0_S2MID[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_0522_ Q_SRAM1 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6 Q_SRAM2
+ _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0453_ Tile_X0Y0_E6END[1] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_E6END[5] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ _0058_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0384_ Q_SRAM5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5 Q_SRAM6
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_1005_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_135_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput41 net41 Tile_X0Y0_FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput30 net30 Tile_X0Y0_FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput52 net52 Tile_X0Y0_FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput6 net6 A_SRAM5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput63 net63 Tile_X0Y0_FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput96 net96 Tile_X0Y0_N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput85 net85 Tile_X0Y0_N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput74 net74 Tile_X0Y0_N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0436_ Tile_X0Y0_E1END[3] Tile_X0Y0_E6END[11] Tile_X0Y0_EE4END[3] Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
+ _0047_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0505_ Q_SRAM1 _0000_ Q_SRAM2 _0005_ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
.ends

