magic
tech gf180mcuD
magscale 1 10
timestamp 1764971299
<< metal1 >>
rect 672 13354 52080 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 52080 13354
rect 672 13268 52080 13302
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 17390 13186 17442 13198
rect 17390 13122 17442 13134
rect 21198 13186 21250 13198
rect 37774 13186 37826 13198
rect 35746 13134 35758 13186
rect 35810 13134 35822 13186
rect 21198 13122 21250 13134
rect 37774 13122 37826 13134
rect 37998 13186 38050 13198
rect 37998 13122 38050 13134
rect 41246 13186 41298 13198
rect 41246 13122 41298 13134
rect 45054 13186 45106 13198
rect 45054 13122 45106 13134
rect 6526 13074 6578 13086
rect 13346 13022 13358 13074
rect 13410 13022 13422 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 15698 13022 15710 13074
rect 15762 13022 15774 13074
rect 22866 13022 22878 13074
rect 22930 13022 22942 13074
rect 25218 13022 25230 13074
rect 25282 13022 25294 13074
rect 40674 13022 40686 13074
rect 40738 13022 40750 13074
rect 43698 13022 43710 13074
rect 43762 13022 43774 13074
rect 6526 13010 6578 13022
rect 35422 12962 35474 12974
rect 42254 12962 42306 12974
rect 50766 12962 50818 12974
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 14130 12910 14142 12962
rect 14194 12910 14206 12962
rect 17938 12910 17950 12962
rect 18002 12910 18014 12962
rect 18386 12910 18398 12962
rect 18450 12910 18462 12962
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 37314 12910 37326 12962
rect 37378 12910 37390 12962
rect 39106 12910 39118 12962
rect 39170 12910 39182 12962
rect 42914 12910 42926 12962
rect 42978 12910 42990 12962
rect 44482 12910 44494 12962
rect 44546 12910 44558 12962
rect 47170 12910 47182 12962
rect 47234 12910 47246 12962
rect 48962 12910 48974 12962
rect 49026 12910 49038 12962
rect 35422 12898 35474 12910
rect 42254 12898 42306 12910
rect 50766 12898 50818 12910
rect 36318 12850 36370 12862
rect 19170 12798 19182 12850
rect 19234 12798 19246 12850
rect 36318 12786 36370 12798
rect 38558 12850 38610 12862
rect 50430 12850 50482 12862
rect 40002 12798 40014 12850
rect 40066 12798 40078 12850
rect 51202 12798 51214 12850
rect 51266 12798 51278 12850
rect 38558 12786 38610 12798
rect 50430 12786 50482 12798
rect 24222 12738 24274 12750
rect 24222 12674 24274 12686
rect 48190 12738 48242 12750
rect 48190 12674 48242 12686
rect 49758 12738 49810 12750
rect 49758 12674 49810 12686
rect 672 12570 52080 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 52080 12570
rect 672 12484 52080 12518
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 18286 12402 18338 12414
rect 18286 12338 18338 12350
rect 21646 12402 21698 12414
rect 21646 12338 21698 12350
rect 22878 12402 22930 12414
rect 22878 12338 22930 12350
rect 36542 12402 36594 12414
rect 36542 12338 36594 12350
rect 38110 12402 38162 12414
rect 38110 12338 38162 12350
rect 40014 12402 40066 12414
rect 40014 12338 40066 12350
rect 41582 12402 41634 12414
rect 41582 12338 41634 12350
rect 48078 12402 48130 12414
rect 48078 12338 48130 12350
rect 14814 12290 14866 12302
rect 26350 12290 26402 12302
rect 28030 12290 28082 12302
rect 49646 12290 49698 12302
rect 6850 12238 6862 12290
rect 6914 12238 6926 12290
rect 7746 12238 7758 12290
rect 7810 12238 7822 12290
rect 9986 12238 9998 12290
rect 10050 12238 10062 12290
rect 19618 12238 19630 12290
rect 19682 12238 19694 12290
rect 27122 12238 27134 12290
rect 27186 12238 27198 12290
rect 28914 12238 28926 12290
rect 28978 12238 28990 12290
rect 14814 12226 14866 12238
rect 26350 12226 26402 12238
rect 28030 12226 28082 12238
rect 49646 12226 49698 12238
rect 51214 12290 51266 12302
rect 51214 12226 51266 12238
rect 6302 12178 6354 12190
rect 26686 12178 26738 12190
rect 15362 12126 15374 12178
rect 15426 12126 15438 12178
rect 15810 12126 15822 12178
rect 15874 12126 15886 12178
rect 17266 12126 17278 12178
rect 17330 12126 17342 12178
rect 20850 12126 20862 12178
rect 20914 12126 20926 12178
rect 23202 12126 23214 12178
rect 23266 12126 23278 12178
rect 6302 12114 6354 12126
rect 26686 12114 26738 12126
rect 28478 12178 28530 12190
rect 42590 12178 42642 12190
rect 39442 12126 39454 12178
rect 39506 12126 39518 12178
rect 41234 12126 41246 12178
rect 41298 12126 41310 12178
rect 48738 12126 48750 12178
rect 48802 12126 48814 12178
rect 28478 12114 28530 12126
rect 42590 12114 42642 12126
rect 2606 12066 2658 12078
rect 2606 12002 2658 12014
rect 5742 12066 5794 12078
rect 12798 12066 12850 12078
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 12226 12014 12238 12066
rect 12290 12014 12302 12066
rect 5742 12002 5794 12014
rect 12798 12002 12850 12014
rect 13358 12066 13410 12078
rect 29934 12066 29986 12078
rect 18834 12014 18846 12066
rect 18898 12014 18910 12066
rect 23762 12014 23774 12066
rect 23826 12014 23838 12066
rect 13358 12002 13410 12014
rect 29934 12002 29986 12014
rect 31166 12066 31218 12078
rect 43150 12066 43202 12078
rect 37538 12014 37550 12066
rect 37602 12014 37614 12066
rect 39106 12014 39118 12066
rect 39170 12014 39182 12066
rect 47058 12014 47070 12066
rect 47122 12014 47134 12066
rect 50194 12014 50206 12066
rect 50258 12014 50270 12066
rect 31166 12002 31218 12014
rect 43150 12002 43202 12014
rect 3166 11954 3218 11966
rect 3166 11890 3218 11902
rect 3502 11954 3554 11966
rect 3502 11890 3554 11902
rect 7310 11954 7362 11966
rect 7310 11890 7362 11902
rect 8206 11954 8258 11966
rect 8206 11890 8258 11902
rect 8542 11954 8594 11966
rect 8542 11890 8594 11902
rect 13694 11954 13746 11966
rect 13694 11890 13746 11902
rect 24334 11954 24386 11966
rect 24334 11890 24386 11902
rect 29374 11954 29426 11966
rect 29374 11890 29426 11902
rect 30382 11954 30434 11966
rect 30382 11890 30434 11902
rect 30606 11954 30658 11966
rect 30606 11890 30658 11902
rect 672 11786 52080 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 52080 11786
rect 672 11700 52080 11734
rect 7086 11618 7138 11630
rect 7086 11554 7138 11566
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 12462 11618 12514 11630
rect 12462 11554 12514 11566
rect 14030 11618 14082 11630
rect 14030 11554 14082 11566
rect 23326 11618 23378 11630
rect 23326 11554 23378 11566
rect 26910 11618 26962 11630
rect 26910 11554 26962 11566
rect 38670 11618 38722 11630
rect 38670 11554 38722 11566
rect 40798 11618 40850 11630
rect 40798 11554 40850 11566
rect 42366 11618 42418 11630
rect 42366 11554 42418 11566
rect 5294 11506 5346 11518
rect 5294 11442 5346 11454
rect 6750 11506 6802 11518
rect 18834 11454 18846 11506
rect 18898 11454 18910 11506
rect 21970 11454 21982 11506
rect 22034 11454 22046 11506
rect 50418 11454 50430 11506
rect 50482 11454 50494 11506
rect 6750 11442 6802 11454
rect 5854 11394 5906 11406
rect 17166 11394 17218 11406
rect 25118 11394 25170 11406
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 13010 11342 13022 11394
rect 13074 11342 13086 11394
rect 14578 11342 14590 11394
rect 14642 11342 14654 11394
rect 16146 11342 16158 11394
rect 16210 11342 16222 11394
rect 18050 11342 18062 11394
rect 18114 11342 18126 11394
rect 19730 11342 19742 11394
rect 19794 11342 19806 11394
rect 21186 11342 21198 11394
rect 21250 11342 21262 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 5854 11330 5906 11342
rect 17166 11330 17218 11342
rect 25118 11330 25170 11342
rect 27918 11394 27970 11406
rect 37762 11342 37774 11394
rect 37826 11342 37838 11394
rect 38098 11342 38110 11394
rect 38162 11342 38174 11394
rect 40450 11342 40462 11394
rect 40514 11342 40526 11394
rect 41794 11342 41806 11394
rect 41858 11342 41870 11394
rect 48850 11342 48862 11394
rect 48914 11342 48926 11394
rect 27918 11330 27970 11342
rect 7646 11282 7698 11294
rect 16830 11282 16882 11294
rect 6290 11230 6302 11282
rect 6354 11230 6366 11282
rect 15474 11230 15486 11282
rect 15538 11230 15550 11282
rect 7646 11218 7698 11230
rect 16830 11218 16882 11230
rect 17726 11282 17778 11294
rect 17726 11218 17778 11230
rect 20190 11282 20242 11294
rect 25342 11282 25394 11294
rect 24658 11230 24670 11282
rect 24722 11230 24734 11282
rect 20190 11218 20242 11230
rect 25342 11218 25394 11230
rect 27582 11282 27634 11294
rect 27582 11218 27634 11230
rect 28478 11282 28530 11294
rect 28478 11218 28530 11230
rect 29038 11282 29090 11294
rect 29038 11218 29090 11230
rect 36766 11282 36818 11294
rect 36766 11218 36818 11230
rect 49870 11282 49922 11294
rect 49870 11218 49922 11230
rect 51438 11170 51490 11182
rect 51438 11106 51490 11118
rect 672 11002 52080 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 52080 11002
rect 672 10916 52080 10950
rect 10446 10834 10498 10846
rect 10446 10770 10498 10782
rect 11678 10834 11730 10846
rect 11678 10770 11730 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 18286 10834 18338 10846
rect 18286 10770 18338 10782
rect 19854 10834 19906 10846
rect 19854 10770 19906 10782
rect 21870 10834 21922 10846
rect 21870 10770 21922 10782
rect 23438 10834 23490 10846
rect 23438 10770 23490 10782
rect 37774 10834 37826 10846
rect 37774 10770 37826 10782
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 40910 10834 40962 10846
rect 40910 10770 40962 10782
rect 42478 10834 42530 10846
rect 42478 10770 42530 10782
rect 49646 10722 49698 10734
rect 1698 10670 1710 10722
rect 1762 10670 1774 10722
rect 14690 10670 14702 10722
rect 14754 10670 14766 10722
rect 26786 10670 26798 10722
rect 26850 10670 26862 10722
rect 49646 10658 49698 10670
rect 27246 10610 27298 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 16930 10558 16942 10610
rect 16994 10558 17006 10610
rect 18834 10558 18846 10610
rect 18898 10558 18910 10610
rect 22866 10558 22878 10610
rect 22930 10558 22942 10610
rect 38770 10558 38782 10610
rect 38834 10558 38846 10610
rect 40562 10558 40574 10610
rect 40626 10558 40638 10610
rect 42018 10558 42030 10610
rect 42082 10558 42094 10610
rect 48738 10558 48750 10610
rect 48802 10558 48814 10610
rect 27246 10546 27298 10558
rect 27806 10498 27858 10510
rect 47518 10498 47570 10510
rect 12226 10446 12238 10498
rect 12290 10446 12302 10498
rect 15362 10446 15374 10498
rect 15426 10446 15438 10498
rect 17266 10446 17278 10498
rect 17330 10446 17342 10498
rect 21298 10446 21310 10498
rect 21362 10446 21374 10498
rect 37202 10446 37214 10498
rect 37266 10446 37278 10498
rect 27806 10434 27858 10446
rect 47518 10434 47570 10446
rect 47742 10498 47794 10510
rect 47742 10434 47794 10446
rect 48302 10498 48354 10510
rect 50194 10446 50206 10498
rect 50258 10446 50270 10498
rect 50978 10446 50990 10498
rect 51042 10446 51054 10498
rect 48302 10434 48354 10446
rect 2158 10386 2210 10398
rect 2158 10322 2210 10334
rect 2494 10386 2546 10398
rect 2494 10322 2546 10334
rect 6078 10386 6130 10398
rect 6078 10322 6130 10334
rect 26126 10386 26178 10398
rect 26126 10322 26178 10334
rect 26350 10386 26402 10398
rect 26350 10322 26402 10334
rect 672 10218 52080 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 52080 10218
rect 672 10132 52080 10166
rect 10446 10050 10498 10062
rect 10446 9986 10498 9998
rect 10670 10050 10722 10062
rect 10670 9986 10722 9998
rect 12462 10050 12514 10062
rect 12462 9986 12514 9998
rect 14030 10050 14082 10062
rect 14030 9986 14082 9998
rect 15598 10050 15650 10062
rect 15598 9986 15650 9998
rect 19294 10050 19346 10062
rect 19294 9986 19346 9998
rect 20862 10050 20914 10062
rect 20862 9986 20914 9998
rect 22318 10050 22370 10062
rect 22318 9986 22370 9998
rect 27358 10050 27410 10062
rect 27358 9986 27410 9998
rect 34190 10050 34242 10062
rect 34190 9986 34242 9998
rect 38894 10050 38946 10062
rect 38894 9986 38946 9998
rect 40798 10050 40850 10062
rect 40798 9986 40850 9998
rect 41806 10050 41858 10062
rect 41806 9986 41858 9998
rect 24558 9938 24610 9950
rect 27682 9886 27694 9938
rect 27746 9886 27758 9938
rect 50418 9886 50430 9938
rect 50482 9886 50494 9938
rect 24558 9874 24610 9886
rect 9438 9826 9490 9838
rect 25118 9826 25170 9838
rect 12786 9774 12798 9826
rect 12850 9774 12862 9826
rect 14578 9774 14590 9826
rect 14642 9774 14654 9826
rect 16146 9774 16158 9826
rect 16210 9774 16222 9826
rect 17042 9774 17054 9826
rect 17106 9774 17118 9826
rect 19842 9774 19854 9826
rect 19906 9774 19918 9826
rect 21410 9774 21422 9826
rect 21474 9774 21486 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 9438 9762 9490 9774
rect 25118 9762 25170 9774
rect 26798 9826 26850 9838
rect 26798 9762 26850 9774
rect 27134 9826 27186 9838
rect 36206 9826 36258 9838
rect 43934 9826 43986 9838
rect 34626 9774 34638 9826
rect 34690 9774 34702 9826
rect 38322 9774 38334 9826
rect 38386 9774 38398 9826
rect 40338 9774 40350 9826
rect 40402 9774 40414 9826
rect 27134 9762 27186 9774
rect 36206 9762 36258 9774
rect 43934 9762 43986 9774
rect 44830 9826 44882 9838
rect 48850 9774 48862 9826
rect 48914 9774 48926 9826
rect 44830 9762 44882 9774
rect 9774 9714 9826 9726
rect 8978 9662 8990 9714
rect 9042 9662 9054 9714
rect 9774 9650 9826 9662
rect 11230 9714 11282 9726
rect 11230 9650 11282 9662
rect 18062 9714 18114 9726
rect 18062 9650 18114 9662
rect 25454 9714 25506 9726
rect 35086 9714 35138 9726
rect 26338 9662 26350 9714
rect 26402 9662 26414 9714
rect 25454 9650 25506 9662
rect 35086 9650 35138 9662
rect 35870 9714 35922 9726
rect 35870 9650 35922 9662
rect 36766 9714 36818 9726
rect 43598 9714 43650 9726
rect 42242 9662 42254 9714
rect 42306 9662 42318 9714
rect 36766 9650 36818 9662
rect 43598 9650 43650 9662
rect 44494 9714 44546 9726
rect 49870 9714 49922 9726
rect 45266 9662 45278 9714
rect 45330 9662 45342 9714
rect 44494 9650 44546 9662
rect 49870 9650 49922 9662
rect 51438 9602 51490 9614
rect 51438 9538 51490 9550
rect 672 9434 52080 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 52080 9434
rect 672 9348 52080 9382
rect 14814 9266 14866 9278
rect 14814 9202 14866 9214
rect 16382 9266 16434 9278
rect 16382 9202 16434 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 20862 9266 20914 9278
rect 20862 9202 20914 9214
rect 40910 9266 40962 9278
rect 40910 9202 40962 9214
rect 49646 9266 49698 9278
rect 49646 9202 49698 9214
rect 22990 9154 23042 9166
rect 8530 9102 8542 9154
rect 8594 9102 8606 9154
rect 11554 9102 11566 9154
rect 11618 9102 11630 9154
rect 17938 9102 17950 9154
rect 18002 9102 18014 9154
rect 22990 9090 23042 9102
rect 25790 9154 25842 9166
rect 25790 9090 25842 9102
rect 27022 9154 27074 9166
rect 27022 9090 27074 9102
rect 38222 9154 38274 9166
rect 38222 9090 38274 9102
rect 41582 9154 41634 9166
rect 41582 9090 41634 9102
rect 44494 9154 44546 9166
rect 44494 9090 44546 9102
rect 22766 9042 22818 9054
rect 21746 8990 21758 9042
rect 21810 8990 21822 9042
rect 22766 8978 22818 8990
rect 23774 9042 23826 9054
rect 23774 8978 23826 8990
rect 24334 9042 24386 9054
rect 24334 8978 24386 8990
rect 38558 9042 38610 9054
rect 48738 8990 48750 9042
rect 48802 8990 48814 9042
rect 38558 8978 38610 8990
rect 13806 8930 13858 8942
rect 22206 8930 22258 8942
rect 12226 8878 12238 8930
rect 12290 8878 12302 8930
rect 15362 8878 15374 8930
rect 15426 8878 15438 8930
rect 16930 8878 16942 8930
rect 16994 8878 17006 8930
rect 17266 8878 17278 8930
rect 17330 8878 17342 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 13806 8866 13858 8878
rect 22206 8866 22258 8878
rect 24894 8930 24946 8942
rect 24894 8866 24946 8878
rect 25230 8930 25282 8942
rect 25230 8866 25282 8878
rect 39118 8930 39170 8942
rect 48302 8930 48354 8942
rect 39890 8878 39902 8930
rect 39954 8878 39966 8930
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 50978 8878 50990 8930
rect 51042 8878 51054 8930
rect 39118 8866 39170 8878
rect 48302 8866 48354 8878
rect 8990 8818 9042 8830
rect 8990 8754 9042 8766
rect 9214 8818 9266 8830
rect 9214 8754 9266 8766
rect 13022 8818 13074 8830
rect 13022 8754 13074 8766
rect 13246 8818 13298 8830
rect 13246 8754 13298 8766
rect 23998 8818 24050 8830
rect 23998 8754 24050 8766
rect 47518 8818 47570 8830
rect 47518 8754 47570 8766
rect 47742 8818 47794 8830
rect 47742 8754 47794 8766
rect 672 8650 52080 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 52080 8650
rect 672 8564 52080 8598
rect 22430 8482 22482 8494
rect 22430 8418 22482 8430
rect 9326 8370 9378 8382
rect 20974 8370 21026 8382
rect 19394 8318 19406 8370
rect 19458 8318 19470 8370
rect 9326 8306 9378 8318
rect 20974 8306 21026 8318
rect 29374 8370 29426 8382
rect 29374 8306 29426 8318
rect 49198 8370 49250 8382
rect 49198 8306 49250 8318
rect 9886 8258 9938 8270
rect 9886 8194 9938 8206
rect 10222 8258 10274 8270
rect 21534 8258 21586 8270
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 14354 8206 14366 8258
rect 14418 8206 14430 8258
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 10222 8194 10274 8206
rect 21534 8194 21586 8206
rect 22430 8258 22482 8270
rect 22430 8194 22482 8206
rect 22766 8258 22818 8270
rect 22766 8194 22818 8206
rect 24894 8258 24946 8270
rect 24894 8194 24946 8206
rect 25454 8258 25506 8270
rect 25454 8194 25506 8206
rect 29934 8258 29986 8270
rect 29934 8194 29986 8206
rect 32398 8258 32450 8270
rect 32398 8194 32450 8206
rect 48638 8258 48690 8270
rect 48638 8194 48690 8206
rect 49534 8258 49586 8270
rect 50418 8206 50430 8258
rect 50482 8206 50494 8258
rect 49534 8194 49586 8206
rect 12238 8146 12290 8158
rect 12238 8082 12290 8094
rect 13022 8146 13074 8158
rect 13022 8082 13074 8094
rect 13582 8146 13634 8158
rect 13582 8082 13634 8094
rect 15150 8146 15202 8158
rect 21870 8146 21922 8158
rect 18498 8094 18510 8146
rect 18562 8094 18574 8146
rect 15150 8082 15202 8094
rect 21870 8082 21922 8094
rect 24670 8146 24722 8158
rect 24670 8082 24722 8094
rect 30158 8146 30210 8158
rect 30158 8082 30210 8094
rect 31838 8146 31890 8158
rect 31838 8082 31890 8094
rect 32958 8146 33010 8158
rect 32958 8082 33010 8094
rect 48190 8146 48242 8158
rect 48190 8082 48242 8094
rect 48302 8146 48354 8158
rect 49970 8094 49982 8146
rect 50034 8094 50046 8146
rect 48302 8082 48354 8094
rect 51438 8034 51490 8046
rect 51438 7970 51490 7982
rect 672 7866 52080 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 52080 7866
rect 672 7780 52080 7814
rect 13022 7698 13074 7710
rect 13022 7634 13074 7646
rect 14590 7698 14642 7710
rect 14590 7634 14642 7646
rect 50878 7698 50930 7710
rect 50878 7634 50930 7646
rect 21870 7586 21922 7598
rect 18498 7534 18510 7586
rect 18562 7534 18574 7586
rect 21870 7522 21922 7534
rect 23326 7586 23378 7598
rect 23326 7522 23378 7534
rect 24110 7586 24162 7598
rect 24110 7522 24162 7534
rect 49646 7586 49698 7598
rect 49646 7522 49698 7534
rect 23886 7474 23938 7486
rect 14018 7422 14030 7474
rect 14082 7422 14094 7474
rect 23886 7410 23938 7422
rect 29934 7474 29986 7486
rect 48738 7422 48750 7474
rect 48802 7422 48814 7474
rect 51314 7422 51326 7474
rect 51378 7422 51390 7474
rect 29934 7410 29986 7422
rect 15586 7310 15598 7362
rect 15650 7310 15662 7362
rect 18958 7250 19010 7262
rect 18958 7186 19010 7198
rect 19294 7250 19346 7262
rect 19294 7186 19346 7198
rect 29150 7250 29202 7262
rect 29150 7186 29202 7198
rect 29374 7250 29426 7262
rect 29374 7186 29426 7198
rect 672 7082 52080 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 52080 7082
rect 672 6996 52080 7030
rect 5854 6690 5906 6702
rect 5854 6626 5906 6638
rect 8990 6690 9042 6702
rect 8990 6626 9042 6638
rect 9550 6690 9602 6702
rect 9550 6626 9602 6638
rect 9886 6690 9938 6702
rect 9886 6626 9938 6638
rect 18734 6690 18786 6702
rect 18734 6626 18786 6638
rect 19294 6690 19346 6702
rect 19294 6626 19346 6638
rect 19630 6690 19682 6702
rect 19630 6626 19682 6638
rect 23326 6690 23378 6702
rect 23326 6626 23378 6638
rect 29374 6690 29426 6702
rect 29374 6626 29426 6638
rect 29934 6690 29986 6702
rect 29934 6626 29986 6638
rect 44606 6690 44658 6702
rect 48850 6638 48862 6690
rect 48914 6638 48926 6690
rect 50418 6638 50430 6690
rect 50482 6638 50494 6690
rect 44606 6626 44658 6638
rect 5518 6578 5570 6590
rect 23662 6578 23714 6590
rect 6290 6526 6302 6578
rect 6354 6526 6366 6578
rect 22866 6526 22878 6578
rect 22930 6526 22942 6578
rect 5518 6514 5570 6526
rect 23662 6514 23714 6526
rect 29038 6578 29090 6590
rect 29038 6514 29090 6526
rect 44382 6578 44434 6590
rect 51438 6578 51490 6590
rect 45042 6526 45054 6578
rect 45106 6526 45118 6578
rect 49746 6526 49758 6578
rect 49810 6526 49822 6578
rect 44382 6514 44434 6526
rect 51438 6514 51490 6526
rect 672 6298 52080 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 52080 6298
rect 672 6212 52080 6246
rect 51214 6130 51266 6142
rect 51214 6066 51266 6078
rect 9550 6018 9602 6030
rect 5058 5966 5070 6018
rect 5122 5966 5134 6018
rect 9550 5954 9602 5966
rect 23774 6018 23826 6030
rect 23774 5954 23826 5966
rect 24558 6018 24610 6030
rect 24558 5954 24610 5966
rect 37550 6018 37602 6030
rect 47742 6018 47794 6030
rect 48974 6018 49026 6030
rect 38210 5966 38222 6018
rect 38274 5966 38286 6018
rect 48514 5966 48526 6018
rect 48578 5966 48590 6018
rect 37550 5954 37602 5966
rect 47742 5954 47794 5966
rect 48974 5954 49026 5966
rect 49870 6018 49922 6030
rect 49870 5954 49922 5966
rect 6750 5906 6802 5918
rect 6750 5842 6802 5854
rect 10110 5906 10162 5918
rect 10110 5842 10162 5854
rect 24334 5906 24386 5918
rect 24334 5842 24386 5854
rect 37774 5906 37826 5918
rect 37774 5842 37826 5854
rect 38670 5906 38722 5918
rect 38670 5842 38722 5854
rect 48078 5906 48130 5918
rect 48078 5842 48130 5854
rect 49310 5906 49362 5918
rect 50194 5854 50206 5906
rect 50258 5854 50270 5906
rect 49310 5842 49362 5854
rect 5518 5794 5570 5806
rect 5518 5730 5570 5742
rect 6414 5794 6466 5806
rect 6414 5730 6466 5742
rect 10446 5794 10498 5806
rect 10446 5730 10498 5742
rect 39230 5794 39282 5806
rect 39230 5730 39282 5742
rect 5854 5682 5906 5694
rect 5854 5618 5906 5630
rect 11006 5682 11058 5694
rect 11006 5618 11058 5630
rect 11230 5682 11282 5694
rect 11230 5618 11282 5630
rect 672 5514 52080 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 52080 5514
rect 672 5428 52080 5462
rect 17614 5346 17666 5358
rect 17614 5282 17666 5294
rect 17838 5346 17890 5358
rect 17838 5282 17890 5294
rect 23102 5346 23154 5358
rect 23102 5282 23154 5294
rect 23438 5346 23490 5358
rect 23438 5282 23490 5294
rect 38334 5346 38386 5358
rect 38334 5282 38386 5294
rect 5966 5234 6018 5246
rect 5966 5170 6018 5182
rect 10446 5234 10498 5246
rect 10446 5170 10498 5182
rect 14254 5234 14306 5246
rect 14254 5170 14306 5182
rect 17054 5234 17106 5246
rect 17054 5170 17106 5182
rect 22542 5234 22594 5246
rect 22542 5170 22594 5182
rect 38670 5234 38722 5246
rect 38670 5170 38722 5182
rect 38894 5234 38946 5246
rect 38894 5170 38946 5182
rect 39454 5234 39506 5246
rect 51202 5182 51214 5234
rect 51266 5182 51278 5234
rect 39454 5170 39506 5182
rect 5518 5122 5570 5134
rect 5518 5058 5570 5070
rect 6526 5122 6578 5134
rect 6526 5058 6578 5070
rect 6750 5122 6802 5134
rect 6750 5058 6802 5070
rect 14814 5122 14866 5134
rect 14814 5058 14866 5070
rect 15150 5122 15202 5134
rect 15150 5058 15202 5070
rect 24558 5122 24610 5134
rect 24558 5058 24610 5070
rect 24894 5122 24946 5134
rect 49074 5070 49086 5122
rect 49138 5070 49150 5122
rect 49634 5070 49646 5122
rect 49698 5070 49710 5122
rect 50530 5070 50542 5122
rect 50594 5070 50606 5122
rect 24894 5058 24946 5070
rect 25454 5010 25506 5022
rect 25454 4946 25506 4958
rect 672 4730 52080 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 52080 4730
rect 672 4644 52080 4678
rect 51214 4562 51266 4574
rect 51214 4498 51266 4510
rect 10894 4450 10946 4462
rect 15598 4450 15650 4462
rect 10210 4398 10222 4450
rect 10274 4398 10286 4450
rect 14914 4398 14926 4450
rect 14978 4398 14990 4450
rect 10894 4386 10946 4398
rect 15598 4386 15650 4398
rect 26126 4450 26178 4462
rect 26126 4386 26178 4398
rect 27022 4450 27074 4462
rect 27022 4386 27074 4398
rect 32286 4450 32338 4462
rect 41918 4450 41970 4462
rect 43598 4450 43650 4462
rect 33058 4398 33070 4450
rect 33122 4398 33134 4450
rect 42690 4398 42702 4450
rect 42754 4398 42766 4450
rect 46834 4398 46846 4450
rect 46898 4398 46910 4450
rect 32286 4386 32338 4398
rect 41918 4386 41970 4398
rect 43598 4386 43650 4398
rect 10670 4338 10722 4350
rect 10670 4274 10722 4286
rect 15374 4338 15426 4350
rect 15374 4274 15426 4286
rect 26462 4338 26514 4350
rect 26462 4274 26514 4286
rect 32622 4338 32674 4350
rect 32622 4274 32674 4286
rect 42254 4338 42306 4350
rect 42254 4274 42306 4286
rect 44158 4338 44210 4350
rect 48738 4286 48750 4338
rect 48802 4286 48814 4338
rect 44158 4274 44210 4286
rect 44718 4226 44770 4238
rect 44718 4162 44770 4174
rect 48302 4226 48354 4238
rect 49410 4174 49422 4226
rect 49474 4174 49486 4226
rect 50194 4174 50206 4226
rect 50258 4174 50270 4226
rect 48302 4162 48354 4174
rect 46174 4114 46226 4126
rect 46174 4050 46226 4062
rect 46398 4114 46450 4126
rect 46398 4050 46450 4062
rect 47406 4114 47458 4126
rect 47406 4050 47458 4062
rect 47742 4114 47794 4126
rect 47742 4050 47794 4062
rect 672 3946 52080 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 52080 3946
rect 672 3860 52080 3894
rect 20302 3778 20354 3790
rect 20302 3714 20354 3726
rect 20638 3778 20690 3790
rect 20638 3714 20690 3726
rect 25118 3778 25170 3790
rect 25118 3714 25170 3726
rect 25342 3778 25394 3790
rect 25342 3714 25394 3726
rect 29038 3778 29090 3790
rect 29038 3714 29090 3726
rect 29262 3778 29314 3790
rect 29262 3714 29314 3726
rect 44494 3778 44546 3790
rect 44494 3714 44546 3726
rect 44718 3778 44770 3790
rect 44718 3714 44770 3726
rect 46734 3778 46786 3790
rect 46734 3714 46786 3726
rect 1822 3666 1874 3678
rect 1822 3602 1874 3614
rect 19742 3666 19794 3678
rect 19742 3602 19794 3614
rect 33518 3666 33570 3678
rect 33518 3602 33570 3614
rect 45278 3666 45330 3678
rect 45278 3602 45330 3614
rect 46398 3666 46450 3678
rect 48850 3614 48862 3666
rect 48914 3614 48926 3666
rect 46398 3602 46450 3614
rect 2382 3554 2434 3566
rect 2382 3490 2434 3502
rect 2718 3554 2770 3566
rect 28030 3554 28082 3566
rect 27682 3502 27694 3554
rect 27746 3502 27758 3554
rect 2718 3490 2770 3502
rect 28030 3490 28082 3502
rect 32958 3554 33010 3566
rect 32958 3490 33010 3502
rect 45614 3554 45666 3566
rect 45614 3490 45666 3502
rect 45838 3554 45890 3566
rect 50418 3502 50430 3554
rect 50482 3502 50494 3554
rect 45838 3490 45890 3502
rect 27246 3442 27298 3454
rect 24658 3390 24670 3442
rect 24722 3390 24734 3442
rect 27246 3378 27298 3390
rect 29822 3442 29874 3454
rect 29822 3378 29874 3390
rect 32734 3442 32786 3454
rect 32734 3378 32786 3390
rect 47294 3442 47346 3454
rect 47294 3378 47346 3390
rect 49870 3442 49922 3454
rect 49870 3378 49922 3390
rect 51438 3442 51490 3454
rect 51438 3378 51490 3390
rect 672 3162 52080 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 52080 3162
rect 672 3076 52080 3110
rect 51214 2994 51266 3006
rect 51214 2930 51266 2942
rect 1262 2882 1314 2894
rect 1262 2818 1314 2830
rect 2158 2882 2210 2894
rect 4846 2882 4898 2894
rect 3938 2830 3950 2882
rect 4002 2830 4014 2882
rect 2158 2818 2210 2830
rect 4846 2818 4898 2830
rect 10782 2882 10834 2894
rect 16830 2882 16882 2894
rect 11778 2830 11790 2882
rect 11842 2830 11854 2882
rect 10782 2818 10834 2830
rect 16830 2818 16882 2830
rect 36766 2882 36818 2894
rect 36766 2818 36818 2830
rect 38558 2882 38610 2894
rect 38558 2818 38610 2830
rect 45166 2882 45218 2894
rect 45166 2818 45218 2830
rect 46510 2882 46562 2894
rect 46510 2818 46562 2830
rect 48078 2882 48130 2894
rect 48078 2818 48130 2830
rect 1598 2770 1650 2782
rect 1598 2706 1650 2718
rect 4398 2770 4450 2782
rect 4398 2706 4450 2718
rect 11342 2770 11394 2782
rect 11342 2706 11394 2718
rect 37102 2770 37154 2782
rect 37102 2706 37154 2718
rect 38894 2770 38946 2782
rect 38894 2706 38946 2718
rect 45390 2770 45442 2782
rect 47058 2718 47070 2770
rect 47122 2718 47134 2770
rect 48738 2718 48750 2770
rect 48802 2718 48814 2770
rect 50306 2718 50318 2770
rect 50370 2718 50382 2770
rect 45390 2706 45442 2718
rect 37662 2658 37714 2670
rect 37662 2594 37714 2606
rect 39454 2658 39506 2670
rect 39454 2594 39506 2606
rect 45950 2658 46002 2670
rect 49410 2606 49422 2658
rect 49474 2606 49486 2658
rect 45950 2594 46002 2606
rect 12238 2546 12290 2558
rect 12238 2482 12290 2494
rect 12686 2546 12738 2558
rect 12686 2482 12738 2494
rect 17390 2546 17442 2558
rect 17390 2482 17442 2494
rect 17614 2546 17666 2558
rect 17614 2482 17666 2494
rect 672 2378 52080 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 52080 2378
rect 672 2292 52080 2326
rect 11678 2210 11730 2222
rect 11678 2146 11730 2158
rect 13694 2210 13746 2222
rect 13694 2146 13746 2158
rect 13918 2210 13970 2222
rect 13918 2146 13970 2158
rect 19518 2210 19570 2222
rect 19518 2146 19570 2158
rect 19854 2210 19906 2222
rect 19854 2146 19906 2158
rect 20750 2210 20802 2222
rect 20750 2146 20802 2158
rect 21086 2210 21138 2222
rect 21086 2146 21138 2158
rect 32622 2210 32674 2222
rect 32622 2146 32674 2158
rect 32846 2210 32898 2222
rect 32846 2146 32898 2158
rect 38894 2210 38946 2222
rect 38894 2146 38946 2158
rect 39118 2210 39170 2222
rect 39118 2146 39170 2158
rect 43598 2210 43650 2222
rect 43598 2146 43650 2158
rect 43822 2210 43874 2222
rect 43822 2146 43874 2158
rect 18958 2098 19010 2110
rect 18958 2034 19010 2046
rect 20190 2098 20242 2110
rect 20190 2034 20242 2046
rect 39678 2098 39730 2110
rect 39678 2034 39730 2046
rect 46734 2098 46786 2110
rect 46734 2034 46786 2046
rect 46958 2098 47010 2110
rect 46958 2034 47010 2046
rect 47518 2098 47570 2110
rect 48850 2046 48862 2098
rect 48914 2046 48926 2098
rect 47518 2034 47570 2046
rect 33406 1986 33458 1998
rect 50642 1934 50654 1986
rect 50706 1934 50718 1986
rect 33406 1922 33458 1934
rect 14478 1874 14530 1886
rect 49870 1874 49922 1886
rect 44258 1822 44270 1874
rect 44322 1822 44334 1874
rect 14478 1810 14530 1822
rect 49870 1810 49922 1822
rect 51438 1874 51490 1886
rect 51438 1810 51490 1822
rect 672 1594 52080 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 52080 1594
rect 672 1508 52080 1542
rect 49758 1426 49810 1438
rect 49758 1362 49810 1374
rect 48190 1314 48242 1326
rect 20402 1262 20414 1314
rect 20466 1262 20478 1314
rect 48190 1250 48242 1262
rect 51326 1314 51378 1326
rect 51326 1250 51378 1262
rect 20862 1202 20914 1214
rect 20862 1138 20914 1150
rect 21086 1202 21138 1214
rect 47170 1150 47182 1202
rect 47234 1150 47246 1202
rect 21086 1138 21138 1150
rect 48738 1038 48750 1090
rect 48802 1038 48814 1090
rect 50430 978 50482 990
rect 50430 914 50482 926
rect 50766 978 50818 990
rect 50766 914 50818 926
rect 672 810 52080 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 52080 810
rect 672 724 52080 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 17390 13134 17442 13186
rect 21198 13134 21250 13186
rect 35758 13134 35810 13186
rect 37774 13134 37826 13186
rect 37998 13134 38050 13186
rect 41246 13134 41298 13186
rect 45054 13134 45106 13186
rect 6526 13022 6578 13074
rect 13358 13022 13410 13074
rect 14926 13022 14978 13074
rect 15710 13022 15762 13074
rect 22878 13022 22930 13074
rect 25230 13022 25282 13074
rect 40686 13022 40738 13074
rect 43710 13022 43762 13074
rect 10334 12910 10386 12962
rect 11902 12910 11954 12962
rect 14142 12910 14194 12962
rect 17950 12910 18002 12962
rect 18398 12910 18450 12962
rect 21758 12910 21810 12962
rect 22094 12910 22146 12962
rect 35422 12910 35474 12962
rect 37326 12910 37378 12962
rect 39118 12910 39170 12962
rect 42254 12910 42306 12962
rect 42926 12910 42978 12962
rect 44494 12910 44546 12962
rect 47182 12910 47234 12962
rect 48974 12910 49026 12962
rect 50766 12910 50818 12962
rect 19182 12798 19234 12850
rect 36318 12798 36370 12850
rect 38558 12798 38610 12850
rect 40014 12798 40066 12850
rect 50430 12798 50482 12850
rect 51214 12798 51266 12850
rect 24222 12686 24274 12738
rect 48190 12686 48242 12738
rect 49758 12686 49810 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 11678 12350 11730 12402
rect 16718 12350 16770 12402
rect 18286 12350 18338 12402
rect 21646 12350 21698 12402
rect 22878 12350 22930 12402
rect 36542 12350 36594 12402
rect 38110 12350 38162 12402
rect 40014 12350 40066 12402
rect 41582 12350 41634 12402
rect 48078 12350 48130 12402
rect 6862 12238 6914 12290
rect 7758 12238 7810 12290
rect 9998 12238 10050 12290
rect 14814 12238 14866 12290
rect 19630 12238 19682 12290
rect 26350 12238 26402 12290
rect 27134 12238 27186 12290
rect 28030 12238 28082 12290
rect 28926 12238 28978 12290
rect 49646 12238 49698 12290
rect 51214 12238 51266 12290
rect 6302 12126 6354 12178
rect 15374 12126 15426 12178
rect 15822 12126 15874 12178
rect 17278 12126 17330 12178
rect 20862 12126 20914 12178
rect 23214 12126 23266 12178
rect 26686 12126 26738 12178
rect 28478 12126 28530 12178
rect 39454 12126 39506 12178
rect 41246 12126 41298 12178
rect 42590 12126 42642 12178
rect 48750 12126 48802 12178
rect 2606 12014 2658 12066
rect 5742 12014 5794 12066
rect 10670 12014 10722 12066
rect 12238 12014 12290 12066
rect 12798 12014 12850 12066
rect 13358 12014 13410 12066
rect 18846 12014 18898 12066
rect 23774 12014 23826 12066
rect 29934 12014 29986 12066
rect 31166 12014 31218 12066
rect 37550 12014 37602 12066
rect 39118 12014 39170 12066
rect 43150 12014 43202 12066
rect 47070 12014 47122 12066
rect 50206 12014 50258 12066
rect 3166 11902 3218 11954
rect 3502 11902 3554 11954
rect 7310 11902 7362 11954
rect 8206 11902 8258 11954
rect 8542 11902 8594 11954
rect 13694 11902 13746 11954
rect 24334 11902 24386 11954
rect 29374 11902 29426 11954
rect 30382 11902 30434 11954
rect 30606 11902 30658 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 7086 11566 7138 11618
rect 10894 11566 10946 11618
rect 12462 11566 12514 11618
rect 14030 11566 14082 11618
rect 23326 11566 23378 11618
rect 26910 11566 26962 11618
rect 38670 11566 38722 11618
rect 40798 11566 40850 11618
rect 42366 11566 42418 11618
rect 5294 11454 5346 11506
rect 6750 11454 6802 11506
rect 18846 11454 18898 11506
rect 21982 11454 22034 11506
rect 50430 11454 50482 11506
rect 5854 11342 5906 11394
rect 11454 11342 11506 11394
rect 13022 11342 13074 11394
rect 14590 11342 14642 11394
rect 16158 11342 16210 11394
rect 17166 11342 17218 11394
rect 18062 11342 18114 11394
rect 19742 11342 19794 11394
rect 21198 11342 21250 11394
rect 22766 11342 22818 11394
rect 25118 11342 25170 11394
rect 27918 11342 27970 11394
rect 37774 11342 37826 11394
rect 38110 11342 38162 11394
rect 40462 11342 40514 11394
rect 41806 11342 41858 11394
rect 48862 11342 48914 11394
rect 6302 11230 6354 11282
rect 7646 11230 7698 11282
rect 15486 11230 15538 11282
rect 16830 11230 16882 11282
rect 17726 11230 17778 11282
rect 20190 11230 20242 11282
rect 24670 11230 24722 11282
rect 25342 11230 25394 11282
rect 27582 11230 27634 11282
rect 28478 11230 28530 11282
rect 29038 11230 29090 11282
rect 36766 11230 36818 11282
rect 49870 11230 49922 11282
rect 51438 11118 51490 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 10446 10782 10498 10834
rect 11678 10782 11730 10834
rect 16382 10782 16434 10834
rect 18286 10782 18338 10834
rect 19854 10782 19906 10834
rect 21870 10782 21922 10834
rect 23438 10782 23490 10834
rect 37774 10782 37826 10834
rect 39342 10782 39394 10834
rect 40910 10782 40962 10834
rect 42478 10782 42530 10834
rect 1710 10670 1762 10722
rect 14702 10670 14754 10722
rect 26798 10670 26850 10722
rect 49646 10670 49698 10722
rect 9550 10558 9602 10610
rect 16942 10558 16994 10610
rect 18846 10558 18898 10610
rect 22878 10558 22930 10610
rect 27246 10558 27298 10610
rect 38782 10558 38834 10610
rect 40574 10558 40626 10610
rect 42030 10558 42082 10610
rect 48750 10558 48802 10610
rect 12238 10446 12290 10498
rect 15374 10446 15426 10498
rect 17278 10446 17330 10498
rect 21310 10446 21362 10498
rect 27806 10446 27858 10498
rect 37214 10446 37266 10498
rect 47518 10446 47570 10498
rect 47742 10446 47794 10498
rect 48302 10446 48354 10498
rect 50206 10446 50258 10498
rect 50990 10446 51042 10498
rect 2158 10334 2210 10386
rect 2494 10334 2546 10386
rect 6078 10334 6130 10386
rect 26126 10334 26178 10386
rect 26350 10334 26402 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 10446 9998 10498 10050
rect 10670 9998 10722 10050
rect 12462 9998 12514 10050
rect 14030 9998 14082 10050
rect 15598 9998 15650 10050
rect 19294 9998 19346 10050
rect 20862 9998 20914 10050
rect 22318 9998 22370 10050
rect 27358 9998 27410 10050
rect 34190 9998 34242 10050
rect 38894 9998 38946 10050
rect 40798 9998 40850 10050
rect 41806 9998 41858 10050
rect 24558 9886 24610 9938
rect 27694 9886 27746 9938
rect 50430 9886 50482 9938
rect 9438 9774 9490 9826
rect 12798 9774 12850 9826
rect 14590 9774 14642 9826
rect 16158 9774 16210 9826
rect 17054 9774 17106 9826
rect 19854 9774 19906 9826
rect 21422 9774 21474 9826
rect 21982 9774 22034 9826
rect 25118 9774 25170 9826
rect 26798 9774 26850 9826
rect 27134 9774 27186 9826
rect 34638 9774 34690 9826
rect 36206 9774 36258 9826
rect 38334 9774 38386 9826
rect 40350 9774 40402 9826
rect 43934 9774 43986 9826
rect 44830 9774 44882 9826
rect 48862 9774 48914 9826
rect 8990 9662 9042 9714
rect 9774 9662 9826 9714
rect 11230 9662 11282 9714
rect 18062 9662 18114 9714
rect 25454 9662 25506 9714
rect 26350 9662 26402 9714
rect 35086 9662 35138 9714
rect 35870 9662 35922 9714
rect 36766 9662 36818 9714
rect 42254 9662 42306 9714
rect 43598 9662 43650 9714
rect 44494 9662 44546 9714
rect 45278 9662 45330 9714
rect 49870 9662 49922 9714
rect 51438 9550 51490 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 14814 9214 14866 9266
rect 16382 9214 16434 9266
rect 19070 9214 19122 9266
rect 20862 9214 20914 9266
rect 40910 9214 40962 9266
rect 49646 9214 49698 9266
rect 8542 9102 8594 9154
rect 11566 9102 11618 9154
rect 17950 9102 18002 9154
rect 22990 9102 23042 9154
rect 25790 9102 25842 9154
rect 27022 9102 27074 9154
rect 38222 9102 38274 9154
rect 41582 9102 41634 9154
rect 44494 9102 44546 9154
rect 21758 8990 21810 9042
rect 22766 8990 22818 9042
rect 23774 8990 23826 9042
rect 24334 8990 24386 9042
rect 38558 8990 38610 9042
rect 48750 8990 48802 9042
rect 12238 8878 12290 8930
rect 13806 8878 13858 8930
rect 15374 8878 15426 8930
rect 16942 8878 16994 8930
rect 17278 8878 17330 8930
rect 20078 8878 20130 8930
rect 22206 8878 22258 8930
rect 24894 8878 24946 8930
rect 25230 8878 25282 8930
rect 39118 8878 39170 8930
rect 39902 8878 39954 8930
rect 48302 8878 48354 8930
rect 50206 8878 50258 8930
rect 50990 8878 51042 8930
rect 8990 8766 9042 8818
rect 9214 8766 9266 8818
rect 13022 8766 13074 8818
rect 13246 8766 13298 8818
rect 23998 8766 24050 8818
rect 47518 8766 47570 8818
rect 47742 8766 47794 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 22430 8430 22482 8482
rect 9326 8318 9378 8370
rect 19406 8318 19458 8370
rect 20974 8318 21026 8370
rect 29374 8318 29426 8370
rect 49198 8318 49250 8370
rect 9886 8206 9938 8258
rect 10222 8206 10274 8258
rect 12574 8206 12626 8258
rect 14366 8206 14418 8258
rect 16158 8206 16210 8258
rect 21534 8206 21586 8258
rect 22430 8206 22482 8258
rect 22766 8206 22818 8258
rect 24894 8206 24946 8258
rect 25454 8206 25506 8258
rect 29934 8206 29986 8258
rect 32398 8206 32450 8258
rect 48638 8206 48690 8258
rect 49534 8206 49586 8258
rect 50430 8206 50482 8258
rect 12238 8094 12290 8146
rect 13022 8094 13074 8146
rect 13582 8094 13634 8146
rect 15150 8094 15202 8146
rect 18510 8094 18562 8146
rect 21870 8094 21922 8146
rect 24670 8094 24722 8146
rect 30158 8094 30210 8146
rect 31838 8094 31890 8146
rect 32958 8094 33010 8146
rect 48190 8094 48242 8146
rect 48302 8094 48354 8146
rect 49982 8094 50034 8146
rect 51438 7982 51490 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 13022 7646 13074 7698
rect 14590 7646 14642 7698
rect 50878 7646 50930 7698
rect 18510 7534 18562 7586
rect 21870 7534 21922 7586
rect 23326 7534 23378 7586
rect 24110 7534 24162 7586
rect 49646 7534 49698 7586
rect 14030 7422 14082 7474
rect 23886 7422 23938 7474
rect 29934 7422 29986 7474
rect 48750 7422 48802 7474
rect 51326 7422 51378 7474
rect 15598 7310 15650 7362
rect 18958 7198 19010 7250
rect 19294 7198 19346 7250
rect 29150 7198 29202 7250
rect 29374 7198 29426 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 5854 6638 5906 6690
rect 8990 6638 9042 6690
rect 9550 6638 9602 6690
rect 9886 6638 9938 6690
rect 18734 6638 18786 6690
rect 19294 6638 19346 6690
rect 19630 6638 19682 6690
rect 23326 6638 23378 6690
rect 29374 6638 29426 6690
rect 29934 6638 29986 6690
rect 44606 6638 44658 6690
rect 48862 6638 48914 6690
rect 50430 6638 50482 6690
rect 5518 6526 5570 6578
rect 6302 6526 6354 6578
rect 22878 6526 22930 6578
rect 23662 6526 23714 6578
rect 29038 6526 29090 6578
rect 44382 6526 44434 6578
rect 45054 6526 45106 6578
rect 49758 6526 49810 6578
rect 51438 6526 51490 6578
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 51214 6078 51266 6130
rect 5070 5966 5122 6018
rect 9550 5966 9602 6018
rect 23774 5966 23826 6018
rect 24558 5966 24610 6018
rect 37550 5966 37602 6018
rect 38222 5966 38274 6018
rect 47742 5966 47794 6018
rect 48526 5966 48578 6018
rect 48974 5966 49026 6018
rect 49870 5966 49922 6018
rect 6750 5854 6802 5906
rect 10110 5854 10162 5906
rect 24334 5854 24386 5906
rect 37774 5854 37826 5906
rect 38670 5854 38722 5906
rect 48078 5854 48130 5906
rect 49310 5854 49362 5906
rect 50206 5854 50258 5906
rect 5518 5742 5570 5794
rect 6414 5742 6466 5794
rect 10446 5742 10498 5794
rect 39230 5742 39282 5794
rect 5854 5630 5906 5682
rect 11006 5630 11058 5682
rect 11230 5630 11282 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 17614 5294 17666 5346
rect 17838 5294 17890 5346
rect 23102 5294 23154 5346
rect 23438 5294 23490 5346
rect 38334 5294 38386 5346
rect 5966 5182 6018 5234
rect 10446 5182 10498 5234
rect 14254 5182 14306 5234
rect 17054 5182 17106 5234
rect 22542 5182 22594 5234
rect 38670 5182 38722 5234
rect 38894 5182 38946 5234
rect 39454 5182 39506 5234
rect 51214 5182 51266 5234
rect 5518 5070 5570 5122
rect 6526 5070 6578 5122
rect 6750 5070 6802 5122
rect 14814 5070 14866 5122
rect 15150 5070 15202 5122
rect 24558 5070 24610 5122
rect 24894 5070 24946 5122
rect 49086 5070 49138 5122
rect 49646 5070 49698 5122
rect 50542 5070 50594 5122
rect 25454 4958 25506 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 51214 4510 51266 4562
rect 10222 4398 10274 4450
rect 10894 4398 10946 4450
rect 14926 4398 14978 4450
rect 15598 4398 15650 4450
rect 26126 4398 26178 4450
rect 27022 4398 27074 4450
rect 32286 4398 32338 4450
rect 33070 4398 33122 4450
rect 41918 4398 41970 4450
rect 42702 4398 42754 4450
rect 43598 4398 43650 4450
rect 46846 4398 46898 4450
rect 10670 4286 10722 4338
rect 15374 4286 15426 4338
rect 26462 4286 26514 4338
rect 32622 4286 32674 4338
rect 42254 4286 42306 4338
rect 44158 4286 44210 4338
rect 48750 4286 48802 4338
rect 44718 4174 44770 4226
rect 48302 4174 48354 4226
rect 49422 4174 49474 4226
rect 50206 4174 50258 4226
rect 46174 4062 46226 4114
rect 46398 4062 46450 4114
rect 47406 4062 47458 4114
rect 47742 4062 47794 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 20302 3726 20354 3778
rect 20638 3726 20690 3778
rect 25118 3726 25170 3778
rect 25342 3726 25394 3778
rect 29038 3726 29090 3778
rect 29262 3726 29314 3778
rect 44494 3726 44546 3778
rect 44718 3726 44770 3778
rect 46734 3726 46786 3778
rect 1822 3614 1874 3666
rect 19742 3614 19794 3666
rect 33518 3614 33570 3666
rect 45278 3614 45330 3666
rect 46398 3614 46450 3666
rect 48862 3614 48914 3666
rect 2382 3502 2434 3554
rect 2718 3502 2770 3554
rect 27694 3502 27746 3554
rect 28030 3502 28082 3554
rect 32958 3502 33010 3554
rect 45614 3502 45666 3554
rect 45838 3502 45890 3554
rect 50430 3502 50482 3554
rect 24670 3390 24722 3442
rect 27246 3390 27298 3442
rect 29822 3390 29874 3442
rect 32734 3390 32786 3442
rect 47294 3390 47346 3442
rect 49870 3390 49922 3442
rect 51438 3390 51490 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 51214 2942 51266 2994
rect 1262 2830 1314 2882
rect 2158 2830 2210 2882
rect 3950 2830 4002 2882
rect 4846 2830 4898 2882
rect 10782 2830 10834 2882
rect 11790 2830 11842 2882
rect 16830 2830 16882 2882
rect 36766 2830 36818 2882
rect 38558 2830 38610 2882
rect 45166 2830 45218 2882
rect 46510 2830 46562 2882
rect 48078 2830 48130 2882
rect 1598 2718 1650 2770
rect 4398 2718 4450 2770
rect 11342 2718 11394 2770
rect 37102 2718 37154 2770
rect 38894 2718 38946 2770
rect 45390 2718 45442 2770
rect 47070 2718 47122 2770
rect 48750 2718 48802 2770
rect 50318 2718 50370 2770
rect 37662 2606 37714 2658
rect 39454 2606 39506 2658
rect 45950 2606 46002 2658
rect 49422 2606 49474 2658
rect 12238 2494 12290 2546
rect 12686 2494 12738 2546
rect 17390 2494 17442 2546
rect 17614 2494 17666 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 11678 2158 11730 2210
rect 13694 2158 13746 2210
rect 13918 2158 13970 2210
rect 19518 2158 19570 2210
rect 19854 2158 19906 2210
rect 20750 2158 20802 2210
rect 21086 2158 21138 2210
rect 32622 2158 32674 2210
rect 32846 2158 32898 2210
rect 38894 2158 38946 2210
rect 39118 2158 39170 2210
rect 43598 2158 43650 2210
rect 43822 2158 43874 2210
rect 18958 2046 19010 2098
rect 20190 2046 20242 2098
rect 39678 2046 39730 2098
rect 46734 2046 46786 2098
rect 46958 2046 47010 2098
rect 47518 2046 47570 2098
rect 48862 2046 48914 2098
rect 33406 1934 33458 1986
rect 50654 1934 50706 1986
rect 14478 1822 14530 1874
rect 44270 1822 44322 1874
rect 49870 1822 49922 1874
rect 51438 1822 51490 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 49758 1374 49810 1426
rect 20414 1262 20466 1314
rect 48190 1262 48242 1314
rect 51326 1262 51378 1314
rect 20862 1150 20914 1202
rect 21086 1150 21138 1202
rect 47182 1150 47234 1202
rect 48750 1038 48802 1090
rect 50430 926 50482 978
rect 50766 926 50818 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 7084 14196 7140 14206
rect 252 13972 308 13982
rect 252 6916 308 13916
rect 5516 13524 5572 13534
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 2268 13076 2324 13086
rect 812 12628 868 12638
rect 812 10500 868 12572
rect 1708 10722 1764 10734
rect 1708 10670 1710 10722
rect 1762 10670 1764 10722
rect 812 10434 868 10444
rect 1148 10612 1204 10622
rect 252 6850 308 6860
rect 1148 6804 1204 10556
rect 1148 6738 1204 6748
rect 1260 9940 1316 9950
rect 1260 2884 1316 9884
rect 1708 9268 1764 10670
rect 2268 10724 2324 13020
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 5180 12180 5236 12190
rect 2268 10658 2324 10668
rect 2604 12066 2660 12078
rect 2604 12014 2606 12066
rect 2658 12014 2660 12066
rect 2156 10388 2212 10398
rect 2492 10388 2548 10398
rect 2156 10386 2548 10388
rect 2156 10334 2158 10386
rect 2210 10334 2494 10386
rect 2546 10334 2548 10386
rect 2156 10332 2548 10334
rect 2156 10322 2212 10332
rect 1708 9202 1764 9212
rect 1596 7700 1652 7710
rect 1596 6692 1652 7644
rect 1596 6626 1652 6636
rect 1820 5796 1876 5806
rect 1820 3666 1876 5740
rect 1820 3614 1822 3666
rect 1874 3614 1876 3666
rect 1820 3602 1876 3614
rect 2380 3556 2436 3566
rect 2380 3462 2436 3500
rect 2156 2884 2212 2894
rect 1260 2882 1652 2884
rect 1260 2830 1262 2882
rect 1314 2830 1652 2882
rect 1260 2828 1652 2830
rect 1260 2818 1316 2828
rect 1596 2770 1652 2828
rect 2156 2790 2212 2828
rect 1596 2718 1598 2770
rect 1650 2718 1652 2770
rect 1596 2706 1652 2718
rect 1596 2212 1652 2222
rect 1596 112 1652 2156
rect 2492 1092 2548 10332
rect 2604 3332 2660 12014
rect 3164 11956 3220 11966
rect 3164 11862 3220 11900
rect 3500 11956 3556 11966
rect 3500 11862 3556 11900
rect 4464 11788 4728 11798
rect 3276 11732 3332 11742
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 2716 10388 2772 10398
rect 2716 7252 2772 10332
rect 3276 9716 3332 11676
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 5068 10948 5124 10958
rect 4956 10724 5012 10734
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 3276 9650 3332 9660
rect 4956 9492 5012 10668
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4956 9426 5012 9436
rect 3804 9370 4068 9380
rect 4464 8652 4728 8662
rect 4284 8596 4340 8606
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 4284 7476 4340 8540
rect 4284 7410 4340 7420
rect 2716 7186 2772 7196
rect 3612 7364 3668 7374
rect 3276 6804 3332 6814
rect 3276 6356 3332 6748
rect 3276 6290 3332 6300
rect 3500 5124 3556 5134
rect 3276 5068 3500 5124
rect 2716 3556 2772 3566
rect 2716 3462 2772 3500
rect 2604 3266 2660 3276
rect 2492 1026 2548 1036
rect 3276 980 3332 5068
rect 3500 5058 3556 5068
rect 3612 3220 3668 7308
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 5068 6018 5124 10892
rect 5180 6356 5236 12124
rect 5292 11844 5348 11854
rect 5292 11506 5348 11788
rect 5292 11454 5294 11506
rect 5346 11454 5348 11506
rect 5292 11442 5348 11454
rect 5516 7812 5572 13468
rect 6524 13076 6580 13086
rect 6300 13020 6524 13076
rect 6300 12178 6356 13020
rect 6524 12982 6580 13020
rect 6860 12290 6916 12302
rect 6860 12238 6862 12290
rect 6914 12238 6916 12290
rect 6300 12126 6302 12178
rect 6354 12126 6356 12178
rect 6300 12114 6356 12126
rect 6524 12180 6580 12190
rect 5740 12066 5796 12078
rect 5740 12014 5742 12066
rect 5794 12014 5796 12066
rect 5740 8596 5796 12014
rect 5852 11394 5908 11406
rect 5852 11342 5854 11394
rect 5906 11342 5908 11394
rect 5852 10388 5908 11342
rect 6300 11282 6356 11294
rect 6300 11230 6302 11282
rect 6354 11230 6356 11282
rect 6188 10500 6244 10510
rect 6076 10388 6132 10398
rect 5852 10386 6132 10388
rect 5852 10334 6078 10386
rect 6130 10334 6132 10386
rect 5852 10332 6132 10334
rect 6076 9940 6132 10332
rect 6076 9874 6132 9884
rect 5740 8530 5796 8540
rect 5516 7746 5572 7756
rect 5964 8148 6020 8158
rect 5852 6690 5908 6702
rect 5852 6638 5854 6690
rect 5906 6638 5908 6690
rect 5516 6580 5572 6590
rect 5852 6580 5908 6638
rect 5516 6578 5908 6580
rect 5516 6526 5518 6578
rect 5570 6526 5908 6578
rect 5516 6524 5908 6526
rect 5516 6514 5572 6524
rect 5180 6300 5348 6356
rect 5068 5966 5070 6018
rect 5122 5966 5124 6018
rect 5068 5954 5124 5966
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4172 4788 4228 4798
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 3612 3154 3668 3164
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3948 2884 4004 2894
rect 4172 2884 4228 4732
rect 5068 4564 5124 4574
rect 4844 4340 4900 4350
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 4844 2884 4900 4284
rect 3948 2882 4228 2884
rect 3948 2830 3950 2882
rect 4002 2830 4228 2882
rect 3948 2828 4228 2830
rect 4396 2882 4900 2884
rect 4396 2830 4846 2882
rect 4898 2830 4900 2882
rect 4396 2828 4900 2830
rect 3948 2818 4004 2828
rect 4396 2770 4452 2828
rect 4844 2818 4900 2828
rect 4396 2718 4398 2770
rect 4450 2718 4452 2770
rect 4396 2706 4452 2718
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 4172 1988 4228 1998
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 3276 914 3332 924
rect 4172 532 4228 1932
rect 5068 1204 5124 4508
rect 5068 1138 5124 1148
rect 5180 3108 5236 3118
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 4172 466 4228 476
rect 4060 420 4116 430
rect 4060 112 4116 364
rect 1568 0 1680 112
rect 4032 0 4144 112
rect 5180 84 5236 3052
rect 5292 2996 5348 6300
rect 5516 5796 5572 5806
rect 5516 5702 5572 5740
rect 5516 5124 5572 5134
rect 5516 5030 5572 5068
rect 5292 2930 5348 2940
rect 5628 1428 5684 6524
rect 5852 5682 5908 5694
rect 5852 5630 5854 5682
rect 5906 5630 5908 5682
rect 5852 5124 5908 5630
rect 5964 5684 6020 8092
rect 5964 5618 6020 5628
rect 5964 5236 6020 5246
rect 5964 5142 6020 5180
rect 5852 5058 5908 5068
rect 6188 4676 6244 10444
rect 6300 7252 6356 11230
rect 6300 7186 6356 7196
rect 6188 4610 6244 4620
rect 6300 6578 6356 6590
rect 6300 6526 6302 6578
rect 6354 6526 6356 6578
rect 6188 3780 6244 3790
rect 6188 2548 6244 3724
rect 6188 2482 6244 2492
rect 6300 1540 6356 6526
rect 6524 5908 6580 12124
rect 6748 11508 6804 11518
rect 6748 11414 6804 11452
rect 6860 10500 6916 12238
rect 7084 11618 7140 14140
rect 12320 14112 12432 14224
rect 12544 14112 12656 14224
rect 12768 14112 12880 14224
rect 12992 14112 13104 14224
rect 13216 14112 13328 14224
rect 13440 14112 13552 14224
rect 13664 14112 13776 14224
rect 13888 14112 14000 14224
rect 14112 14112 14224 14224
rect 14336 14112 14448 14224
rect 14560 14112 14672 14224
rect 14784 14112 14896 14224
rect 15008 14112 15120 14224
rect 15232 14112 15344 14224
rect 15456 14112 15568 14224
rect 15680 14112 15792 14224
rect 15904 14112 16016 14224
rect 16128 14112 16240 14224
rect 16352 14112 16464 14224
rect 16576 14112 16688 14224
rect 16800 14112 16912 14224
rect 17024 14112 17136 14224
rect 17248 14112 17360 14224
rect 17472 14112 17584 14224
rect 17696 14112 17808 14224
rect 17920 14112 18032 14224
rect 18144 14112 18256 14224
rect 18368 14112 18480 14224
rect 18592 14112 18704 14224
rect 18816 14112 18928 14224
rect 19040 14112 19152 14224
rect 19264 14112 19376 14224
rect 19488 14112 19600 14224
rect 19712 14112 19824 14224
rect 19936 14112 20048 14224
rect 20160 14112 20272 14224
rect 20384 14112 20496 14224
rect 20608 14112 20720 14224
rect 20832 14112 20944 14224
rect 21056 14112 21168 14224
rect 21280 14112 21392 14224
rect 21504 14112 21616 14224
rect 21728 14112 21840 14224
rect 21952 14112 22064 14224
rect 22176 14112 22288 14224
rect 22400 14112 22512 14224
rect 22624 14112 22736 14224
rect 22848 14112 22960 14224
rect 23072 14112 23184 14224
rect 23296 14112 23408 14224
rect 23520 14112 23632 14224
rect 23744 14112 23856 14224
rect 23968 14112 24080 14224
rect 24192 14112 24304 14224
rect 24416 14112 24528 14224
rect 24640 14112 24752 14224
rect 24864 14112 24976 14224
rect 25088 14112 25200 14224
rect 25312 14112 25424 14224
rect 25536 14112 25648 14224
rect 25760 14112 25872 14224
rect 25984 14112 26096 14224
rect 26208 14112 26320 14224
rect 26432 14112 26544 14224
rect 26656 14112 26768 14224
rect 26880 14112 26992 14224
rect 27104 14112 27216 14224
rect 27328 14112 27440 14224
rect 27552 14112 27664 14224
rect 27776 14112 27888 14224
rect 28000 14112 28112 14224
rect 28224 14112 28336 14224
rect 28448 14112 28560 14224
rect 28672 14112 28784 14224
rect 28896 14112 29008 14224
rect 29120 14112 29232 14224
rect 29344 14112 29456 14224
rect 29568 14112 29680 14224
rect 29792 14112 29904 14224
rect 30016 14112 30128 14224
rect 30240 14112 30352 14224
rect 30464 14112 30576 14224
rect 30688 14112 30800 14224
rect 30912 14112 31024 14224
rect 31136 14112 31248 14224
rect 31360 14112 31472 14224
rect 31584 14112 31696 14224
rect 31808 14112 31920 14224
rect 32032 14112 32144 14224
rect 32256 14112 32368 14224
rect 32480 14112 32592 14224
rect 32704 14112 32816 14224
rect 32928 14112 33040 14224
rect 33152 14112 33264 14224
rect 33376 14112 33488 14224
rect 33600 14112 33712 14224
rect 33824 14112 33936 14224
rect 34048 14112 34160 14224
rect 34272 14112 34384 14224
rect 34496 14112 34608 14224
rect 34720 14112 34832 14224
rect 34944 14112 35056 14224
rect 35168 14112 35280 14224
rect 35392 14112 35504 14224
rect 35616 14112 35728 14224
rect 35840 14112 35952 14224
rect 36064 14112 36176 14224
rect 36288 14112 36400 14224
rect 36512 14112 36624 14224
rect 36736 14112 36848 14224
rect 36960 14112 37072 14224
rect 37184 14112 37296 14224
rect 37408 14112 37520 14224
rect 37632 14112 37744 14224
rect 37856 14112 37968 14224
rect 38080 14112 38192 14224
rect 38304 14112 38416 14224
rect 38528 14112 38640 14224
rect 38752 14112 38864 14224
rect 38976 14112 39088 14224
rect 39200 14112 39312 14224
rect 39424 14112 39536 14224
rect 39648 14112 39760 14224
rect 39872 14112 39984 14224
rect 40096 14112 40208 14224
rect 41692 14196 41748 14206
rect 11564 14084 11620 14094
rect 9996 13636 10052 13646
rect 9772 13412 9828 13422
rect 9772 13186 9828 13356
rect 9772 13134 9774 13186
rect 9826 13134 9828 13186
rect 9772 13122 9828 13134
rect 7756 12292 7812 12302
rect 7756 12290 7924 12292
rect 7756 12238 7758 12290
rect 7810 12238 7924 12290
rect 7756 12236 7924 12238
rect 7756 12226 7812 12236
rect 7084 11566 7086 11618
rect 7138 11566 7140 11618
rect 7084 11508 7140 11566
rect 7084 11442 7140 11452
rect 7308 11954 7364 11966
rect 7308 11902 7310 11954
rect 7362 11902 7364 11954
rect 7308 11284 7364 11902
rect 7644 11284 7700 11294
rect 7308 11282 7700 11284
rect 7308 11230 7646 11282
rect 7698 11230 7700 11282
rect 7308 11228 7700 11230
rect 6860 10434 6916 10444
rect 7420 9940 7476 9950
rect 6524 5842 6580 5852
rect 6636 9492 6692 9502
rect 6412 5794 6468 5806
rect 6412 5742 6414 5794
rect 6466 5742 6468 5794
rect 6412 4564 6468 5742
rect 6524 5124 6580 5134
rect 6524 5030 6580 5068
rect 6412 4498 6468 4508
rect 6636 3388 6692 9436
rect 6972 9380 7028 9390
rect 6748 5908 6804 5918
rect 6748 5814 6804 5852
rect 6748 5124 6804 5134
rect 6748 5030 6804 5068
rect 6972 4788 7028 9324
rect 6972 4722 7028 4732
rect 6972 3444 7028 3454
rect 6636 3332 6804 3388
rect 6300 1474 6356 1484
rect 6524 1652 6580 1662
rect 5628 1362 5684 1372
rect 6524 112 6580 1596
rect 6748 532 6804 3332
rect 6972 2884 7028 3388
rect 6972 2818 7028 2828
rect 6748 466 6804 476
rect 7420 196 7476 9884
rect 7644 9940 7700 11228
rect 7644 9874 7700 9884
rect 7756 10836 7812 10846
rect 7644 8484 7700 8494
rect 7532 7140 7588 7150
rect 7532 5572 7588 7084
rect 7532 5506 7588 5516
rect 7532 4564 7588 4574
rect 7532 2884 7588 4508
rect 7644 3108 7700 8428
rect 7756 5796 7812 10780
rect 7756 5730 7812 5740
rect 7868 4564 7924 12236
rect 9996 12290 10052 13580
rect 11340 13524 11396 13534
rect 11004 13300 11060 13310
rect 9996 12238 9998 12290
rect 10050 12238 10052 12290
rect 9996 12226 10052 12238
rect 10332 12962 10388 12974
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 8204 11956 8260 11966
rect 8204 11862 8260 11900
rect 8540 11956 8596 11966
rect 8540 11862 8596 11900
rect 9324 11956 9380 11966
rect 8092 10388 8148 10398
rect 7980 9268 8036 9278
rect 7980 6132 8036 9212
rect 8092 8820 8148 10332
rect 8764 10276 8820 10286
rect 8204 10164 8260 10174
rect 8204 9044 8260 10108
rect 8652 9940 8708 9950
rect 8204 8978 8260 8988
rect 8316 9604 8372 9614
rect 8092 8754 8148 8764
rect 8316 8372 8372 9548
rect 8540 9156 8596 9166
rect 8540 9062 8596 9100
rect 8316 8306 8372 8316
rect 8652 8036 8708 9884
rect 8764 9716 8820 10220
rect 8764 9650 8820 9660
rect 8988 9716 9044 9726
rect 8988 9622 9044 9660
rect 9324 9604 9380 11900
rect 9548 10610 9604 10622
rect 9548 10558 9550 10610
rect 9602 10558 9604 10610
rect 9548 10388 9604 10558
rect 9548 10322 9604 10332
rect 10332 10388 10388 12910
rect 10668 12068 10724 12078
rect 10668 12066 10836 12068
rect 10668 12014 10670 12066
rect 10722 12014 10836 12066
rect 10668 12012 10836 12014
rect 10668 12002 10724 12012
rect 10444 10836 10500 10846
rect 10444 10742 10500 10780
rect 10332 10322 10388 10332
rect 10444 10052 10500 10062
rect 10444 9958 10500 9996
rect 10668 10052 10724 10062
rect 10668 9958 10724 9996
rect 9436 9826 9492 9838
rect 9436 9774 9438 9826
rect 9490 9774 9492 9826
rect 9436 9716 9492 9774
rect 9772 9716 9828 9726
rect 9436 9714 9828 9716
rect 9436 9662 9774 9714
rect 9826 9662 9828 9714
rect 9436 9660 9828 9662
rect 9324 9548 9492 9604
rect 8652 7970 8708 7980
rect 8876 9268 8932 9278
rect 7980 6066 8036 6076
rect 8092 7252 8148 7262
rect 8092 5572 8148 7196
rect 8316 6916 8372 6926
rect 8316 6020 8372 6860
rect 8876 6692 8932 9212
rect 9324 9044 9380 9054
rect 8988 8820 9044 8830
rect 9212 8820 9268 8830
rect 8988 8818 9268 8820
rect 8988 8766 8990 8818
rect 9042 8766 9214 8818
rect 9266 8766 9268 8818
rect 8988 8764 9268 8766
rect 8988 8754 9044 8764
rect 9212 7924 9268 8764
rect 9324 8370 9380 8988
rect 9324 8318 9326 8370
rect 9378 8318 9380 8370
rect 9324 8306 9380 8318
rect 9212 7858 9268 7868
rect 9212 7588 9268 7598
rect 9212 6804 9268 7532
rect 9212 6738 9268 6748
rect 8988 6692 9044 6702
rect 8876 6690 9044 6692
rect 8876 6638 8990 6690
rect 9042 6638 9044 6690
rect 8876 6636 9044 6638
rect 8988 6626 9044 6636
rect 8316 5954 8372 5964
rect 8092 5506 8148 5516
rect 8204 5684 8260 5694
rect 7868 4498 7924 4508
rect 8092 4116 8148 4126
rect 8092 3220 8148 4060
rect 8092 3154 8148 3164
rect 7644 3042 7700 3052
rect 7532 2818 7588 2828
rect 8204 2436 8260 5628
rect 8316 5236 8372 5246
rect 8316 3892 8372 5180
rect 8316 3826 8372 3836
rect 8764 4900 8820 4910
rect 8204 2370 8260 2380
rect 8764 2100 8820 4844
rect 8764 2034 8820 2044
rect 7420 130 7476 140
rect 8988 1652 9044 1662
rect 8988 112 9044 1596
rect 5180 18 5236 28
rect 6496 0 6608 112
rect 8960 0 9072 112
rect 9436 84 9492 9548
rect 9772 8148 9828 9660
rect 10108 9604 10164 9614
rect 9884 8260 9940 8270
rect 9884 8166 9940 8204
rect 9772 8082 9828 8092
rect 10108 6804 10164 9548
rect 10220 8260 10276 8270
rect 10220 8166 10276 8204
rect 9996 6748 10164 6804
rect 10556 8036 10612 8046
rect 9548 6692 9604 6702
rect 9548 6598 9604 6636
rect 9884 6692 9940 6702
rect 9884 6598 9940 6636
rect 9548 6244 9604 6254
rect 9548 6018 9604 6188
rect 9548 5966 9550 6018
rect 9602 5966 9604 6018
rect 9548 5954 9604 5966
rect 9772 5124 9828 5134
rect 9772 2548 9828 5068
rect 9884 4676 9940 4686
rect 9884 2660 9940 4620
rect 9884 2594 9940 2604
rect 9772 2482 9828 2492
rect 9996 2212 10052 6748
rect 10108 6244 10164 6254
rect 10108 5908 10164 6188
rect 10108 5906 10388 5908
rect 10108 5854 10110 5906
rect 10162 5854 10388 5906
rect 10108 5852 10388 5854
rect 10108 5842 10164 5852
rect 10332 5236 10388 5852
rect 10444 5794 10500 5806
rect 10444 5742 10446 5794
rect 10498 5742 10500 5794
rect 10444 5460 10500 5742
rect 10444 5394 10500 5404
rect 10444 5236 10500 5246
rect 10332 5234 10500 5236
rect 10332 5182 10446 5234
rect 10498 5182 10500 5234
rect 10332 5180 10500 5182
rect 10444 5170 10500 5180
rect 10220 4452 10276 4462
rect 10220 4358 10276 4396
rect 10556 2436 10612 7980
rect 10780 7028 10836 12012
rect 10892 11844 10948 11854
rect 10892 11618 10948 11788
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 10780 6962 10836 6972
rect 11004 6020 11060 13244
rect 11340 13186 11396 13468
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 11452 11394 11508 11406
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11228 9714 11284 9726
rect 11228 9662 11230 9714
rect 11282 9662 11284 9714
rect 11228 6804 11284 9662
rect 11228 6738 11284 6748
rect 10892 5964 11060 6020
rect 10892 5460 10948 5964
rect 11004 5684 11060 5694
rect 11228 5684 11284 5694
rect 11004 5682 11284 5684
rect 11004 5630 11006 5682
rect 11058 5630 11230 5682
rect 11282 5630 11284 5682
rect 11004 5628 11284 5630
rect 11004 5618 11060 5628
rect 10892 5404 11060 5460
rect 10892 5236 10948 5246
rect 10892 4452 10948 5180
rect 10668 4450 10948 4452
rect 10668 4398 10894 4450
rect 10946 4398 10948 4450
rect 10668 4396 10948 4398
rect 10668 4338 10724 4396
rect 10892 4386 10948 4396
rect 10668 4286 10670 4338
rect 10722 4286 10724 4338
rect 10668 4274 10724 4286
rect 11004 3388 11060 5404
rect 11228 4788 11284 5628
rect 11228 4722 11284 4732
rect 11452 4676 11508 11342
rect 11564 9154 11620 14028
rect 12348 14084 12404 14112
rect 12348 14018 12404 14028
rect 11900 12964 11956 12974
rect 11900 12870 11956 12908
rect 11900 12740 11956 12750
rect 11676 12404 11732 12414
rect 11676 12310 11732 12348
rect 11788 12292 11844 12302
rect 11788 11732 11844 12236
rect 11676 11676 11844 11732
rect 11676 10834 11732 11676
rect 11900 11396 11956 12684
rect 12460 12628 12516 12638
rect 12236 12066 12292 12078
rect 12236 12014 12238 12066
rect 12290 12014 12292 12066
rect 12236 11508 12292 12014
rect 12460 11618 12516 12572
rect 12460 11566 12462 11618
rect 12514 11566 12516 11618
rect 12460 11554 12516 11566
rect 12236 11442 12292 11452
rect 11676 10782 11678 10834
rect 11730 10782 11732 10834
rect 11676 10770 11732 10782
rect 11788 11340 11956 11396
rect 11788 10388 11844 11340
rect 12012 11284 12068 11294
rect 11564 9102 11566 9154
rect 11618 9102 11620 9154
rect 11564 9090 11620 9102
rect 11676 10332 11844 10388
rect 11900 11172 11956 11182
rect 11564 7700 11620 7710
rect 11564 6692 11620 7644
rect 11676 7140 11732 10332
rect 11676 7074 11732 7084
rect 11788 10164 11844 10174
rect 11788 6804 11844 10108
rect 11900 9156 11956 11116
rect 11900 9090 11956 9100
rect 11900 8372 11956 8382
rect 11900 8148 11956 8316
rect 11900 8082 11956 8092
rect 11564 6626 11620 6636
rect 11676 6748 11844 6804
rect 11676 5878 11732 6748
rect 11452 4610 11508 4620
rect 11564 5822 11732 5878
rect 11788 6468 11844 6478
rect 10780 3332 11060 3388
rect 11340 3668 11396 3678
rect 10780 2882 10836 3332
rect 10780 2830 10782 2882
rect 10834 2830 10836 2882
rect 10780 2818 10836 2830
rect 11228 3220 11284 3230
rect 10556 2370 10612 2380
rect 9996 2146 10052 2156
rect 11228 1652 11284 3164
rect 11340 2770 11396 3612
rect 11564 3388 11620 5822
rect 11676 5684 11732 5694
rect 11676 4228 11732 5628
rect 11788 4452 11844 6412
rect 11788 4386 11844 4396
rect 11676 4162 11732 4172
rect 11340 2718 11342 2770
rect 11394 2718 11396 2770
rect 11340 2706 11396 2718
rect 11452 3332 11620 3388
rect 11676 3668 11732 3678
rect 11228 1586 11284 1596
rect 11452 112 11508 3332
rect 11564 2772 11620 2782
rect 11564 1652 11620 2716
rect 11676 2210 11732 3612
rect 12012 3388 12068 11228
rect 12572 10836 12628 14112
rect 12572 10770 12628 10780
rect 12684 12852 12740 12862
rect 12236 10498 12292 10510
rect 12236 10446 12238 10498
rect 12290 10446 12292 10498
rect 12236 9492 12292 10446
rect 12460 10052 12516 10062
rect 12460 9958 12516 9996
rect 12236 9426 12292 9436
rect 12124 9156 12180 9166
rect 12124 8484 12180 9100
rect 12236 8932 12292 8942
rect 12236 8838 12292 8876
rect 12124 8418 12180 8428
rect 12572 8258 12628 8270
rect 12572 8206 12574 8258
rect 12626 8206 12628 8258
rect 12236 8148 12292 8158
rect 12572 8148 12628 8206
rect 12236 8146 12628 8148
rect 12236 8094 12238 8146
rect 12290 8094 12628 8146
rect 12236 8092 12628 8094
rect 12236 8082 12292 8092
rect 12572 6916 12628 8092
rect 12572 6850 12628 6860
rect 12684 6132 12740 12796
rect 12796 12292 12852 14112
rect 12796 12236 12964 12292
rect 12796 12066 12852 12078
rect 12796 12014 12798 12066
rect 12850 12014 12852 12066
rect 12796 11956 12852 12014
rect 12796 11890 12852 11900
rect 12572 6076 12740 6132
rect 12796 9826 12852 9838
rect 12796 9774 12798 9826
rect 12850 9774 12852 9826
rect 12572 5908 12628 6076
rect 12572 5842 12628 5852
rect 12796 5908 12852 9774
rect 12908 7700 12964 12236
rect 13020 11844 13076 14112
rect 13244 12292 13300 14112
rect 13356 13188 13412 13198
rect 13356 13074 13412 13132
rect 13356 13022 13358 13074
rect 13410 13022 13412 13074
rect 13356 13010 13412 13022
rect 13244 12226 13300 12236
rect 13356 12068 13412 12078
rect 13356 11974 13412 12012
rect 13020 11778 13076 11788
rect 13020 11396 13076 11406
rect 13020 11302 13076 11340
rect 13020 8820 13076 8830
rect 13244 8820 13300 8830
rect 13020 8818 13300 8820
rect 13020 8766 13022 8818
rect 13074 8766 13246 8818
rect 13298 8766 13300 8818
rect 13020 8764 13300 8766
rect 13020 8754 13076 8764
rect 13020 8146 13076 8158
rect 13020 8094 13022 8146
rect 13074 8094 13076 8146
rect 13020 8036 13076 8094
rect 13020 7970 13076 7980
rect 13020 7700 13076 7710
rect 12908 7698 13076 7700
rect 12908 7646 13022 7698
rect 13074 7646 13076 7698
rect 12908 7644 13076 7646
rect 13020 7634 13076 7644
rect 13244 7252 13300 8764
rect 13468 8148 13524 14112
rect 13692 12292 13748 14112
rect 13916 13636 13972 14112
rect 13916 13570 13972 13580
rect 14140 13188 14196 14112
rect 14364 13412 14420 14112
rect 14364 13346 14420 13356
rect 14140 13132 14532 13188
rect 13580 12236 13748 12292
rect 14140 12962 14196 12974
rect 14140 12910 14142 12962
rect 14194 12910 14196 12962
rect 13580 10052 13636 12236
rect 13692 12068 13748 12078
rect 13692 11954 13748 12012
rect 13692 11902 13694 11954
rect 13746 11902 13748 11954
rect 13692 10724 13748 11902
rect 14028 12068 14084 12078
rect 14028 11618 14084 12012
rect 14028 11566 14030 11618
rect 14082 11566 14084 11618
rect 14028 11554 14084 11566
rect 13916 11396 13972 11406
rect 13692 10658 13748 10668
rect 13804 11284 13860 11294
rect 13580 9986 13636 9996
rect 13804 9268 13860 11228
rect 13804 9202 13860 9212
rect 13804 8930 13860 8942
rect 13804 8878 13806 8930
rect 13858 8878 13860 8930
rect 13580 8148 13636 8158
rect 13468 8146 13636 8148
rect 13468 8094 13582 8146
rect 13634 8094 13636 8146
rect 13468 8092 13636 8094
rect 13580 8082 13636 8092
rect 13804 7364 13860 8878
rect 13804 7298 13860 7308
rect 13244 7186 13300 7196
rect 13804 6804 13860 6814
rect 12796 5842 12852 5852
rect 13692 6692 13748 6702
rect 11900 3332 12068 3388
rect 13356 5796 13412 5806
rect 13356 3388 13412 5740
rect 13692 4452 13748 6636
rect 13692 4386 13748 4396
rect 13356 3332 13748 3388
rect 11788 3108 11844 3118
rect 11788 2882 11844 3052
rect 11788 2830 11790 2882
rect 11842 2830 11844 2882
rect 11788 2818 11844 2830
rect 11676 2158 11678 2210
rect 11730 2158 11732 2210
rect 11676 2146 11732 2158
rect 11564 1586 11620 1596
rect 11900 532 11956 3332
rect 12460 2772 12516 2782
rect 12236 2546 12292 2558
rect 12236 2494 12238 2546
rect 12290 2494 12292 2546
rect 12236 2324 12292 2494
rect 12236 2258 12292 2268
rect 12460 1876 12516 2716
rect 12684 2546 12740 2558
rect 12684 2494 12686 2546
rect 12738 2494 12740 2546
rect 12460 1810 12516 1820
rect 12572 2436 12628 2446
rect 12572 980 12628 2380
rect 12572 914 12628 924
rect 12684 2324 12740 2494
rect 11900 466 11956 476
rect 12684 420 12740 2268
rect 13692 2212 13748 3332
rect 13804 2660 13860 6748
rect 13916 6692 13972 11340
rect 14140 11060 14196 12910
rect 14140 10994 14196 11004
rect 14364 12740 14420 12750
rect 14252 10948 14308 10958
rect 14028 10050 14084 10062
rect 14028 9998 14030 10050
rect 14082 9998 14084 10050
rect 14028 9940 14084 9998
rect 14028 9874 14084 9884
rect 14028 7476 14084 7486
rect 14028 7382 14084 7420
rect 13916 6626 13972 6636
rect 14252 5234 14308 10892
rect 14364 10164 14420 12684
rect 14364 10098 14420 10108
rect 14364 8258 14420 8270
rect 14364 8206 14366 8258
rect 14418 8206 14420 8258
rect 14364 5796 14420 8206
rect 14476 7700 14532 13132
rect 14588 12404 14644 14112
rect 14700 13860 14756 13870
rect 14700 12740 14756 13804
rect 14700 12674 14756 12684
rect 14812 12628 14868 14112
rect 14924 13300 14980 13310
rect 14924 13074 14980 13244
rect 14924 13022 14926 13074
rect 14978 13022 14980 13074
rect 14924 13010 14980 13022
rect 14812 12562 14868 12572
rect 14588 12338 14644 12348
rect 14700 12516 14756 12526
rect 14588 11396 14644 11406
rect 14588 11302 14644 11340
rect 14700 10722 14756 12460
rect 14812 12292 14868 12302
rect 14812 12198 14868 12236
rect 14700 10670 14702 10722
rect 14754 10670 14756 10722
rect 14700 10658 14756 10670
rect 15036 10612 15092 14112
rect 15148 13636 15204 13646
rect 15148 12068 15204 13580
rect 15148 12002 15204 12012
rect 15036 10556 15204 10612
rect 14924 10164 14980 10174
rect 14588 9828 14644 9838
rect 14588 9734 14644 9772
rect 14812 9268 14868 9278
rect 14812 9174 14868 9212
rect 14588 7700 14644 7710
rect 14476 7698 14644 7700
rect 14476 7646 14590 7698
rect 14642 7646 14644 7698
rect 14476 7644 14644 7646
rect 14588 7634 14644 7644
rect 14588 7140 14644 7150
rect 14364 5730 14420 5740
rect 14476 6580 14532 6590
rect 14252 5182 14254 5234
rect 14306 5182 14308 5234
rect 14252 5170 14308 5182
rect 14252 4788 14308 4798
rect 13804 2594 13860 2604
rect 14140 2996 14196 3006
rect 14140 2660 14196 2940
rect 14140 2594 14196 2604
rect 13916 2212 13972 2222
rect 13692 2210 13972 2212
rect 13692 2158 13694 2210
rect 13746 2158 13918 2210
rect 13970 2158 13972 2210
rect 13692 2156 13972 2158
rect 13692 2146 13748 2156
rect 13916 2146 13972 2156
rect 14252 2100 14308 4732
rect 14476 4788 14532 6524
rect 14476 4722 14532 4732
rect 14588 3108 14644 7084
rect 14700 5908 14756 5918
rect 14700 4228 14756 5852
rect 14812 5124 14868 5134
rect 14812 5030 14868 5068
rect 14924 4450 14980 10108
rect 15148 8146 15204 10556
rect 15260 9940 15316 14112
rect 15484 13860 15540 14112
rect 15484 13804 15652 13860
rect 15484 13636 15540 13646
rect 15372 12180 15428 12190
rect 15372 12086 15428 12124
rect 15372 11620 15428 11630
rect 15372 11060 15428 11564
rect 15484 11282 15540 13580
rect 15596 12740 15652 13804
rect 15708 13524 15764 14112
rect 15932 13748 15988 14112
rect 15932 13682 15988 13692
rect 15708 13458 15764 13468
rect 15708 13076 15764 13086
rect 15708 13074 15988 13076
rect 15708 13022 15710 13074
rect 15762 13022 15988 13074
rect 15708 13020 15988 13022
rect 15708 13010 15764 13020
rect 15820 12852 15876 12862
rect 15596 12684 15764 12740
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15484 11218 15540 11230
rect 15596 12404 15652 12414
rect 15372 11004 15540 11060
rect 15372 10498 15428 10510
rect 15372 10446 15374 10498
rect 15426 10446 15428 10498
rect 15372 10388 15428 10446
rect 15372 10322 15428 10332
rect 15484 10276 15540 11004
rect 15484 10210 15540 10220
rect 15596 10050 15652 12348
rect 15596 9998 15598 10050
rect 15650 9998 15652 10050
rect 15596 9986 15652 9998
rect 15260 9874 15316 9884
rect 15708 9268 15764 12684
rect 15820 12178 15876 12796
rect 15820 12126 15822 12178
rect 15874 12126 15876 12178
rect 15820 12114 15876 12126
rect 15932 11732 15988 13020
rect 16156 12404 16212 14112
rect 16380 12628 16436 14112
rect 16380 12562 16436 12572
rect 16156 12338 16212 12348
rect 16380 12404 16436 12414
rect 15932 11666 15988 11676
rect 16044 11396 16100 11406
rect 15932 10612 15988 10622
rect 15932 10276 15988 10556
rect 15932 10210 15988 10220
rect 15932 9268 15988 9278
rect 15708 9202 15764 9212
rect 15820 9212 15932 9268
rect 15484 9156 15540 9166
rect 15372 8930 15428 8942
rect 15372 8878 15374 8930
rect 15426 8878 15428 8930
rect 15148 8094 15150 8146
rect 15202 8094 15204 8146
rect 15148 8082 15204 8094
rect 15260 8372 15316 8382
rect 15148 7700 15204 7710
rect 15260 7700 15316 8316
rect 15204 7644 15316 7700
rect 15372 7700 15428 8878
rect 15148 7634 15204 7644
rect 15372 7634 15428 7644
rect 15372 7364 15428 7374
rect 15372 5460 15428 7308
rect 15484 6244 15540 9100
rect 15596 7364 15652 7374
rect 15596 7270 15652 7308
rect 15484 6178 15540 6188
rect 15596 5460 15652 5470
rect 15372 5404 15596 5460
rect 15596 5394 15652 5404
rect 15148 5124 15204 5134
rect 15820 5124 15876 9212
rect 15932 9202 15988 9212
rect 16044 6244 16100 11340
rect 16156 11394 16212 11406
rect 16156 11342 16158 11394
rect 16210 11342 16212 11394
rect 16156 10612 16212 11342
rect 16380 10834 16436 12348
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10770 16436 10782
rect 16156 10546 16212 10556
rect 16492 10724 16548 10734
rect 16492 9940 16548 10668
rect 16492 9874 16548 9884
rect 16156 9828 16212 9838
rect 16156 9826 16324 9828
rect 16156 9774 16158 9826
rect 16210 9774 16324 9826
rect 16156 9772 16324 9774
rect 16156 9762 16212 9772
rect 16044 6178 16100 6188
rect 16156 8258 16212 8270
rect 16156 8206 16158 8258
rect 16210 8206 16212 8258
rect 15148 5030 15204 5068
rect 15372 5068 15876 5124
rect 15372 4900 15428 5068
rect 15372 4834 15428 4844
rect 15596 4900 15652 4910
rect 15596 4452 15652 4844
rect 14924 4398 14926 4450
rect 14978 4398 14980 4450
rect 14924 4386 14980 4398
rect 15372 4450 15652 4452
rect 15372 4398 15598 4450
rect 15650 4398 15652 4450
rect 15372 4396 15652 4398
rect 15372 4338 15428 4396
rect 15596 4386 15652 4396
rect 15372 4286 15374 4338
rect 15426 4286 15428 4338
rect 15372 4274 15428 4286
rect 14700 4172 14980 4228
rect 14924 4004 14980 4172
rect 15092 4004 15204 4116
rect 14924 3948 15204 4004
rect 14588 3042 14644 3052
rect 15148 2996 15204 3948
rect 15820 3892 15876 3902
rect 15148 2930 15204 2940
rect 15372 3780 15428 3790
rect 15372 2324 15428 3724
rect 15820 3668 15876 3836
rect 15820 3602 15876 3612
rect 16156 2884 16212 8206
rect 16268 3556 16324 9772
rect 16380 9268 16436 9278
rect 16604 9268 16660 14112
rect 16828 13188 16884 14112
rect 16828 13122 16884 13132
rect 16716 12516 16772 12526
rect 16716 12402 16772 12460
rect 16716 12350 16718 12402
rect 16770 12350 16772 12402
rect 16716 12338 16772 12350
rect 17052 12404 17108 14112
rect 17164 13748 17220 13758
rect 17164 13300 17220 13692
rect 17276 13636 17332 14112
rect 17276 13570 17332 13580
rect 17164 13234 17220 13244
rect 17276 13412 17332 13422
rect 17052 12338 17108 12348
rect 17276 12178 17332 13356
rect 17388 13300 17444 13310
rect 17388 13186 17444 13244
rect 17388 13134 17390 13186
rect 17442 13134 17444 13186
rect 17388 13122 17444 13134
rect 17276 12126 17278 12178
rect 17330 12126 17332 12178
rect 17276 12114 17332 12126
rect 17388 12404 17444 12414
rect 16380 9266 16660 9268
rect 16380 9214 16382 9266
rect 16434 9214 16660 9266
rect 16380 9212 16660 9214
rect 16716 11508 16772 11518
rect 16380 9202 16436 9212
rect 16716 6468 16772 11452
rect 17164 11394 17220 11406
rect 17164 11342 17166 11394
rect 17218 11342 17220 11394
rect 16828 11284 16884 11294
rect 17164 11284 17220 11342
rect 16828 11282 17220 11284
rect 16828 11230 16830 11282
rect 16882 11230 17220 11282
rect 16828 11228 17220 11230
rect 16828 7588 16884 11228
rect 16940 10724 16996 10734
rect 16940 10610 16996 10668
rect 16940 10558 16942 10610
rect 16994 10558 16996 10610
rect 16940 10546 16996 10558
rect 17276 10500 17332 10510
rect 17276 10406 17332 10444
rect 17052 9826 17108 9838
rect 17052 9774 17054 9826
rect 17106 9774 17108 9826
rect 17052 9044 17108 9774
rect 17052 8978 17108 8988
rect 17164 9604 17220 9614
rect 16828 7522 16884 7532
rect 16940 8930 16996 8942
rect 16940 8878 16942 8930
rect 16994 8878 16996 8930
rect 16716 6402 16772 6412
rect 16380 6020 16436 6030
rect 16436 5964 16772 6020
rect 16380 5954 16436 5964
rect 16716 5012 16772 5964
rect 16940 5572 16996 8878
rect 17052 8820 17108 8830
rect 17052 7252 17108 8764
rect 17052 7186 17108 7196
rect 17164 7028 17220 9548
rect 17276 8930 17332 8942
rect 17276 8878 17278 8930
rect 17330 8878 17332 8930
rect 17276 8596 17332 8878
rect 17276 8530 17332 8540
rect 17164 6962 17220 6972
rect 17388 6804 17444 12348
rect 17500 12292 17556 14112
rect 17500 12226 17556 12236
rect 17612 12628 17668 12638
rect 17500 12068 17556 12078
rect 17500 10164 17556 12012
rect 17500 10098 17556 10108
rect 16940 5506 16996 5516
rect 17052 6748 17444 6804
rect 17052 5234 17108 6748
rect 17612 5348 17668 12572
rect 17724 11508 17780 14112
rect 17836 13636 17892 13646
rect 17836 12404 17892 13580
rect 17948 13188 18004 14112
rect 17948 13122 18004 13132
rect 17836 12338 17892 12348
rect 17948 12962 18004 12974
rect 17948 12910 17950 12962
rect 18002 12910 18004 12962
rect 17948 12180 18004 12910
rect 17948 12114 18004 12124
rect 17724 11452 18004 11508
rect 17724 11282 17780 11294
rect 17724 11230 17726 11282
rect 17778 11230 17780 11282
rect 17724 9268 17780 11230
rect 17724 9202 17780 9212
rect 17948 9154 18004 11452
rect 18060 11394 18116 11406
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18060 11284 18116 11342
rect 18060 11218 18116 11228
rect 18060 9716 18116 9726
rect 18172 9716 18228 14112
rect 18396 13748 18452 14112
rect 18396 13682 18452 13692
rect 18508 13188 18564 13198
rect 18396 12962 18452 12974
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18284 12404 18340 12414
rect 18284 12310 18340 12348
rect 18396 11508 18452 12910
rect 18396 11442 18452 11452
rect 18284 11396 18340 11406
rect 18284 10834 18340 11340
rect 18284 10782 18286 10834
rect 18338 10782 18340 10834
rect 18284 10770 18340 10782
rect 18396 11284 18452 11294
rect 18060 9714 18228 9716
rect 18060 9662 18062 9714
rect 18114 9662 18228 9714
rect 18060 9660 18228 9662
rect 18284 10500 18340 10510
rect 18060 9650 18116 9660
rect 18284 9380 18340 10444
rect 18284 9314 18340 9324
rect 17948 9102 17950 9154
rect 18002 9102 18004 9154
rect 17948 9090 18004 9102
rect 17724 8372 17780 8382
rect 17724 6916 17780 8316
rect 18396 8036 18452 11228
rect 18508 8146 18564 13132
rect 18620 11396 18676 14112
rect 18620 11330 18676 11340
rect 18732 13188 18788 13198
rect 18732 9156 18788 13132
rect 18844 12516 18900 14112
rect 18844 12450 18900 12460
rect 18844 12068 18900 12078
rect 18844 11974 18900 12012
rect 18844 11508 18900 11518
rect 18844 11414 18900 11452
rect 18956 11396 19012 11406
rect 18844 10948 18900 10958
rect 18844 10610 18900 10892
rect 18844 10558 18846 10610
rect 18898 10558 18900 10610
rect 18844 10546 18900 10558
rect 18732 9090 18788 9100
rect 18844 9940 18900 9950
rect 18844 8932 18900 9884
rect 18956 9716 19012 11340
rect 18956 9650 19012 9660
rect 19068 9266 19124 14112
rect 19180 12852 19236 12862
rect 19180 12758 19236 12796
rect 19292 10050 19348 14112
rect 19516 12404 19572 14112
rect 19516 12338 19572 12348
rect 19628 12292 19684 12302
rect 19740 12292 19796 14112
rect 19740 12236 19908 12292
rect 19628 12198 19684 12236
rect 19292 9998 19294 10050
rect 19346 9998 19348 10050
rect 19292 9986 19348 9998
rect 19740 11394 19796 11406
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19068 9214 19070 9266
rect 19122 9214 19124 9266
rect 19068 9202 19124 9214
rect 18508 8094 18510 8146
rect 18562 8094 18564 8146
rect 18508 8082 18564 8094
rect 18732 8876 18900 8932
rect 19404 9156 19460 9166
rect 17948 7980 18452 8036
rect 17948 7140 18004 7980
rect 18396 7812 18452 7822
rect 17948 7074 18004 7084
rect 18060 7364 18116 7374
rect 17724 6860 18004 6916
rect 17724 6468 17780 6478
rect 17724 6020 17780 6412
rect 17724 5954 17780 5964
rect 17836 5348 17892 5358
rect 17612 5346 17892 5348
rect 17612 5294 17614 5346
rect 17666 5294 17838 5346
rect 17890 5294 17892 5346
rect 17612 5292 17892 5294
rect 17612 5282 17668 5292
rect 17836 5282 17892 5292
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 16716 4946 16772 4956
rect 16940 5124 16996 5134
rect 16268 3490 16324 3500
rect 16156 2818 16212 2828
rect 16828 2884 16884 2894
rect 16828 2790 16884 2828
rect 15372 2258 15428 2268
rect 16716 2548 16772 2558
rect 14252 2034 14308 2044
rect 13468 1988 13524 1998
rect 13356 1764 13412 1774
rect 13356 1540 13412 1708
rect 13356 1474 13412 1484
rect 13468 1428 13524 1932
rect 13468 1362 13524 1372
rect 13916 1876 13972 1886
rect 12684 354 12740 364
rect 13916 112 13972 1820
rect 14476 1874 14532 1886
rect 14476 1822 14478 1874
rect 14530 1822 14532 1874
rect 14476 1316 14532 1822
rect 14476 1250 14532 1260
rect 16380 1652 16436 1662
rect 16380 112 16436 1596
rect 16716 532 16772 2492
rect 16940 2212 16996 5068
rect 17276 4116 17332 4126
rect 17164 4004 17220 4014
rect 17164 3668 17220 3948
rect 17164 3602 17220 3612
rect 16940 2146 16996 2156
rect 17164 3220 17220 3230
rect 17164 1988 17220 3164
rect 17276 1988 17332 4060
rect 17948 4116 18004 6860
rect 18060 5460 18116 7308
rect 18396 6468 18452 7756
rect 18508 7586 18564 7598
rect 18508 7534 18510 7586
rect 18562 7534 18564 7586
rect 18508 7252 18564 7534
rect 18508 7186 18564 7196
rect 18732 6916 18788 8876
rect 19404 8370 19460 9100
rect 19404 8318 19406 8370
rect 19458 8318 19460 8370
rect 19404 8306 19460 8318
rect 19628 7588 19684 7598
rect 18956 7250 19012 7262
rect 18956 7198 18958 7250
rect 19010 7198 19012 7250
rect 18956 7140 19012 7198
rect 18956 7074 19012 7084
rect 19292 7250 19348 7262
rect 19292 7198 19294 7250
rect 19346 7198 19348 7250
rect 19292 7140 19348 7198
rect 19628 7140 19684 7532
rect 19292 7074 19348 7084
rect 19404 7084 19684 7140
rect 18732 6850 18788 6860
rect 19180 6916 19236 6926
rect 18732 6692 18788 6702
rect 18732 6598 18788 6636
rect 18396 6402 18452 6412
rect 18060 5394 18116 5404
rect 18284 5348 18340 5358
rect 17948 4050 18004 4060
rect 18060 4564 18116 4574
rect 18060 3780 18116 4508
rect 18284 4564 18340 5292
rect 18508 5348 18564 5358
rect 18508 4788 18564 5292
rect 18508 4722 18564 4732
rect 18284 4498 18340 4508
rect 18060 3714 18116 3724
rect 18620 4004 18676 4014
rect 18284 3332 18340 3342
rect 17388 2548 17444 2558
rect 17612 2548 17668 2558
rect 17388 2546 17668 2548
rect 17388 2494 17390 2546
rect 17442 2494 17614 2546
rect 17666 2494 17668 2546
rect 17388 2492 17668 2494
rect 17388 2482 17444 2492
rect 17388 1988 17444 1998
rect 17276 1932 17388 1988
rect 17164 1922 17220 1932
rect 17388 1922 17444 1932
rect 17612 644 17668 2492
rect 18284 1988 18340 3276
rect 18284 1922 18340 1932
rect 18620 1652 18676 3948
rect 19180 3388 19236 6860
rect 19292 6692 19348 6702
rect 19404 6692 19460 7084
rect 19292 6690 19460 6692
rect 19292 6638 19294 6690
rect 19346 6638 19460 6690
rect 19292 6636 19460 6638
rect 19628 6690 19684 7084
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19292 6626 19348 6636
rect 19628 6626 19684 6638
rect 19740 3666 19796 11342
rect 19852 10834 19908 12236
rect 19964 11508 20020 14112
rect 20188 13300 20244 14112
rect 20188 13234 20244 13244
rect 20300 13748 20356 13758
rect 20300 12628 20356 13692
rect 19964 11442 20020 11452
rect 20188 12572 20356 12628
rect 20188 11282 20244 12572
rect 20300 12180 20356 12190
rect 20300 11732 20356 12124
rect 20300 11666 20356 11676
rect 20412 11638 20468 14112
rect 20636 12292 20692 14112
rect 20748 13300 20804 13310
rect 20860 13300 20916 14112
rect 21084 13748 21140 14112
rect 21084 13682 21140 13692
rect 20804 13244 20916 13300
rect 20748 13234 20804 13244
rect 21196 13188 21252 13198
rect 21196 13094 21252 13132
rect 21308 12852 21364 14112
rect 21308 12786 21364 12796
rect 21420 13748 21476 13758
rect 20636 12236 20804 12292
rect 20748 12068 20804 12236
rect 20860 12180 20916 12190
rect 21084 12180 21140 12190
rect 20860 12178 21084 12180
rect 20860 12126 20862 12178
rect 20914 12126 21084 12178
rect 20860 12124 21084 12126
rect 20860 12114 20916 12124
rect 21084 12114 21140 12124
rect 20636 12012 20804 12068
rect 20636 11844 20692 12012
rect 21308 11956 21364 11966
rect 21196 11844 21252 11854
rect 20636 11788 20916 11844
rect 20412 11582 20804 11638
rect 20188 11230 20190 11282
rect 20242 11230 20244 11282
rect 20188 11218 20244 11230
rect 19852 10782 19854 10834
rect 19906 10782 19908 10834
rect 19852 10770 19908 10782
rect 20076 10164 20132 10174
rect 20076 10018 20132 10108
rect 20076 9962 20244 10018
rect 19852 9828 19908 9838
rect 19852 9734 19908 9772
rect 19964 9044 20020 9054
rect 19740 3614 19742 3666
rect 19794 3614 19796 3666
rect 19740 3602 19796 3614
rect 19852 7476 19908 7486
rect 19852 3388 19908 7420
rect 19964 6804 20020 8988
rect 20076 8930 20132 8942
rect 20076 8878 20078 8930
rect 20130 8878 20132 8930
rect 20076 8372 20132 8878
rect 20076 8306 20132 8316
rect 20188 8036 20244 9962
rect 20748 9268 20804 11582
rect 20860 10050 20916 11788
rect 20860 9998 20862 10050
rect 20914 9998 20916 10050
rect 20860 9986 20916 9998
rect 20972 11788 21196 11844
rect 20860 9268 20916 9278
rect 20748 9266 20916 9268
rect 20748 9214 20862 9266
rect 20914 9214 20916 9266
rect 20748 9212 20916 9214
rect 20860 9202 20916 9212
rect 20972 8596 21028 11788
rect 21196 11778 21252 11788
rect 21196 11396 21252 11406
rect 21196 11302 21252 11340
rect 21308 11060 21364 11900
rect 20972 8530 21028 8540
rect 21084 11004 21364 11060
rect 20972 8372 21028 8382
rect 20972 8278 21028 8316
rect 20188 7970 20244 7980
rect 21084 7700 21140 11004
rect 21308 10500 21364 10510
rect 21308 10406 21364 10444
rect 21420 10052 21476 13692
rect 21532 11732 21588 14112
rect 21756 13188 21812 14112
rect 21756 13132 21924 13188
rect 21756 12962 21812 12974
rect 21756 12910 21758 12962
rect 21810 12910 21812 12962
rect 21644 12404 21700 12414
rect 21644 12310 21700 12348
rect 21532 11666 21588 11676
rect 21644 12180 21700 12190
rect 21644 11508 21700 12124
rect 21308 9996 21476 10052
rect 21532 11452 21700 11508
rect 21196 8372 21252 8382
rect 21196 7924 21252 8316
rect 21196 7858 21252 7868
rect 20412 7644 21140 7700
rect 20412 7476 20468 7644
rect 21308 7588 21364 9996
rect 21308 7522 21364 7532
rect 21420 9826 21476 9838
rect 21420 9774 21422 9826
rect 21474 9774 21476 9826
rect 20412 7410 20468 7420
rect 20636 7476 20692 7486
rect 19964 6738 20020 6748
rect 20188 6580 20244 6590
rect 19180 3332 19460 3388
rect 19852 3332 20020 3388
rect 18956 2996 19012 3006
rect 18956 2098 19012 2940
rect 18956 2046 18958 2098
rect 19010 2046 19012 2098
rect 18956 2034 19012 2046
rect 19180 2996 19236 3006
rect 18620 1586 18676 1596
rect 17612 578 17668 588
rect 18844 1540 18900 1550
rect 16716 466 16772 476
rect 18844 112 18900 1484
rect 19180 1428 19236 2940
rect 19404 1652 19460 3332
rect 19516 3220 19572 3230
rect 19516 2772 19572 3164
rect 19516 2706 19572 2716
rect 19516 2212 19572 2222
rect 19516 2118 19572 2156
rect 19852 2212 19908 2222
rect 19852 2118 19908 2156
rect 19964 1988 20020 3332
rect 20076 2772 20132 2782
rect 20076 2548 20132 2716
rect 20076 2482 20132 2492
rect 20188 2098 20244 6524
rect 20300 3780 20356 3790
rect 20636 3780 20692 7420
rect 20972 6132 21028 6142
rect 20300 3778 20692 3780
rect 20300 3726 20302 3778
rect 20354 3726 20638 3778
rect 20690 3726 20692 3778
rect 20300 3724 20692 3726
rect 20300 3714 20356 3724
rect 20636 3714 20692 3724
rect 20748 5796 20804 5806
rect 20748 2436 20804 5740
rect 20860 5684 20916 5694
rect 20860 3668 20916 5628
rect 20972 3892 21028 6076
rect 21420 5796 21476 9774
rect 21532 9716 21588 11452
rect 21644 10836 21700 10846
rect 21644 9940 21700 10780
rect 21756 10052 21812 12910
rect 21868 10834 21924 13132
rect 21980 11506 22036 14112
rect 21980 11454 21982 11506
rect 22034 11454 22036 11506
rect 21980 11442 22036 11454
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 21868 10782 21870 10834
rect 21922 10782 21924 10834
rect 21868 10770 21924 10782
rect 21756 9996 21924 10052
rect 21644 9874 21700 9884
rect 21532 9660 21700 9716
rect 21532 8260 21588 8270
rect 21532 8166 21588 8204
rect 21420 5730 21476 5740
rect 21532 8036 21588 8046
rect 21308 5124 21364 5134
rect 21364 5068 21476 5124
rect 21308 5058 21364 5068
rect 20972 3826 21028 3836
rect 21084 4564 21140 4574
rect 20860 3602 20916 3612
rect 20188 2046 20190 2098
rect 20242 2046 20244 2098
rect 20188 2034 20244 2046
rect 20412 2380 20804 2436
rect 19404 1586 19460 1596
rect 19852 1932 20020 1988
rect 19180 1362 19236 1372
rect 19852 308 19908 1932
rect 20188 1428 20244 1438
rect 19964 980 20020 990
rect 20188 980 20244 1372
rect 20412 1314 20468 2380
rect 20748 2212 20804 2222
rect 21084 2212 21140 4508
rect 20748 2210 21140 2212
rect 20748 2158 20750 2210
rect 20802 2158 21086 2210
rect 21138 2158 21140 2210
rect 20748 2156 21140 2158
rect 20748 2146 20804 2156
rect 21084 2146 21140 2156
rect 21196 4228 21252 4238
rect 20412 1262 20414 1314
rect 20466 1262 20468 1314
rect 20412 1250 20468 1262
rect 20860 1204 20916 1214
rect 20860 1110 20916 1148
rect 21084 1204 21140 1214
rect 21084 1110 21140 1148
rect 20020 924 20244 980
rect 19964 914 20020 924
rect 21196 756 21252 4172
rect 21420 4228 21476 5068
rect 21420 4162 21476 4172
rect 21308 3668 21364 3678
rect 21308 2996 21364 3612
rect 21308 2930 21364 2940
rect 21532 1876 21588 7980
rect 21644 2212 21700 9660
rect 21756 9042 21812 9054
rect 21756 8990 21758 9042
rect 21810 8990 21812 9042
rect 21756 5012 21812 8990
rect 21868 8596 21924 9996
rect 21868 8530 21924 8540
rect 21980 9826 22036 9838
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21868 8146 21924 8158
rect 21868 8094 21870 8146
rect 21922 8094 21924 8146
rect 21868 8036 21924 8094
rect 21868 7970 21924 7980
rect 21868 7588 21924 7598
rect 21868 7494 21924 7532
rect 21756 4946 21812 4956
rect 21868 7140 21924 7150
rect 21756 4676 21812 4686
rect 21756 2996 21812 4620
rect 21868 4116 21924 7084
rect 21980 6580 22036 9774
rect 22092 9118 22148 12910
rect 22204 12404 22260 14112
rect 22428 13188 22484 14112
rect 22428 13122 22484 13132
rect 22540 13524 22596 13534
rect 22204 12338 22260 12348
rect 22428 12740 22484 12750
rect 22316 11732 22372 11742
rect 22204 11620 22260 11630
rect 22204 9716 22260 11564
rect 22316 10050 22372 11676
rect 22316 9998 22318 10050
rect 22370 9998 22372 10050
rect 22316 9986 22372 9998
rect 22204 9650 22260 9660
rect 22092 9062 22372 9118
rect 22204 8932 22260 8942
rect 22204 8838 22260 8876
rect 22092 8820 22148 8830
rect 22092 8260 22148 8764
rect 22092 7588 22148 8204
rect 22092 7522 22148 7532
rect 22204 8036 22260 8046
rect 21980 6514 22036 6524
rect 22092 6692 22148 6702
rect 21868 4050 21924 4060
rect 21756 2930 21812 2940
rect 21756 2436 21812 2446
rect 21812 2380 21924 2436
rect 21756 2370 21812 2380
rect 21644 2146 21700 2156
rect 21532 1810 21588 1820
rect 21196 690 21252 700
rect 21308 1652 21364 1662
rect 19852 242 19908 252
rect 21308 112 21364 1596
rect 21532 1652 21588 1662
rect 21532 1428 21588 1596
rect 21532 1362 21588 1372
rect 21868 1428 21924 2380
rect 22092 2212 22148 6636
rect 22204 5124 22260 7980
rect 22316 6356 22372 9062
rect 22428 8482 22484 12684
rect 22540 10612 22596 13468
rect 22652 10836 22708 14112
rect 22876 13748 22932 14112
rect 22764 13692 22932 13748
rect 22764 11620 22820 13692
rect 22876 13524 22932 13534
rect 22876 13074 22932 13468
rect 22876 13022 22878 13074
rect 22930 13022 22932 13074
rect 22876 13010 22932 13022
rect 22876 12404 22932 12414
rect 23100 12404 23156 14112
rect 23324 13524 23380 14112
rect 23324 13458 23380 13468
rect 22876 12402 23156 12404
rect 22876 12350 22878 12402
rect 22930 12350 23156 12402
rect 22876 12348 23156 12350
rect 23324 12404 23380 12414
rect 23380 12348 23492 12404
rect 22876 12338 22932 12348
rect 23324 12338 23380 12348
rect 23212 12178 23268 12190
rect 23212 12126 23214 12178
rect 23266 12126 23268 12178
rect 22764 11554 22820 11564
rect 22988 11956 23044 11966
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 11284 22820 11342
rect 22764 11218 22820 11228
rect 22652 10770 22708 10780
rect 22876 11060 22932 11070
rect 22540 10556 22820 10612
rect 22428 8430 22430 8482
rect 22482 8430 22484 8482
rect 22428 8418 22484 8430
rect 22540 10164 22596 10174
rect 22428 8260 22484 8270
rect 22428 8166 22484 8204
rect 22316 6290 22372 6300
rect 22428 7924 22484 7934
rect 22428 5158 22484 7868
rect 22540 5234 22596 10108
rect 22764 10164 22820 10556
rect 22876 10610 22932 11004
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22876 10546 22932 10558
rect 22764 10098 22820 10108
rect 22988 9156 23044 11900
rect 23212 9940 23268 12126
rect 23324 11620 23380 11630
rect 23324 11526 23380 11564
rect 23436 11284 23492 12348
rect 23548 12292 23604 14112
rect 23772 12740 23828 14112
rect 23996 13188 24052 14112
rect 24220 13412 24276 14112
rect 24444 13524 24500 14112
rect 24220 13346 24276 13356
rect 24332 13468 24500 13524
rect 24668 13524 24724 14112
rect 24892 13748 24948 14112
rect 24892 13682 24948 13692
rect 25116 13636 25172 14112
rect 25116 13570 25172 13580
rect 25340 13636 25396 14112
rect 25340 13570 25396 13580
rect 25564 13524 25620 14112
rect 24668 13468 24948 13524
rect 24332 13300 24388 13468
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24332 13234 24388 13244
rect 23996 13122 24052 13132
rect 24892 13076 24948 13468
rect 25564 13458 25620 13468
rect 25676 13748 25732 13758
rect 24444 13020 24948 13076
rect 25004 13132 25228 13188
rect 24220 12740 24276 12750
rect 23772 12738 24276 12740
rect 23772 12686 24222 12738
rect 24274 12686 24276 12738
rect 23772 12684 24276 12686
rect 24220 12674 24276 12684
rect 23660 12628 23716 12638
rect 24444 12628 24500 13020
rect 23660 12404 23716 12572
rect 23804 12572 24068 12582
rect 24444 12572 24724 12628
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 24556 12404 24612 12414
rect 23660 12348 24556 12404
rect 24556 12338 24612 12348
rect 23548 12236 24388 12292
rect 23772 12066 23828 12078
rect 23772 12014 23774 12066
rect 23826 12014 23828 12066
rect 23772 11844 23828 12014
rect 24332 11954 24388 12236
rect 24332 11902 24334 11954
rect 24386 11902 24388 11954
rect 24332 11890 24388 11902
rect 24668 11956 24724 12572
rect 24668 11890 24724 11900
rect 23772 11778 23828 11788
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24668 11284 24724 11294
rect 23436 11228 24388 11284
rect 23660 11116 24276 11172
rect 23660 11060 23716 11116
rect 24220 11060 24276 11116
rect 23660 10994 23716 11004
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24220 10994 24276 11004
rect 23804 10938 24068 10948
rect 24332 10948 24388 11228
rect 24668 11190 24724 11228
rect 24332 10882 24388 10892
rect 23436 10836 23492 10846
rect 23436 10742 23492 10780
rect 23212 9874 23268 9884
rect 23436 10500 23492 10510
rect 22764 9154 23044 9156
rect 22764 9102 22990 9154
rect 23042 9102 23044 9154
rect 22764 9100 23044 9102
rect 22764 9042 22820 9100
rect 22988 9090 23044 9100
rect 23212 9380 23268 9390
rect 22764 8990 22766 9042
rect 22818 8990 22820 9042
rect 22764 8978 22820 8990
rect 22876 8596 22932 8606
rect 22764 8260 22820 8270
rect 22764 8166 22820 8204
rect 22876 6578 22932 8540
rect 23212 8260 23268 9324
rect 23212 8194 23268 8204
rect 23436 7924 23492 10444
rect 24108 10332 24948 10388
rect 24108 10276 24164 10332
rect 24108 10210 24164 10220
rect 24464 10220 24728 10230
rect 24332 10164 24388 10174
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24332 9380 24388 10108
rect 24556 9940 24612 9950
rect 24556 9846 24612 9884
rect 24892 9940 24948 10332
rect 25004 10276 25060 13132
rect 25172 13086 25228 13132
rect 25172 13074 25284 13086
rect 25172 13022 25230 13074
rect 25282 13022 25284 13074
rect 25172 13020 25284 13022
rect 25228 13010 25284 13020
rect 25564 12852 25620 12862
rect 25172 12796 25564 12852
rect 25172 12628 25228 12796
rect 25564 12786 25620 12796
rect 25116 12572 25228 12628
rect 25116 11732 25172 12572
rect 25452 12404 25508 12414
rect 25676 12404 25732 13692
rect 25452 12180 25508 12348
rect 25452 12114 25508 12124
rect 25564 12348 25732 12404
rect 25116 11666 25172 11676
rect 25116 11394 25172 11406
rect 25116 11342 25118 11394
rect 25170 11342 25172 11394
rect 25116 11284 25172 11342
rect 25340 11284 25396 11294
rect 25116 11282 25396 11284
rect 25116 11230 25342 11282
rect 25394 11230 25396 11282
rect 25116 11228 25396 11230
rect 25340 10836 25396 11228
rect 25340 10770 25396 10780
rect 25564 10500 25620 12348
rect 25564 10434 25620 10444
rect 25676 12180 25732 12190
rect 25004 10210 25060 10220
rect 24892 9874 24948 9884
rect 25116 9826 25172 9838
rect 25116 9774 25118 9826
rect 25170 9774 25172 9826
rect 25116 9716 25172 9774
rect 25116 9650 25172 9660
rect 25452 9716 25508 9726
rect 25452 9622 25508 9660
rect 24332 9314 24388 9324
rect 25004 9380 25060 9390
rect 25060 9324 25508 9380
rect 25004 9314 25060 9324
rect 25340 9156 25396 9166
rect 23772 9044 23828 9054
rect 23772 8950 23828 8988
rect 24332 9044 24388 9054
rect 24332 8950 24388 8988
rect 24556 9044 24612 9054
rect 23996 8932 24052 8942
rect 23996 8818 24052 8876
rect 24556 8820 24612 8988
rect 24892 8932 24948 8942
rect 25228 8932 25284 8942
rect 24892 8930 25060 8932
rect 24892 8878 24894 8930
rect 24946 8878 25060 8930
rect 24892 8876 25060 8878
rect 24892 8866 24948 8876
rect 23996 8766 23998 8818
rect 24050 8766 24052 8818
rect 23996 8708 24052 8766
rect 23996 8642 24052 8652
rect 24332 8764 24612 8820
rect 24332 8596 24388 8764
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24332 8530 24388 8540
rect 24892 8258 24948 8270
rect 24892 8206 24894 8258
rect 24946 8206 24948 8258
rect 24668 8148 24724 8158
rect 24892 8148 24948 8206
rect 24668 8146 24948 8148
rect 24668 8094 24670 8146
rect 24722 8094 24948 8146
rect 24668 8092 24948 8094
rect 24668 8036 24724 8092
rect 24668 7970 24724 7980
rect 24220 7924 24276 7934
rect 23436 7858 23492 7868
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 23324 7700 23380 7710
rect 23324 7586 23380 7644
rect 24108 7588 24164 7598
rect 23324 7534 23326 7586
rect 23378 7534 23380 7586
rect 23324 7522 23380 7534
rect 23884 7532 24108 7588
rect 23884 7474 23940 7532
rect 24108 7494 24164 7532
rect 23884 7422 23886 7474
rect 23938 7422 23940 7474
rect 23884 7410 23940 7422
rect 24108 7140 24164 7150
rect 22988 6916 23044 6926
rect 22988 6692 23044 6860
rect 23436 6916 23492 6926
rect 22988 6626 23044 6636
rect 23324 6690 23380 6702
rect 23324 6638 23326 6690
rect 23378 6638 23380 6690
rect 22876 6526 22878 6578
rect 22930 6526 22932 6578
rect 22876 6514 22932 6526
rect 23324 6468 23380 6638
rect 23324 6402 23380 6412
rect 23100 5348 23156 5358
rect 23436 5348 23492 6860
rect 23660 6578 23716 6590
rect 23660 6526 23662 6578
rect 23714 6526 23716 6578
rect 23660 6468 23716 6526
rect 24108 6468 24164 7084
rect 24220 7028 24276 7868
rect 25004 7140 25060 8876
rect 25228 8838 25284 8876
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 25004 7074 25060 7084
rect 25228 8260 25284 8270
rect 24464 7018 24728 7028
rect 24892 7028 24948 7038
rect 24220 6962 24276 6972
rect 24444 6468 24500 6478
rect 24108 6412 24444 6468
rect 23660 6402 23716 6412
rect 24444 6402 24500 6412
rect 23804 6300 24068 6310
rect 23660 6244 23716 6254
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 23660 6020 23716 6188
rect 23772 6020 23828 6030
rect 24556 6020 24612 6030
rect 23660 6018 23828 6020
rect 23660 5966 23774 6018
rect 23826 5966 23828 6018
rect 23660 5964 23828 5966
rect 23772 5954 23828 5964
rect 24332 5964 24556 6020
rect 24332 5906 24388 5964
rect 24556 5926 24612 5964
rect 24332 5854 24334 5906
rect 24386 5854 24388 5906
rect 24332 5842 24388 5854
rect 23100 5346 23492 5348
rect 23100 5294 23102 5346
rect 23154 5294 23438 5346
rect 23490 5294 23492 5346
rect 23100 5292 23492 5294
rect 24332 5572 24388 5582
rect 24332 5348 24388 5516
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24892 5348 24948 6972
rect 24332 5292 24500 5348
rect 23100 5282 23156 5292
rect 23436 5282 23492 5292
rect 22540 5182 22542 5234
rect 22594 5182 22596 5234
rect 22540 5170 22596 5182
rect 22204 5058 22260 5068
rect 22316 5102 22484 5158
rect 23212 5124 23268 5134
rect 22316 3388 22372 5102
rect 22652 5012 22708 5022
rect 22092 2146 22148 2156
rect 22204 3332 22372 3388
rect 22540 4228 22596 4238
rect 22204 1652 22260 3332
rect 22204 1586 22260 1596
rect 22540 1652 22596 4172
rect 22652 3444 22708 4956
rect 23212 3388 23268 5068
rect 23660 4844 24388 4900
rect 23660 4788 23716 4844
rect 24332 4788 24388 4844
rect 23660 4722 23716 4732
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24332 4722 24388 4732
rect 23804 4666 24068 4676
rect 24220 4676 24276 4686
rect 24220 4004 24276 4620
rect 24444 4228 24500 5292
rect 24668 5292 24948 5348
rect 25004 6804 25060 6814
rect 24556 5124 24612 5134
rect 24556 5030 24612 5068
rect 24668 4452 24724 5292
rect 24892 5124 24948 5134
rect 24892 5030 24948 5068
rect 24780 4788 24836 4798
rect 24780 4564 24836 4732
rect 25004 4788 25060 6748
rect 25228 5796 25284 8204
rect 25228 5730 25284 5740
rect 25340 5348 25396 9100
rect 25452 8932 25508 9324
rect 25452 8866 25508 8876
rect 25452 8260 25508 8270
rect 25452 8166 25508 8204
rect 25452 7812 25508 7822
rect 25452 6692 25508 7756
rect 25676 7588 25732 12124
rect 25788 11060 25844 14112
rect 25900 13860 25956 13870
rect 25900 11732 25956 13804
rect 26012 12404 26068 14112
rect 26012 12338 26068 12348
rect 25900 11666 25956 11676
rect 25788 10994 25844 11004
rect 25900 11396 25956 11406
rect 25900 10500 25956 11340
rect 25900 10434 25956 10444
rect 26124 10386 26180 10398
rect 26124 10334 26126 10386
rect 26178 10334 26180 10386
rect 26124 10164 26180 10334
rect 26124 10098 26180 10108
rect 26124 9604 26180 9614
rect 25788 9156 25844 9166
rect 25788 9062 25844 9100
rect 25788 8932 25844 8942
rect 25788 7812 25844 8876
rect 25788 7746 25844 7756
rect 25676 7522 25732 7532
rect 25452 6626 25508 6636
rect 25340 5282 25396 5292
rect 25452 5012 25508 5022
rect 25452 4918 25508 4956
rect 25004 4722 25060 4732
rect 24780 4508 25956 4564
rect 24668 4386 24724 4396
rect 24444 4172 25284 4228
rect 24892 4004 24948 4014
rect 24220 3938 24276 3948
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 22652 3378 22708 3388
rect 22540 1586 22596 1596
rect 23100 3332 23268 3388
rect 24220 3780 24276 3790
rect 23884 3332 23940 3342
rect 23100 1540 23156 3332
rect 23660 3276 23884 3332
rect 23660 3220 23716 3276
rect 23884 3266 23940 3276
rect 23660 3154 23716 3164
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24220 2212 24276 3724
rect 24332 3556 24388 3566
rect 24892 3556 24948 3948
rect 25116 3780 25172 3818
rect 25116 3714 25172 3724
rect 24332 3332 24388 3500
rect 24780 3500 24948 3556
rect 25228 3556 25284 4172
rect 25340 3780 25396 3790
rect 25340 3686 25396 3724
rect 24668 3444 24724 3454
rect 24780 3444 24836 3500
rect 25228 3490 25284 3500
rect 25452 3668 25508 3678
rect 24668 3442 24836 3444
rect 24668 3390 24670 3442
rect 24722 3390 24836 3442
rect 24668 3388 24836 3390
rect 24668 3378 24724 3388
rect 24444 3332 24500 3342
rect 24332 3276 24444 3332
rect 24444 3266 24500 3276
rect 25340 3332 25396 3342
rect 25452 3332 25508 3612
rect 25396 3276 25508 3332
rect 25340 3266 25396 3276
rect 24892 3220 24948 3230
rect 24332 3108 24388 3118
rect 24332 2436 24388 3052
rect 24892 2436 24948 3164
rect 24332 2370 24388 2380
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24892 2370 24948 2380
rect 25788 3220 25844 3230
rect 24464 2314 24728 2324
rect 24220 2156 24948 2212
rect 23660 1708 24500 1764
rect 23660 1652 23716 1708
rect 23660 1586 23716 1596
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 24220 1540 24276 1550
rect 23100 1474 23156 1484
rect 21868 1362 21924 1372
rect 24220 980 24276 1484
rect 23324 924 24276 980
rect 24444 980 24500 1708
rect 24780 1652 24836 1662
rect 24892 1652 24948 2156
rect 25788 2100 25844 3164
rect 25900 3108 25956 4508
rect 26124 4452 26180 9548
rect 26236 5572 26292 14112
rect 26348 13188 26404 13198
rect 26348 12292 26404 13132
rect 26460 12740 26516 14112
rect 26460 12674 26516 12684
rect 26684 12404 26740 14112
rect 26684 12348 26852 12404
rect 26348 12290 26740 12292
rect 26348 12238 26350 12290
rect 26402 12238 26740 12290
rect 26348 12236 26740 12238
rect 26348 12226 26404 12236
rect 26684 12178 26740 12236
rect 26684 12126 26686 12178
rect 26738 12126 26740 12178
rect 26684 12114 26740 12126
rect 26796 11844 26852 12348
rect 26572 11788 26852 11844
rect 26460 11396 26516 11406
rect 26348 10386 26404 10398
rect 26348 10334 26350 10386
rect 26402 10334 26404 10386
rect 26348 10052 26404 10334
rect 26348 9986 26404 9996
rect 26348 9828 26404 9838
rect 26348 9714 26404 9772
rect 26348 9662 26350 9714
rect 26402 9662 26404 9714
rect 26348 9650 26404 9662
rect 26460 6020 26516 11340
rect 26572 9604 26628 11788
rect 26908 11620 26964 14112
rect 27132 12852 27188 14112
rect 27356 12964 27412 14112
rect 27580 13188 27636 14112
rect 27580 13122 27636 13132
rect 27356 12908 27636 12964
rect 27132 12796 27524 12852
rect 27132 12628 27188 12638
rect 27132 12290 27188 12572
rect 27132 12238 27134 12290
rect 27186 12238 27188 12290
rect 27132 12226 27188 12238
rect 26908 11618 27300 11620
rect 26908 11566 26910 11618
rect 26962 11566 27300 11618
rect 26908 11564 27300 11566
rect 26908 11554 26964 11564
rect 26796 10724 26852 10734
rect 26572 9538 26628 9548
rect 26684 10722 26852 10724
rect 26684 10670 26798 10722
rect 26850 10670 26852 10722
rect 26684 10668 26852 10670
rect 26460 5954 26516 5964
rect 26572 8820 26628 8830
rect 26236 5506 26292 5516
rect 26572 5236 26628 8764
rect 26684 8260 26740 10668
rect 26796 10658 26852 10668
rect 27244 10610 27300 11564
rect 27244 10558 27246 10610
rect 27298 10558 27300 10610
rect 27244 10546 27300 10558
rect 27356 11172 27412 11182
rect 27356 10052 27412 11116
rect 27020 10050 27412 10052
rect 27020 9998 27358 10050
rect 27410 9998 27412 10050
rect 27020 9996 27412 9998
rect 26796 9828 26852 9838
rect 26796 9734 26852 9772
rect 27020 9154 27076 9996
rect 27356 9986 27412 9996
rect 27132 9828 27188 9838
rect 27132 9734 27188 9772
rect 27020 9102 27022 9154
rect 27074 9102 27076 9154
rect 27020 9090 27076 9102
rect 27132 8932 27188 8942
rect 26684 8194 26740 8204
rect 26908 8596 26964 8606
rect 26908 5908 26964 8540
rect 26572 5170 26628 5180
rect 26684 5852 26964 5908
rect 26124 4450 26516 4452
rect 26124 4398 26126 4450
rect 26178 4398 26516 4450
rect 26124 4396 26516 4398
rect 26124 4386 26180 4396
rect 26460 4338 26516 4396
rect 26460 4286 26462 4338
rect 26514 4286 26516 4338
rect 26460 4274 26516 4286
rect 26124 4116 26180 4126
rect 26012 3108 26068 3118
rect 25900 3052 26012 3108
rect 26012 3042 26068 3052
rect 25788 2034 25844 2044
rect 25228 1876 25284 1886
rect 25004 1652 25060 1662
rect 24892 1596 25004 1652
rect 24780 1428 24836 1596
rect 25004 1586 25060 1596
rect 25228 1540 25284 1820
rect 26124 1876 26180 4060
rect 26124 1810 26180 1820
rect 26348 4116 26404 4126
rect 25228 1474 25284 1484
rect 24780 1372 25172 1428
rect 24444 924 24948 980
rect 22540 756 22596 766
rect 22764 756 22820 766
rect 22540 420 22596 700
rect 22540 354 22596 364
rect 22652 700 22764 756
rect 22316 308 22372 318
rect 22316 196 22372 252
rect 22652 196 22708 700
rect 22764 690 22820 700
rect 22876 532 22932 542
rect 22876 308 22932 476
rect 23324 420 23380 924
rect 24332 868 24388 878
rect 23212 364 23380 420
rect 23996 756 24052 766
rect 23212 308 23268 364
rect 22876 252 23268 308
rect 22316 140 22708 196
rect 23772 196 23828 206
rect 23772 112 23828 140
rect 23996 196 24052 700
rect 24332 532 24388 812
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24892 756 24948 924
rect 25116 868 25172 1372
rect 26348 1204 26404 4060
rect 26684 2884 26740 5852
rect 27132 4788 27188 8876
rect 27356 6356 27412 6366
rect 27356 6020 27412 6300
rect 27356 5954 27412 5964
rect 26908 4732 27188 4788
rect 27356 5684 27412 5694
rect 26908 4564 26964 4732
rect 26908 4498 26964 4508
rect 27132 4564 27188 4574
rect 27020 4452 27076 4462
rect 27020 4358 27076 4396
rect 27132 4228 27188 4508
rect 26908 4172 27188 4228
rect 26796 3556 26852 3566
rect 26796 2996 26852 3500
rect 26796 2930 26852 2940
rect 26684 2818 26740 2828
rect 26460 2772 26516 2782
rect 26460 2436 26516 2716
rect 26908 2436 26964 4172
rect 27244 3444 27300 3482
rect 27244 3378 27300 3388
rect 27356 2996 27412 5628
rect 27468 3556 27524 12796
rect 27580 11508 27636 12908
rect 27804 12180 27860 14112
rect 28028 14084 28084 14112
rect 28028 14018 28084 14028
rect 28140 13636 28196 13646
rect 28140 12628 28196 13580
rect 28140 12562 28196 12572
rect 28140 12404 28196 12414
rect 28028 12292 28084 12302
rect 28028 12198 28084 12236
rect 27804 12114 27860 12124
rect 27580 11442 27636 11452
rect 27804 11844 27860 11854
rect 27804 11508 27860 11788
rect 27804 11442 27860 11452
rect 28028 11844 28084 11854
rect 27916 11394 27972 11406
rect 27916 11342 27918 11394
rect 27970 11342 27972 11394
rect 27580 11284 27636 11294
rect 27916 11284 27972 11342
rect 27580 11282 27972 11284
rect 27580 11230 27582 11282
rect 27634 11230 27972 11282
rect 27580 11228 27972 11230
rect 27580 6244 27636 11228
rect 27804 10498 27860 10510
rect 27804 10446 27806 10498
rect 27858 10446 27860 10498
rect 27804 10388 27860 10446
rect 27804 10322 27860 10332
rect 27804 10164 27860 10174
rect 27580 6178 27636 6188
rect 27692 9938 27748 9950
rect 27692 9886 27694 9938
rect 27746 9886 27748 9938
rect 27692 5684 27748 9886
rect 27804 6468 27860 10108
rect 27804 6402 27860 6412
rect 28028 6132 28084 11788
rect 28140 9828 28196 12348
rect 28140 9762 28196 9772
rect 28028 6066 28084 6076
rect 27692 5618 27748 5628
rect 27692 3556 27748 3566
rect 28028 3556 28084 3566
rect 27468 3554 28084 3556
rect 27468 3502 27694 3554
rect 27746 3502 28030 3554
rect 28082 3502 28084 3554
rect 27468 3500 28084 3502
rect 27692 3490 27748 3500
rect 28028 3490 28084 3500
rect 28252 3388 28308 14112
rect 28476 12516 28532 14112
rect 28700 13300 28756 14112
rect 28700 13234 28756 13244
rect 28924 12516 28980 14112
rect 28364 12460 28532 12516
rect 28588 12460 28980 12516
rect 28364 6916 28420 12460
rect 28476 12292 28532 12302
rect 28476 12178 28532 12236
rect 28476 12126 28478 12178
rect 28530 12126 28532 12178
rect 28476 12114 28532 12126
rect 28476 11282 28532 11294
rect 28476 11230 28478 11282
rect 28530 11230 28532 11282
rect 28476 10836 28532 11230
rect 28476 10770 28532 10780
rect 28588 8596 28644 12460
rect 28924 12290 28980 12302
rect 28924 12238 28926 12290
rect 28978 12238 28980 12290
rect 28588 8530 28644 8540
rect 28700 12180 28756 12190
rect 28700 8148 28756 12124
rect 28700 8082 28756 8092
rect 28812 9940 28868 9950
rect 28364 6850 28420 6860
rect 28812 4116 28868 9884
rect 28924 7364 28980 12238
rect 29148 11844 29204 14112
rect 29372 12180 29428 14112
rect 29372 12124 29540 12180
rect 29148 11778 29204 11788
rect 29372 11954 29428 11966
rect 29372 11902 29374 11954
rect 29426 11902 29428 11954
rect 28924 7298 28980 7308
rect 29036 11284 29092 11294
rect 29372 11284 29428 11902
rect 29484 11732 29540 12124
rect 29484 11666 29540 11676
rect 29036 11282 29428 11284
rect 29036 11230 29038 11282
rect 29090 11230 29428 11282
rect 29036 11228 29428 11230
rect 29484 11508 29540 11518
rect 29036 7140 29092 11228
rect 29260 9940 29316 9950
rect 29148 9604 29204 9614
rect 29148 7588 29204 9548
rect 29148 7522 29204 7532
rect 29260 7476 29316 9884
rect 29372 9604 29428 9614
rect 29372 8370 29428 9548
rect 29372 8318 29374 8370
rect 29426 8318 29428 8370
rect 29372 8306 29428 8318
rect 29260 7410 29316 7420
rect 28924 7084 29092 7140
rect 29148 7252 29204 7262
rect 29372 7252 29428 7262
rect 29148 7250 29428 7252
rect 29148 7198 29150 7250
rect 29202 7198 29374 7250
rect 29426 7198 29428 7250
rect 29148 7196 29428 7198
rect 28924 5572 28980 7084
rect 29148 6804 29204 7196
rect 29372 7186 29428 7196
rect 29484 7140 29540 11452
rect 29596 8708 29652 14112
rect 29820 13860 29876 14112
rect 29820 13794 29876 13804
rect 30044 13748 30100 14112
rect 30268 13860 30324 14112
rect 30268 13794 30324 13804
rect 30044 13682 30100 13692
rect 29820 13636 29876 13646
rect 29820 11284 29876 13580
rect 30044 12628 30100 12638
rect 29932 12066 29988 12078
rect 29932 12014 29934 12066
rect 29986 12014 29988 12066
rect 29932 11508 29988 12014
rect 29932 11442 29988 11452
rect 29820 11218 29876 11228
rect 29596 8642 29652 8652
rect 29708 11172 29764 11182
rect 29708 8484 29764 11116
rect 30044 9828 30100 12572
rect 30156 12292 30212 12302
rect 30156 11620 30212 12236
rect 30492 12180 30548 14112
rect 30716 12898 30772 14112
rect 30940 13076 30996 14112
rect 30940 13010 30996 13020
rect 30716 12842 30996 12898
rect 30828 12740 30884 12750
rect 30492 12114 30548 12124
rect 30716 12628 30772 12638
rect 30380 11956 30436 11966
rect 30604 11956 30660 11966
rect 30380 11954 30660 11956
rect 30380 11902 30382 11954
rect 30434 11902 30606 11954
rect 30658 11902 30660 11954
rect 30380 11900 30660 11902
rect 30156 11554 30212 11564
rect 30268 11844 30324 11854
rect 30044 9762 30100 9772
rect 30156 11396 30212 11406
rect 30156 9492 30212 11340
rect 30156 9426 30212 9436
rect 29484 7074 29540 7084
rect 29596 8428 29764 8484
rect 29148 6738 29204 6748
rect 29596 6804 29652 8428
rect 29932 8258 29988 8270
rect 29932 8206 29934 8258
rect 29986 8206 29988 8258
rect 29932 8148 29988 8206
rect 30156 8148 30212 8158
rect 29932 8092 30156 8148
rect 30156 8054 30212 8092
rect 29596 6738 29652 6748
rect 29708 8036 29764 8046
rect 29372 6690 29428 6702
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 28924 5506 28980 5516
rect 29036 6580 29092 6590
rect 29372 6580 29428 6638
rect 29036 6578 29428 6580
rect 29036 6526 29038 6578
rect 29090 6526 29428 6578
rect 29036 6524 29428 6526
rect 29036 4340 29092 6524
rect 29708 5572 29764 7980
rect 30268 7924 30324 11788
rect 30380 9380 30436 11900
rect 30604 11890 30660 11900
rect 30380 9314 30436 9324
rect 30604 10052 30660 10062
rect 30044 7868 30324 7924
rect 30380 9044 30436 9054
rect 29932 7476 29988 7486
rect 29932 7382 29988 7420
rect 29708 5506 29764 5516
rect 29820 6916 29876 6926
rect 29820 5460 29876 6860
rect 29932 6692 29988 6702
rect 29932 6598 29988 6636
rect 29820 5394 29876 5404
rect 29036 4274 29092 4284
rect 29596 4900 29652 4910
rect 28812 4060 29092 4116
rect 29036 3780 29092 4060
rect 29260 3780 29316 3790
rect 29036 3778 29316 3780
rect 29036 3726 29038 3778
rect 29090 3726 29262 3778
rect 29314 3726 29316 3778
rect 29036 3724 29316 3726
rect 29036 3714 29092 3724
rect 29260 3714 29316 3724
rect 27356 2930 27412 2940
rect 27692 3332 28308 3388
rect 26460 2370 26516 2380
rect 26796 2380 26964 2436
rect 26348 1138 26404 1148
rect 26796 1092 26852 2380
rect 26796 1026 26852 1036
rect 27692 868 27748 3332
rect 29596 2884 29652 4844
rect 29820 3444 29876 3482
rect 29820 3378 29876 3388
rect 30044 3388 30100 7868
rect 30156 6244 30212 6254
rect 30156 4452 30212 6188
rect 30380 6020 30436 8988
rect 30380 5954 30436 5964
rect 30604 6020 30660 9996
rect 30716 9940 30772 12572
rect 30716 9874 30772 9884
rect 30828 7028 30884 12684
rect 30940 11284 30996 12842
rect 31164 12852 31220 14112
rect 31164 12786 31220 12796
rect 31388 12180 31444 14112
rect 31612 13636 31668 14112
rect 31836 13636 31892 14112
rect 31612 13570 31668 13580
rect 31724 13580 31892 13636
rect 31388 12114 31444 12124
rect 31612 13188 31668 13198
rect 30940 11218 30996 11228
rect 31164 12066 31220 12078
rect 31164 12014 31166 12066
rect 31218 12014 31220 12066
rect 30828 6962 30884 6972
rect 30940 10388 30996 10398
rect 30940 6132 30996 10332
rect 31164 10388 31220 12014
rect 31164 10322 31220 10332
rect 31052 10052 31108 10062
rect 31052 8932 31108 9996
rect 31052 8866 31108 8876
rect 31500 9828 31556 9838
rect 30940 6066 30996 6076
rect 31164 8148 31220 8158
rect 30604 5954 30660 5964
rect 30156 4386 30212 4396
rect 30268 5684 30324 5694
rect 30044 3332 30212 3388
rect 30156 3220 30212 3332
rect 30268 3332 30324 5628
rect 30268 3266 30324 3276
rect 30380 3444 30436 3454
rect 30156 3154 30212 3164
rect 29596 2818 29652 2828
rect 28812 2660 28868 2670
rect 25116 812 26964 868
rect 24892 700 25396 756
rect 25228 532 25284 542
rect 24332 476 25228 532
rect 25228 466 25284 476
rect 25340 420 25396 700
rect 26796 420 26852 430
rect 25340 364 26796 420
rect 26796 354 26852 364
rect 23996 130 24052 140
rect 26236 196 26292 206
rect 26236 112 26292 140
rect 9660 84 9716 94
rect 9436 28 9660 84
rect 9660 18 9716 28
rect 11424 0 11536 112
rect 13888 0 14000 112
rect 16352 0 16464 112
rect 18816 0 18928 112
rect 21280 0 21392 112
rect 23744 0 23856 112
rect 26208 0 26320 112
rect 26908 84 26964 812
rect 27692 802 27748 812
rect 28700 1876 28756 1886
rect 28700 112 28756 1820
rect 28812 1428 28868 2604
rect 28812 1362 28868 1372
rect 30044 2548 30100 2558
rect 30044 756 30100 2492
rect 30380 2436 30436 3388
rect 30380 2370 30436 2380
rect 30604 2996 30660 3006
rect 30604 2436 30660 2940
rect 30604 2370 30660 2380
rect 30828 1988 30884 1998
rect 30156 1764 30212 1774
rect 30156 1092 30212 1708
rect 30828 1540 30884 1932
rect 30828 1474 30884 1484
rect 30156 1026 30212 1036
rect 30044 690 30100 700
rect 31164 112 31220 8092
rect 31500 4228 31556 9772
rect 31612 8932 31668 13132
rect 31724 12404 31780 13580
rect 31724 12338 31780 12348
rect 31836 13412 31892 13422
rect 31836 10612 31892 13356
rect 31836 10546 31892 10556
rect 31612 8866 31668 8876
rect 31836 8148 31892 8158
rect 31724 6468 31780 6478
rect 31724 4452 31780 6412
rect 31724 4386 31780 4396
rect 31500 4162 31556 4172
rect 31836 4004 31892 8092
rect 32060 7476 32116 14112
rect 32284 14084 32340 14112
rect 32284 14018 32340 14028
rect 32284 13076 32340 13086
rect 32284 7700 32340 13020
rect 32396 12964 32452 12974
rect 32396 11620 32452 12908
rect 32508 11844 32564 14112
rect 32508 11778 32564 11788
rect 32396 11554 32452 11564
rect 32508 10500 32564 10510
rect 32508 9492 32564 10444
rect 32732 9716 32788 14112
rect 32956 13972 33012 14112
rect 32956 13906 33012 13916
rect 33068 13188 33124 13198
rect 33068 10052 33124 13132
rect 33068 9986 33124 9996
rect 32732 9650 32788 9660
rect 32508 9426 32564 9436
rect 32508 8820 32564 8830
rect 32396 8258 32452 8270
rect 32396 8206 32398 8258
rect 32450 8206 32452 8258
rect 32396 8148 32452 8206
rect 32396 8082 32452 8092
rect 32284 7634 32340 7644
rect 32060 7420 32340 7476
rect 31948 6916 32004 6926
rect 31948 6468 32004 6860
rect 31948 6402 32004 6412
rect 32284 4452 32340 7420
rect 32508 5124 32564 8764
rect 33180 8596 33236 14112
rect 33180 8530 33236 8540
rect 33292 10836 33348 10846
rect 32732 8484 32788 8494
rect 32732 6356 32788 8428
rect 32956 8146 33012 8158
rect 32956 8094 32958 8146
rect 33010 8094 33012 8146
rect 32956 8036 33012 8094
rect 32956 7970 33012 7980
rect 32732 6290 32788 6300
rect 32956 7588 33012 7598
rect 32508 5058 32564 5068
rect 32844 5460 32900 5470
rect 32844 4564 32900 5404
rect 32844 4498 32900 4508
rect 32284 4450 32676 4452
rect 32284 4398 32286 4450
rect 32338 4398 32676 4450
rect 32284 4396 32676 4398
rect 32284 4386 32340 4396
rect 32620 4338 32676 4396
rect 32620 4286 32622 4338
rect 32674 4286 32676 4338
rect 32620 4274 32676 4286
rect 32956 4228 33012 7532
rect 33180 5572 33236 5582
rect 33068 4452 33124 4462
rect 33068 4358 33124 4396
rect 32956 4172 33124 4228
rect 31836 3938 31892 3948
rect 32620 3556 32676 3566
rect 31948 3108 32004 3118
rect 31948 2660 32004 3052
rect 31948 2594 32004 2604
rect 32620 2212 32676 3500
rect 32956 3554 33012 3566
rect 32956 3502 32958 3554
rect 33010 3502 33012 3554
rect 32732 3444 32788 3482
rect 32956 3444 33012 3502
rect 32788 3388 33012 3444
rect 33068 3388 33124 4172
rect 33180 3556 33236 5516
rect 33292 4004 33348 10780
rect 33404 10612 33460 14112
rect 33628 12740 33684 14112
rect 33628 12674 33684 12684
rect 33628 12516 33684 12526
rect 33628 10836 33684 12460
rect 33628 10770 33684 10780
rect 33740 12068 33796 12078
rect 33852 12068 33908 14112
rect 34076 13076 34132 14112
rect 34300 13188 34356 14112
rect 34300 13122 34356 13132
rect 34076 13010 34132 13020
rect 33852 12012 34020 12068
rect 33404 10556 33572 10612
rect 33404 10388 33460 10398
rect 33404 5684 33460 10332
rect 33516 9044 33572 10556
rect 33516 8978 33572 8988
rect 33628 10052 33684 10062
rect 33516 8820 33572 8830
rect 33516 5796 33572 8764
rect 33628 6804 33684 9996
rect 33740 9716 33796 12012
rect 33740 9650 33796 9660
rect 33852 11844 33908 11854
rect 33852 9156 33908 11788
rect 33852 9090 33908 9100
rect 33740 9044 33796 9054
rect 33740 7812 33796 8988
rect 33964 8708 34020 12012
rect 34300 11732 34356 11742
rect 34188 10164 34244 10174
rect 34188 10050 34244 10108
rect 34188 9998 34190 10050
rect 34242 9998 34244 10050
rect 34188 9986 34244 9998
rect 33964 8642 34020 8652
rect 34076 9380 34132 9390
rect 34076 8148 34132 9324
rect 34076 8082 34132 8092
rect 33740 7746 33796 7756
rect 33964 7924 34020 7934
rect 33852 7700 33908 7710
rect 33628 6738 33684 6748
rect 33740 6916 33796 6926
rect 33740 6132 33796 6860
rect 33740 6066 33796 6076
rect 33516 5730 33572 5740
rect 33852 5796 33908 7644
rect 33852 5730 33908 5740
rect 33404 5618 33460 5628
rect 33292 3938 33348 3948
rect 33404 5236 33460 5246
rect 33180 3490 33236 3500
rect 32732 3378 32788 3388
rect 33068 3332 33236 3388
rect 33180 2996 33236 3332
rect 33404 3108 33460 5180
rect 33628 5124 33684 5134
rect 33516 4564 33572 4574
rect 33516 3666 33572 4508
rect 33516 3614 33518 3666
rect 33570 3614 33572 3666
rect 33516 3602 33572 3614
rect 33628 3388 33684 5068
rect 33964 4676 34020 7868
rect 34300 7812 34356 11676
rect 34524 9940 34580 14112
rect 34748 12628 34804 14112
rect 34748 12562 34804 12572
rect 34524 9874 34580 9884
rect 34636 10164 34692 10174
rect 34636 9826 34692 10108
rect 34636 9774 34638 9826
rect 34690 9774 34692 9826
rect 34636 9762 34692 9774
rect 34972 8596 35028 14112
rect 35196 13188 35252 14112
rect 35196 13122 35252 13132
rect 35308 13860 35364 13870
rect 35308 11060 35364 13804
rect 35420 13412 35476 14112
rect 35420 13346 35476 13356
rect 35532 13300 35588 13310
rect 35308 10994 35364 11004
rect 35420 12962 35476 12974
rect 35420 12910 35422 12962
rect 35474 12910 35476 12962
rect 35084 9716 35140 9726
rect 35084 9714 35364 9716
rect 35084 9662 35086 9714
rect 35138 9662 35364 9714
rect 35084 9660 35364 9662
rect 35084 9650 35140 9660
rect 34972 8530 35028 8540
rect 35308 8260 35364 9660
rect 35308 8194 35364 8204
rect 34300 7746 34356 7756
rect 35308 7252 35364 7262
rect 35308 5908 35364 7196
rect 35308 5842 35364 5852
rect 35308 5572 35364 5582
rect 35308 4788 35364 5516
rect 35308 4722 35364 4732
rect 33964 4610 34020 4620
rect 35308 4228 35364 4238
rect 35308 3388 35364 4172
rect 33404 3042 33460 3052
rect 33516 3332 33684 3388
rect 35196 3332 35364 3388
rect 35420 3332 35476 12910
rect 35532 12898 35588 13244
rect 35644 13188 35700 14112
rect 35756 13188 35812 13198
rect 35644 13186 35812 13188
rect 35644 13134 35758 13186
rect 35810 13134 35812 13186
rect 35644 13132 35812 13134
rect 35756 13122 35812 13132
rect 35532 12842 35812 12898
rect 35532 12740 35588 12750
rect 35532 10388 35588 12684
rect 35532 10322 35588 10332
rect 35644 11284 35700 11294
rect 35532 10052 35588 10062
rect 35532 8484 35588 9996
rect 35532 8418 35588 8428
rect 35532 6692 35588 6702
rect 35532 4340 35588 6636
rect 35644 6468 35700 11228
rect 35756 8596 35812 12842
rect 35868 12852 35924 14112
rect 36092 13076 36148 14112
rect 36316 13076 36372 14112
rect 36540 13300 36596 14112
rect 36764 13748 36820 14112
rect 36764 13682 36820 13692
rect 36540 13234 36596 13244
rect 36876 13412 36932 13422
rect 36540 13076 36596 13086
rect 36316 13020 36484 13076
rect 36092 13010 36148 13020
rect 36316 12852 36372 12862
rect 35868 12850 36372 12852
rect 35868 12798 36318 12850
rect 36370 12798 36372 12850
rect 35868 12796 36372 12798
rect 36316 12786 36372 12796
rect 36316 12180 36372 12190
rect 36204 9826 36260 9838
rect 36204 9774 36206 9826
rect 36258 9774 36260 9826
rect 35756 8530 35812 8540
rect 35868 9716 35924 9726
rect 36204 9716 36260 9774
rect 35868 9714 36260 9716
rect 35868 9662 35870 9714
rect 35922 9662 36260 9714
rect 35868 9660 36260 9662
rect 35644 6402 35700 6412
rect 35868 5012 35924 9660
rect 36316 9156 36372 12124
rect 36428 11284 36484 13020
rect 36540 12402 36596 13020
rect 36540 12350 36542 12402
rect 36594 12350 36596 12402
rect 36540 12338 36596 12350
rect 36764 11284 36820 11294
rect 36428 11282 36820 11284
rect 36428 11230 36766 11282
rect 36818 11230 36820 11282
rect 36428 11228 36820 11230
rect 36764 11218 36820 11228
rect 36764 9714 36820 9726
rect 36764 9662 36766 9714
rect 36818 9662 36820 9714
rect 36316 9090 36372 9100
rect 36652 9380 36708 9390
rect 36652 8372 36708 9324
rect 36764 8484 36820 9662
rect 36764 8418 36820 8428
rect 36652 8306 36708 8316
rect 35868 4946 35924 4956
rect 35980 6356 36036 6366
rect 35532 4274 35588 4284
rect 35756 4788 35812 4798
rect 33180 2930 33236 2940
rect 32844 2212 32900 2222
rect 32620 2210 32900 2212
rect 32620 2158 32622 2210
rect 32674 2158 32846 2210
rect 32898 2158 32900 2210
rect 32620 2156 32900 2158
rect 32620 2146 32676 2156
rect 32844 2146 32900 2156
rect 33404 1988 33460 1998
rect 33404 1894 33460 1932
rect 32732 1764 32788 1774
rect 32732 196 32788 1708
rect 33516 868 33572 3332
rect 33516 802 33572 812
rect 33628 2212 33684 2222
rect 32732 130 32788 140
rect 33628 112 33684 2156
rect 35196 1652 35252 3332
rect 35420 3266 35476 3276
rect 35756 3220 35812 4732
rect 35980 4676 36036 6300
rect 35980 4610 36036 4620
rect 36092 6020 36148 6030
rect 35756 3154 35812 3164
rect 35196 1586 35252 1596
rect 35308 3108 35364 3118
rect 35308 1316 35364 3052
rect 35308 1250 35364 1260
rect 36092 112 36148 5964
rect 36652 3668 36708 3678
rect 36652 1204 36708 3612
rect 36764 2884 36820 2894
rect 36876 2884 36932 13356
rect 36988 10836 37044 14112
rect 37100 12852 37156 12862
rect 37100 11620 37156 12796
rect 37212 12740 37268 14112
rect 37324 12962 37380 12974
rect 37324 12910 37326 12962
rect 37378 12910 37380 12962
rect 37324 12852 37380 12910
rect 37324 12786 37380 12796
rect 37212 12674 37268 12684
rect 37436 12516 37492 14112
rect 37660 13412 37716 14112
rect 37660 13346 37716 13356
rect 37772 13188 37828 13198
rect 37772 13094 37828 13132
rect 37436 12450 37492 12460
rect 37884 12404 37940 14112
rect 38108 13524 38164 14112
rect 38108 13468 38276 13524
rect 38108 13300 38164 13310
rect 37996 13188 38052 13198
rect 37996 13094 38052 13132
rect 37884 12338 37940 12348
rect 38108 12402 38164 13244
rect 38108 12350 38110 12402
rect 38162 12350 38164 12402
rect 38108 12338 38164 12350
rect 37100 11554 37156 11564
rect 37548 12066 37604 12078
rect 37548 12014 37550 12066
rect 37602 12014 37604 12066
rect 37548 11284 37604 12014
rect 38220 11732 38276 13468
rect 38332 13076 38388 14112
rect 38556 13412 38612 14112
rect 38332 13010 38388 13020
rect 38444 13356 38612 13412
rect 38668 13524 38724 13534
rect 38444 12628 38500 13356
rect 38668 13300 38724 13468
rect 38668 13234 38724 13244
rect 38444 12562 38500 12572
rect 38556 12850 38612 12862
rect 38556 12798 38558 12850
rect 38610 12798 38612 12850
rect 38220 11666 38276 11676
rect 37772 11396 37828 11406
rect 38108 11396 38164 11406
rect 37772 11394 37940 11396
rect 37772 11342 37774 11394
rect 37826 11342 37940 11394
rect 37772 11340 37940 11342
rect 37772 11330 37828 11340
rect 37548 11218 37604 11228
rect 37772 10836 37828 10846
rect 36988 10834 37828 10836
rect 36988 10782 37774 10834
rect 37826 10782 37828 10834
rect 36988 10780 37828 10782
rect 37772 10770 37828 10780
rect 37212 10498 37268 10510
rect 37212 10446 37214 10498
rect 37266 10446 37268 10498
rect 37212 10164 37268 10446
rect 37772 10388 37828 10398
rect 37212 10098 37268 10108
rect 37548 10276 37604 10286
rect 36988 9268 37044 9278
rect 36988 5012 37044 9212
rect 36988 4946 37044 4956
rect 37100 7812 37156 7822
rect 37100 3444 37156 7756
rect 37548 6020 37604 10220
rect 37772 9716 37828 10332
rect 37884 9940 37940 11340
rect 37884 9874 37940 9884
rect 37996 11394 38164 11396
rect 37996 11342 38110 11394
rect 38162 11342 38164 11394
rect 37996 11340 38164 11342
rect 37772 9660 37940 9716
rect 37548 6018 37828 6020
rect 37548 5966 37550 6018
rect 37602 5966 37828 6018
rect 37548 5964 37828 5966
rect 37548 5954 37604 5964
rect 37772 5906 37828 5964
rect 37772 5854 37774 5906
rect 37826 5854 37828 5906
rect 37772 5842 37828 5854
rect 37660 5796 37716 5806
rect 37100 3378 37156 3388
rect 37548 4676 37604 4686
rect 36764 2882 37156 2884
rect 36764 2830 36766 2882
rect 36818 2830 37156 2882
rect 36764 2828 37156 2830
rect 36764 2818 36820 2828
rect 37100 2770 37156 2828
rect 37100 2718 37102 2770
rect 37154 2718 37156 2770
rect 37100 2706 37156 2718
rect 36652 1138 36708 1148
rect 36988 2100 37044 2110
rect 36988 532 37044 2044
rect 36988 466 37044 476
rect 37548 308 37604 4620
rect 37660 4452 37716 5740
rect 37884 4676 37940 9660
rect 37996 5572 38052 11340
rect 38108 11330 38164 11340
rect 38332 9828 38388 9838
rect 38332 9734 38388 9772
rect 38556 9380 38612 12798
rect 38668 12740 38724 12750
rect 38668 11618 38724 12684
rect 38780 12180 38836 14112
rect 39004 13524 39060 14112
rect 39004 13458 39060 13468
rect 39116 12964 39172 12974
rect 38780 12114 38836 12124
rect 39004 12962 39172 12964
rect 39004 12910 39118 12962
rect 39170 12910 39172 12962
rect 39004 12908 39172 12910
rect 38668 11566 38670 11618
rect 38722 11566 38724 11618
rect 38668 11554 38724 11566
rect 38892 11732 38948 11742
rect 38780 11172 38836 11182
rect 38780 10610 38836 11116
rect 38780 10558 38782 10610
rect 38834 10558 38836 10610
rect 38780 10546 38836 10558
rect 38668 10164 38724 10174
rect 38668 9604 38724 10108
rect 38780 10052 38836 10062
rect 38780 9716 38836 9996
rect 38892 10050 38948 11676
rect 38892 9998 38894 10050
rect 38946 9998 38948 10050
rect 38892 9986 38948 9998
rect 38780 9650 38836 9660
rect 38668 9538 38724 9548
rect 38332 9324 38612 9380
rect 38220 9156 38276 9166
rect 38220 9062 38276 9100
rect 38332 7028 38388 9324
rect 38556 9156 38612 9166
rect 38556 9042 38612 9100
rect 38556 8990 38558 9042
rect 38610 8990 38612 9042
rect 38556 8978 38612 8990
rect 38668 9044 38724 9054
rect 38668 8596 38724 8988
rect 38668 8530 38724 8540
rect 39004 8428 39060 12908
rect 39116 12898 39172 12908
rect 39228 12740 39284 14112
rect 39228 12674 39284 12684
rect 39452 12516 39508 14112
rect 39452 12460 39620 12516
rect 39340 12404 39396 12414
rect 39116 12066 39172 12078
rect 39116 12014 39118 12066
rect 39170 12014 39172 12066
rect 39116 10276 39172 12014
rect 39340 10834 39396 12348
rect 39452 12292 39508 12302
rect 39452 12178 39508 12236
rect 39452 12126 39454 12178
rect 39506 12126 39508 12178
rect 39452 12114 39508 12126
rect 39340 10782 39342 10834
rect 39394 10782 39396 10834
rect 39340 10770 39396 10782
rect 39116 10210 39172 10220
rect 39564 10052 39620 12460
rect 39676 11508 39732 14112
rect 39676 11452 39844 11508
rect 39564 9986 39620 9996
rect 39676 10836 39732 10846
rect 38780 8372 39060 8428
rect 39116 8930 39172 8942
rect 39116 8878 39118 8930
rect 39170 8878 39172 8930
rect 38780 7476 38836 8372
rect 38780 7410 38836 7420
rect 38332 6962 38388 6972
rect 38444 6916 38500 6926
rect 38500 6860 38612 6916
rect 38444 6850 38500 6860
rect 37996 5506 38052 5516
rect 38108 6692 38164 6702
rect 37884 4610 37940 4620
rect 37660 4396 38052 4452
rect 37884 3892 37940 3902
rect 37660 2658 37716 2670
rect 37660 2606 37662 2658
rect 37714 2606 37716 2658
rect 37660 2548 37716 2606
rect 37660 2482 37716 2492
rect 37884 1428 37940 3836
rect 37884 1362 37940 1372
rect 37548 242 37604 252
rect 37996 196 38052 4396
rect 38108 1316 38164 6636
rect 38556 6590 38612 6860
rect 38444 6580 38500 6590
rect 38556 6580 38668 6590
rect 38556 6524 38612 6580
rect 38444 6418 38500 6524
rect 38612 6514 38668 6524
rect 39116 6580 39172 8878
rect 39116 6514 39172 6524
rect 39564 8820 39620 8830
rect 38444 6362 38724 6418
rect 38220 6018 38276 6030
rect 38220 5966 38222 6018
rect 38274 5966 38276 6018
rect 38220 2772 38276 5966
rect 38332 5348 38388 5358
rect 38444 5348 38500 6362
rect 38668 5906 38724 6362
rect 38668 5854 38670 5906
rect 38722 5854 38724 5906
rect 38668 5842 38724 5854
rect 38332 5346 38500 5348
rect 38332 5294 38334 5346
rect 38386 5294 38500 5346
rect 38332 5292 38500 5294
rect 39228 5794 39284 5806
rect 39228 5742 39230 5794
rect 39282 5742 39284 5794
rect 38332 5282 38388 5292
rect 38668 5236 38724 5246
rect 38668 5142 38724 5180
rect 38892 5236 38948 5246
rect 38892 5142 38948 5180
rect 38780 5124 38836 5134
rect 38780 3332 38836 5068
rect 38780 3266 38836 3276
rect 38556 2996 38612 3006
rect 38556 2882 38612 2940
rect 38556 2830 38558 2882
rect 38610 2830 38612 2882
rect 38556 2818 38612 2830
rect 38892 2996 38948 3006
rect 38220 2706 38276 2716
rect 38892 2770 38948 2940
rect 38892 2718 38894 2770
rect 38946 2718 38948 2770
rect 38892 2706 38948 2718
rect 38668 2548 38724 2558
rect 38668 2324 38724 2492
rect 38668 2258 38724 2268
rect 39228 2324 39284 5742
rect 39452 5236 39508 5246
rect 39452 5142 39508 5180
rect 39452 2658 39508 2670
rect 39452 2606 39454 2658
rect 39506 2606 39508 2658
rect 39452 2436 39508 2606
rect 39564 2548 39620 8764
rect 39676 4340 39732 10780
rect 39788 9604 39844 11452
rect 39900 10836 39956 14112
rect 40012 13748 40068 13758
rect 40012 12850 40068 13692
rect 40124 13188 40180 14112
rect 40684 13636 40740 13646
rect 40124 13122 40180 13132
rect 40236 13300 40292 13310
rect 40236 12964 40292 13244
rect 40684 13074 40740 13580
rect 41244 13412 41300 13422
rect 41244 13186 41300 13356
rect 41244 13134 41246 13186
rect 41298 13134 41300 13186
rect 41244 13122 41300 13134
rect 40684 13022 40686 13074
rect 40738 13022 40740 13074
rect 40684 13010 40740 13022
rect 41580 13076 41636 13086
rect 40012 12798 40014 12850
rect 40066 12798 40068 12850
rect 40012 12786 40068 12798
rect 40124 12908 40292 12964
rect 40012 12516 40068 12526
rect 40012 12402 40068 12460
rect 40012 12350 40014 12402
rect 40066 12350 40068 12402
rect 40012 12338 40068 12350
rect 39900 10770 39956 10780
rect 40012 11620 40068 11630
rect 40012 10612 40068 11564
rect 39788 9538 39844 9548
rect 39900 10556 40068 10612
rect 39900 9380 39956 10556
rect 39788 9324 39956 9380
rect 40012 9492 40068 9502
rect 39788 5124 39844 9324
rect 39900 8930 39956 8942
rect 39900 8878 39902 8930
rect 39954 8878 39956 8930
rect 39900 6804 39956 8878
rect 39900 6738 39956 6748
rect 39788 5058 39844 5068
rect 40012 5012 40068 9436
rect 40124 6132 40180 12908
rect 40796 12628 40852 12638
rect 40796 11618 40852 12572
rect 41580 12402 41636 13020
rect 41580 12350 41582 12402
rect 41634 12350 41636 12402
rect 41580 12338 41636 12350
rect 40796 11566 40798 11618
rect 40850 11566 40852 11618
rect 40796 11554 40852 11566
rect 40908 12180 40964 12190
rect 40460 11394 40516 11406
rect 40460 11342 40462 11394
rect 40514 11342 40516 11394
rect 40348 9828 40404 9838
rect 40348 9734 40404 9772
rect 40460 9268 40516 11342
rect 40908 10834 40964 12124
rect 41132 12180 41188 12190
rect 40908 10782 40910 10834
rect 40962 10782 40964 10834
rect 40908 10770 40964 10782
rect 41020 11844 41076 11854
rect 40572 10612 40628 10622
rect 40572 10610 40740 10612
rect 40572 10558 40574 10610
rect 40626 10558 40740 10610
rect 40572 10556 40740 10558
rect 40572 10546 40628 10556
rect 40684 9380 40740 10556
rect 40908 10500 40964 10510
rect 40796 10052 40852 10062
rect 40796 9958 40852 9996
rect 40908 9828 40964 10444
rect 41020 10052 41076 11788
rect 41020 9986 41076 9996
rect 40908 9772 41076 9828
rect 40908 9604 40964 9614
rect 40684 9324 40852 9380
rect 40460 9212 40740 9268
rect 40460 8932 40516 8942
rect 40236 8596 40292 8606
rect 40236 7476 40292 8540
rect 40460 8148 40516 8876
rect 40460 8082 40516 8092
rect 40236 7410 40292 7420
rect 40124 6066 40180 6076
rect 40572 6580 40628 6590
rect 40012 4956 40516 5012
rect 39676 4284 39844 4340
rect 39564 2482 39620 2492
rect 39452 2370 39508 2380
rect 39228 2258 39284 2268
rect 38892 2212 38948 2222
rect 38892 2118 38948 2156
rect 39116 2212 39172 2222
rect 39116 2118 39172 2156
rect 39676 2100 39732 2110
rect 39676 2006 39732 2044
rect 38108 1250 38164 1260
rect 37996 130 38052 140
rect 38556 196 38612 206
rect 38556 112 38612 140
rect 39788 196 39844 4284
rect 40348 3668 40404 3678
rect 40348 1764 40404 3612
rect 40460 2884 40516 4956
rect 40572 4900 40628 6524
rect 40572 4834 40628 4844
rect 40684 4788 40740 9212
rect 40684 4722 40740 4732
rect 40460 2818 40516 2828
rect 40796 2660 40852 9324
rect 40908 9266 40964 9548
rect 40908 9214 40910 9266
rect 40962 9214 40964 9266
rect 40908 9202 40964 9214
rect 41020 8428 41076 9772
rect 40908 8372 41076 8428
rect 40908 7588 40964 8372
rect 40908 7522 40964 7532
rect 41132 6244 41188 12124
rect 41244 12178 41300 12190
rect 41244 12126 41246 12178
rect 41298 12126 41300 12178
rect 41244 10164 41300 12126
rect 41468 10388 41524 10398
rect 41244 10098 41300 10108
rect 41356 10276 41412 10286
rect 41356 8372 41412 10220
rect 41356 8306 41412 8316
rect 41132 6178 41188 6188
rect 40796 2594 40852 2604
rect 41020 5460 41076 5470
rect 40236 1708 40404 1764
rect 40236 1540 40292 1708
rect 40236 1474 40292 1484
rect 39788 130 39844 140
rect 41020 112 41076 5404
rect 41468 2100 41524 10332
rect 41692 10052 41748 14140
rect 51100 13972 51156 13982
rect 42588 13860 42644 13870
rect 42252 12964 42308 12974
rect 42588 12964 42644 13804
rect 43708 13524 43764 13534
rect 43708 13074 43764 13468
rect 50876 13524 50932 13534
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 45052 13188 45108 13198
rect 45052 13094 45108 13132
rect 43708 13022 43710 13074
rect 43762 13022 43764 13074
rect 43708 13010 43764 13022
rect 48076 13076 48132 13086
rect 42252 12962 42644 12964
rect 42252 12910 42254 12962
rect 42306 12910 42644 12962
rect 42252 12908 42644 12910
rect 42252 12898 42308 12908
rect 42364 12740 42420 12750
rect 42364 11618 42420 12684
rect 42588 12178 42644 12908
rect 42588 12126 42590 12178
rect 42642 12126 42644 12178
rect 42588 12114 42644 12126
rect 42924 12962 42980 12974
rect 44492 12964 44548 12974
rect 42924 12910 42926 12962
rect 42978 12910 42980 12962
rect 42924 11956 42980 12910
rect 44268 12962 44548 12964
rect 44268 12910 44494 12962
rect 44546 12910 44548 12962
rect 44268 12908 44548 12910
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 42924 11890 42980 11900
rect 43036 12068 43092 12078
rect 42364 11566 42366 11618
rect 42418 11566 42420 11618
rect 42364 11554 42420 11566
rect 41804 11396 41860 11406
rect 41804 11302 41860 11340
rect 42476 10836 42532 10846
rect 42476 10742 42532 10780
rect 42028 10612 42084 10622
rect 42028 10518 42084 10556
rect 41804 10052 41860 10062
rect 41692 10050 41860 10052
rect 41692 9998 41806 10050
rect 41858 9998 41860 10050
rect 41692 9996 41860 9998
rect 41580 9156 41636 9166
rect 41692 9156 41748 9996
rect 41804 9986 41860 9996
rect 41916 9940 41972 9950
rect 41580 9154 41748 9156
rect 41580 9102 41582 9154
rect 41634 9102 41748 9154
rect 41580 9100 41748 9102
rect 41804 9604 41860 9614
rect 41580 9090 41636 9100
rect 41804 7924 41860 9548
rect 41804 7858 41860 7868
rect 41916 4900 41972 9884
rect 42140 9940 42196 9950
rect 42140 9380 42196 9884
rect 42252 9716 42308 9726
rect 42252 9622 42308 9660
rect 42140 9314 42196 9324
rect 42364 9156 42420 9166
rect 42140 8708 42196 8718
rect 42140 6804 42196 8652
rect 42140 6738 42196 6748
rect 41916 4834 41972 4844
rect 41916 4676 41972 4686
rect 41916 4452 41972 4620
rect 41916 4450 42308 4452
rect 41916 4398 41918 4450
rect 41970 4398 42308 4450
rect 41916 4396 42308 4398
rect 41916 4386 41972 4396
rect 42252 4338 42308 4396
rect 42252 4286 42254 4338
rect 42306 4286 42308 4338
rect 42252 4274 42308 4286
rect 42364 2996 42420 9100
rect 42700 5012 42756 5022
rect 42700 4450 42756 4956
rect 42700 4398 42702 4450
rect 42754 4398 42756 4450
rect 42700 4386 42756 4398
rect 43036 3108 43092 12012
rect 43148 12066 43204 12078
rect 43148 12014 43150 12066
rect 43202 12014 43204 12066
rect 43148 6580 43204 12014
rect 43148 6514 43204 6524
rect 43260 11732 43316 11742
rect 43036 3042 43092 3052
rect 42364 2930 42420 2940
rect 41468 2034 41524 2044
rect 43260 868 43316 11676
rect 44268 11732 44324 12908
rect 44492 12898 44548 12908
rect 45164 12964 45220 12974
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44268 11666 44324 11676
rect 44940 11508 44996 11518
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 43932 9826 43988 9838
rect 44828 9828 44884 9838
rect 43932 9774 43934 9826
rect 43986 9774 43988 9826
rect 43596 9714 43652 9726
rect 43596 9662 43598 9714
rect 43650 9662 43652 9714
rect 43596 9604 43652 9662
rect 43932 9716 43988 9774
rect 44604 9826 44884 9828
rect 44604 9774 44830 9826
rect 44882 9774 44884 9826
rect 44604 9772 44884 9774
rect 43932 9650 43988 9660
rect 44492 9716 44548 9726
rect 44492 9622 44548 9660
rect 43596 9538 43652 9548
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 43596 9268 43652 9278
rect 43260 802 43316 812
rect 43484 6916 43540 6926
rect 43484 112 43540 6860
rect 43596 4450 43652 9212
rect 44492 9156 44548 9166
rect 44604 9156 44660 9772
rect 44828 9762 44884 9772
rect 44940 9828 44996 11452
rect 44940 9762 44996 9772
rect 44492 9154 44660 9156
rect 44492 9102 44494 9154
rect 44546 9102 44660 9154
rect 44492 9100 44660 9102
rect 45164 9156 45220 12908
rect 47180 12964 47236 12974
rect 47180 12870 47236 12908
rect 45276 12404 45332 12414
rect 45276 11620 45332 12348
rect 48076 12402 48132 13020
rect 48972 12964 49028 12974
rect 48972 12962 50148 12964
rect 48972 12910 48974 12962
rect 49026 12910 50148 12962
rect 48972 12908 50148 12910
rect 48972 12898 49028 12908
rect 48188 12738 48244 12750
rect 48188 12686 48190 12738
rect 48242 12686 48244 12738
rect 48188 12628 48244 12686
rect 48188 12562 48244 12572
rect 49756 12738 49812 12750
rect 49756 12686 49758 12738
rect 49810 12686 49812 12738
rect 48076 12350 48078 12402
rect 48130 12350 48132 12402
rect 48076 12338 48132 12350
rect 49644 12290 49700 12302
rect 49644 12238 49646 12290
rect 49698 12238 49700 12290
rect 48748 12180 48804 12190
rect 48748 12086 48804 12124
rect 47068 12066 47124 12078
rect 47068 12014 47070 12066
rect 47122 12014 47124 12066
rect 45276 11564 45780 11620
rect 45612 11396 45668 11406
rect 45276 11172 45332 11182
rect 45276 9714 45332 11116
rect 45276 9662 45278 9714
rect 45330 9662 45332 9714
rect 45276 9650 45332 9662
rect 44492 8932 44548 9100
rect 45164 9090 45220 9100
rect 44492 8866 44548 8876
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 45388 8484 45444 8494
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44268 6804 44324 6814
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 43596 4398 43598 4450
rect 43650 4398 43652 4450
rect 43596 4340 43652 4398
rect 43596 4274 43652 4284
rect 44156 4340 44212 4350
rect 44156 4246 44212 4284
rect 44268 3780 44324 6748
rect 44604 6690 44660 6702
rect 44604 6638 44606 6690
rect 44658 6638 44660 6690
rect 44380 6580 44436 6590
rect 44604 6580 44660 6638
rect 44380 6578 44660 6580
rect 44380 6526 44382 6578
rect 44434 6526 44660 6578
rect 44380 6524 44660 6526
rect 45052 6578 45108 6590
rect 45052 6526 45054 6578
rect 45106 6526 45108 6578
rect 44380 6468 44436 6524
rect 44380 6402 44436 6412
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 45052 5348 45108 6526
rect 45052 5282 45108 5292
rect 45388 4340 45444 8428
rect 45612 4564 45668 11340
rect 45724 6020 45780 11564
rect 47068 10052 47124 12014
rect 49644 11844 49700 12238
rect 49756 12180 49812 12686
rect 49756 12114 49812 12124
rect 49644 11778 49700 11788
rect 48860 11396 48916 11406
rect 48860 11302 48916 11340
rect 49868 11284 49924 11294
rect 49868 11190 49924 11228
rect 48748 10836 48804 10846
rect 47852 10724 47908 10734
rect 47516 10500 47572 10510
rect 47516 10406 47572 10444
rect 47740 10500 47796 10510
rect 47740 10406 47796 10444
rect 47068 9986 47124 9996
rect 47516 8820 47572 8830
rect 47740 8820 47796 8830
rect 47516 8818 47796 8820
rect 47516 8766 47518 8818
rect 47570 8766 47742 8818
rect 47794 8766 47796 8818
rect 47516 8764 47796 8766
rect 45724 5954 45780 5964
rect 46172 8036 46228 8046
rect 46172 4788 46228 7980
rect 46732 5124 46788 5134
rect 46172 4722 46228 4732
rect 46508 5012 46564 5022
rect 45612 4498 45668 4508
rect 45388 4274 45444 4284
rect 44716 4228 44772 4238
rect 44716 4134 44772 4172
rect 46172 4116 46228 4126
rect 46396 4116 46452 4126
rect 46172 4114 46452 4116
rect 46172 4062 46174 4114
rect 46226 4062 46398 4114
rect 46450 4062 46452 4114
rect 46172 4060 46452 4062
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 45276 3892 45332 3902
rect 44492 3780 44548 3790
rect 44716 3780 44772 3790
rect 44268 3778 44772 3780
rect 44268 3726 44494 3778
rect 44546 3726 44718 3778
rect 44770 3726 44772 3778
rect 44268 3724 44772 3726
rect 44492 3714 44548 3724
rect 44716 3714 44772 3724
rect 45276 3666 45332 3836
rect 45276 3614 45278 3666
rect 45330 3614 45332 3666
rect 45276 3602 45332 3614
rect 45612 3556 45668 3566
rect 45612 3462 45668 3500
rect 45836 3556 45892 3566
rect 45836 3462 45892 3500
rect 43596 3444 43652 3454
rect 43596 2212 43652 3388
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 45164 2884 45220 2894
rect 45220 2828 45444 2884
rect 45164 2790 45220 2828
rect 45388 2770 45444 2828
rect 45388 2718 45390 2770
rect 45442 2718 45444 2770
rect 45388 2706 45444 2718
rect 45948 2660 46004 2670
rect 45948 2566 46004 2604
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 43820 2212 43876 2222
rect 43596 2210 43876 2212
rect 43596 2158 43598 2210
rect 43650 2158 43822 2210
rect 43874 2158 43876 2210
rect 43596 2156 43876 2158
rect 43596 2118 43652 2156
rect 43820 2146 43876 2156
rect 44268 1876 44324 1886
rect 44268 1782 44324 1820
rect 46172 1764 46228 4060
rect 46396 4050 46452 4060
rect 46396 3668 46452 3678
rect 46508 3668 46564 4956
rect 46732 3780 46788 5068
rect 46844 4900 46900 4910
rect 46844 4450 46900 4844
rect 46844 4398 46846 4450
rect 46898 4398 46900 4450
rect 46844 4386 46900 4398
rect 47404 4116 47460 4126
rect 47404 4022 47460 4060
rect 46396 3666 46564 3668
rect 46396 3614 46398 3666
rect 46450 3614 46564 3666
rect 46396 3612 46564 3614
rect 46620 3778 46788 3780
rect 46620 3726 46734 3778
rect 46786 3726 46788 3778
rect 46620 3724 46788 3726
rect 46396 3602 46452 3612
rect 46508 2884 46564 2894
rect 46620 2884 46676 3724
rect 46732 3714 46788 3724
rect 46508 2882 46676 2884
rect 46508 2830 46510 2882
rect 46562 2830 46676 2882
rect 46508 2828 46676 2830
rect 47292 3442 47348 3454
rect 47292 3390 47294 3442
rect 47346 3390 47348 3442
rect 46508 2818 46564 2828
rect 47068 2772 47124 2782
rect 47068 2678 47124 2716
rect 46732 2100 46788 2110
rect 46732 2006 46788 2044
rect 46956 2100 47012 2110
rect 46956 2006 47012 2044
rect 46172 1698 46228 1708
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 45948 1428 46004 1438
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 45948 112 46004 1372
rect 47180 1204 47236 1214
rect 47180 1110 47236 1148
rect 47292 644 47348 3390
rect 47516 3332 47572 8764
rect 47740 8754 47796 8764
rect 47852 6244 47908 10668
rect 48748 10610 48804 10780
rect 48748 10558 48750 10610
rect 48802 10558 48804 10610
rect 48748 10546 48804 10558
rect 49644 10722 49700 10734
rect 49644 10670 49646 10722
rect 49698 10670 49700 10722
rect 48300 10498 48356 10510
rect 48300 10446 48302 10498
rect 48354 10446 48356 10498
rect 48300 10164 48356 10446
rect 49644 10388 49700 10670
rect 49644 10322 49700 10332
rect 48300 10098 48356 10108
rect 48860 9826 48916 9838
rect 48860 9774 48862 9826
rect 48914 9774 48916 9826
rect 48076 9044 48132 9054
rect 47852 6178 47908 6188
rect 47964 8708 48020 8718
rect 47740 6020 47796 6030
rect 47740 5926 47796 5964
rect 47964 5684 48020 8652
rect 48076 6692 48132 8988
rect 48748 9042 48804 9054
rect 48748 8990 48750 9042
rect 48802 8990 48804 9042
rect 48300 8932 48356 8942
rect 48300 8838 48356 8876
rect 48748 8820 48804 8990
rect 48748 8754 48804 8764
rect 48636 8258 48692 8270
rect 48636 8206 48638 8258
rect 48690 8206 48692 8258
rect 48188 8148 48244 8158
rect 48188 7252 48244 8092
rect 48300 8148 48356 8158
rect 48636 8148 48692 8206
rect 48300 8146 48692 8148
rect 48300 8094 48302 8146
rect 48354 8094 48692 8146
rect 48300 8092 48692 8094
rect 48300 7476 48356 8092
rect 48300 7410 48356 7420
rect 48748 7474 48804 7486
rect 48748 7422 48750 7474
rect 48802 7422 48804 7474
rect 48748 7364 48804 7422
rect 48748 7298 48804 7308
rect 48188 7186 48244 7196
rect 48860 6916 48916 9774
rect 48076 6626 48132 6636
rect 48748 6860 48916 6916
rect 48972 9828 49028 9838
rect 48972 6916 49028 9772
rect 48524 6580 48580 6590
rect 48076 6020 48132 6030
rect 48076 5906 48132 5964
rect 48524 6018 48580 6524
rect 48524 5966 48526 6018
rect 48578 5966 48580 6018
rect 48524 5954 48580 5966
rect 48076 5854 48078 5906
rect 48130 5854 48132 5906
rect 48076 5842 48132 5854
rect 47964 5618 48020 5628
rect 48748 5012 48804 6860
rect 48972 6850 49028 6860
rect 49084 9716 49140 9726
rect 48860 6690 48916 6702
rect 48860 6638 48862 6690
rect 48914 6638 48916 6690
rect 48860 5012 48916 6638
rect 48972 6132 49028 6142
rect 48972 6018 49028 6076
rect 48972 5966 48974 6018
rect 49026 5966 49028 6018
rect 48972 5954 49028 5966
rect 49084 5122 49140 9660
rect 49868 9716 49924 9726
rect 49868 9622 49924 9660
rect 49644 9268 49700 9278
rect 49644 9174 49700 9212
rect 49196 8372 49252 8382
rect 49196 8278 49252 8316
rect 49532 8258 49588 8270
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 8148 49588 8206
rect 49532 8082 49588 8092
rect 49980 8146 50036 8158
rect 49980 8094 49982 8146
rect 50034 8094 50036 8146
rect 49644 7586 49700 7598
rect 49644 7534 49646 7586
rect 49698 7534 49700 7586
rect 49644 6804 49700 7534
rect 49980 7588 50036 8094
rect 49980 7522 50036 7532
rect 49644 6738 49700 6748
rect 49756 6578 49812 6590
rect 49756 6526 49758 6578
rect 49810 6526 49812 6578
rect 49308 6132 49364 6142
rect 49308 5906 49364 6076
rect 49308 5854 49310 5906
rect 49362 5854 49364 5906
rect 49308 5842 49364 5854
rect 49756 5908 49812 6526
rect 49868 6244 49924 6254
rect 49868 6018 49924 6188
rect 49868 5966 49870 6018
rect 49922 5966 49924 6018
rect 49868 5954 49924 5966
rect 49756 5842 49812 5852
rect 50092 5236 50148 12908
rect 50764 12962 50820 12974
rect 50764 12910 50766 12962
rect 50818 12910 50820 12962
rect 50428 12852 50484 12862
rect 50764 12852 50820 12910
rect 50428 12850 50820 12852
rect 50428 12798 50430 12850
rect 50482 12798 50820 12850
rect 50428 12796 50820 12798
rect 50428 12786 50484 12796
rect 50204 12068 50260 12078
rect 50204 11974 50260 12012
rect 50428 11620 50484 11630
rect 50428 11506 50484 11564
rect 50428 11454 50430 11506
rect 50482 11454 50484 11506
rect 50428 11442 50484 11454
rect 50204 10500 50260 10510
rect 50204 10406 50260 10444
rect 50540 10164 50596 10174
rect 50428 9940 50484 9950
rect 50428 9846 50484 9884
rect 50204 8930 50260 8942
rect 50204 8878 50206 8930
rect 50258 8878 50260 8930
rect 50204 8708 50260 8878
rect 50204 8642 50260 8652
rect 50316 8932 50372 8942
rect 50204 6692 50260 6702
rect 50204 5906 50260 6636
rect 50204 5854 50206 5906
rect 50258 5854 50260 5906
rect 50204 5842 50260 5854
rect 50092 5170 50148 5180
rect 49084 5070 49086 5122
rect 49138 5070 49140 5122
rect 49084 5058 49140 5070
rect 49644 5124 49700 5134
rect 49644 5030 49700 5068
rect 48860 4956 49028 5012
rect 48748 4946 48804 4956
rect 48860 4788 48916 4798
rect 48748 4340 48804 4350
rect 48748 4246 48804 4284
rect 48300 4226 48356 4238
rect 48300 4174 48302 4226
rect 48354 4174 48356 4226
rect 47740 4116 47796 4126
rect 47740 4022 47796 4060
rect 48300 3668 48356 4174
rect 48300 3602 48356 3612
rect 48860 3666 48916 4732
rect 48860 3614 48862 3666
rect 48914 3614 48916 3666
rect 48860 3602 48916 3614
rect 47516 3266 47572 3276
rect 48076 2884 48132 2894
rect 48076 2790 48132 2828
rect 48748 2770 48804 2782
rect 48748 2718 48750 2770
rect 48802 2718 48804 2770
rect 47516 2548 47572 2558
rect 47516 2098 47572 2492
rect 48748 2212 48804 2718
rect 48748 2146 48804 2156
rect 48860 2660 48916 2670
rect 47516 2046 47518 2098
rect 47570 2046 47572 2098
rect 47516 2034 47572 2046
rect 48860 2098 48916 2604
rect 48860 2046 48862 2098
rect 48914 2046 48916 2098
rect 48860 2034 48916 2046
rect 48972 1988 49028 4956
rect 49420 4226 49476 4238
rect 49420 4174 49422 4226
rect 49474 4174 49476 4226
rect 49420 3668 49476 4174
rect 50204 4226 50260 4238
rect 50204 4174 50206 4226
rect 50258 4174 50260 4226
rect 50204 3780 50260 4174
rect 50204 3714 50260 3724
rect 49420 3602 49476 3612
rect 49868 3444 49924 3454
rect 49868 3350 49924 3388
rect 50316 2770 50372 8876
rect 50428 8260 50484 8270
rect 50428 8166 50484 8204
rect 50428 6690 50484 6702
rect 50428 6638 50430 6690
rect 50482 6638 50484 6690
rect 50428 3892 50484 6638
rect 50540 5122 50596 10108
rect 50540 5070 50542 5122
rect 50594 5070 50596 5122
rect 50540 5058 50596 5070
rect 50652 6916 50708 6926
rect 50428 3826 50484 3836
rect 50316 2718 50318 2770
rect 50370 2718 50372 2770
rect 50316 2706 50372 2718
rect 50428 3554 50484 3566
rect 50428 3502 50430 3554
rect 50482 3502 50484 3554
rect 49420 2660 49476 2670
rect 49420 2566 49476 2604
rect 50428 2548 50484 3502
rect 50428 2482 50484 2492
rect 50540 2884 50596 2894
rect 48972 1922 49028 1932
rect 49868 1876 49924 1886
rect 49868 1782 49924 1820
rect 49756 1428 49812 1438
rect 49756 1334 49812 1372
rect 48188 1314 48244 1326
rect 48188 1262 48190 1314
rect 48242 1262 48244 1314
rect 48188 868 48244 1262
rect 48748 1092 48804 1102
rect 48748 998 48804 1036
rect 50428 980 50484 990
rect 50428 886 50484 924
rect 48188 802 48244 812
rect 47292 578 47348 588
rect 50540 532 50596 2828
rect 50652 1986 50708 6860
rect 50764 6020 50820 12796
rect 50876 9716 50932 13468
rect 50876 9650 50932 9660
rect 50988 10498 51044 10510
rect 50988 10446 50990 10498
rect 51042 10446 51044 10498
rect 50988 9492 51044 10446
rect 50988 9426 51044 9436
rect 51100 9268 51156 13916
rect 51212 12852 51268 12862
rect 51212 12758 51268 12796
rect 51212 12290 51268 12302
rect 51212 12238 51214 12290
rect 51266 12238 51268 12290
rect 51212 10836 51268 12238
rect 51212 10770 51268 10780
rect 51436 11170 51492 11182
rect 51436 11118 51438 11170
rect 51490 11118 51492 11170
rect 51436 9940 51492 11118
rect 51436 9874 51492 9884
rect 51100 9202 51156 9212
rect 51436 9602 51492 9614
rect 51436 9550 51438 9602
rect 51490 9550 51492 9602
rect 51436 9044 51492 9550
rect 51436 8978 51492 8988
rect 50988 8930 51044 8942
rect 50988 8878 50990 8930
rect 51042 8878 51044 8930
rect 50988 8596 51044 8878
rect 50988 8530 51044 8540
rect 50876 8148 50932 8158
rect 50876 7698 50932 8092
rect 50876 7646 50878 7698
rect 50930 7646 50932 7698
rect 50876 7634 50932 7646
rect 51436 8034 51492 8046
rect 51436 7982 51438 8034
rect 51490 7982 51492 8034
rect 51436 7700 51492 7982
rect 51436 7634 51492 7644
rect 51324 7474 51380 7486
rect 51324 7422 51326 7474
rect 51378 7422 51380 7474
rect 51212 6356 51268 6366
rect 51212 6130 51268 6300
rect 51212 6078 51214 6130
rect 51266 6078 51268 6130
rect 51212 6066 51268 6078
rect 50764 5954 50820 5964
rect 51212 5460 51268 5470
rect 51212 5234 51268 5404
rect 51212 5182 51214 5234
rect 51266 5182 51268 5234
rect 51212 5170 51268 5182
rect 51100 5124 51156 5134
rect 51100 4564 51156 5068
rect 51100 4498 51156 4508
rect 51212 5012 51268 5022
rect 51212 4562 51268 4956
rect 51212 4510 51214 4562
rect 51266 4510 51268 4562
rect 51212 4498 51268 4510
rect 51100 3444 51156 3454
rect 51100 2772 51156 3388
rect 51212 3220 51268 3230
rect 51212 2994 51268 3164
rect 51212 2942 51214 2994
rect 51266 2942 51268 2994
rect 51212 2930 51268 2942
rect 51100 2706 51156 2716
rect 50652 1934 50654 1986
rect 50706 1934 50708 1986
rect 50652 1922 50708 1934
rect 51324 1314 51380 7422
rect 51436 7252 51492 7262
rect 51436 6578 51492 7196
rect 51436 6526 51438 6578
rect 51490 6526 51492 6578
rect 51436 6514 51492 6526
rect 51436 4116 51492 4126
rect 51436 3442 51492 4060
rect 51436 3390 51438 3442
rect 51490 3390 51492 3442
rect 51436 3378 51492 3390
rect 51548 2660 51604 2670
rect 51436 2324 51492 2334
rect 51436 1874 51492 2268
rect 51436 1822 51438 1874
rect 51490 1822 51492 1874
rect 51436 1810 51492 1822
rect 51324 1262 51326 1314
rect 51378 1262 51380 1314
rect 51324 1250 51380 1262
rect 50764 980 50820 990
rect 50764 886 50820 924
rect 50540 466 50596 476
rect 50876 308 50932 318
rect 48412 196 48468 206
rect 48412 112 48468 140
rect 50876 112 50932 252
rect 26908 18 26964 28
rect 28672 0 28784 112
rect 31136 0 31248 112
rect 33600 0 33712 112
rect 36064 0 36176 112
rect 38528 0 38640 112
rect 40992 0 41104 112
rect 43456 0 43568 112
rect 45920 0 46032 112
rect 48384 0 48496 112
rect 50848 0 50960 112
rect 51548 84 51604 2604
rect 51548 18 51604 28
<< via2 >>
rect 7084 14140 7140 14196
rect 252 13916 308 13972
rect 5516 13468 5572 13524
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 2268 13020 2324 13076
rect 812 12572 868 12628
rect 812 10444 868 10500
rect 1148 10556 1204 10612
rect 252 6860 308 6916
rect 1148 6748 1204 6804
rect 1260 9884 1316 9940
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 5180 12124 5236 12180
rect 2268 10668 2324 10724
rect 1708 9212 1764 9268
rect 1596 7644 1652 7700
rect 1596 6636 1652 6692
rect 1820 5740 1876 5796
rect 2380 3554 2436 3556
rect 2380 3502 2382 3554
rect 2382 3502 2434 3554
rect 2434 3502 2436 3554
rect 2380 3500 2436 3502
rect 2156 2882 2212 2884
rect 2156 2830 2158 2882
rect 2158 2830 2210 2882
rect 2210 2830 2212 2882
rect 2156 2828 2212 2830
rect 1596 2156 1652 2212
rect 3164 11954 3220 11956
rect 3164 11902 3166 11954
rect 3166 11902 3218 11954
rect 3218 11902 3220 11954
rect 3164 11900 3220 11902
rect 3500 11954 3556 11956
rect 3500 11902 3502 11954
rect 3502 11902 3554 11954
rect 3554 11902 3556 11954
rect 3500 11900 3556 11902
rect 4464 11786 4520 11788
rect 3276 11676 3332 11732
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 2716 10332 2772 10388
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 5068 10892 5124 10948
rect 4956 10668 5012 10724
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 3276 9660 3332 9716
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4956 9436 5012 9492
rect 4012 9380 4068 9382
rect 4464 8650 4520 8652
rect 4284 8540 4340 8596
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4284 7420 4340 7476
rect 2716 7196 2772 7252
rect 3612 7308 3668 7364
rect 3276 6748 3332 6804
rect 3276 6300 3332 6356
rect 3500 5068 3556 5124
rect 2716 3554 2772 3556
rect 2716 3502 2718 3554
rect 2718 3502 2770 3554
rect 2770 3502 2772 3554
rect 2716 3500 2772 3502
rect 2604 3276 2660 3332
rect 2492 1036 2548 1092
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 5292 11788 5348 11844
rect 6524 13074 6580 13076
rect 6524 13022 6526 13074
rect 6526 13022 6578 13074
rect 6578 13022 6580 13074
rect 6524 13020 6580 13022
rect 6524 12124 6580 12180
rect 6188 10444 6244 10500
rect 6076 9884 6132 9940
rect 5740 8540 5796 8596
rect 5516 7756 5572 7812
rect 5964 8092 6020 8148
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4172 4732 4228 4788
rect 3612 3164 3668 3220
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 5068 4508 5124 4564
rect 4844 4284 4900 4340
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 4172 1932 4228 1988
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 3276 924 3332 980
rect 5068 1148 5124 1204
rect 5180 3052 5236 3108
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 4172 476 4228 532
rect 4060 364 4116 420
rect 5516 5794 5572 5796
rect 5516 5742 5518 5794
rect 5518 5742 5570 5794
rect 5570 5742 5572 5794
rect 5516 5740 5572 5742
rect 5516 5122 5572 5124
rect 5516 5070 5518 5122
rect 5518 5070 5570 5122
rect 5570 5070 5572 5122
rect 5516 5068 5572 5070
rect 5292 2940 5348 2996
rect 5964 5628 6020 5684
rect 5964 5234 6020 5236
rect 5964 5182 5966 5234
rect 5966 5182 6018 5234
rect 6018 5182 6020 5234
rect 5964 5180 6020 5182
rect 5852 5068 5908 5124
rect 6300 7196 6356 7252
rect 6188 4620 6244 4676
rect 6188 3724 6244 3780
rect 6188 2492 6244 2548
rect 6748 11506 6804 11508
rect 6748 11454 6750 11506
rect 6750 11454 6802 11506
rect 6802 11454 6804 11506
rect 6748 11452 6804 11454
rect 41692 14140 41748 14196
rect 11564 14028 11620 14084
rect 9996 13580 10052 13636
rect 9772 13356 9828 13412
rect 7084 11452 7140 11508
rect 6860 10444 6916 10500
rect 7420 9884 7476 9940
rect 6524 5852 6580 5908
rect 6636 9436 6692 9492
rect 6524 5122 6580 5124
rect 6524 5070 6526 5122
rect 6526 5070 6578 5122
rect 6578 5070 6580 5122
rect 6524 5068 6580 5070
rect 6412 4508 6468 4564
rect 6972 9324 7028 9380
rect 6748 5906 6804 5908
rect 6748 5854 6750 5906
rect 6750 5854 6802 5906
rect 6802 5854 6804 5906
rect 6748 5852 6804 5854
rect 6748 5122 6804 5124
rect 6748 5070 6750 5122
rect 6750 5070 6802 5122
rect 6802 5070 6804 5122
rect 6748 5068 6804 5070
rect 6972 4732 7028 4788
rect 6972 3388 7028 3444
rect 6300 1484 6356 1540
rect 6524 1596 6580 1652
rect 5628 1372 5684 1428
rect 6972 2828 7028 2884
rect 6748 476 6804 532
rect 7644 9884 7700 9940
rect 7756 10780 7812 10836
rect 7644 8428 7700 8484
rect 7532 7084 7588 7140
rect 7532 5516 7588 5572
rect 7532 4508 7588 4564
rect 7756 5740 7812 5796
rect 11340 13468 11396 13524
rect 11004 13244 11060 13300
rect 8204 11954 8260 11956
rect 8204 11902 8206 11954
rect 8206 11902 8258 11954
rect 8258 11902 8260 11954
rect 8204 11900 8260 11902
rect 8540 11954 8596 11956
rect 8540 11902 8542 11954
rect 8542 11902 8594 11954
rect 8594 11902 8596 11954
rect 8540 11900 8596 11902
rect 9324 11900 9380 11956
rect 8092 10332 8148 10388
rect 7980 9212 8036 9268
rect 8764 10220 8820 10276
rect 8204 10108 8260 10164
rect 8652 9884 8708 9940
rect 8204 8988 8260 9044
rect 8316 9548 8372 9604
rect 8092 8764 8148 8820
rect 8540 9154 8596 9156
rect 8540 9102 8542 9154
rect 8542 9102 8594 9154
rect 8594 9102 8596 9154
rect 8540 9100 8596 9102
rect 8316 8316 8372 8372
rect 8764 9660 8820 9716
rect 8988 9714 9044 9716
rect 8988 9662 8990 9714
rect 8990 9662 9042 9714
rect 9042 9662 9044 9714
rect 8988 9660 9044 9662
rect 9548 10332 9604 10388
rect 10444 10834 10500 10836
rect 10444 10782 10446 10834
rect 10446 10782 10498 10834
rect 10498 10782 10500 10834
rect 10444 10780 10500 10782
rect 10332 10332 10388 10388
rect 10444 10050 10500 10052
rect 10444 9998 10446 10050
rect 10446 9998 10498 10050
rect 10498 9998 10500 10050
rect 10444 9996 10500 9998
rect 10668 10050 10724 10052
rect 10668 9998 10670 10050
rect 10670 9998 10722 10050
rect 10722 9998 10724 10050
rect 10668 9996 10724 9998
rect 8652 7980 8708 8036
rect 8876 9212 8932 9268
rect 7980 6076 8036 6132
rect 8092 7196 8148 7252
rect 8316 6860 8372 6916
rect 9324 8988 9380 9044
rect 9212 7868 9268 7924
rect 9212 7532 9268 7588
rect 9212 6748 9268 6804
rect 8316 5964 8372 6020
rect 8092 5516 8148 5572
rect 8204 5628 8260 5684
rect 7868 4508 7924 4564
rect 8092 4060 8148 4116
rect 8092 3164 8148 3220
rect 7644 3052 7700 3108
rect 7532 2828 7588 2884
rect 8316 5180 8372 5236
rect 8316 3836 8372 3892
rect 8764 4844 8820 4900
rect 8204 2380 8260 2436
rect 8764 2044 8820 2100
rect 7420 140 7476 196
rect 8988 1596 9044 1652
rect 5180 28 5236 84
rect 10108 9548 10164 9604
rect 9884 8258 9940 8260
rect 9884 8206 9886 8258
rect 9886 8206 9938 8258
rect 9938 8206 9940 8258
rect 9884 8204 9940 8206
rect 9772 8092 9828 8148
rect 10220 8258 10276 8260
rect 10220 8206 10222 8258
rect 10222 8206 10274 8258
rect 10274 8206 10276 8258
rect 10220 8204 10276 8206
rect 10556 7980 10612 8036
rect 9548 6690 9604 6692
rect 9548 6638 9550 6690
rect 9550 6638 9602 6690
rect 9602 6638 9604 6690
rect 9548 6636 9604 6638
rect 9884 6690 9940 6692
rect 9884 6638 9886 6690
rect 9886 6638 9938 6690
rect 9938 6638 9940 6690
rect 9884 6636 9940 6638
rect 9548 6188 9604 6244
rect 9772 5068 9828 5124
rect 9884 4620 9940 4676
rect 9884 2604 9940 2660
rect 9772 2492 9828 2548
rect 10108 6188 10164 6244
rect 10444 5404 10500 5460
rect 10220 4450 10276 4452
rect 10220 4398 10222 4450
rect 10222 4398 10274 4450
rect 10274 4398 10276 4450
rect 10220 4396 10276 4398
rect 10892 11788 10948 11844
rect 10780 6972 10836 7028
rect 11228 6748 11284 6804
rect 10892 5180 10948 5236
rect 11228 4732 11284 4788
rect 12348 14028 12404 14084
rect 11900 12962 11956 12964
rect 11900 12910 11902 12962
rect 11902 12910 11954 12962
rect 11954 12910 11956 12962
rect 11900 12908 11956 12910
rect 11900 12684 11956 12740
rect 11676 12402 11732 12404
rect 11676 12350 11678 12402
rect 11678 12350 11730 12402
rect 11730 12350 11732 12402
rect 11676 12348 11732 12350
rect 11788 12236 11844 12292
rect 12460 12572 12516 12628
rect 12236 11452 12292 11508
rect 12012 11228 12068 11284
rect 11900 11116 11956 11172
rect 11564 7644 11620 7700
rect 11676 7084 11732 7140
rect 11788 10108 11844 10164
rect 11900 9100 11956 9156
rect 11900 8316 11956 8372
rect 11900 8092 11956 8148
rect 11564 6636 11620 6692
rect 11452 4620 11508 4676
rect 11788 6412 11844 6468
rect 11340 3612 11396 3668
rect 11228 3164 11284 3220
rect 10556 2380 10612 2436
rect 9996 2156 10052 2212
rect 11676 5628 11732 5684
rect 11788 4396 11844 4452
rect 11676 4172 11732 4228
rect 11676 3612 11732 3668
rect 11228 1596 11284 1652
rect 11564 2716 11620 2772
rect 12572 10780 12628 10836
rect 12684 12796 12740 12852
rect 12460 10050 12516 10052
rect 12460 9998 12462 10050
rect 12462 9998 12514 10050
rect 12514 9998 12516 10050
rect 12460 9996 12516 9998
rect 12236 9436 12292 9492
rect 12124 9100 12180 9156
rect 12236 8930 12292 8932
rect 12236 8878 12238 8930
rect 12238 8878 12290 8930
rect 12290 8878 12292 8930
rect 12236 8876 12292 8878
rect 12124 8428 12180 8484
rect 12572 6860 12628 6916
rect 12796 11900 12852 11956
rect 12572 5852 12628 5908
rect 13356 13132 13412 13188
rect 13244 12236 13300 12292
rect 13356 12066 13412 12068
rect 13356 12014 13358 12066
rect 13358 12014 13410 12066
rect 13410 12014 13412 12066
rect 13356 12012 13412 12014
rect 13020 11788 13076 11844
rect 13020 11394 13076 11396
rect 13020 11342 13022 11394
rect 13022 11342 13074 11394
rect 13074 11342 13076 11394
rect 13020 11340 13076 11342
rect 13020 7980 13076 8036
rect 13916 13580 13972 13636
rect 14364 13356 14420 13412
rect 13692 12012 13748 12068
rect 14028 12012 14084 12068
rect 13916 11340 13972 11396
rect 13692 10668 13748 10724
rect 13804 11228 13860 11284
rect 13580 9996 13636 10052
rect 13804 9212 13860 9268
rect 13804 7308 13860 7364
rect 13244 7196 13300 7252
rect 13804 6748 13860 6804
rect 12796 5852 12852 5908
rect 13692 6636 13748 6692
rect 13356 5740 13412 5796
rect 13692 4396 13748 4452
rect 11788 3052 11844 3108
rect 11564 1596 11620 1652
rect 12460 2716 12516 2772
rect 12236 2268 12292 2324
rect 12460 1820 12516 1876
rect 12572 2380 12628 2436
rect 12572 924 12628 980
rect 12684 2268 12740 2324
rect 11900 476 11956 532
rect 14140 11004 14196 11060
rect 14364 12684 14420 12740
rect 14252 10892 14308 10948
rect 14028 9884 14084 9940
rect 14028 7474 14084 7476
rect 14028 7422 14030 7474
rect 14030 7422 14082 7474
rect 14082 7422 14084 7474
rect 14028 7420 14084 7422
rect 13916 6636 13972 6692
rect 14364 10108 14420 10164
rect 14700 13804 14756 13860
rect 14700 12684 14756 12740
rect 14924 13244 14980 13300
rect 14812 12572 14868 12628
rect 14588 12348 14644 12404
rect 14700 12460 14756 12516
rect 14588 11394 14644 11396
rect 14588 11342 14590 11394
rect 14590 11342 14642 11394
rect 14642 11342 14644 11394
rect 14588 11340 14644 11342
rect 14812 12290 14868 12292
rect 14812 12238 14814 12290
rect 14814 12238 14866 12290
rect 14866 12238 14868 12290
rect 14812 12236 14868 12238
rect 15148 13580 15204 13636
rect 15148 12012 15204 12068
rect 14924 10108 14980 10164
rect 14588 9826 14644 9828
rect 14588 9774 14590 9826
rect 14590 9774 14642 9826
rect 14642 9774 14644 9826
rect 14588 9772 14644 9774
rect 14812 9266 14868 9268
rect 14812 9214 14814 9266
rect 14814 9214 14866 9266
rect 14866 9214 14868 9266
rect 14812 9212 14868 9214
rect 14588 7084 14644 7140
rect 14364 5740 14420 5796
rect 14476 6524 14532 6580
rect 14252 4732 14308 4788
rect 13804 2604 13860 2660
rect 14140 2940 14196 2996
rect 14140 2604 14196 2660
rect 14476 4732 14532 4788
rect 14700 5852 14756 5908
rect 14812 5122 14868 5124
rect 14812 5070 14814 5122
rect 14814 5070 14866 5122
rect 14866 5070 14868 5122
rect 14812 5068 14868 5070
rect 15484 13580 15540 13636
rect 15372 12178 15428 12180
rect 15372 12126 15374 12178
rect 15374 12126 15426 12178
rect 15426 12126 15428 12178
rect 15372 12124 15428 12126
rect 15372 11564 15428 11620
rect 15932 13692 15988 13748
rect 15708 13468 15764 13524
rect 15820 12796 15876 12852
rect 15596 12348 15652 12404
rect 15372 10332 15428 10388
rect 15484 10220 15540 10276
rect 15260 9884 15316 9940
rect 16380 12572 16436 12628
rect 16156 12348 16212 12404
rect 16380 12348 16436 12404
rect 15932 11676 15988 11732
rect 16044 11340 16100 11396
rect 15932 10556 15988 10612
rect 15932 10220 15988 10276
rect 15708 9212 15764 9268
rect 15932 9212 15988 9268
rect 15484 9100 15540 9156
rect 15260 8316 15316 8372
rect 15148 7644 15204 7700
rect 15372 7644 15428 7700
rect 15372 7308 15428 7364
rect 15596 7362 15652 7364
rect 15596 7310 15598 7362
rect 15598 7310 15650 7362
rect 15650 7310 15652 7362
rect 15596 7308 15652 7310
rect 15484 6188 15540 6244
rect 15596 5404 15652 5460
rect 16156 10556 16212 10612
rect 16492 10668 16548 10724
rect 16492 9884 16548 9940
rect 16044 6188 16100 6244
rect 15148 5122 15204 5124
rect 15148 5070 15150 5122
rect 15150 5070 15202 5122
rect 15202 5070 15204 5122
rect 15148 5068 15204 5070
rect 15372 4844 15428 4900
rect 15596 4844 15652 4900
rect 14588 3052 14644 3108
rect 15820 3836 15876 3892
rect 15148 2940 15204 2996
rect 15372 3724 15428 3780
rect 15820 3612 15876 3668
rect 16828 13132 16884 13188
rect 16716 12460 16772 12516
rect 17164 13692 17220 13748
rect 17276 13580 17332 13636
rect 17164 13244 17220 13300
rect 17276 13356 17332 13412
rect 17052 12348 17108 12404
rect 17388 13244 17444 13300
rect 17388 12348 17444 12404
rect 16716 11452 16772 11508
rect 16940 10668 16996 10724
rect 17276 10498 17332 10500
rect 17276 10446 17278 10498
rect 17278 10446 17330 10498
rect 17330 10446 17332 10498
rect 17276 10444 17332 10446
rect 17052 8988 17108 9044
rect 17164 9548 17220 9604
rect 16828 7532 16884 7588
rect 16716 6412 16772 6468
rect 16380 5964 16436 6020
rect 17052 8764 17108 8820
rect 17052 7196 17108 7252
rect 17276 8540 17332 8596
rect 17164 6972 17220 7028
rect 17500 12236 17556 12292
rect 17612 12572 17668 12628
rect 17500 12012 17556 12068
rect 17500 10108 17556 10164
rect 16940 5516 16996 5572
rect 17836 13580 17892 13636
rect 17948 13132 18004 13188
rect 17836 12348 17892 12404
rect 17948 12124 18004 12180
rect 17724 9212 17780 9268
rect 18060 11228 18116 11284
rect 18396 13692 18452 13748
rect 18508 13132 18564 13188
rect 18284 12402 18340 12404
rect 18284 12350 18286 12402
rect 18286 12350 18338 12402
rect 18338 12350 18340 12402
rect 18284 12348 18340 12350
rect 18396 11452 18452 11508
rect 18284 11340 18340 11396
rect 18396 11228 18452 11284
rect 18284 10444 18340 10500
rect 18284 9324 18340 9380
rect 17724 8316 17780 8372
rect 18620 11340 18676 11396
rect 18732 13132 18788 13188
rect 18844 12460 18900 12516
rect 18844 12066 18900 12068
rect 18844 12014 18846 12066
rect 18846 12014 18898 12066
rect 18898 12014 18900 12066
rect 18844 12012 18900 12014
rect 18844 11506 18900 11508
rect 18844 11454 18846 11506
rect 18846 11454 18898 11506
rect 18898 11454 18900 11506
rect 18844 11452 18900 11454
rect 18956 11340 19012 11396
rect 18844 10892 18900 10948
rect 18732 9100 18788 9156
rect 18844 9884 18900 9940
rect 18956 9660 19012 9716
rect 19180 12850 19236 12852
rect 19180 12798 19182 12850
rect 19182 12798 19234 12850
rect 19234 12798 19236 12850
rect 19180 12796 19236 12798
rect 19516 12348 19572 12404
rect 19628 12290 19684 12292
rect 19628 12238 19630 12290
rect 19630 12238 19682 12290
rect 19682 12238 19684 12290
rect 19628 12236 19684 12238
rect 19404 9100 19460 9156
rect 18396 7756 18452 7812
rect 17948 7084 18004 7140
rect 18060 7308 18116 7364
rect 17724 6412 17780 6468
rect 17724 5964 17780 6020
rect 16716 4956 16772 5012
rect 16940 5068 16996 5124
rect 16268 3500 16324 3556
rect 16156 2828 16212 2884
rect 16828 2882 16884 2884
rect 16828 2830 16830 2882
rect 16830 2830 16882 2882
rect 16882 2830 16884 2882
rect 16828 2828 16884 2830
rect 15372 2268 15428 2324
rect 16716 2492 16772 2548
rect 14252 2044 14308 2100
rect 13468 1932 13524 1988
rect 13356 1708 13412 1764
rect 13356 1484 13412 1540
rect 13468 1372 13524 1428
rect 13916 1820 13972 1876
rect 12684 364 12740 420
rect 14476 1260 14532 1316
rect 16380 1596 16436 1652
rect 17276 4060 17332 4116
rect 17164 3948 17220 4004
rect 17164 3612 17220 3668
rect 16940 2156 16996 2212
rect 17164 3164 17220 3220
rect 17164 1932 17220 1988
rect 18508 7196 18564 7252
rect 19628 7532 19684 7588
rect 18956 7084 19012 7140
rect 19292 7084 19348 7140
rect 18732 6860 18788 6916
rect 19180 6860 19236 6916
rect 18732 6690 18788 6692
rect 18732 6638 18734 6690
rect 18734 6638 18786 6690
rect 18786 6638 18788 6690
rect 18732 6636 18788 6638
rect 18396 6412 18452 6468
rect 18060 5404 18116 5460
rect 18284 5292 18340 5348
rect 17948 4060 18004 4116
rect 18060 4508 18116 4564
rect 18508 5292 18564 5348
rect 18508 4732 18564 4788
rect 18284 4508 18340 4564
rect 18060 3724 18116 3780
rect 18620 3948 18676 4004
rect 18284 3276 18340 3332
rect 17388 1932 17444 1988
rect 18284 1932 18340 1988
rect 20188 13244 20244 13300
rect 20300 13692 20356 13748
rect 19964 11452 20020 11508
rect 20300 12124 20356 12180
rect 20300 11676 20356 11732
rect 21084 13692 21140 13748
rect 20748 13244 20804 13300
rect 21196 13186 21252 13188
rect 21196 13134 21198 13186
rect 21198 13134 21250 13186
rect 21250 13134 21252 13186
rect 21196 13132 21252 13134
rect 21308 12796 21364 12852
rect 21420 13692 21476 13748
rect 21084 12124 21140 12180
rect 21308 11900 21364 11956
rect 20076 10108 20132 10164
rect 19852 9826 19908 9828
rect 19852 9774 19854 9826
rect 19854 9774 19906 9826
rect 19906 9774 19908 9826
rect 19852 9772 19908 9774
rect 19964 8988 20020 9044
rect 19852 7420 19908 7476
rect 20076 8316 20132 8372
rect 21196 11788 21252 11844
rect 21196 11394 21252 11396
rect 21196 11342 21198 11394
rect 21198 11342 21250 11394
rect 21250 11342 21252 11394
rect 21196 11340 21252 11342
rect 20972 8540 21028 8596
rect 20972 8370 21028 8372
rect 20972 8318 20974 8370
rect 20974 8318 21026 8370
rect 21026 8318 21028 8370
rect 20972 8316 21028 8318
rect 20188 7980 20244 8036
rect 21308 10498 21364 10500
rect 21308 10446 21310 10498
rect 21310 10446 21362 10498
rect 21362 10446 21364 10498
rect 21308 10444 21364 10446
rect 21644 12402 21700 12404
rect 21644 12350 21646 12402
rect 21646 12350 21698 12402
rect 21698 12350 21700 12402
rect 21644 12348 21700 12350
rect 21532 11676 21588 11732
rect 21644 12124 21700 12180
rect 21196 8316 21252 8372
rect 21196 7868 21252 7924
rect 21308 7532 21364 7588
rect 20412 7420 20468 7476
rect 20636 7420 20692 7476
rect 19964 6748 20020 6804
rect 20188 6524 20244 6580
rect 18956 2940 19012 2996
rect 19180 2940 19236 2996
rect 18620 1596 18676 1652
rect 17612 588 17668 644
rect 18844 1484 18900 1540
rect 16716 476 16772 532
rect 19516 3164 19572 3220
rect 19516 2716 19572 2772
rect 19516 2210 19572 2212
rect 19516 2158 19518 2210
rect 19518 2158 19570 2210
rect 19570 2158 19572 2210
rect 19516 2156 19572 2158
rect 19852 2210 19908 2212
rect 19852 2158 19854 2210
rect 19854 2158 19906 2210
rect 19906 2158 19908 2210
rect 19852 2156 19908 2158
rect 20076 2716 20132 2772
rect 20076 2492 20132 2548
rect 20972 6076 21028 6132
rect 20748 5740 20804 5796
rect 20860 5628 20916 5684
rect 21644 10780 21700 10836
rect 21644 9884 21700 9940
rect 21532 8258 21588 8260
rect 21532 8206 21534 8258
rect 21534 8206 21586 8258
rect 21586 8206 21588 8258
rect 21532 8204 21588 8206
rect 21420 5740 21476 5796
rect 21532 7980 21588 8036
rect 21308 5068 21364 5124
rect 20972 3836 21028 3892
rect 21084 4508 21140 4564
rect 20860 3612 20916 3668
rect 19404 1596 19460 1652
rect 19180 1372 19236 1428
rect 20188 1372 20244 1428
rect 21196 4172 21252 4228
rect 20860 1202 20916 1204
rect 20860 1150 20862 1202
rect 20862 1150 20914 1202
rect 20914 1150 20916 1202
rect 20860 1148 20916 1150
rect 21084 1202 21140 1204
rect 21084 1150 21086 1202
rect 21086 1150 21138 1202
rect 21138 1150 21140 1202
rect 21084 1148 21140 1150
rect 19964 924 20020 980
rect 21420 4172 21476 4228
rect 21308 3612 21364 3668
rect 21308 2940 21364 2996
rect 21868 8540 21924 8596
rect 21868 7980 21924 8036
rect 21868 7586 21924 7588
rect 21868 7534 21870 7586
rect 21870 7534 21922 7586
rect 21922 7534 21924 7586
rect 21868 7532 21924 7534
rect 21756 4956 21812 5012
rect 21868 7084 21924 7140
rect 21756 4620 21812 4676
rect 22428 13132 22484 13188
rect 22540 13468 22596 13524
rect 22204 12348 22260 12404
rect 22428 12684 22484 12740
rect 22316 11676 22372 11732
rect 22204 11564 22260 11620
rect 22204 9660 22260 9716
rect 22204 8930 22260 8932
rect 22204 8878 22206 8930
rect 22206 8878 22258 8930
rect 22258 8878 22260 8930
rect 22204 8876 22260 8878
rect 22092 8764 22148 8820
rect 22092 8204 22148 8260
rect 22092 7532 22148 7588
rect 22204 7980 22260 8036
rect 21980 6524 22036 6580
rect 22092 6636 22148 6692
rect 21868 4060 21924 4116
rect 21756 2940 21812 2996
rect 21756 2380 21812 2436
rect 21644 2156 21700 2212
rect 21532 1820 21588 1876
rect 21196 700 21252 756
rect 21308 1596 21364 1652
rect 19852 252 19908 308
rect 21532 1596 21588 1652
rect 21532 1372 21588 1428
rect 22876 13468 22932 13524
rect 23324 13468 23380 13524
rect 23324 12348 23380 12404
rect 22764 11564 22820 11620
rect 22988 11900 23044 11956
rect 22764 11228 22820 11284
rect 22652 10780 22708 10836
rect 22876 11004 22932 11060
rect 22540 10108 22596 10164
rect 22428 8258 22484 8260
rect 22428 8206 22430 8258
rect 22430 8206 22482 8258
rect 22482 8206 22484 8258
rect 22428 8204 22484 8206
rect 22316 6300 22372 6356
rect 22428 7868 22484 7924
rect 22764 10108 22820 10164
rect 23324 11618 23380 11620
rect 23324 11566 23326 11618
rect 23326 11566 23378 11618
rect 23378 11566 23380 11618
rect 23324 11564 23380 11566
rect 24220 13356 24276 13412
rect 24892 13692 24948 13748
rect 25116 13580 25172 13636
rect 25340 13580 25396 13636
rect 24332 13244 24388 13300
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 23996 13132 24052 13188
rect 25564 13468 25620 13524
rect 25676 13692 25732 13748
rect 23660 12572 23716 12628
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 24556 12348 24612 12404
rect 24668 11900 24724 11956
rect 23772 11788 23828 11844
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 23660 11004 23716 11060
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24220 11004 24276 11060
rect 24012 10948 24068 10950
rect 24668 11282 24724 11284
rect 24668 11230 24670 11282
rect 24670 11230 24722 11282
rect 24722 11230 24724 11282
rect 24668 11228 24724 11230
rect 24332 10892 24388 10948
rect 23436 10834 23492 10836
rect 23436 10782 23438 10834
rect 23438 10782 23490 10834
rect 23490 10782 23492 10834
rect 23436 10780 23492 10782
rect 23212 9884 23268 9940
rect 23436 10444 23492 10500
rect 23212 9324 23268 9380
rect 22876 8540 22932 8596
rect 22764 8258 22820 8260
rect 22764 8206 22766 8258
rect 22766 8206 22818 8258
rect 22818 8206 22820 8258
rect 22764 8204 22820 8206
rect 23212 8204 23268 8260
rect 24108 10220 24164 10276
rect 24464 10218 24520 10220
rect 24332 10108 24388 10164
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24556 9938 24612 9940
rect 24556 9886 24558 9938
rect 24558 9886 24610 9938
rect 24610 9886 24612 9938
rect 24556 9884 24612 9886
rect 25564 12796 25620 12852
rect 25452 12348 25508 12404
rect 25452 12124 25508 12180
rect 25116 11676 25172 11732
rect 25340 10780 25396 10836
rect 25564 10444 25620 10500
rect 25676 12124 25732 12180
rect 25004 10220 25060 10276
rect 24892 9884 24948 9940
rect 25116 9660 25172 9716
rect 25452 9714 25508 9716
rect 25452 9662 25454 9714
rect 25454 9662 25506 9714
rect 25506 9662 25508 9714
rect 25452 9660 25508 9662
rect 24332 9324 24388 9380
rect 25004 9324 25060 9380
rect 25340 9100 25396 9156
rect 23772 9042 23828 9044
rect 23772 8990 23774 9042
rect 23774 8990 23826 9042
rect 23826 8990 23828 9042
rect 23772 8988 23828 8990
rect 24332 9042 24388 9044
rect 24332 8990 24334 9042
rect 24334 8990 24386 9042
rect 24386 8990 24388 9042
rect 24332 8988 24388 8990
rect 24556 8988 24612 9044
rect 23996 8876 24052 8932
rect 23996 8652 24052 8708
rect 24332 8540 24388 8596
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24668 7980 24724 8036
rect 23436 7868 23492 7924
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24220 7868 24276 7924
rect 23324 7644 23380 7700
rect 24108 7586 24164 7588
rect 24108 7534 24110 7586
rect 24110 7534 24162 7586
rect 24162 7534 24164 7586
rect 24108 7532 24164 7534
rect 24108 7084 24164 7140
rect 22988 6860 23044 6916
rect 23436 6860 23492 6916
rect 22988 6636 23044 6692
rect 23324 6412 23380 6468
rect 23660 6412 23716 6468
rect 25228 8930 25284 8932
rect 25228 8878 25230 8930
rect 25230 8878 25282 8930
rect 25282 8878 25284 8930
rect 25228 8876 25284 8878
rect 24220 6972 24276 7028
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 25004 7084 25060 7140
rect 25228 8204 25284 8260
rect 24672 7028 24728 7030
rect 24892 6972 24948 7028
rect 24444 6412 24500 6468
rect 23804 6298 23860 6300
rect 23660 6188 23716 6244
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24556 6018 24612 6020
rect 24556 5966 24558 6018
rect 24558 5966 24610 6018
rect 24610 5966 24612 6018
rect 24556 5964 24612 5966
rect 24332 5516 24388 5572
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 22204 5068 22260 5124
rect 23212 5068 23268 5124
rect 22652 4956 22708 5012
rect 22092 2156 22148 2212
rect 22540 4172 22596 4228
rect 22204 1596 22260 1652
rect 22652 3388 22708 3444
rect 23660 4732 23716 4788
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24332 4732 24388 4788
rect 24012 4676 24068 4678
rect 24220 4620 24276 4676
rect 25004 6748 25060 6804
rect 24556 5122 24612 5124
rect 24556 5070 24558 5122
rect 24558 5070 24610 5122
rect 24610 5070 24612 5122
rect 24556 5068 24612 5070
rect 24892 5122 24948 5124
rect 24892 5070 24894 5122
rect 24894 5070 24946 5122
rect 24946 5070 24948 5122
rect 24892 5068 24948 5070
rect 24780 4732 24836 4788
rect 25228 5740 25284 5796
rect 25452 8876 25508 8932
rect 25452 8258 25508 8260
rect 25452 8206 25454 8258
rect 25454 8206 25506 8258
rect 25506 8206 25508 8258
rect 25452 8204 25508 8206
rect 25452 7756 25508 7812
rect 25900 13804 25956 13860
rect 26012 12348 26068 12404
rect 25900 11676 25956 11732
rect 25788 11004 25844 11060
rect 25900 11340 25956 11396
rect 25900 10444 25956 10500
rect 26124 10108 26180 10164
rect 26124 9548 26180 9604
rect 25788 9154 25844 9156
rect 25788 9102 25790 9154
rect 25790 9102 25842 9154
rect 25842 9102 25844 9154
rect 25788 9100 25844 9102
rect 25788 8876 25844 8932
rect 25788 7756 25844 7812
rect 25676 7532 25732 7588
rect 25452 6636 25508 6692
rect 25340 5292 25396 5348
rect 25452 5010 25508 5012
rect 25452 4958 25454 5010
rect 25454 4958 25506 5010
rect 25506 4958 25508 5010
rect 25452 4956 25508 4958
rect 25004 4732 25060 4788
rect 24668 4396 24724 4452
rect 24220 3948 24276 4004
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 24892 3948 24948 4004
rect 22540 1596 22596 1652
rect 24220 3724 24276 3780
rect 23884 3276 23940 3332
rect 23660 3164 23716 3220
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 25116 3778 25172 3780
rect 25116 3726 25118 3778
rect 25118 3726 25170 3778
rect 25170 3726 25172 3778
rect 25116 3724 25172 3726
rect 24332 3500 24388 3556
rect 25340 3778 25396 3780
rect 25340 3726 25342 3778
rect 25342 3726 25394 3778
rect 25394 3726 25396 3778
rect 25340 3724 25396 3726
rect 25228 3500 25284 3556
rect 25452 3612 25508 3668
rect 24444 3276 24500 3332
rect 25340 3276 25396 3332
rect 24892 3164 24948 3220
rect 24332 3052 24388 3108
rect 24332 2380 24388 2436
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24892 2380 24948 2436
rect 25788 3164 25844 3220
rect 24672 2324 24728 2326
rect 23660 1596 23716 1652
rect 23804 1594 23860 1596
rect 23100 1484 23156 1540
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24220 1484 24276 1540
rect 21868 1372 21924 1428
rect 24780 1596 24836 1652
rect 26348 13132 26404 13188
rect 26460 12684 26516 12740
rect 26460 11340 26516 11396
rect 26348 9996 26404 10052
rect 26348 9772 26404 9828
rect 27580 13132 27636 13188
rect 27132 12572 27188 12628
rect 26572 9548 26628 9604
rect 26460 5964 26516 6020
rect 26572 8764 26628 8820
rect 26236 5516 26292 5572
rect 27356 11116 27412 11172
rect 26796 9826 26852 9828
rect 26796 9774 26798 9826
rect 26798 9774 26850 9826
rect 26850 9774 26852 9826
rect 26796 9772 26852 9774
rect 27132 9826 27188 9828
rect 27132 9774 27134 9826
rect 27134 9774 27186 9826
rect 27186 9774 27188 9826
rect 27132 9772 27188 9774
rect 27132 8876 27188 8932
rect 26684 8204 26740 8260
rect 26908 8540 26964 8596
rect 26572 5180 26628 5236
rect 26124 4060 26180 4116
rect 26012 3052 26068 3108
rect 25788 2044 25844 2100
rect 25228 1820 25284 1876
rect 25004 1596 25060 1652
rect 26124 1820 26180 1876
rect 26348 4060 26404 4116
rect 25228 1484 25284 1540
rect 22540 700 22596 756
rect 22540 364 22596 420
rect 22764 700 22820 756
rect 22316 252 22372 308
rect 22876 476 22932 532
rect 24332 812 24388 868
rect 23996 700 24052 756
rect 23772 140 23828 196
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 27356 6300 27412 6356
rect 27356 5964 27412 6020
rect 27356 5628 27412 5684
rect 26908 4508 26964 4564
rect 27132 4508 27188 4564
rect 27020 4450 27076 4452
rect 27020 4398 27022 4450
rect 27022 4398 27074 4450
rect 27074 4398 27076 4450
rect 27020 4396 27076 4398
rect 26796 3500 26852 3556
rect 26796 2940 26852 2996
rect 26684 2828 26740 2884
rect 26460 2716 26516 2772
rect 27244 3442 27300 3444
rect 27244 3390 27246 3442
rect 27246 3390 27298 3442
rect 27298 3390 27300 3442
rect 27244 3388 27300 3390
rect 28028 14028 28084 14084
rect 28140 13580 28196 13636
rect 28140 12572 28196 12628
rect 28140 12348 28196 12404
rect 28028 12290 28084 12292
rect 28028 12238 28030 12290
rect 28030 12238 28082 12290
rect 28082 12238 28084 12290
rect 28028 12236 28084 12238
rect 27804 12124 27860 12180
rect 27580 11452 27636 11508
rect 27804 11788 27860 11844
rect 27804 11452 27860 11508
rect 28028 11788 28084 11844
rect 27804 10332 27860 10388
rect 27804 10108 27860 10164
rect 27580 6188 27636 6244
rect 27804 6412 27860 6468
rect 28140 9772 28196 9828
rect 28028 6076 28084 6132
rect 27692 5628 27748 5684
rect 28700 13244 28756 13300
rect 28476 12236 28532 12292
rect 28476 10780 28532 10836
rect 28588 8540 28644 8596
rect 28700 12124 28756 12180
rect 28700 8092 28756 8148
rect 28812 9884 28868 9940
rect 28364 6860 28420 6916
rect 29148 11788 29204 11844
rect 28924 7308 28980 7364
rect 29484 11676 29540 11732
rect 29484 11452 29540 11508
rect 29260 9884 29316 9940
rect 29148 9548 29204 9604
rect 29148 7532 29204 7588
rect 29372 9548 29428 9604
rect 29260 7420 29316 7476
rect 29820 13804 29876 13860
rect 30268 13804 30324 13860
rect 30044 13692 30100 13748
rect 29820 13580 29876 13636
rect 30044 12572 30100 12628
rect 29932 11452 29988 11508
rect 29820 11228 29876 11284
rect 29596 8652 29652 8708
rect 29708 11116 29764 11172
rect 30156 12236 30212 12292
rect 30940 13020 30996 13076
rect 30828 12684 30884 12740
rect 30492 12124 30548 12180
rect 30716 12572 30772 12628
rect 30156 11564 30212 11620
rect 30268 11788 30324 11844
rect 30044 9772 30100 9828
rect 30156 11340 30212 11396
rect 30156 9436 30212 9492
rect 29484 7084 29540 7140
rect 29148 6748 29204 6804
rect 30156 8146 30212 8148
rect 30156 8094 30158 8146
rect 30158 8094 30210 8146
rect 30210 8094 30212 8146
rect 30156 8092 30212 8094
rect 29596 6748 29652 6804
rect 29708 7980 29764 8036
rect 28924 5516 28980 5572
rect 30380 9324 30436 9380
rect 30604 9996 30660 10052
rect 30380 8988 30436 9044
rect 29932 7474 29988 7476
rect 29932 7422 29934 7474
rect 29934 7422 29986 7474
rect 29986 7422 29988 7474
rect 29932 7420 29988 7422
rect 29708 5516 29764 5572
rect 29820 6860 29876 6916
rect 29932 6690 29988 6692
rect 29932 6638 29934 6690
rect 29934 6638 29986 6690
rect 29986 6638 29988 6690
rect 29932 6636 29988 6638
rect 29820 5404 29876 5460
rect 29036 4284 29092 4340
rect 29596 4844 29652 4900
rect 27356 2940 27412 2996
rect 26460 2380 26516 2436
rect 26348 1148 26404 1204
rect 26796 1036 26852 1092
rect 29820 3442 29876 3444
rect 29820 3390 29822 3442
rect 29822 3390 29874 3442
rect 29874 3390 29876 3442
rect 29820 3388 29876 3390
rect 30156 6188 30212 6244
rect 30380 5964 30436 6020
rect 30716 9884 30772 9940
rect 31164 12796 31220 12852
rect 31612 13580 31668 13636
rect 31388 12124 31444 12180
rect 31612 13132 31668 13188
rect 30940 11228 30996 11284
rect 30828 6972 30884 7028
rect 30940 10332 30996 10388
rect 31164 10332 31220 10388
rect 31052 9996 31108 10052
rect 31052 8876 31108 8932
rect 31500 9772 31556 9828
rect 30940 6076 30996 6132
rect 31164 8092 31220 8148
rect 30604 5964 30660 6020
rect 30156 4396 30212 4452
rect 30268 5628 30324 5684
rect 30268 3276 30324 3332
rect 30380 3388 30436 3444
rect 30156 3164 30212 3220
rect 29596 2828 29652 2884
rect 28812 2604 28868 2660
rect 25228 476 25284 532
rect 26796 364 26852 420
rect 23996 140 24052 196
rect 26236 140 26292 196
rect 9660 28 9716 84
rect 27692 812 27748 868
rect 28700 1820 28756 1876
rect 28812 1372 28868 1428
rect 30044 2492 30100 2548
rect 30380 2380 30436 2436
rect 30604 2940 30660 2996
rect 30604 2380 30660 2436
rect 30828 1932 30884 1988
rect 30156 1708 30212 1764
rect 30828 1484 30884 1540
rect 30156 1036 30212 1092
rect 30044 700 30100 756
rect 31724 12348 31780 12404
rect 31836 13356 31892 13412
rect 31836 10556 31892 10612
rect 31612 8876 31668 8932
rect 31836 8146 31892 8148
rect 31836 8094 31838 8146
rect 31838 8094 31890 8146
rect 31890 8094 31892 8146
rect 31836 8092 31892 8094
rect 31724 6412 31780 6468
rect 31724 4396 31780 4452
rect 31500 4172 31556 4228
rect 32284 14028 32340 14084
rect 32284 13020 32340 13076
rect 32396 12908 32452 12964
rect 32508 11788 32564 11844
rect 32396 11564 32452 11620
rect 32508 10444 32564 10500
rect 32956 13916 33012 13972
rect 33068 13132 33124 13188
rect 33068 9996 33124 10052
rect 32732 9660 32788 9716
rect 32508 9436 32564 9492
rect 32508 8764 32564 8820
rect 32396 8092 32452 8148
rect 32284 7644 32340 7700
rect 31948 6860 32004 6916
rect 31948 6412 32004 6468
rect 33180 8540 33236 8596
rect 33292 10780 33348 10836
rect 32732 8428 32788 8484
rect 32956 7980 33012 8036
rect 32732 6300 32788 6356
rect 32956 7532 33012 7588
rect 32508 5068 32564 5124
rect 32844 5404 32900 5460
rect 32844 4508 32900 4564
rect 33180 5516 33236 5572
rect 33068 4450 33124 4452
rect 33068 4398 33070 4450
rect 33070 4398 33122 4450
rect 33122 4398 33124 4450
rect 33068 4396 33124 4398
rect 31836 3948 31892 4004
rect 32620 3500 32676 3556
rect 31948 3052 32004 3108
rect 31948 2604 32004 2660
rect 32732 3442 32788 3444
rect 32732 3390 32734 3442
rect 32734 3390 32786 3442
rect 32786 3390 32788 3442
rect 32732 3388 32788 3390
rect 33628 12684 33684 12740
rect 33628 12460 33684 12516
rect 33628 10780 33684 10836
rect 33740 12012 33796 12068
rect 34300 13132 34356 13188
rect 34076 13020 34132 13076
rect 33404 10332 33460 10388
rect 33516 8988 33572 9044
rect 33628 9996 33684 10052
rect 33516 8764 33572 8820
rect 33740 9660 33796 9716
rect 33852 11788 33908 11844
rect 33852 9100 33908 9156
rect 33740 8988 33796 9044
rect 34300 11676 34356 11732
rect 34188 10108 34244 10164
rect 33964 8652 34020 8708
rect 34076 9324 34132 9380
rect 34076 8092 34132 8148
rect 33740 7756 33796 7812
rect 33964 7868 34020 7924
rect 33852 7644 33908 7700
rect 33628 6748 33684 6804
rect 33740 6860 33796 6916
rect 33740 6076 33796 6132
rect 33516 5740 33572 5796
rect 33852 5740 33908 5796
rect 33404 5628 33460 5684
rect 33292 3948 33348 4004
rect 33404 5180 33460 5236
rect 33180 3500 33236 3556
rect 33628 5068 33684 5124
rect 33516 4508 33572 4564
rect 34748 12572 34804 12628
rect 34524 9884 34580 9940
rect 34636 10108 34692 10164
rect 35196 13132 35252 13188
rect 35308 13804 35364 13860
rect 35420 13356 35476 13412
rect 35532 13244 35588 13300
rect 35308 11004 35364 11060
rect 34972 8540 35028 8596
rect 35308 8204 35364 8260
rect 34300 7756 34356 7812
rect 35308 7196 35364 7252
rect 35308 5852 35364 5908
rect 35308 5516 35364 5572
rect 35308 4732 35364 4788
rect 33964 4620 34020 4676
rect 35308 4172 35364 4228
rect 33404 3052 33460 3108
rect 35532 12684 35588 12740
rect 35532 10332 35588 10388
rect 35644 11228 35700 11284
rect 35532 9996 35588 10052
rect 35532 8428 35588 8484
rect 35532 6636 35588 6692
rect 36092 13020 36148 13076
rect 36764 13692 36820 13748
rect 36540 13244 36596 13300
rect 36876 13356 36932 13412
rect 36316 12124 36372 12180
rect 35756 8540 35812 8596
rect 35644 6412 35700 6468
rect 36540 13020 36596 13076
rect 36316 9100 36372 9156
rect 36652 9324 36708 9380
rect 36764 8428 36820 8484
rect 36652 8316 36708 8372
rect 35868 4956 35924 5012
rect 35980 6300 36036 6356
rect 35532 4284 35588 4340
rect 35756 4732 35812 4788
rect 33180 2940 33236 2996
rect 33404 1986 33460 1988
rect 33404 1934 33406 1986
rect 33406 1934 33458 1986
rect 33458 1934 33460 1986
rect 33404 1932 33460 1934
rect 32732 1708 32788 1764
rect 33516 812 33572 868
rect 33628 2156 33684 2212
rect 32732 140 32788 196
rect 35420 3276 35476 3332
rect 35980 4620 36036 4676
rect 36092 5964 36148 6020
rect 35756 3164 35812 3220
rect 35196 1596 35252 1652
rect 35308 3052 35364 3108
rect 35308 1260 35364 1316
rect 36652 3612 36708 3668
rect 37100 12796 37156 12852
rect 37324 12796 37380 12852
rect 37212 12684 37268 12740
rect 37660 13356 37716 13412
rect 37772 13186 37828 13188
rect 37772 13134 37774 13186
rect 37774 13134 37826 13186
rect 37826 13134 37828 13186
rect 37772 13132 37828 13134
rect 37436 12460 37492 12516
rect 38108 13244 38164 13300
rect 37996 13186 38052 13188
rect 37996 13134 37998 13186
rect 37998 13134 38050 13186
rect 38050 13134 38052 13186
rect 37996 13132 38052 13134
rect 37884 12348 37940 12404
rect 37100 11564 37156 11620
rect 38332 13020 38388 13076
rect 38668 13468 38724 13524
rect 38668 13244 38724 13300
rect 38444 12572 38500 12628
rect 38220 11676 38276 11732
rect 37548 11228 37604 11284
rect 37772 10332 37828 10388
rect 37212 10108 37268 10164
rect 37548 10220 37604 10276
rect 36988 9212 37044 9268
rect 36988 4956 37044 5012
rect 37100 7756 37156 7812
rect 37884 9884 37940 9940
rect 37660 5740 37716 5796
rect 37100 3388 37156 3444
rect 37548 4620 37604 4676
rect 36652 1148 36708 1204
rect 36988 2044 37044 2100
rect 36988 476 37044 532
rect 38332 9826 38388 9828
rect 38332 9774 38334 9826
rect 38334 9774 38386 9826
rect 38386 9774 38388 9826
rect 38332 9772 38388 9774
rect 38668 12684 38724 12740
rect 39004 13468 39060 13524
rect 38780 12124 38836 12180
rect 38892 11676 38948 11732
rect 38780 11116 38836 11172
rect 38668 10108 38724 10164
rect 38780 9996 38836 10052
rect 38780 9660 38836 9716
rect 38668 9548 38724 9604
rect 38220 9154 38276 9156
rect 38220 9102 38222 9154
rect 38222 9102 38274 9154
rect 38274 9102 38276 9154
rect 38220 9100 38276 9102
rect 38556 9100 38612 9156
rect 38668 8988 38724 9044
rect 38668 8540 38724 8596
rect 39228 12684 39284 12740
rect 39340 12348 39396 12404
rect 39452 12236 39508 12292
rect 39116 10220 39172 10276
rect 39564 9996 39620 10052
rect 39676 10780 39732 10836
rect 38780 7420 38836 7476
rect 38332 6972 38388 7028
rect 38444 6860 38500 6916
rect 37996 5516 38052 5572
rect 38108 6636 38164 6692
rect 37884 4620 37940 4676
rect 37884 3836 37940 3892
rect 37660 2492 37716 2548
rect 37884 1372 37940 1428
rect 37548 252 37604 308
rect 38444 6524 38500 6580
rect 38612 6524 38668 6580
rect 39116 6524 39172 6580
rect 39564 8764 39620 8820
rect 38668 5234 38724 5236
rect 38668 5182 38670 5234
rect 38670 5182 38722 5234
rect 38722 5182 38724 5234
rect 38668 5180 38724 5182
rect 38892 5234 38948 5236
rect 38892 5182 38894 5234
rect 38894 5182 38946 5234
rect 38946 5182 38948 5234
rect 38892 5180 38948 5182
rect 38780 5068 38836 5124
rect 38780 3276 38836 3332
rect 38556 2940 38612 2996
rect 38892 2940 38948 2996
rect 38220 2716 38276 2772
rect 38668 2492 38724 2548
rect 38668 2268 38724 2324
rect 39452 5234 39508 5236
rect 39452 5182 39454 5234
rect 39454 5182 39506 5234
rect 39506 5182 39508 5234
rect 39452 5180 39508 5182
rect 40012 13692 40068 13748
rect 40684 13580 40740 13636
rect 40124 13132 40180 13188
rect 40236 13244 40292 13300
rect 41244 13356 41300 13412
rect 41580 13020 41636 13076
rect 40012 12460 40068 12516
rect 39900 10780 39956 10836
rect 40012 11564 40068 11620
rect 39788 9548 39844 9604
rect 40012 9436 40068 9492
rect 39900 6748 39956 6804
rect 39788 5068 39844 5124
rect 40796 12572 40852 12628
rect 40908 12124 40964 12180
rect 40348 9826 40404 9828
rect 40348 9774 40350 9826
rect 40350 9774 40402 9826
rect 40402 9774 40404 9826
rect 40348 9772 40404 9774
rect 41132 12124 41188 12180
rect 41020 11788 41076 11844
rect 40908 10444 40964 10500
rect 40796 10050 40852 10052
rect 40796 9998 40798 10050
rect 40798 9998 40850 10050
rect 40850 9998 40852 10050
rect 40796 9996 40852 9998
rect 41020 9996 41076 10052
rect 40908 9548 40964 9604
rect 40460 8876 40516 8932
rect 40236 8540 40292 8596
rect 40460 8092 40516 8148
rect 40236 7420 40292 7476
rect 40124 6076 40180 6132
rect 40572 6524 40628 6580
rect 39564 2492 39620 2548
rect 39452 2380 39508 2436
rect 39228 2268 39284 2324
rect 38892 2210 38948 2212
rect 38892 2158 38894 2210
rect 38894 2158 38946 2210
rect 38946 2158 38948 2210
rect 38892 2156 38948 2158
rect 39116 2210 39172 2212
rect 39116 2158 39118 2210
rect 39118 2158 39170 2210
rect 39170 2158 39172 2210
rect 39116 2156 39172 2158
rect 39676 2098 39732 2100
rect 39676 2046 39678 2098
rect 39678 2046 39730 2098
rect 39730 2046 39732 2098
rect 39676 2044 39732 2046
rect 38108 1260 38164 1316
rect 37996 140 38052 196
rect 38556 140 38612 196
rect 40348 3612 40404 3668
rect 40572 4844 40628 4900
rect 40684 4732 40740 4788
rect 40460 2828 40516 2884
rect 40908 7532 40964 7588
rect 41468 10332 41524 10388
rect 41244 10108 41300 10164
rect 41356 10220 41412 10276
rect 41356 8316 41412 8372
rect 41132 6188 41188 6244
rect 40796 2604 40852 2660
rect 41020 5404 41076 5460
rect 40236 1484 40292 1540
rect 39788 140 39844 196
rect 51100 13916 51156 13972
rect 42588 13804 42644 13860
rect 43708 13468 43764 13524
rect 50876 13468 50932 13524
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 45052 13186 45108 13188
rect 45052 13134 45054 13186
rect 45054 13134 45106 13186
rect 45106 13134 45108 13186
rect 45052 13132 45108 13134
rect 48076 13020 48132 13076
rect 42364 12684 42420 12740
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 42924 11900 42980 11956
rect 43036 12012 43092 12068
rect 41804 11394 41860 11396
rect 41804 11342 41806 11394
rect 41806 11342 41858 11394
rect 41858 11342 41860 11394
rect 41804 11340 41860 11342
rect 42476 10834 42532 10836
rect 42476 10782 42478 10834
rect 42478 10782 42530 10834
rect 42530 10782 42532 10834
rect 42476 10780 42532 10782
rect 42028 10610 42084 10612
rect 42028 10558 42030 10610
rect 42030 10558 42082 10610
rect 42082 10558 42084 10610
rect 42028 10556 42084 10558
rect 41916 9884 41972 9940
rect 41804 9548 41860 9604
rect 41804 7868 41860 7924
rect 42140 9884 42196 9940
rect 42252 9714 42308 9716
rect 42252 9662 42254 9714
rect 42254 9662 42306 9714
rect 42306 9662 42308 9714
rect 42252 9660 42308 9662
rect 42140 9324 42196 9380
rect 42364 9100 42420 9156
rect 42140 8652 42196 8708
rect 42140 6748 42196 6804
rect 41916 4844 41972 4900
rect 41916 4620 41972 4676
rect 42700 4956 42756 5012
rect 43148 6524 43204 6580
rect 43260 11676 43316 11732
rect 43036 3052 43092 3108
rect 42364 2940 42420 2996
rect 41468 2044 41524 2100
rect 45164 12908 45220 12964
rect 44268 11676 44324 11732
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44940 11452 44996 11508
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 43932 9660 43988 9716
rect 44492 9714 44548 9716
rect 44492 9662 44494 9714
rect 44494 9662 44546 9714
rect 44546 9662 44548 9714
rect 44492 9660 44548 9662
rect 43596 9548 43652 9604
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 43596 9212 43652 9268
rect 43260 812 43316 868
rect 43484 6860 43540 6916
rect 44940 9772 44996 9828
rect 47180 12962 47236 12964
rect 47180 12910 47182 12962
rect 47182 12910 47234 12962
rect 47234 12910 47236 12962
rect 47180 12908 47236 12910
rect 45276 12348 45332 12404
rect 48188 12572 48244 12628
rect 48748 12178 48804 12180
rect 48748 12126 48750 12178
rect 48750 12126 48802 12178
rect 48802 12126 48804 12178
rect 48748 12124 48804 12126
rect 45612 11340 45668 11396
rect 45276 11116 45332 11172
rect 45164 9100 45220 9156
rect 44492 8876 44548 8932
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 45388 8428 45444 8484
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44268 6748 44324 6804
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 43596 4284 43652 4340
rect 44156 4338 44212 4340
rect 44156 4286 44158 4338
rect 44158 4286 44210 4338
rect 44210 4286 44212 4338
rect 44156 4284 44212 4286
rect 44380 6412 44436 6468
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 45052 5292 45108 5348
rect 49756 12124 49812 12180
rect 49644 11788 49700 11844
rect 48860 11394 48916 11396
rect 48860 11342 48862 11394
rect 48862 11342 48914 11394
rect 48914 11342 48916 11394
rect 48860 11340 48916 11342
rect 49868 11282 49924 11284
rect 49868 11230 49870 11282
rect 49870 11230 49922 11282
rect 49922 11230 49924 11282
rect 49868 11228 49924 11230
rect 48748 10780 48804 10836
rect 47852 10668 47908 10724
rect 47516 10498 47572 10500
rect 47516 10446 47518 10498
rect 47518 10446 47570 10498
rect 47570 10446 47572 10498
rect 47516 10444 47572 10446
rect 47740 10498 47796 10500
rect 47740 10446 47742 10498
rect 47742 10446 47794 10498
rect 47794 10446 47796 10498
rect 47740 10444 47796 10446
rect 47068 9996 47124 10052
rect 45724 5964 45780 6020
rect 46172 7980 46228 8036
rect 46732 5068 46788 5124
rect 46172 4732 46228 4788
rect 46508 4956 46564 5012
rect 45612 4508 45668 4564
rect 45388 4284 45444 4340
rect 44716 4226 44772 4228
rect 44716 4174 44718 4226
rect 44718 4174 44770 4226
rect 44770 4174 44772 4226
rect 44716 4172 44772 4174
rect 44464 3946 44520 3948
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 45276 3836 45332 3892
rect 45612 3554 45668 3556
rect 45612 3502 45614 3554
rect 45614 3502 45666 3554
rect 45666 3502 45668 3554
rect 45612 3500 45668 3502
rect 45836 3554 45892 3556
rect 45836 3502 45838 3554
rect 45838 3502 45890 3554
rect 45890 3502 45892 3554
rect 45836 3500 45892 3502
rect 43596 3388 43652 3444
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 45164 2882 45220 2884
rect 45164 2830 45166 2882
rect 45166 2830 45218 2882
rect 45218 2830 45220 2882
rect 45164 2828 45220 2830
rect 45948 2658 46004 2660
rect 45948 2606 45950 2658
rect 45950 2606 46002 2658
rect 46002 2606 46004 2658
rect 45948 2604 46004 2606
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 44268 1874 44324 1876
rect 44268 1822 44270 1874
rect 44270 1822 44322 1874
rect 44322 1822 44324 1874
rect 44268 1820 44324 1822
rect 46844 4844 46900 4900
rect 47404 4114 47460 4116
rect 47404 4062 47406 4114
rect 47406 4062 47458 4114
rect 47458 4062 47460 4114
rect 47404 4060 47460 4062
rect 47068 2770 47124 2772
rect 47068 2718 47070 2770
rect 47070 2718 47122 2770
rect 47122 2718 47124 2770
rect 47068 2716 47124 2718
rect 46732 2098 46788 2100
rect 46732 2046 46734 2098
rect 46734 2046 46786 2098
rect 46786 2046 46788 2098
rect 46732 2044 46788 2046
rect 46956 2098 47012 2100
rect 46956 2046 46958 2098
rect 46958 2046 47010 2098
rect 47010 2046 47012 2098
rect 46956 2044 47012 2046
rect 46172 1708 46228 1764
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 45948 1372 46004 1428
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 47180 1202 47236 1204
rect 47180 1150 47182 1202
rect 47182 1150 47234 1202
rect 47234 1150 47236 1202
rect 47180 1148 47236 1150
rect 49644 10332 49700 10388
rect 48300 10108 48356 10164
rect 48076 8988 48132 9044
rect 47852 6188 47908 6244
rect 47964 8652 48020 8708
rect 47740 6018 47796 6020
rect 47740 5966 47742 6018
rect 47742 5966 47794 6018
rect 47794 5966 47796 6018
rect 47740 5964 47796 5966
rect 48300 8930 48356 8932
rect 48300 8878 48302 8930
rect 48302 8878 48354 8930
rect 48354 8878 48356 8930
rect 48300 8876 48356 8878
rect 48748 8764 48804 8820
rect 48188 8146 48244 8148
rect 48188 8094 48190 8146
rect 48190 8094 48242 8146
rect 48242 8094 48244 8146
rect 48188 8092 48244 8094
rect 48300 7420 48356 7476
rect 48748 7308 48804 7364
rect 48188 7196 48244 7252
rect 48076 6636 48132 6692
rect 48972 9772 49028 9828
rect 48972 6860 49028 6916
rect 48524 6524 48580 6580
rect 48076 5964 48132 6020
rect 47964 5628 48020 5684
rect 49084 9660 49140 9716
rect 48748 4956 48804 5012
rect 48972 6076 49028 6132
rect 49868 9714 49924 9716
rect 49868 9662 49870 9714
rect 49870 9662 49922 9714
rect 49922 9662 49924 9714
rect 49868 9660 49924 9662
rect 49644 9266 49700 9268
rect 49644 9214 49646 9266
rect 49646 9214 49698 9266
rect 49698 9214 49700 9266
rect 49644 9212 49700 9214
rect 49196 8370 49252 8372
rect 49196 8318 49198 8370
rect 49198 8318 49250 8370
rect 49250 8318 49252 8370
rect 49196 8316 49252 8318
rect 49532 8092 49588 8148
rect 49980 7532 50036 7588
rect 49644 6748 49700 6804
rect 49308 6076 49364 6132
rect 49868 6188 49924 6244
rect 49756 5852 49812 5908
rect 50204 12066 50260 12068
rect 50204 12014 50206 12066
rect 50206 12014 50258 12066
rect 50258 12014 50260 12066
rect 50204 12012 50260 12014
rect 50428 11564 50484 11620
rect 50204 10498 50260 10500
rect 50204 10446 50206 10498
rect 50206 10446 50258 10498
rect 50258 10446 50260 10498
rect 50204 10444 50260 10446
rect 50540 10108 50596 10164
rect 50428 9938 50484 9940
rect 50428 9886 50430 9938
rect 50430 9886 50482 9938
rect 50482 9886 50484 9938
rect 50428 9884 50484 9886
rect 50204 8652 50260 8708
rect 50316 8876 50372 8932
rect 50204 6636 50260 6692
rect 50092 5180 50148 5236
rect 49644 5122 49700 5124
rect 49644 5070 49646 5122
rect 49646 5070 49698 5122
rect 49698 5070 49700 5122
rect 49644 5068 49700 5070
rect 48860 4732 48916 4788
rect 48748 4338 48804 4340
rect 48748 4286 48750 4338
rect 48750 4286 48802 4338
rect 48802 4286 48804 4338
rect 48748 4284 48804 4286
rect 47740 4114 47796 4116
rect 47740 4062 47742 4114
rect 47742 4062 47794 4114
rect 47794 4062 47796 4114
rect 47740 4060 47796 4062
rect 48300 3612 48356 3668
rect 47516 3276 47572 3332
rect 48076 2882 48132 2884
rect 48076 2830 48078 2882
rect 48078 2830 48130 2882
rect 48130 2830 48132 2882
rect 48076 2828 48132 2830
rect 47516 2492 47572 2548
rect 48748 2156 48804 2212
rect 48860 2604 48916 2660
rect 50204 3724 50260 3780
rect 49420 3612 49476 3668
rect 49868 3442 49924 3444
rect 49868 3390 49870 3442
rect 49870 3390 49922 3442
rect 49922 3390 49924 3442
rect 49868 3388 49924 3390
rect 50428 8258 50484 8260
rect 50428 8206 50430 8258
rect 50430 8206 50482 8258
rect 50482 8206 50484 8258
rect 50428 8204 50484 8206
rect 50652 6860 50708 6916
rect 50428 3836 50484 3892
rect 49420 2658 49476 2660
rect 49420 2606 49422 2658
rect 49422 2606 49474 2658
rect 49474 2606 49476 2658
rect 49420 2604 49476 2606
rect 50428 2492 50484 2548
rect 50540 2828 50596 2884
rect 48972 1932 49028 1988
rect 49868 1874 49924 1876
rect 49868 1822 49870 1874
rect 49870 1822 49922 1874
rect 49922 1822 49924 1874
rect 49868 1820 49924 1822
rect 49756 1426 49812 1428
rect 49756 1374 49758 1426
rect 49758 1374 49810 1426
rect 49810 1374 49812 1426
rect 49756 1372 49812 1374
rect 48748 1090 48804 1092
rect 48748 1038 48750 1090
rect 48750 1038 48802 1090
rect 48802 1038 48804 1090
rect 48748 1036 48804 1038
rect 50428 978 50484 980
rect 50428 926 50430 978
rect 50430 926 50482 978
rect 50482 926 50484 978
rect 50428 924 50484 926
rect 48188 812 48244 868
rect 47292 588 47348 644
rect 50876 9660 50932 9716
rect 50988 9436 51044 9492
rect 51212 12850 51268 12852
rect 51212 12798 51214 12850
rect 51214 12798 51266 12850
rect 51266 12798 51268 12850
rect 51212 12796 51268 12798
rect 51212 10780 51268 10836
rect 51436 9884 51492 9940
rect 51100 9212 51156 9268
rect 51436 8988 51492 9044
rect 50988 8540 51044 8596
rect 50876 8092 50932 8148
rect 51436 7644 51492 7700
rect 51212 6300 51268 6356
rect 50764 5964 50820 6020
rect 51212 5404 51268 5460
rect 51100 5068 51156 5124
rect 51100 4508 51156 4564
rect 51212 4956 51268 5012
rect 51100 3388 51156 3444
rect 51212 3164 51268 3220
rect 51100 2716 51156 2772
rect 51436 7196 51492 7252
rect 51436 4060 51492 4116
rect 51548 2604 51604 2660
rect 51436 2268 51492 2324
rect 50764 978 50820 980
rect 50764 926 50766 978
rect 50766 926 50818 978
rect 50818 926 50820 978
rect 50764 924 50820 926
rect 50540 476 50596 532
rect 50876 252 50932 308
rect 48412 140 48468 196
rect 26908 28 26964 84
rect 51548 28 51604 84
<< metal3 >>
rect 7074 14140 7084 14196
rect 7140 14140 32340 14196
rect 32284 14084 32340 14140
rect 38612 14140 41692 14196
rect 41748 14140 41758 14196
rect 11554 14028 11564 14084
rect 11620 14028 12348 14084
rect 12404 14028 12414 14084
rect 14700 14028 16156 14084
rect 16212 14028 16222 14084
rect 16370 14028 16380 14084
rect 16436 14028 26684 14084
rect 26740 14028 26750 14084
rect 28018 14028 28028 14084
rect 28084 14028 32060 14084
rect 32116 14028 32126 14084
rect 32274 14028 32284 14084
rect 32340 14028 32350 14084
rect 0 13972 112 14000
rect 0 13916 252 13972
rect 308 13916 318 13972
rect 0 13888 112 13916
rect 14700 13860 14756 14028
rect 38612 13972 38668 14140
rect 52640 13972 52752 14000
rect 14914 13916 14924 13972
rect 14980 13916 21420 13972
rect 21476 13916 21486 13972
rect 22866 13916 22876 13972
rect 22932 13916 32956 13972
rect 33012 13916 33022 13972
rect 34524 13916 38668 13972
rect 51090 13916 51100 13972
rect 51156 13916 52752 13972
rect 34524 13860 34580 13916
rect 52640 13888 52752 13916
rect 14690 13804 14700 13860
rect 14756 13804 14766 13860
rect 15092 13804 25900 13860
rect 25956 13804 25966 13860
rect 29362 13804 29372 13860
rect 29428 13804 29820 13860
rect 29876 13804 29886 13860
rect 30258 13804 30268 13860
rect 30324 13804 34580 13860
rect 35298 13804 35308 13860
rect 35364 13804 42588 13860
rect 42644 13804 42654 13860
rect 15092 13748 15148 13804
rect 13570 13692 13580 13748
rect 13636 13692 15148 13748
rect 15260 13692 15932 13748
rect 15988 13692 15998 13748
rect 17154 13692 17164 13748
rect 17220 13692 18396 13748
rect 18452 13692 18462 13748
rect 20290 13692 20300 13748
rect 20356 13692 21084 13748
rect 21140 13692 21150 13748
rect 21410 13692 21420 13748
rect 21476 13692 24892 13748
rect 24948 13692 24958 13748
rect 25666 13692 25676 13748
rect 25732 13692 30044 13748
rect 30100 13692 30110 13748
rect 30268 13692 34692 13748
rect 36754 13692 36764 13748
rect 36820 13692 40012 13748
rect 40068 13692 40078 13748
rect 15260 13636 15316 13692
rect 30268 13636 30324 13692
rect 34636 13636 34692 13692
rect 9986 13580 9996 13636
rect 10052 13580 13916 13636
rect 13972 13580 13982 13636
rect 15138 13580 15148 13636
rect 15204 13580 15316 13636
rect 15474 13580 15484 13636
rect 15540 13580 17276 13636
rect 17332 13580 17342 13636
rect 17826 13580 17836 13636
rect 17892 13580 24892 13636
rect 24948 13580 24958 13636
rect 25106 13580 25116 13636
rect 25172 13580 25210 13636
rect 25330 13580 25340 13636
rect 25396 13580 28140 13636
rect 28196 13580 28206 13636
rect 29810 13580 29820 13636
rect 29876 13580 30324 13636
rect 31602 13580 31612 13636
rect 31668 13580 34580 13636
rect 34636 13580 40684 13636
rect 40740 13580 40750 13636
rect 0 13524 112 13552
rect 34524 13524 34580 13580
rect 52640 13524 52752 13552
rect 0 13468 5516 13524
rect 5572 13468 5582 13524
rect 11330 13468 11340 13524
rect 11396 13468 15708 13524
rect 15764 13468 15774 13524
rect 16146 13468 16156 13524
rect 16212 13468 22540 13524
rect 22596 13468 22606 13524
rect 22866 13468 22876 13524
rect 22932 13468 23324 13524
rect 23380 13468 23390 13524
rect 23548 13468 25172 13524
rect 25554 13468 25564 13524
rect 25620 13468 32732 13524
rect 32788 13468 32798 13524
rect 34524 13468 38668 13524
rect 38724 13468 38734 13524
rect 38994 13468 39004 13524
rect 39060 13468 43708 13524
rect 43764 13468 43774 13524
rect 50866 13468 50876 13524
rect 50932 13468 52752 13524
rect 0 13440 112 13468
rect 23548 13412 23604 13468
rect 25116 13412 25172 13468
rect 52640 13440 52752 13468
rect 9762 13356 9772 13412
rect 9828 13356 14364 13412
rect 14420 13356 14430 13412
rect 14588 13356 17276 13412
rect 17332 13356 17342 13412
rect 18722 13356 18732 13412
rect 18788 13356 21868 13412
rect 21924 13356 21934 13412
rect 22194 13356 22204 13412
rect 22260 13356 23604 13412
rect 24182 13356 24220 13412
rect 24276 13356 24286 13412
rect 25116 13356 26460 13412
rect 26516 13356 26526 13412
rect 26684 13356 31836 13412
rect 31892 13356 31902 13412
rect 32050 13356 32060 13412
rect 32116 13356 33852 13412
rect 33908 13356 33918 13412
rect 35410 13356 35420 13412
rect 35476 13356 36876 13412
rect 36932 13356 36942 13412
rect 37650 13356 37660 13412
rect 37716 13356 41244 13412
rect 41300 13356 41310 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 14588 13300 14644 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 26684 13300 26740 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 10994 13244 11004 13300
rect 11060 13244 14644 13300
rect 14914 13244 14924 13300
rect 14980 13244 17164 13300
rect 17220 13244 17230 13300
rect 17378 13244 17388 13300
rect 17444 13244 20188 13300
rect 20244 13244 20254 13300
rect 20710 13244 20748 13300
rect 20804 13244 20814 13300
rect 20972 13244 24332 13300
rect 24388 13244 24398 13300
rect 24882 13244 24892 13300
rect 24948 13244 26740 13300
rect 26898 13244 26908 13300
rect 26964 13244 28700 13300
rect 28756 13244 28766 13300
rect 30930 13244 30940 13300
rect 30996 13244 35532 13300
rect 35588 13244 35598 13300
rect 36530 13244 36540 13300
rect 36596 13244 38108 13300
rect 38164 13244 38174 13300
rect 38658 13244 38668 13300
rect 38724 13244 40236 13300
rect 40292 13244 40302 13300
rect 20972 13188 21028 13244
rect 13346 13132 13356 13188
rect 13412 13132 16828 13188
rect 16884 13132 16894 13188
rect 17938 13132 17948 13188
rect 18004 13132 18508 13188
rect 18564 13132 18574 13188
rect 18722 13132 18732 13188
rect 18788 13132 21028 13188
rect 21186 13132 21196 13188
rect 21252 13132 22428 13188
rect 22484 13132 22494 13188
rect 23650 13132 23660 13188
rect 23716 13132 23996 13188
rect 24052 13132 24062 13188
rect 24210 13132 24220 13188
rect 24276 13132 26348 13188
rect 26404 13132 26414 13188
rect 27570 13132 27580 13188
rect 27636 13132 31612 13188
rect 31668 13132 31678 13188
rect 33058 13132 33068 13188
rect 33124 13132 34300 13188
rect 34356 13132 34366 13188
rect 35186 13132 35196 13188
rect 35252 13132 37772 13188
rect 37828 13132 37996 13188
rect 38052 13132 38062 13188
rect 40114 13132 40124 13188
rect 40180 13132 45052 13188
rect 45108 13132 45118 13188
rect 0 13076 112 13104
rect 52640 13076 52752 13104
rect 0 13020 2268 13076
rect 2324 13020 2334 13076
rect 6514 13020 6524 13076
rect 6580 13020 30940 13076
rect 30996 13020 31006 13076
rect 31154 13020 31164 13076
rect 31220 13020 32284 13076
rect 32340 13020 32350 13076
rect 33618 13020 33628 13076
rect 33684 13020 34076 13076
rect 34132 13020 34142 13076
rect 36082 13020 36092 13076
rect 36148 13020 36540 13076
rect 36596 13020 36606 13076
rect 38322 13020 38332 13076
rect 38388 13020 41580 13076
rect 41636 13020 41646 13076
rect 48066 13020 48076 13076
rect 48132 13020 52752 13076
rect 0 12992 112 13020
rect 52640 12992 52752 13020
rect 11890 12908 11900 12964
rect 11956 12908 13244 12964
rect 13300 12908 13310 12964
rect 13468 12908 26908 12964
rect 28242 12908 28252 12964
rect 28308 12908 32396 12964
rect 32452 12908 32462 12964
rect 32722 12908 32732 12964
rect 32788 12908 39564 12964
rect 39620 12908 39630 12964
rect 45154 12908 45164 12964
rect 45220 12908 47180 12964
rect 47236 12908 47246 12964
rect 13468 12852 13524 12908
rect 26852 12852 26908 12908
rect 12674 12796 12684 12852
rect 12740 12796 13524 12852
rect 13580 12796 15820 12852
rect 15876 12796 15886 12852
rect 16044 12796 18732 12852
rect 18788 12796 18798 12852
rect 19170 12796 19180 12852
rect 19236 12796 21308 12852
rect 21364 12796 21374 12852
rect 21532 12796 25340 12852
rect 25396 12796 25406 12852
rect 25554 12796 25564 12852
rect 25620 12796 26740 12852
rect 26852 12796 30940 12852
rect 30996 12796 31006 12852
rect 31154 12796 31164 12852
rect 31220 12796 37100 12852
rect 37156 12796 37166 12852
rect 37314 12796 37324 12852
rect 37380 12796 51212 12852
rect 51268 12796 51278 12852
rect 13580 12740 13636 12796
rect 16044 12740 16100 12796
rect 21532 12740 21588 12796
rect 26684 12740 26740 12796
rect 11890 12684 11900 12740
rect 11956 12684 13636 12740
rect 14354 12684 14364 12740
rect 14420 12684 14700 12740
rect 14756 12684 14766 12740
rect 15138 12684 15148 12740
rect 15204 12684 16100 12740
rect 16482 12684 16492 12740
rect 16548 12684 21588 12740
rect 22418 12684 22428 12740
rect 22484 12684 26460 12740
rect 26516 12684 26526 12740
rect 26684 12684 30604 12740
rect 30660 12684 30670 12740
rect 30818 12684 30828 12740
rect 30884 12684 33628 12740
rect 33684 12684 33694 12740
rect 33842 12684 33852 12740
rect 33908 12684 35532 12740
rect 35588 12684 35598 12740
rect 37202 12684 37212 12740
rect 37268 12684 38668 12740
rect 38724 12684 38734 12740
rect 39218 12684 39228 12740
rect 39284 12684 42364 12740
rect 42420 12684 42430 12740
rect 0 12628 112 12656
rect 52640 12628 52752 12656
rect 0 12572 812 12628
rect 868 12572 878 12628
rect 12450 12572 12460 12628
rect 12516 12572 14812 12628
rect 14868 12572 14878 12628
rect 16370 12572 16380 12628
rect 16436 12572 16446 12628
rect 17602 12572 17612 12628
rect 17668 12572 19124 12628
rect 19282 12572 19292 12628
rect 19348 12572 23660 12628
rect 23716 12572 23726 12628
rect 24210 12572 24220 12628
rect 24276 12572 27132 12628
rect 27188 12572 27198 12628
rect 28130 12572 28140 12628
rect 28196 12572 30044 12628
rect 30100 12572 30110 12628
rect 30706 12572 30716 12628
rect 30772 12572 34748 12628
rect 34804 12572 34814 12628
rect 38434 12572 38444 12628
rect 38500 12572 40796 12628
rect 40852 12572 40862 12628
rect 48178 12572 48188 12628
rect 48244 12572 52752 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 16380 12516 16436 12572
rect 19068 12516 19124 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 52640 12544 52752 12572
rect 14690 12460 14700 12516
rect 14756 12460 16436 12516
rect 16706 12460 16716 12516
rect 16772 12460 18844 12516
rect 18900 12460 18910 12516
rect 19068 12460 23604 12516
rect 23548 12404 23604 12460
rect 24332 12460 33628 12516
rect 33684 12460 33694 12516
rect 37426 12460 37436 12516
rect 37492 12460 40012 12516
rect 40068 12460 40078 12516
rect 24332 12404 24388 12460
rect 11666 12348 11676 12404
rect 11732 12348 14588 12404
rect 14644 12348 14654 12404
rect 15586 12348 15596 12404
rect 15652 12348 16156 12404
rect 16212 12348 16222 12404
rect 16370 12348 16380 12404
rect 16436 12348 17052 12404
rect 17108 12348 17118 12404
rect 17378 12348 17388 12404
rect 17444 12348 17836 12404
rect 17892 12348 17902 12404
rect 18274 12348 18284 12404
rect 18340 12348 19516 12404
rect 19572 12348 19582 12404
rect 19730 12348 19740 12404
rect 19796 12348 21140 12404
rect 21634 12348 21644 12404
rect 21700 12348 22204 12404
rect 22260 12348 22270 12404
rect 22428 12348 23324 12404
rect 23380 12348 23390 12404
rect 23548 12348 24388 12404
rect 24546 12348 24556 12404
rect 24612 12348 24892 12404
rect 24948 12348 24958 12404
rect 25442 12348 25452 12404
rect 25508 12348 26012 12404
rect 26068 12348 26078 12404
rect 28130 12348 28140 12404
rect 28196 12348 31724 12404
rect 31780 12348 31790 12404
rect 31938 12348 31948 12404
rect 32004 12348 33964 12404
rect 34020 12348 34030 12404
rect 37874 12348 37884 12404
rect 37940 12348 39340 12404
rect 39396 12348 39406 12404
rect 39554 12348 39564 12404
rect 39620 12348 45276 12404
rect 45332 12348 45342 12404
rect 21084 12292 21140 12348
rect 22428 12292 22484 12348
rect 11778 12236 11788 12292
rect 11844 12236 13244 12292
rect 13300 12236 13310 12292
rect 14802 12236 14812 12292
rect 14868 12236 17500 12292
rect 17556 12236 17566 12292
rect 17714 12236 17724 12292
rect 17780 12236 19404 12292
rect 19460 12236 19470 12292
rect 19618 12236 19628 12292
rect 19684 12236 20748 12292
rect 20804 12236 20814 12292
rect 21084 12236 22484 12292
rect 23426 12236 23436 12292
rect 23492 12236 28028 12292
rect 28084 12236 28476 12292
rect 28532 12236 28542 12292
rect 30146 12236 30156 12292
rect 30212 12236 39452 12292
rect 39508 12236 39518 12292
rect 0 12180 112 12208
rect 52640 12180 52752 12208
rect 0 12124 5180 12180
rect 5236 12124 5246 12180
rect 6514 12124 6524 12180
rect 6580 12124 15148 12180
rect 15204 12124 15214 12180
rect 15362 12124 15372 12180
rect 15428 12124 17612 12180
rect 17668 12124 17678 12180
rect 17938 12124 17948 12180
rect 18004 12124 20300 12180
rect 20356 12124 20366 12180
rect 20514 12124 20524 12180
rect 20580 12124 21084 12180
rect 21140 12124 21150 12180
rect 21634 12124 21644 12180
rect 21700 12124 25452 12180
rect 25508 12124 25518 12180
rect 25666 12124 25676 12180
rect 25732 12124 27804 12180
rect 27860 12124 27870 12180
rect 28690 12124 28700 12180
rect 28756 12124 30492 12180
rect 30548 12124 30558 12180
rect 31378 12124 31388 12180
rect 31444 12124 36316 12180
rect 36372 12124 36382 12180
rect 38770 12124 38780 12180
rect 38836 12124 40908 12180
rect 40964 12124 40974 12180
rect 41122 12124 41132 12180
rect 41188 12124 48748 12180
rect 48804 12124 48814 12180
rect 49746 12124 49756 12180
rect 49812 12124 52752 12180
rect 0 12096 112 12124
rect 52640 12096 52752 12124
rect 13346 12012 13356 12068
rect 13412 12012 13692 12068
rect 13748 12012 13758 12068
rect 14018 12012 14028 12068
rect 14084 12012 15148 12068
rect 15204 12012 15214 12068
rect 17490 12012 17500 12068
rect 17556 12012 18844 12068
rect 18900 12012 18910 12068
rect 19068 12012 26348 12068
rect 26404 12012 26414 12068
rect 26572 12012 28252 12068
rect 28308 12012 28318 12068
rect 28466 12012 28476 12068
rect 28532 12012 33740 12068
rect 33796 12012 33806 12068
rect 33954 12012 33964 12068
rect 34020 12012 39116 12068
rect 39172 12012 39182 12068
rect 43026 12012 43036 12068
rect 43092 12012 50204 12068
rect 50260 12012 50270 12068
rect 19068 11956 19124 12012
rect 26572 11956 26628 12012
rect 3154 11900 3164 11956
rect 3220 11900 3500 11956
rect 3556 11900 7364 11956
rect 8194 11900 8204 11956
rect 8260 11900 8540 11956
rect 8596 11900 9324 11956
rect 9380 11900 9390 11956
rect 12786 11900 12796 11956
rect 12852 11900 17948 11956
rect 18004 11900 18014 11956
rect 18610 11900 18620 11956
rect 18676 11900 19124 11956
rect 21298 11900 21308 11956
rect 21364 11900 22316 11956
rect 22372 11900 22382 11956
rect 22978 11900 22988 11956
rect 23044 11900 24668 11956
rect 24724 11900 24734 11956
rect 24882 11900 24892 11956
rect 24948 11900 26628 11956
rect 26786 11900 26796 11956
rect 26852 11900 42924 11956
rect 42980 11900 42990 11956
rect 5282 11788 5292 11844
rect 5348 11788 6804 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 0 11676 3276 11732
rect 3332 11676 3342 11732
rect 0 11648 112 11676
rect 6748 11620 6804 11788
rect 7308 11732 7364 11900
rect 10882 11788 10892 11844
rect 10948 11788 13020 11844
rect 13076 11788 13086 11844
rect 13458 11788 13468 11844
rect 13524 11788 14924 11844
rect 14980 11788 14990 11844
rect 15708 11788 18060 11844
rect 18116 11788 18126 11844
rect 18722 11788 18732 11844
rect 18788 11788 18798 11844
rect 20076 11788 20188 11844
rect 20244 11788 20254 11844
rect 21186 11788 21196 11844
rect 21252 11788 23772 11844
rect 23828 11788 23838 11844
rect 25106 11788 25116 11844
rect 25172 11788 27804 11844
rect 27860 11788 27870 11844
rect 28018 11788 28028 11844
rect 28084 11788 29148 11844
rect 29204 11788 29214 11844
rect 30258 11788 30268 11844
rect 30324 11788 32508 11844
rect 32564 11788 32574 11844
rect 33842 11788 33852 11844
rect 33908 11788 41020 11844
rect 41076 11788 41086 11844
rect 49634 11788 49644 11844
rect 49700 11788 51044 11844
rect 15708 11732 15764 11788
rect 18732 11732 18788 11788
rect 20076 11732 20132 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 50988 11732 51044 11788
rect 52640 11732 52752 11760
rect 7308 11676 15764 11732
rect 15922 11676 15932 11732
rect 15988 11676 18508 11732
rect 18564 11676 18574 11732
rect 18732 11676 20132 11732
rect 20290 11676 20300 11732
rect 20356 11676 20394 11732
rect 21522 11676 21532 11732
rect 21588 11676 22316 11732
rect 22372 11676 22382 11732
rect 22530 11676 22540 11732
rect 22596 11676 24220 11732
rect 24276 11676 24286 11732
rect 24882 11676 24892 11732
rect 24948 11676 25116 11732
rect 25172 11676 25182 11732
rect 25890 11676 25900 11732
rect 25956 11676 28476 11732
rect 28532 11676 28542 11732
rect 29474 11676 29484 11732
rect 29540 11676 34300 11732
rect 34356 11676 34366 11732
rect 38210 11676 38220 11732
rect 38276 11676 38892 11732
rect 38948 11676 38958 11732
rect 43250 11676 43260 11732
rect 43316 11676 44268 11732
rect 44324 11676 44334 11732
rect 50988 11676 52752 11732
rect 52640 11648 52752 11676
rect 6748 11564 13468 11620
rect 13524 11564 13534 11620
rect 15362 11564 15372 11620
rect 15428 11564 22204 11620
rect 22260 11564 22270 11620
rect 22754 11564 22764 11620
rect 22820 11564 23324 11620
rect 23380 11564 23390 11620
rect 23548 11564 30156 11620
rect 30212 11564 30222 11620
rect 32386 11564 32396 11620
rect 32452 11564 35532 11620
rect 35588 11564 35598 11620
rect 37090 11564 37100 11620
rect 37156 11564 40012 11620
rect 40068 11564 40078 11620
rect 41794 11564 41804 11620
rect 41860 11564 50428 11620
rect 50484 11564 50494 11620
rect 23548 11508 23604 11564
rect 6738 11452 6748 11508
rect 6804 11452 7084 11508
rect 7140 11452 7150 11508
rect 12226 11452 12236 11508
rect 12292 11452 16492 11508
rect 16548 11452 16558 11508
rect 16706 11452 16716 11508
rect 16772 11452 18396 11508
rect 18452 11452 18462 11508
rect 18834 11452 18844 11508
rect 18900 11452 19964 11508
rect 20020 11452 20030 11508
rect 20178 11452 20188 11508
rect 20244 11452 23604 11508
rect 23660 11452 27356 11508
rect 27412 11452 27422 11508
rect 27570 11452 27580 11508
rect 27636 11452 27646 11508
rect 27794 11452 27804 11508
rect 27860 11452 29484 11508
rect 29540 11452 29550 11508
rect 29922 11452 29932 11508
rect 29988 11452 44940 11508
rect 44996 11452 45006 11508
rect 23660 11396 23716 11452
rect 27580 11396 27636 11452
rect 13010 11340 13020 11396
rect 13076 11340 13916 11396
rect 13972 11340 13982 11396
rect 14578 11340 14588 11396
rect 14644 11340 16044 11396
rect 16100 11340 16110 11396
rect 16258 11340 16268 11396
rect 16324 11340 17724 11396
rect 17780 11340 17790 11396
rect 18274 11340 18284 11396
rect 18340 11340 18620 11396
rect 18676 11340 18686 11396
rect 18946 11340 18956 11396
rect 19012 11340 21196 11396
rect 21252 11340 21262 11396
rect 21410 11340 21420 11396
rect 21476 11340 23716 11396
rect 23772 11340 25900 11396
rect 25956 11340 25966 11396
rect 26450 11340 26460 11396
rect 26516 11340 27636 11396
rect 30146 11340 30156 11396
rect 30212 11340 41804 11396
rect 41860 11340 41870 11396
rect 45602 11340 45612 11396
rect 45668 11340 48860 11396
rect 48916 11340 48926 11396
rect 0 11284 112 11312
rect 23772 11284 23828 11340
rect 52640 11284 52752 11312
rect 0 11228 12012 11284
rect 12068 11228 12078 11284
rect 13794 11228 13804 11284
rect 13860 11228 18060 11284
rect 18116 11228 18126 11284
rect 18386 11228 18396 11284
rect 18452 11228 22764 11284
rect 22820 11228 22830 11284
rect 22978 11228 22988 11284
rect 23044 11228 23828 11284
rect 24658 11228 24668 11284
rect 24724 11228 26348 11284
rect 26404 11228 26414 11284
rect 27346 11228 27356 11284
rect 27412 11228 29820 11284
rect 29876 11228 29886 11284
rect 30930 11228 30940 11284
rect 30996 11228 35644 11284
rect 35700 11228 35710 11284
rect 37538 11228 37548 11284
rect 37604 11228 43708 11284
rect 49858 11228 49868 11284
rect 49924 11228 52752 11284
rect 0 11200 112 11228
rect 43652 11172 43708 11228
rect 52640 11200 52752 11228
rect 11890 11116 11900 11172
rect 11956 11116 16548 11172
rect 16706 11116 16716 11172
rect 16772 11116 27356 11172
rect 27412 11116 27422 11172
rect 28242 11116 28252 11172
rect 28308 11116 29708 11172
rect 29764 11116 29774 11172
rect 29922 11116 29932 11172
rect 29988 11116 38780 11172
rect 38836 11116 38846 11172
rect 43652 11116 45276 11172
rect 45332 11116 45342 11172
rect 16492 11060 16548 11116
rect 14130 11004 14140 11060
rect 14196 11004 16324 11060
rect 16492 11004 22876 11060
rect 22932 11004 22942 11060
rect 23090 11004 23100 11060
rect 23156 11004 23660 11060
rect 23716 11004 23726 11060
rect 24210 11004 24220 11060
rect 24276 11004 24892 11060
rect 24948 11004 24958 11060
rect 25778 11004 25788 11060
rect 25844 11004 35308 11060
rect 35364 11004 35374 11060
rect 38612 11004 43708 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 5058 10892 5068 10948
rect 5124 10892 13580 10948
rect 13636 10892 13646 10948
rect 14242 10892 14252 10948
rect 14308 10892 16044 10948
rect 16100 10892 16110 10948
rect 0 10836 112 10864
rect 16268 10836 16324 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 38612 10948 38668 11004
rect 16482 10892 16492 10948
rect 16548 10892 18844 10948
rect 18900 10892 18910 10948
rect 19058 10892 19068 10948
rect 19124 10892 23716 10948
rect 24322 10892 24332 10948
rect 24388 10892 26796 10948
rect 26852 10892 26862 10948
rect 27010 10892 27020 10948
rect 27076 10892 31500 10948
rect 31556 10892 31566 10948
rect 34178 10892 34188 10948
rect 34244 10892 38668 10948
rect 23660 10836 23716 10892
rect 43652 10836 43708 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 52640 10836 52752 10864
rect 0 10780 7756 10836
rect 7812 10780 7822 10836
rect 10434 10780 10444 10836
rect 10500 10780 12572 10836
rect 12628 10780 12638 10836
rect 13468 10780 15932 10836
rect 15988 10780 15998 10836
rect 16268 10780 21644 10836
rect 21700 10780 21710 10836
rect 21858 10780 21868 10836
rect 21924 10780 22428 10836
rect 22484 10780 22494 10836
rect 22642 10780 22652 10836
rect 22708 10780 23436 10836
rect 23492 10780 23502 10836
rect 23660 10780 24220 10836
rect 24276 10780 24286 10836
rect 25330 10780 25340 10836
rect 25396 10780 28252 10836
rect 28308 10780 28318 10836
rect 28466 10780 28476 10836
rect 28532 10780 33292 10836
rect 33348 10780 33358 10836
rect 33618 10780 33628 10836
rect 33684 10780 39676 10836
rect 39732 10780 39742 10836
rect 39890 10780 39900 10836
rect 39956 10780 42476 10836
rect 42532 10780 42542 10836
rect 43652 10780 48748 10836
rect 48804 10780 48814 10836
rect 51202 10780 51212 10836
rect 51268 10780 52752 10836
rect 0 10752 112 10780
rect 13468 10724 13524 10780
rect 52640 10752 52752 10780
rect 2258 10668 2268 10724
rect 2324 10668 4956 10724
rect 5012 10668 5022 10724
rect 8978 10668 8988 10724
rect 9044 10668 13524 10724
rect 13682 10668 13692 10724
rect 13748 10668 16492 10724
rect 16548 10668 16558 10724
rect 16930 10668 16940 10724
rect 16996 10668 47852 10724
rect 47908 10668 47918 10724
rect 1138 10556 1148 10612
rect 1204 10556 15932 10612
rect 15988 10556 15998 10612
rect 16146 10556 16156 10612
rect 16212 10556 26684 10612
rect 26740 10556 26750 10612
rect 26898 10556 26908 10612
rect 26964 10556 29932 10612
rect 29988 10556 29998 10612
rect 31826 10556 31836 10612
rect 31892 10556 42028 10612
rect 42084 10556 42094 10612
rect 802 10444 812 10500
rect 868 10444 6188 10500
rect 6244 10444 6254 10500
rect 6850 10444 6860 10500
rect 6916 10444 17276 10500
rect 17332 10444 17342 10500
rect 18274 10444 18284 10500
rect 18340 10444 21308 10500
rect 21364 10444 21374 10500
rect 21522 10444 21532 10500
rect 21588 10444 23100 10500
rect 23156 10444 23166 10500
rect 23426 10444 23436 10500
rect 23492 10444 25564 10500
rect 25620 10444 25630 10500
rect 25890 10444 25900 10500
rect 25956 10444 32508 10500
rect 32564 10444 32574 10500
rect 33506 10444 33516 10500
rect 33572 10444 40908 10500
rect 40964 10444 40974 10500
rect 41132 10444 47516 10500
rect 47572 10444 47740 10500
rect 47796 10444 47806 10500
rect 47964 10444 50204 10500
rect 50260 10444 50270 10500
rect 0 10388 112 10416
rect 41132 10388 41188 10444
rect 47964 10388 48020 10444
rect 52640 10388 52752 10416
rect 0 10332 1652 10388
rect 2706 10332 2716 10388
rect 2772 10332 8092 10388
rect 8148 10332 8158 10388
rect 9510 10332 9548 10388
rect 9604 10332 9614 10388
rect 10322 10332 10332 10388
rect 10388 10332 14028 10388
rect 14084 10332 14094 10388
rect 15362 10332 15372 10388
rect 15428 10332 27804 10388
rect 27860 10332 27870 10388
rect 28252 10332 30940 10388
rect 30996 10332 31006 10388
rect 31154 10332 31164 10388
rect 31220 10332 33404 10388
rect 33460 10332 33470 10388
rect 35522 10332 35532 10388
rect 35588 10332 37772 10388
rect 37828 10332 37838 10388
rect 39218 10332 39228 10388
rect 39284 10332 41188 10388
rect 41458 10332 41468 10388
rect 41524 10332 48020 10388
rect 49634 10332 49644 10388
rect 49700 10332 52752 10388
rect 0 10304 112 10332
rect 1596 10052 1652 10332
rect 28252 10276 28308 10332
rect 52640 10304 52752 10332
rect 8754 10220 8764 10276
rect 8820 10220 15484 10276
rect 15540 10220 15550 10276
rect 15922 10220 15932 10276
rect 15988 10220 23436 10276
rect 23492 10220 23502 10276
rect 23650 10220 23660 10276
rect 23716 10220 24108 10276
rect 24164 10220 24174 10276
rect 24994 10220 25004 10276
rect 25060 10220 26404 10276
rect 26674 10220 26684 10276
rect 26740 10220 28308 10276
rect 28466 10220 28476 10276
rect 28532 10220 37548 10276
rect 37604 10220 37614 10276
rect 39106 10220 39116 10276
rect 39172 10220 41356 10276
rect 41412 10220 41422 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 26348 10164 26404 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 8194 10108 8204 10164
rect 8260 10108 10948 10164
rect 11778 10108 11788 10164
rect 11844 10108 14364 10164
rect 14420 10108 14430 10164
rect 14914 10108 14924 10164
rect 14980 10108 17500 10164
rect 17556 10108 17566 10164
rect 17714 10108 17724 10164
rect 17780 10108 19068 10164
rect 19124 10108 19134 10164
rect 20038 10108 20076 10164
rect 20132 10108 20142 10164
rect 20290 10108 20300 10164
rect 20356 10108 22540 10164
rect 22596 10108 22606 10164
rect 22754 10108 22764 10164
rect 22820 10108 24332 10164
rect 24388 10108 24398 10164
rect 26114 10108 26124 10164
rect 26180 10108 26190 10164
rect 26348 10108 27804 10164
rect 27860 10108 27870 10164
rect 28914 10108 28924 10164
rect 28980 10108 34188 10164
rect 34244 10108 34636 10164
rect 34692 10108 34702 10164
rect 35308 10108 37212 10164
rect 37268 10108 37278 10164
rect 38658 10108 38668 10164
rect 38724 10108 41244 10164
rect 41300 10108 41310 10164
rect 48290 10108 48300 10164
rect 48356 10108 50540 10164
rect 50596 10108 50606 10164
rect 1596 9996 10444 10052
rect 10500 9996 10668 10052
rect 10724 9996 10734 10052
rect 0 9940 112 9968
rect 10892 9940 10948 10108
rect 26124 10052 26180 10108
rect 35308 10052 35364 10108
rect 12450 9996 12460 10052
rect 12516 9996 13580 10052
rect 13636 9996 13646 10052
rect 13804 9996 26348 10052
rect 26404 9996 26414 10052
rect 26562 9996 26572 10052
rect 26628 9996 30604 10052
rect 30660 9996 30670 10052
rect 31042 9996 31052 10052
rect 31108 9996 33068 10052
rect 33124 9996 33134 10052
rect 33618 9996 33628 10052
rect 33684 9996 35364 10052
rect 35522 9996 35532 10052
rect 35588 9996 38780 10052
rect 38836 9996 38846 10052
rect 39554 9996 39564 10052
rect 39620 9996 40796 10052
rect 40852 9996 40862 10052
rect 41010 9996 41020 10052
rect 41076 9996 47068 10052
rect 47124 9996 47134 10052
rect 13804 9940 13860 9996
rect 52640 9940 52752 9968
rect 0 9884 1260 9940
rect 1316 9884 1326 9940
rect 6066 9884 6076 9940
rect 6132 9884 7420 9940
rect 7476 9884 7486 9940
rect 7634 9884 7644 9940
rect 7700 9884 8652 9940
rect 8708 9884 8718 9940
rect 10892 9884 13860 9940
rect 14018 9884 14028 9940
rect 14084 9884 15260 9940
rect 15316 9884 15326 9940
rect 16482 9884 16492 9940
rect 16548 9884 18844 9940
rect 18900 9884 18910 9940
rect 19058 9884 19068 9940
rect 19124 9884 21252 9940
rect 21634 9884 21644 9940
rect 21700 9884 23044 9940
rect 23202 9884 23212 9940
rect 23268 9884 24556 9940
rect 24612 9884 24622 9940
rect 24882 9884 24892 9940
rect 24948 9884 28812 9940
rect 28868 9884 28878 9940
rect 29250 9884 29260 9940
rect 29316 9884 30716 9940
rect 30772 9884 30782 9940
rect 30930 9884 30940 9940
rect 30996 9884 34524 9940
rect 34580 9884 34590 9940
rect 37874 9884 37884 9940
rect 37940 9884 41916 9940
rect 41972 9884 41982 9940
rect 42130 9884 42140 9940
rect 42196 9884 50428 9940
rect 50484 9884 50494 9940
rect 51426 9884 51436 9940
rect 51492 9884 52752 9940
rect 0 9856 112 9884
rect 21196 9828 21252 9884
rect 22988 9828 23044 9884
rect 52640 9856 52752 9884
rect 14578 9772 14588 9828
rect 14644 9772 19684 9828
rect 19842 9772 19852 9828
rect 19908 9772 20972 9828
rect 21028 9772 21038 9828
rect 21196 9772 22652 9828
rect 22708 9772 22718 9828
rect 22988 9772 26348 9828
rect 26404 9772 26414 9828
rect 26786 9772 26796 9828
rect 26852 9772 27132 9828
rect 27188 9772 28140 9828
rect 28196 9772 28206 9828
rect 30034 9772 30044 9828
rect 30100 9772 31500 9828
rect 31556 9772 31566 9828
rect 31714 9772 31724 9828
rect 31780 9772 38332 9828
rect 38388 9772 38398 9828
rect 38612 9772 40348 9828
rect 40404 9772 40414 9828
rect 44930 9772 44940 9828
rect 44996 9772 48972 9828
rect 49028 9772 49038 9828
rect 19628 9716 19684 9772
rect 38612 9716 38668 9772
rect 3266 9660 3276 9716
rect 3332 9660 8764 9716
rect 8820 9660 8830 9716
rect 8978 9660 8988 9716
rect 9044 9660 18956 9716
rect 19012 9660 19022 9716
rect 19628 9660 21868 9716
rect 21924 9660 21934 9716
rect 22194 9660 22204 9716
rect 22260 9660 24948 9716
rect 25106 9660 25116 9716
rect 25172 9660 25452 9716
rect 25508 9660 32732 9716
rect 32788 9660 32798 9716
rect 33730 9660 33740 9716
rect 33796 9660 38668 9716
rect 38770 9660 38780 9716
rect 38836 9660 42252 9716
rect 42308 9660 42318 9716
rect 43596 9660 43932 9716
rect 43988 9660 43998 9716
rect 44482 9660 44492 9716
rect 44548 9660 49084 9716
rect 49140 9660 49150 9716
rect 49858 9660 49868 9716
rect 49924 9660 50876 9716
rect 50932 9660 50942 9716
rect 24892 9604 24948 9660
rect 43596 9604 43652 9660
rect 3332 9548 8316 9604
rect 8372 9548 8382 9604
rect 10098 9548 10108 9604
rect 10164 9548 16716 9604
rect 16772 9548 16782 9604
rect 17154 9548 17164 9604
rect 17220 9548 24276 9604
rect 24892 9548 26124 9604
rect 26180 9548 26190 9604
rect 26562 9548 26572 9604
rect 26628 9548 29148 9604
rect 29204 9548 29214 9604
rect 29362 9548 29372 9604
rect 29428 9548 38668 9604
rect 38724 9548 38734 9604
rect 39778 9548 39788 9604
rect 39844 9548 40908 9604
rect 40964 9548 40974 9604
rect 41794 9548 41804 9604
rect 41860 9548 43596 9604
rect 43652 9548 43662 9604
rect 0 9492 112 9520
rect 3332 9492 3388 9548
rect 24220 9492 24276 9548
rect 52640 9492 52752 9520
rect 0 9436 3388 9492
rect 4946 9436 4956 9492
rect 5012 9436 6636 9492
rect 6692 9436 6702 9492
rect 12226 9436 12236 9492
rect 12292 9436 21532 9492
rect 21588 9436 21598 9492
rect 21756 9436 22988 9492
rect 23044 9436 23054 9492
rect 24220 9436 30156 9492
rect 30212 9436 30222 9492
rect 32498 9436 32508 9492
rect 32564 9436 40012 9492
rect 40068 9436 40078 9492
rect 50978 9436 50988 9492
rect 51044 9436 52752 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 21756 9380 21812 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 52640 9408 52752 9436
rect 6962 9324 6972 9380
rect 7028 9324 18284 9380
rect 18340 9324 18350 9380
rect 18498 9324 18508 9380
rect 18564 9324 21812 9380
rect 21868 9324 23212 9380
rect 23268 9324 23278 9380
rect 24322 9324 24332 9380
rect 24388 9324 25004 9380
rect 25060 9324 25070 9380
rect 25218 9324 25228 9380
rect 25284 9324 30380 9380
rect 30436 9324 30446 9380
rect 31490 9324 31500 9380
rect 31556 9324 34076 9380
rect 34132 9324 34142 9380
rect 36642 9324 36652 9380
rect 36708 9324 42140 9380
rect 42196 9324 42206 9380
rect 21868 9268 21924 9324
rect 1698 9212 1708 9268
rect 1764 9212 7980 9268
rect 8036 9212 8046 9268
rect 8866 9212 8876 9268
rect 8932 9212 13804 9268
rect 13860 9212 13870 9268
rect 14802 9212 14812 9268
rect 14868 9212 15708 9268
rect 15764 9212 15774 9268
rect 15922 9212 15932 9268
rect 15988 9212 17276 9268
rect 17332 9212 17342 9268
rect 17714 9212 17724 9268
rect 17780 9212 21924 9268
rect 22082 9212 22092 9268
rect 22148 9212 36988 9268
rect 37044 9212 37054 9268
rect 37202 9212 37212 9268
rect 37268 9212 43596 9268
rect 43652 9212 43662 9268
rect 49634 9212 49644 9268
rect 49700 9212 51100 9268
rect 51156 9212 51166 9268
rect 8530 9100 8540 9156
rect 8596 9100 11900 9156
rect 11956 9100 11966 9156
rect 12114 9100 12124 9156
rect 12180 9100 15148 9156
rect 15204 9100 15214 9156
rect 15474 9100 15484 9156
rect 15540 9100 18732 9156
rect 18788 9100 18798 9156
rect 19394 9100 19404 9156
rect 19460 9100 25340 9156
rect 25396 9100 25406 9156
rect 25778 9100 25788 9156
rect 25844 9100 33852 9156
rect 33908 9100 33918 9156
rect 36306 9100 36316 9156
rect 36372 9100 38220 9156
rect 38276 9100 38556 9156
rect 38612 9100 38622 9156
rect 42354 9100 42364 9156
rect 42420 9100 45164 9156
rect 45220 9100 45230 9156
rect 0 9044 112 9072
rect 52640 9044 52752 9072
rect 0 8988 8204 9044
rect 8260 8988 8270 9044
rect 9314 8988 9324 9044
rect 9380 8988 17052 9044
rect 17108 8988 17118 9044
rect 17266 8988 17276 9044
rect 17332 8988 19292 9044
rect 19348 8988 19358 9044
rect 19954 8988 19964 9044
rect 20020 8988 23772 9044
rect 23828 8988 24332 9044
rect 24388 8988 24398 9044
rect 24546 8988 24556 9044
rect 24612 8988 28476 9044
rect 28532 8988 28542 9044
rect 30370 8988 30380 9044
rect 30436 8988 33516 9044
rect 33572 8988 33582 9044
rect 33730 8988 33740 9044
rect 33796 8988 38668 9044
rect 38724 8988 38734 9044
rect 39116 8988 48076 9044
rect 48132 8988 48142 9044
rect 51426 8988 51436 9044
rect 51492 8988 52752 9044
rect 0 8960 112 8988
rect 12226 8876 12236 8932
rect 12292 8876 22204 8932
rect 22260 8876 22270 8932
rect 22418 8876 22428 8932
rect 22484 8876 23100 8932
rect 23156 8876 23166 8932
rect 23986 8876 23996 8932
rect 24052 8876 25228 8932
rect 25284 8876 25294 8932
rect 25442 8876 25452 8932
rect 25508 8876 25788 8932
rect 25844 8876 25854 8932
rect 26012 8876 26908 8932
rect 26964 8876 26974 8932
rect 27122 8876 27132 8932
rect 27188 8876 31052 8932
rect 31108 8876 31118 8932
rect 31602 8876 31612 8932
rect 31668 8876 37212 8932
rect 37268 8876 37278 8932
rect 26012 8820 26068 8876
rect 39116 8820 39172 8988
rect 52640 8960 52752 8988
rect 40450 8876 40460 8932
rect 40516 8876 44492 8932
rect 44548 8876 44558 8932
rect 48290 8876 48300 8932
rect 48356 8876 50316 8932
rect 50372 8876 50382 8932
rect 8082 8764 8092 8820
rect 8148 8764 16828 8820
rect 16884 8764 16894 8820
rect 17042 8764 17052 8820
rect 17108 8764 19964 8820
rect 20020 8764 20030 8820
rect 20178 8764 20188 8820
rect 20244 8764 21868 8820
rect 21924 8764 21934 8820
rect 22082 8764 22092 8820
rect 22148 8764 24948 8820
rect 25554 8764 25564 8820
rect 25620 8764 26068 8820
rect 26562 8764 26572 8820
rect 26628 8764 30940 8820
rect 30996 8764 31006 8820
rect 32498 8764 32508 8820
rect 32564 8764 33292 8820
rect 33348 8764 33358 8820
rect 33506 8764 33516 8820
rect 33572 8764 39172 8820
rect 39554 8764 39564 8820
rect 39620 8764 48748 8820
rect 48804 8764 48814 8820
rect 24892 8708 24948 8764
rect 11666 8652 11676 8708
rect 11732 8652 20076 8708
rect 20132 8652 20142 8708
rect 20402 8652 20412 8708
rect 20468 8652 23996 8708
rect 24052 8652 24062 8708
rect 24892 8652 29596 8708
rect 29652 8652 29662 8708
rect 29820 8652 33964 8708
rect 34020 8652 34030 8708
rect 34850 8652 34860 8708
rect 34916 8652 42140 8708
rect 42196 8652 42206 8708
rect 47954 8652 47964 8708
rect 48020 8652 50204 8708
rect 50260 8652 50270 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 0 8540 4284 8596
rect 4340 8540 4350 8596
rect 5730 8540 5740 8596
rect 5796 8540 17276 8596
rect 17332 8540 17342 8596
rect 17490 8540 17500 8596
rect 17556 8540 20972 8596
rect 21028 8540 21038 8596
rect 21858 8540 21868 8596
rect 21924 8540 22876 8596
rect 22932 8540 22942 8596
rect 23090 8540 23100 8596
rect 23156 8540 24332 8596
rect 24388 8540 24398 8596
rect 26898 8540 26908 8596
rect 26964 8540 28588 8596
rect 28644 8540 28654 8596
rect 0 8512 112 8540
rect 29820 8484 29876 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 52640 8596 52752 8624
rect 7634 8428 7644 8484
rect 7700 8428 12124 8484
rect 12180 8428 12190 8484
rect 15092 8428 29876 8484
rect 29932 8540 33180 8596
rect 33236 8540 33246 8596
rect 33394 8540 33404 8596
rect 33460 8540 34972 8596
rect 35028 8540 35038 8596
rect 35746 8540 35756 8596
rect 35812 8540 38444 8596
rect 38500 8540 38510 8596
rect 38658 8540 38668 8596
rect 38724 8540 40236 8596
rect 40292 8540 40302 8596
rect 50978 8540 50988 8596
rect 51044 8540 52752 8596
rect 15092 8372 15148 8428
rect 29932 8372 29988 8540
rect 52640 8512 52752 8540
rect 32722 8428 32732 8484
rect 32788 8428 35532 8484
rect 35588 8428 35598 8484
rect 36754 8428 36764 8484
rect 36820 8428 45388 8484
rect 45444 8428 45454 8484
rect 8306 8316 8316 8372
rect 8372 8316 11676 8372
rect 11732 8316 11742 8372
rect 11890 8316 11900 8372
rect 11956 8316 15148 8372
rect 15250 8316 15260 8372
rect 15316 8316 15820 8372
rect 15876 8316 15886 8372
rect 16594 8316 16604 8372
rect 16660 8316 17724 8372
rect 17780 8316 17790 8372
rect 20066 8316 20076 8372
rect 20132 8316 20972 8372
rect 21028 8316 21038 8372
rect 21186 8316 21196 8372
rect 21252 8316 29988 8372
rect 32732 8316 36652 8372
rect 36708 8316 36718 8372
rect 41346 8316 41356 8372
rect 41412 8316 49196 8372
rect 49252 8316 49262 8372
rect 32732 8260 32788 8316
rect 9874 8204 9884 8260
rect 9940 8204 10220 8260
rect 10276 8204 21028 8260
rect 21522 8204 21532 8260
rect 21588 8204 22092 8260
rect 22148 8204 22158 8260
rect 22418 8204 22428 8260
rect 22484 8204 22764 8260
rect 22820 8204 22830 8260
rect 23202 8204 23212 8260
rect 23268 8204 25228 8260
rect 25284 8204 25294 8260
rect 25442 8204 25452 8260
rect 25508 8204 25676 8260
rect 25732 8204 25742 8260
rect 26674 8204 26684 8260
rect 26740 8204 32788 8260
rect 35298 8204 35308 8260
rect 35364 8204 50428 8260
rect 50484 8204 50494 8260
rect 0 8148 112 8176
rect 20972 8148 21028 8204
rect 52640 8148 52752 8176
rect 0 8092 5964 8148
rect 6020 8092 6030 8148
rect 9762 8092 9772 8148
rect 9828 8092 11900 8148
rect 11956 8092 11966 8148
rect 14018 8092 14028 8148
rect 14084 8092 16604 8148
rect 16660 8092 16670 8148
rect 16818 8092 16828 8148
rect 16884 8092 20804 8148
rect 20972 8092 28700 8148
rect 28756 8092 28766 8148
rect 30146 8092 30156 8148
rect 30212 8092 31164 8148
rect 31220 8092 31230 8148
rect 31826 8092 31836 8148
rect 31892 8092 32396 8148
rect 32452 8092 32462 8148
rect 34066 8092 34076 8148
rect 34132 8092 40460 8148
rect 40516 8092 40526 8148
rect 48178 8092 48188 8148
rect 48244 8092 49532 8148
rect 49588 8092 49598 8148
rect 50866 8092 50876 8148
rect 50932 8092 52752 8148
rect 0 8064 112 8092
rect 20748 8036 20804 8092
rect 52640 8064 52752 8092
rect 8642 7980 8652 8036
rect 8708 7980 10556 8036
rect 10612 7980 10622 8036
rect 13010 7980 13020 8036
rect 13076 7980 20188 8036
rect 20244 7980 20254 8036
rect 20748 7980 21532 8036
rect 21588 7980 21598 8036
rect 21830 7980 21868 8036
rect 21924 7980 21934 8036
rect 22194 7980 22204 8036
rect 22260 7980 24668 8036
rect 24724 7980 24734 8036
rect 24892 7980 29708 8036
rect 29764 7980 29774 8036
rect 32946 7980 32956 8036
rect 33012 7980 46172 8036
rect 46228 7980 46238 8036
rect 24892 7924 24948 7980
rect 9202 7868 9212 7924
rect 9268 7868 21196 7924
rect 21252 7868 21262 7924
rect 22418 7868 22428 7924
rect 22484 7868 23436 7924
rect 23492 7868 23502 7924
rect 24210 7868 24220 7924
rect 24276 7868 24948 7924
rect 25330 7868 25340 7924
rect 25396 7868 33516 7924
rect 33572 7868 33582 7924
rect 33954 7868 33964 7924
rect 34020 7868 41804 7924
rect 41860 7868 41870 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 5506 7756 5516 7812
rect 5572 7756 9996 7812
rect 10052 7756 10062 7812
rect 15138 7756 15148 7812
rect 15204 7756 18396 7812
rect 18452 7756 18462 7812
rect 20066 7756 20076 7812
rect 20132 7756 23604 7812
rect 24210 7756 24220 7812
rect 24276 7756 25452 7812
rect 25508 7756 25518 7812
rect 25778 7756 25788 7812
rect 25844 7756 33740 7812
rect 33796 7756 33806 7812
rect 34290 7756 34300 7812
rect 34356 7756 37100 7812
rect 37156 7756 37166 7812
rect 0 7700 112 7728
rect 23548 7700 23604 7756
rect 52640 7700 52752 7728
rect 0 7644 1596 7700
rect 1652 7644 1662 7700
rect 11554 7644 11564 7700
rect 11620 7644 15148 7700
rect 15204 7644 15214 7700
rect 15362 7644 15372 7700
rect 15428 7644 23324 7700
rect 23380 7644 23390 7700
rect 23548 7644 31948 7700
rect 32004 7644 32014 7700
rect 32274 7644 32284 7700
rect 32340 7644 33852 7700
rect 33908 7644 33918 7700
rect 51426 7644 51436 7700
rect 51492 7644 52752 7700
rect 0 7616 112 7644
rect 52640 7616 52752 7644
rect 9202 7532 9212 7588
rect 9268 7532 16828 7588
rect 16884 7532 16894 7588
rect 17388 7532 19404 7588
rect 19460 7532 19470 7588
rect 19618 7532 19628 7588
rect 19684 7532 21308 7588
rect 21364 7532 21374 7588
rect 21858 7532 21868 7588
rect 21924 7532 22092 7588
rect 22148 7532 22158 7588
rect 22306 7532 22316 7588
rect 22372 7532 22876 7588
rect 22932 7532 22942 7588
rect 24098 7532 24108 7588
rect 24164 7532 25676 7588
rect 25732 7532 25742 7588
rect 26562 7532 26572 7588
rect 26628 7532 28924 7588
rect 28980 7532 28990 7588
rect 29138 7532 29148 7588
rect 29204 7532 32956 7588
rect 33012 7532 33022 7588
rect 40898 7532 40908 7588
rect 40964 7532 49980 7588
rect 50036 7532 50046 7588
rect 17388 7476 17444 7532
rect 4274 7420 4284 7476
rect 4340 7420 13804 7476
rect 13860 7420 13870 7476
rect 14018 7420 14028 7476
rect 14084 7420 17444 7476
rect 17602 7420 17612 7476
rect 17668 7420 19852 7476
rect 19908 7420 19918 7476
rect 20066 7420 20076 7476
rect 20132 7420 20412 7476
rect 20468 7420 20478 7476
rect 20626 7420 20636 7476
rect 20692 7420 29260 7476
rect 29316 7420 29326 7476
rect 29922 7420 29932 7476
rect 29988 7420 38780 7476
rect 38836 7420 38846 7476
rect 40226 7420 40236 7476
rect 40292 7420 48300 7476
rect 48356 7420 48366 7476
rect 3602 7308 3612 7364
rect 3668 7308 13356 7364
rect 13412 7308 13422 7364
rect 13794 7308 13804 7364
rect 13860 7308 15372 7364
rect 15428 7308 15438 7364
rect 15586 7308 15596 7364
rect 15652 7308 18060 7364
rect 18116 7308 18126 7364
rect 18284 7308 28476 7364
rect 28532 7308 28542 7364
rect 28914 7308 28924 7364
rect 28980 7308 48748 7364
rect 48804 7308 48814 7364
rect 0 7252 112 7280
rect 0 7196 2716 7252
rect 2772 7196 2782 7252
rect 6290 7196 6300 7252
rect 6356 7196 8092 7252
rect 8148 7196 8158 7252
rect 13234 7196 13244 7252
rect 13300 7196 15932 7252
rect 15988 7196 15998 7252
rect 16146 7196 16156 7252
rect 16212 7196 17052 7252
rect 17108 7196 17118 7252
rect 0 7168 112 7196
rect 7522 7084 7532 7140
rect 7588 7084 11676 7140
rect 11732 7084 11742 7140
rect 14578 7084 14588 7140
rect 14644 7084 17948 7140
rect 18004 7084 18014 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 10770 6972 10780 7028
rect 10836 6972 15484 7028
rect 15540 6972 15550 7028
rect 15698 6972 15708 7028
rect 15764 6972 17164 7028
rect 17220 6972 17230 7028
rect 18284 6916 18340 7308
rect 52640 7252 52752 7280
rect 18498 7196 18508 7252
rect 18564 7196 26908 7252
rect 27010 7196 27020 7252
rect 27076 7196 28140 7252
rect 28196 7196 28206 7252
rect 28364 7196 31724 7252
rect 31780 7196 31790 7252
rect 35298 7196 35308 7252
rect 35364 7196 39228 7252
rect 39284 7196 39294 7252
rect 43652 7196 48188 7252
rect 48244 7196 48254 7252
rect 51426 7196 51436 7252
rect 51492 7196 52752 7252
rect 26852 7140 26908 7196
rect 28364 7140 28420 7196
rect 43652 7140 43708 7196
rect 52640 7168 52752 7196
rect 18946 7084 18956 7140
rect 19012 7084 19292 7140
rect 19348 7084 21868 7140
rect 21924 7084 21934 7140
rect 22754 7084 22764 7140
rect 22820 7084 24108 7140
rect 24164 7084 24174 7140
rect 24994 7084 25004 7140
rect 25060 7084 26684 7140
rect 26740 7084 26750 7140
rect 26852 7084 28420 7140
rect 29474 7084 29484 7140
rect 29540 7084 43708 7140
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 18498 6972 18508 7028
rect 18564 6972 19852 7028
rect 19908 6972 19918 7028
rect 20066 6972 20076 7028
rect 20132 6972 24220 7028
rect 24276 6972 24286 7028
rect 24882 6972 24892 7028
rect 24948 6972 28252 7028
rect 28308 6972 28318 7028
rect 28466 6972 28476 7028
rect 28532 6972 30828 7028
rect 30884 6972 30894 7028
rect 31052 6972 38332 7028
rect 38388 6972 38398 7028
rect 38546 6972 38556 7028
rect 31052 6916 31108 6972
rect 38612 6916 38668 7028
rect 242 6860 252 6916
rect 308 6860 8316 6916
rect 8372 6860 8382 6916
rect 12562 6860 12572 6916
rect 12628 6860 18340 6916
rect 18722 6860 18732 6916
rect 18788 6860 19180 6916
rect 19236 6860 19246 6916
rect 19394 6860 19404 6916
rect 19460 6860 22988 6916
rect 23044 6860 23054 6916
rect 23426 6860 23436 6916
rect 23492 6860 28364 6916
rect 28420 6860 28430 6916
rect 29810 6860 29820 6916
rect 29876 6860 31108 6916
rect 31612 6860 31948 6916
rect 32004 6860 32014 6916
rect 33730 6860 33740 6916
rect 33796 6860 38444 6916
rect 38500 6860 38510 6916
rect 38612 6860 43484 6916
rect 43540 6860 43550 6916
rect 48962 6860 48972 6916
rect 49028 6860 50652 6916
rect 50708 6860 50718 6916
rect 0 6804 112 6832
rect 31612 6804 31668 6860
rect 52640 6804 52752 6832
rect 0 6748 1148 6804
rect 1204 6748 1214 6804
rect 3266 6748 3276 6804
rect 3332 6748 9212 6804
rect 9268 6748 9278 6804
rect 11218 6748 11228 6804
rect 11284 6748 13188 6804
rect 13794 6748 13804 6804
rect 13860 6748 19964 6804
rect 20020 6748 20030 6804
rect 20132 6748 22820 6804
rect 23202 6748 23212 6804
rect 23268 6748 25004 6804
rect 25060 6748 25070 6804
rect 25228 6748 29148 6804
rect 29204 6748 29214 6804
rect 29586 6748 29596 6804
rect 29652 6748 31668 6804
rect 31836 6748 33628 6804
rect 33684 6748 33694 6804
rect 36988 6748 39900 6804
rect 39956 6748 39966 6804
rect 42130 6748 42140 6804
rect 42196 6748 44268 6804
rect 44324 6748 44334 6804
rect 49634 6748 49644 6804
rect 49700 6748 52752 6804
rect 0 6720 112 6748
rect 13132 6692 13188 6748
rect 20132 6692 20188 6748
rect 22764 6692 22820 6748
rect 25228 6692 25284 6748
rect 31836 6692 31892 6748
rect 36988 6692 37044 6748
rect 52640 6720 52752 6748
rect 1586 6636 1596 6692
rect 1652 6636 3388 6692
rect 9538 6636 9548 6692
rect 9604 6636 9884 6692
rect 9940 6636 11564 6692
rect 11620 6636 11630 6692
rect 13132 6636 13692 6692
rect 13748 6636 13758 6692
rect 13906 6636 13916 6692
rect 13972 6636 18732 6692
rect 18788 6636 18798 6692
rect 18956 6636 20188 6692
rect 20962 6636 20972 6692
rect 21028 6636 22092 6692
rect 22148 6636 22158 6692
rect 22754 6636 22764 6692
rect 22820 6636 22830 6692
rect 22978 6636 22988 6692
rect 23044 6636 25284 6692
rect 25442 6636 25452 6692
rect 25508 6636 29708 6692
rect 29764 6636 29774 6692
rect 29922 6636 29932 6692
rect 29988 6636 31892 6692
rect 35522 6636 35532 6692
rect 35588 6636 37044 6692
rect 38098 6636 38108 6692
rect 38164 6636 43708 6692
rect 48066 6636 48076 6692
rect 48132 6636 50204 6692
rect 50260 6636 50270 6692
rect 3332 6580 3388 6636
rect 18956 6580 19012 6636
rect 43652 6580 43708 6636
rect 3332 6524 14476 6580
rect 14532 6524 14542 6580
rect 14690 6524 14700 6580
rect 14756 6524 15708 6580
rect 15764 6524 15774 6580
rect 15922 6524 15932 6580
rect 15988 6524 19012 6580
rect 20178 6524 20188 6580
rect 20244 6524 21980 6580
rect 22036 6524 22046 6580
rect 22204 6524 38444 6580
rect 38500 6524 38510 6580
rect 38602 6524 38612 6580
rect 38668 6524 39116 6580
rect 39172 6524 39182 6580
rect 40562 6524 40572 6580
rect 40628 6524 43148 6580
rect 43204 6524 43214 6580
rect 43652 6524 48524 6580
rect 48580 6524 48590 6580
rect 22204 6468 22260 6524
rect 11778 6412 11788 6468
rect 11844 6412 16716 6468
rect 16772 6412 16782 6468
rect 16930 6412 16940 6468
rect 16996 6412 17724 6468
rect 17780 6412 17790 6468
rect 18386 6412 18396 6468
rect 18452 6412 22260 6468
rect 23314 6412 23324 6468
rect 23380 6412 23660 6468
rect 23716 6412 24276 6468
rect 24434 6412 24444 6468
rect 24500 6412 25452 6468
rect 25508 6412 25518 6468
rect 27794 6412 27804 6468
rect 27860 6412 31724 6468
rect 31780 6412 31790 6468
rect 31938 6412 31948 6468
rect 32004 6412 33012 6468
rect 35634 6412 35644 6468
rect 35700 6412 44380 6468
rect 44436 6412 44446 6468
rect 0 6356 112 6384
rect 24220 6356 24276 6412
rect 32956 6356 33012 6412
rect 52640 6356 52752 6384
rect 0 6300 3276 6356
rect 3332 6300 3342 6356
rect 13794 6300 13804 6356
rect 13860 6300 16604 6356
rect 16660 6300 16670 6356
rect 17042 6300 17052 6356
rect 17108 6300 22316 6356
rect 22372 6300 22382 6356
rect 24220 6300 27356 6356
rect 27412 6300 27422 6356
rect 29698 6300 29708 6356
rect 29764 6300 32732 6356
rect 32788 6300 32798 6356
rect 32956 6300 35980 6356
rect 36036 6300 36046 6356
rect 51202 6300 51212 6356
rect 51268 6300 52752 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 52640 6272 52752 6300
rect 9510 6188 9548 6244
rect 9604 6188 9614 6244
rect 10098 6188 10108 6244
rect 10164 6188 15484 6244
rect 15540 6188 15550 6244
rect 16034 6188 16044 6244
rect 16100 6188 23660 6244
rect 23716 6188 23726 6244
rect 24210 6188 24220 6244
rect 24276 6188 25004 6244
rect 25060 6188 25070 6244
rect 25218 6188 25228 6244
rect 25284 6188 27580 6244
rect 27636 6188 27646 6244
rect 28130 6188 28140 6244
rect 28196 6188 29932 6244
rect 29988 6188 29998 6244
rect 30146 6188 30156 6244
rect 30212 6188 41132 6244
rect 41188 6188 41198 6244
rect 47842 6188 47852 6244
rect 47908 6188 49868 6244
rect 49924 6188 49934 6244
rect 7970 6076 7980 6132
rect 8036 6076 14700 6132
rect 14756 6076 14766 6132
rect 15026 6076 15036 6132
rect 15092 6076 17500 6132
rect 17556 6076 17566 6132
rect 20962 6076 20972 6132
rect 21028 6076 28028 6132
rect 28084 6076 28094 6132
rect 30930 6076 30940 6132
rect 30996 6076 33740 6132
rect 33796 6076 33806 6132
rect 40114 6076 40124 6132
rect 40180 6076 48972 6132
rect 49028 6076 49308 6132
rect 49364 6076 49374 6132
rect 8306 5964 8316 6020
rect 8372 5964 16380 6020
rect 16436 5964 16446 6020
rect 17714 5964 17724 6020
rect 17780 5964 24220 6020
rect 24276 5964 24286 6020
rect 24546 5964 24556 6020
rect 24612 5964 26460 6020
rect 26516 5964 26526 6020
rect 27346 5964 27356 6020
rect 27412 5964 30380 6020
rect 30436 5964 30446 6020
rect 30594 5964 30604 6020
rect 30660 5964 36092 6020
rect 36148 5964 36158 6020
rect 45714 5964 45724 6020
rect 45780 5964 47740 6020
rect 47796 5964 48076 6020
rect 48132 5964 48142 6020
rect 48300 5964 50764 6020
rect 50820 5964 50830 6020
rect 0 5908 112 5936
rect 48300 5908 48356 5964
rect 52640 5908 52752 5936
rect 0 5852 6524 5908
rect 6580 5852 6590 5908
rect 6738 5852 6748 5908
rect 6804 5852 12572 5908
rect 12628 5852 12638 5908
rect 12786 5852 12796 5908
rect 12852 5852 14700 5908
rect 14756 5852 14766 5908
rect 16258 5852 16268 5908
rect 16324 5852 27020 5908
rect 27076 5852 27086 5908
rect 28242 5852 28252 5908
rect 28308 5852 35308 5908
rect 35364 5852 35374 5908
rect 35522 5852 35532 5908
rect 35588 5852 48356 5908
rect 49746 5852 49756 5908
rect 49812 5852 52752 5908
rect 0 5824 112 5852
rect 6748 5796 6804 5852
rect 52640 5824 52752 5852
rect 1810 5740 1820 5796
rect 1876 5740 5348 5796
rect 5506 5740 5516 5796
rect 5572 5740 6804 5796
rect 7746 5740 7756 5796
rect 7812 5740 13356 5796
rect 13412 5740 13422 5796
rect 14354 5740 14364 5796
rect 14420 5740 20748 5796
rect 20804 5740 20814 5796
rect 21410 5740 21420 5796
rect 21476 5740 24892 5796
rect 24948 5740 24958 5796
rect 25218 5740 25228 5796
rect 25284 5740 33516 5796
rect 33572 5740 33582 5796
rect 33842 5740 33852 5796
rect 33908 5740 37660 5796
rect 37716 5740 37726 5796
rect 5292 5572 5348 5740
rect 5954 5628 5964 5684
rect 6020 5628 8204 5684
rect 8260 5628 8270 5684
rect 11666 5628 11676 5684
rect 11732 5628 20636 5684
rect 20692 5628 20702 5684
rect 20850 5628 20860 5684
rect 20916 5628 21588 5684
rect 21746 5628 21756 5684
rect 21812 5628 27356 5684
rect 27412 5628 27422 5684
rect 27682 5628 27692 5684
rect 27748 5628 30268 5684
rect 30324 5628 30334 5684
rect 33394 5628 33404 5684
rect 33460 5628 47964 5684
rect 48020 5628 48030 5684
rect 21532 5572 21588 5628
rect 5292 5516 7532 5572
rect 7588 5516 7598 5572
rect 8082 5516 8092 5572
rect 8148 5516 15036 5572
rect 15092 5516 15102 5572
rect 15260 5516 16716 5572
rect 16772 5516 16782 5572
rect 16930 5516 16940 5572
rect 16996 5516 21308 5572
rect 21364 5516 21374 5572
rect 21532 5516 24332 5572
rect 24388 5516 24398 5572
rect 24994 5516 25004 5572
rect 25060 5516 26236 5572
rect 26292 5516 26302 5572
rect 26450 5516 26460 5572
rect 26516 5516 28924 5572
rect 28980 5516 28990 5572
rect 29698 5516 29708 5572
rect 29764 5516 33180 5572
rect 33236 5516 33246 5572
rect 35298 5516 35308 5572
rect 35364 5516 37996 5572
rect 38052 5516 38062 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 15260 5460 15316 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 52640 5460 52752 5488
rect 0 5404 3332 5460
rect 10434 5404 10444 5460
rect 10500 5404 15316 5460
rect 15586 5404 15596 5460
rect 15652 5404 17836 5460
rect 17892 5404 17902 5460
rect 18050 5404 18060 5460
rect 18116 5404 23436 5460
rect 23492 5404 23502 5460
rect 24882 5404 24892 5460
rect 24948 5404 29820 5460
rect 29876 5404 29886 5460
rect 32834 5404 32844 5460
rect 32900 5404 41020 5460
rect 41076 5404 41086 5460
rect 51202 5404 51212 5460
rect 51268 5404 52752 5460
rect 0 5376 112 5404
rect 0 5012 112 5040
rect 3276 5012 3332 5404
rect 52640 5376 52752 5404
rect 11666 5292 11676 5348
rect 11732 5292 18284 5348
rect 18340 5292 18350 5348
rect 18498 5292 18508 5348
rect 18564 5292 25116 5348
rect 25172 5292 25182 5348
rect 25330 5292 25340 5348
rect 25396 5292 45052 5348
rect 45108 5292 45118 5348
rect 5954 5180 5964 5236
rect 6020 5180 8316 5236
rect 8372 5180 8382 5236
rect 10882 5180 10892 5236
rect 10948 5180 26572 5236
rect 26628 5180 26638 5236
rect 27794 5180 27804 5236
rect 27860 5180 33236 5236
rect 33394 5180 33404 5236
rect 33460 5180 38668 5236
rect 38724 5180 38892 5236
rect 38948 5180 38958 5236
rect 39442 5180 39452 5236
rect 39508 5180 50092 5236
rect 50148 5180 50158 5236
rect 3490 5068 3500 5124
rect 3556 5068 5516 5124
rect 5572 5068 5852 5124
rect 5908 5068 5918 5124
rect 6514 5068 6524 5124
rect 6580 5068 6748 5124
rect 6804 5068 9772 5124
rect 9828 5068 9838 5124
rect 9986 5068 9996 5124
rect 10052 5068 12068 5124
rect 14802 5068 14812 5124
rect 14868 5068 15148 5124
rect 15204 5068 16940 5124
rect 16996 5068 17006 5124
rect 17826 5068 17836 5124
rect 17892 5068 18732 5124
rect 18788 5068 18798 5124
rect 18946 5068 18956 5124
rect 19012 5068 21308 5124
rect 21364 5068 21374 5124
rect 21532 5068 22204 5124
rect 22260 5068 22270 5124
rect 22428 5068 22988 5124
rect 23044 5068 23054 5124
rect 23202 5068 23212 5124
rect 23268 5068 24556 5124
rect 24612 5068 24892 5124
rect 24948 5068 24958 5124
rect 25106 5068 25116 5124
rect 25172 5068 26572 5124
rect 26628 5068 26638 5124
rect 26908 5102 27188 5158
rect 33180 5124 33236 5180
rect 12012 5012 12068 5068
rect 21532 5012 21588 5068
rect 22428 5012 22484 5068
rect 26908 5012 26964 5102
rect 0 4956 3220 5012
rect 3276 4956 11676 5012
rect 11732 4956 11742 5012
rect 12012 4956 16492 5012
rect 16548 4956 16558 5012
rect 16706 4956 16716 5012
rect 16772 4956 21588 5012
rect 21746 4956 21756 5012
rect 21812 4956 22484 5012
rect 22642 4956 22652 5012
rect 22708 4956 25228 5012
rect 25284 4956 25294 5012
rect 25442 4956 25452 5012
rect 25508 4956 26964 5012
rect 27132 5012 27188 5102
rect 28578 5068 28588 5124
rect 28644 5068 32508 5124
rect 32564 5068 32574 5124
rect 33180 5068 33404 5124
rect 33460 5068 33470 5124
rect 33618 5068 33628 5124
rect 33684 5068 38780 5124
rect 38836 5068 38846 5124
rect 39778 5068 39788 5124
rect 39844 5068 46732 5124
rect 46788 5068 46798 5124
rect 49634 5068 49644 5124
rect 49700 5068 51100 5124
rect 51156 5068 51166 5124
rect 52640 5012 52752 5040
rect 27132 4956 29428 5012
rect 29586 4956 29596 5012
rect 29652 4956 35868 5012
rect 35924 4956 35934 5012
rect 36978 4956 36988 5012
rect 37044 4956 42700 5012
rect 42756 4956 42766 5012
rect 46498 4956 46508 5012
rect 46564 4956 48748 5012
rect 48804 4956 48814 5012
rect 51202 4956 51212 5012
rect 51268 4956 52752 5012
rect 0 4928 112 4956
rect 3164 4900 3220 4956
rect 3164 4844 8764 4900
rect 8820 4844 8830 4900
rect 8988 4844 15372 4900
rect 15428 4844 15438 4900
rect 15586 4844 15596 4900
rect 15652 4844 26852 4900
rect 26908 4844 26918 4900
rect 8988 4788 9044 4844
rect 29372 4788 29428 4956
rect 52640 4928 52752 4956
rect 29586 4844 29596 4900
rect 29652 4844 40572 4900
rect 40628 4844 40638 4900
rect 41906 4844 41916 4900
rect 41972 4844 46844 4900
rect 46900 4844 46910 4900
rect 4162 4732 4172 4788
rect 4228 4732 6972 4788
rect 7028 4732 7038 4788
rect 8306 4732 8316 4788
rect 8372 4732 9044 4788
rect 11218 4732 11228 4788
rect 11284 4732 14252 4788
rect 14308 4732 14318 4788
rect 14466 4732 14476 4788
rect 14532 4732 18508 4788
rect 18564 4732 18574 4788
rect 18722 4732 18732 4788
rect 18788 4732 23660 4788
rect 23716 4732 23726 4788
rect 24322 4732 24332 4788
rect 24388 4732 24780 4788
rect 24836 4732 24846 4788
rect 24994 4732 25004 4788
rect 25060 4732 29148 4788
rect 29204 4732 29214 4788
rect 29372 4732 35308 4788
rect 35364 4732 35374 4788
rect 35746 4732 35756 4788
rect 35812 4732 40684 4788
rect 40740 4732 40750 4788
rect 46162 4732 46172 4788
rect 46228 4732 48860 4788
rect 48916 4732 48926 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 6178 4620 6188 4676
rect 6244 4620 9884 4676
rect 9940 4620 9950 4676
rect 11442 4620 11452 4676
rect 11508 4620 21756 4676
rect 21812 4620 21822 4676
rect 24210 4620 24220 4676
rect 24276 4620 25900 4676
rect 25956 4620 25966 4676
rect 26898 4620 26908 4676
rect 26964 4620 33964 4676
rect 34020 4620 34030 4676
rect 35970 4620 35980 4676
rect 36036 4620 37548 4676
rect 37604 4620 37614 4676
rect 37874 4620 37884 4676
rect 37940 4620 41916 4676
rect 41972 4620 41982 4676
rect 0 4564 112 4592
rect 52640 4564 52752 4592
rect 0 4508 5068 4564
rect 5124 4508 5134 4564
rect 6402 4508 6412 4564
rect 6468 4508 7532 4564
rect 7588 4508 7598 4564
rect 7858 4508 7868 4564
rect 7924 4508 13020 4564
rect 13076 4508 13086 4564
rect 13234 4508 13244 4564
rect 13300 4508 18060 4564
rect 18116 4508 18126 4564
rect 18274 4508 18284 4564
rect 18340 4508 20916 4564
rect 21074 4508 21084 4564
rect 21140 4508 26908 4564
rect 26964 4508 26974 4564
rect 27122 4508 27132 4564
rect 27188 4508 32844 4564
rect 32900 4508 32910 4564
rect 33506 4508 33516 4564
rect 33572 4508 45612 4564
rect 45668 4508 45678 4564
rect 51090 4508 51100 4564
rect 51156 4508 52752 4564
rect 0 4480 112 4508
rect 20860 4452 20916 4508
rect 52640 4480 52752 4508
rect 10210 4396 10220 4452
rect 10276 4396 11788 4452
rect 11844 4396 11854 4452
rect 13682 4396 13692 4452
rect 13748 4396 14700 4452
rect 14756 4396 14766 4452
rect 15250 4396 15260 4452
rect 15316 4396 20356 4452
rect 20860 4396 24668 4452
rect 24724 4396 24734 4452
rect 24882 4396 24892 4452
rect 24948 4396 26796 4452
rect 26852 4396 26862 4452
rect 27010 4396 27020 4452
rect 27076 4396 30156 4452
rect 30212 4396 30222 4452
rect 31714 4396 31724 4452
rect 31780 4396 33068 4452
rect 33124 4396 33134 4452
rect 20300 4340 20356 4396
rect 4834 4284 4844 4340
rect 4900 4284 16268 4340
rect 16324 4284 16334 4340
rect 16482 4284 16492 4340
rect 16548 4284 20076 4340
rect 20132 4284 20142 4340
rect 20300 4284 25564 4340
rect 25620 4284 25630 4340
rect 25890 4284 25900 4340
rect 25956 4284 29036 4340
rect 29092 4284 29102 4340
rect 29932 4284 35532 4340
rect 35588 4284 35598 4340
rect 43586 4284 43596 4340
rect 43652 4284 44156 4340
rect 44212 4284 44222 4340
rect 45378 4284 45388 4340
rect 45444 4284 48748 4340
rect 48804 4284 48814 4340
rect 29932 4228 29988 4284
rect 3332 4172 11676 4228
rect 11732 4172 11742 4228
rect 15138 4172 15148 4228
rect 15204 4172 21196 4228
rect 21252 4172 21262 4228
rect 21410 4172 21420 4228
rect 21476 4172 22540 4228
rect 22596 4172 22606 4228
rect 23650 4172 23660 4228
rect 23716 4172 26460 4228
rect 26516 4172 26526 4228
rect 26796 4172 29988 4228
rect 31490 4172 31500 4228
rect 31556 4172 34692 4228
rect 35298 4172 35308 4228
rect 35364 4172 44716 4228
rect 44772 4172 44782 4228
rect 0 4116 112 4144
rect 3332 4116 3388 4172
rect 0 4060 3388 4116
rect 8082 4060 8092 4116
rect 8148 4060 17276 4116
rect 17332 4060 17342 4116
rect 17938 4060 17948 4116
rect 18004 4060 21196 4116
rect 21252 4060 21262 4116
rect 21858 4060 21868 4116
rect 21924 4060 26124 4116
rect 26180 4060 26190 4116
rect 26338 4060 26348 4116
rect 26404 4060 26442 4116
rect 0 4032 112 4060
rect 26796 4004 26852 4172
rect 34636 4116 34692 4172
rect 52640 4116 52752 4144
rect 27010 4060 27020 4116
rect 27076 4060 30380 4116
rect 30436 4060 30446 4116
rect 34636 4060 47404 4116
rect 47460 4060 47740 4116
rect 47796 4060 47806 4116
rect 51426 4060 51436 4116
rect 51492 4060 52752 4116
rect 52640 4032 52752 4060
rect 13010 3948 13020 4004
rect 13076 3948 15260 4004
rect 15316 3948 15326 4004
rect 15484 3948 16380 4004
rect 16436 3948 16446 4004
rect 17154 3948 17164 4004
rect 17220 3948 17612 4004
rect 17668 3948 17678 4004
rect 18610 3948 18620 4004
rect 18676 3948 24220 4004
rect 24276 3948 24286 4004
rect 24882 3948 24892 4004
rect 24948 3948 26852 4004
rect 27020 3948 31836 4004
rect 31892 3948 31902 4004
rect 33282 3948 33292 4004
rect 33348 3948 43708 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 15484 3892 15540 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 27020 3898 27076 3948
rect 26908 3892 27076 3898
rect 8306 3836 8316 3892
rect 8372 3836 15540 3892
rect 15810 3836 15820 3892
rect 15876 3836 20972 3892
rect 21028 3836 21038 3892
rect 21186 3836 21196 3892
rect 21252 3836 24220 3892
rect 24276 3836 24286 3892
rect 25218 3836 25228 3892
rect 25284 3842 27076 3892
rect 25284 3836 26964 3842
rect 27132 3836 37884 3892
rect 37940 3836 37950 3892
rect 27132 3780 27188 3836
rect 43652 3780 43708 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 45266 3836 45276 3892
rect 45332 3836 50428 3892
rect 50484 3836 50494 3892
rect 6178 3724 6188 3780
rect 6244 3724 15372 3780
rect 15428 3724 15438 3780
rect 16818 3724 16828 3780
rect 16884 3724 17444 3780
rect 18050 3724 18060 3780
rect 18116 3724 24220 3780
rect 24276 3724 24286 3780
rect 25106 3724 25116 3780
rect 25172 3724 25340 3780
rect 25396 3724 27188 3780
rect 27468 3724 29372 3780
rect 29428 3724 29438 3780
rect 43652 3724 50204 3780
rect 50260 3724 50270 3780
rect 0 3668 112 3696
rect 17388 3668 17444 3724
rect 27468 3668 27524 3724
rect 52640 3668 52752 3696
rect 0 3612 2212 3668
rect 11330 3612 11340 3668
rect 11396 3612 11676 3668
rect 11732 3612 15820 3668
rect 15876 3612 15886 3668
rect 16044 3612 17164 3668
rect 17220 3612 17230 3668
rect 17388 3612 20860 3668
rect 20916 3612 20926 3668
rect 21298 3612 21308 3668
rect 21364 3612 25228 3668
rect 25284 3612 25294 3668
rect 25442 3612 25452 3668
rect 25508 3612 27524 3668
rect 28690 3612 28700 3668
rect 28756 3612 36652 3668
rect 36708 3612 36718 3668
rect 40338 3612 40348 3668
rect 40404 3612 48300 3668
rect 48356 3612 48366 3668
rect 49410 3612 49420 3668
rect 49476 3612 52752 3668
rect 0 3584 112 3612
rect 2156 3444 2212 3612
rect 16044 3556 16100 3612
rect 52640 3584 52752 3612
rect 2370 3500 2380 3556
rect 2436 3500 2716 3556
rect 2772 3500 16100 3556
rect 16258 3500 16268 3556
rect 16324 3500 17052 3556
rect 17108 3500 17118 3556
rect 17388 3500 18844 3556
rect 18900 3500 18910 3556
rect 19068 3500 24332 3556
rect 24388 3500 24398 3556
rect 25218 3500 25228 3556
rect 25284 3500 26572 3556
rect 26628 3500 26638 3556
rect 26786 3500 26796 3556
rect 26852 3500 28420 3556
rect 17388 3444 17444 3500
rect 19068 3444 19124 3500
rect 28364 3444 28420 3500
rect 30044 3500 32620 3556
rect 32676 3500 32686 3556
rect 33170 3500 33180 3556
rect 33236 3500 45612 3556
rect 45668 3500 45836 3556
rect 45892 3500 45902 3556
rect 2156 3388 6804 3444
rect 6962 3388 6972 3444
rect 7028 3388 17444 3444
rect 17602 3388 17612 3444
rect 17668 3388 19124 3444
rect 19282 3388 19292 3444
rect 19348 3388 22652 3444
rect 22708 3388 22718 3444
rect 23548 3388 27244 3444
rect 27300 3388 27310 3444
rect 28364 3388 29820 3444
rect 29876 3388 29886 3444
rect 6748 3332 6804 3388
rect 23548 3332 23604 3388
rect 30044 3332 30100 3500
rect 30370 3388 30380 3444
rect 30436 3388 32732 3444
rect 32788 3388 32798 3444
rect 37090 3388 37100 3444
rect 37156 3388 43596 3444
rect 43652 3388 43662 3444
rect 49858 3388 49868 3444
rect 49924 3388 51100 3444
rect 51156 3388 51166 3444
rect 2594 3276 2604 3332
rect 2660 3276 5236 3332
rect 6748 3276 18284 3332
rect 18340 3276 18350 3332
rect 18610 3276 18620 3332
rect 18676 3276 22428 3332
rect 22484 3276 22494 3332
rect 23538 3276 23548 3332
rect 23604 3276 23614 3332
rect 23874 3276 23884 3332
rect 23940 3276 24276 3332
rect 24434 3276 24444 3332
rect 24500 3276 25340 3332
rect 25396 3276 25406 3332
rect 25554 3276 25564 3332
rect 25620 3276 30100 3332
rect 30258 3276 30268 3332
rect 30324 3276 35420 3332
rect 35476 3276 35486 3332
rect 38770 3276 38780 3332
rect 38836 3276 47516 3332
rect 47572 3276 47582 3332
rect 0 3220 112 3248
rect 5180 3220 5236 3276
rect 24220 3220 24276 3276
rect 52640 3220 52752 3248
rect 0 3164 3612 3220
rect 3668 3164 3678 3220
rect 5180 3164 8092 3220
rect 8148 3164 8158 3220
rect 11218 3164 11228 3220
rect 11284 3164 16940 3220
rect 16996 3164 17006 3220
rect 17154 3164 17164 3220
rect 17220 3164 19292 3220
rect 19348 3164 19358 3220
rect 19506 3164 19516 3220
rect 19572 3164 23660 3220
rect 23716 3164 23726 3220
rect 24220 3164 24892 3220
rect 24948 3164 24958 3220
rect 25778 3164 25788 3220
rect 25844 3164 26796 3220
rect 26852 3164 26862 3220
rect 27010 3164 27020 3220
rect 27076 3164 30156 3220
rect 30212 3164 30222 3220
rect 30380 3164 35756 3220
rect 35812 3164 35822 3220
rect 51202 3164 51212 3220
rect 51268 3164 52752 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 30380 3108 30436 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 52640 3136 52752 3164
rect 5170 3052 5180 3108
rect 5236 3052 7644 3108
rect 7700 3052 7710 3108
rect 11778 3052 11788 3108
rect 11844 3052 14588 3108
rect 14644 3052 14654 3108
rect 17154 3052 17164 3108
rect 17220 3052 23548 3108
rect 23604 3052 23614 3108
rect 24322 3052 24332 3108
rect 24388 3052 25788 3108
rect 25844 3052 25854 3108
rect 26002 3052 26012 3108
rect 26068 3052 30436 3108
rect 31938 3052 31948 3108
rect 32004 3052 33404 3108
rect 33460 3052 33470 3108
rect 35298 3052 35308 3108
rect 35364 3052 43036 3108
rect 43092 3052 43102 3108
rect 5282 2940 5292 2996
rect 5348 2940 14140 2996
rect 14196 2940 14206 2996
rect 15138 2940 15148 2996
rect 15204 2940 18956 2996
rect 19012 2940 19022 2996
rect 19170 2940 19180 2996
rect 19236 2940 21308 2996
rect 21364 2940 21374 2996
rect 21746 2940 21756 2996
rect 21812 2940 26796 2996
rect 26852 2940 26862 2996
rect 27346 2940 27356 2996
rect 27412 2940 30604 2996
rect 30660 2940 30670 2996
rect 33170 2940 33180 2996
rect 33236 2940 38556 2996
rect 38612 2940 38892 2996
rect 38948 2940 38958 2996
rect 39116 2940 42364 2996
rect 42420 2940 42430 2996
rect 39116 2884 39172 2940
rect 2146 2828 2156 2884
rect 2212 2828 6972 2884
rect 7028 2828 7038 2884
rect 7522 2828 7532 2884
rect 7588 2828 14140 2884
rect 14196 2828 14206 2884
rect 16146 2828 16156 2884
rect 16212 2828 16828 2884
rect 16884 2828 16894 2884
rect 17042 2828 17052 2884
rect 17108 2828 22204 2884
rect 22260 2828 22270 2884
rect 22418 2828 22428 2884
rect 22484 2828 26684 2884
rect 26740 2828 26750 2884
rect 26898 2828 26908 2884
rect 26964 2828 29596 2884
rect 29652 2828 29662 2884
rect 29922 2828 29932 2884
rect 29988 2828 39172 2884
rect 40450 2828 40460 2884
rect 40516 2828 45164 2884
rect 45220 2828 45230 2884
rect 48066 2828 48076 2884
rect 48132 2828 50540 2884
rect 50596 2828 50606 2884
rect 0 2772 112 2800
rect 52640 2772 52752 2800
rect 0 2716 11564 2772
rect 11620 2716 11630 2772
rect 12450 2716 12460 2772
rect 12516 2716 18396 2772
rect 18452 2716 18462 2772
rect 18722 2716 18732 2772
rect 18788 2716 19516 2772
rect 19572 2716 19582 2772
rect 20066 2716 20076 2772
rect 20132 2716 26236 2772
rect 26292 2716 26302 2772
rect 26450 2716 26460 2772
rect 26516 2716 32788 2772
rect 38210 2716 38220 2772
rect 38276 2716 47068 2772
rect 47124 2716 47134 2772
rect 51090 2716 51100 2772
rect 51156 2716 52752 2772
rect 0 2688 112 2716
rect 32732 2660 32788 2716
rect 52640 2688 52752 2716
rect 9874 2604 9884 2660
rect 9940 2604 13804 2660
rect 13860 2604 13870 2660
rect 14130 2604 14140 2660
rect 14196 2604 22148 2660
rect 23426 2604 23436 2660
rect 23492 2604 28812 2660
rect 28868 2604 28878 2660
rect 29820 2604 31948 2660
rect 32004 2604 32014 2660
rect 32732 2604 40796 2660
rect 40852 2604 40862 2660
rect 45938 2604 45948 2660
rect 46004 2604 48860 2660
rect 48916 2604 48926 2660
rect 49410 2604 49420 2660
rect 49476 2604 51548 2660
rect 51604 2604 51614 2660
rect 22092 2548 22148 2604
rect 29820 2548 29876 2604
rect 4172 2492 6188 2548
rect 6244 2492 6254 2548
rect 9762 2492 9772 2548
rect 9828 2492 16156 2548
rect 16212 2492 16222 2548
rect 16706 2492 16716 2548
rect 16772 2492 20076 2548
rect 20132 2492 20142 2548
rect 20290 2492 20300 2548
rect 20356 2492 22036 2548
rect 22092 2492 29876 2548
rect 30034 2492 30044 2548
rect 30100 2492 37660 2548
rect 37716 2492 37726 2548
rect 38658 2492 38668 2548
rect 38724 2492 39564 2548
rect 39620 2492 39630 2548
rect 47506 2492 47516 2548
rect 47572 2492 50428 2548
rect 50484 2492 50494 2548
rect 0 2324 112 2352
rect 4172 2324 4228 2492
rect 21980 2436 22036 2492
rect 8194 2380 8204 2436
rect 8260 2380 10388 2436
rect 10546 2380 10556 2436
rect 10612 2380 12572 2436
rect 12628 2380 12638 2436
rect 14130 2380 14140 2436
rect 14196 2380 21756 2436
rect 21812 2380 21822 2436
rect 21980 2380 24332 2436
rect 24388 2380 24398 2436
rect 24882 2380 24892 2436
rect 24948 2380 26460 2436
rect 26516 2380 26526 2436
rect 28578 2380 28588 2436
rect 28644 2380 30380 2436
rect 30436 2380 30446 2436
rect 30594 2380 30604 2436
rect 30660 2380 39452 2436
rect 39508 2380 39518 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 0 2268 4228 2324
rect 0 2240 112 2268
rect 10332 2212 10388 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 52640 2324 52752 2352
rect 12226 2268 12236 2324
rect 12292 2268 12684 2324
rect 12740 2268 12750 2324
rect 15362 2268 15372 2324
rect 15428 2268 23660 2324
rect 23716 2268 23726 2324
rect 25666 2268 25676 2324
rect 25732 2268 38668 2324
rect 38724 2268 38734 2324
rect 39218 2268 39228 2324
rect 39284 2268 43708 2324
rect 51426 2268 51436 2324
rect 51492 2268 52752 2324
rect 43652 2212 43708 2268
rect 52640 2240 52752 2268
rect 1586 2156 1596 2212
rect 1652 2156 9996 2212
rect 10052 2156 10062 2212
rect 10332 2156 16716 2212
rect 16772 2156 16782 2212
rect 16930 2156 16940 2212
rect 16996 2156 18620 2212
rect 18676 2156 18686 2212
rect 19506 2156 19516 2212
rect 19572 2156 19852 2212
rect 19908 2156 21644 2212
rect 21700 2156 21710 2212
rect 22082 2156 22092 2212
rect 22148 2156 26068 2212
rect 26226 2156 26236 2212
rect 26292 2156 28588 2212
rect 28644 2156 28654 2212
rect 29138 2156 29148 2212
rect 29204 2156 33628 2212
rect 33684 2156 33694 2212
rect 38882 2156 38892 2212
rect 38948 2156 39116 2212
rect 39172 2156 39182 2212
rect 39340 2156 41748 2212
rect 43652 2156 48748 2212
rect 48804 2156 48814 2212
rect 26012 2100 26068 2156
rect 39340 2100 39396 2156
rect 41692 2100 41748 2156
rect 8754 2044 8764 2100
rect 8820 2044 13748 2100
rect 14242 2044 14252 2100
rect 14308 2044 25788 2100
rect 25844 2044 25854 2100
rect 26012 2044 32620 2100
rect 32676 2044 32686 2100
rect 32844 2044 34860 2100
rect 34916 2044 34926 2100
rect 36978 2044 36988 2100
rect 37044 2044 39396 2100
rect 39666 2044 39676 2100
rect 39732 2044 41468 2100
rect 41524 2044 41534 2100
rect 41692 2044 46732 2100
rect 46788 2044 46956 2100
rect 47012 2044 47022 2100
rect 13692 1988 13748 2044
rect 32844 1988 32900 2044
rect 4162 1932 4172 1988
rect 4228 1932 13468 1988
rect 13524 1932 13534 1988
rect 13692 1932 17164 1988
rect 17220 1932 17230 1988
rect 17378 1932 17388 1988
rect 17444 1932 18060 1988
rect 18116 1932 18126 1988
rect 18274 1932 18284 1988
rect 18340 1932 29596 1988
rect 29652 1932 29662 1988
rect 30818 1932 30828 1988
rect 30884 1932 32900 1988
rect 33394 1932 33404 1988
rect 33460 1932 48972 1988
rect 49028 1932 49038 1988
rect 0 1876 112 1904
rect 52640 1876 52752 1904
rect 0 1820 12460 1876
rect 12516 1820 12526 1876
rect 13906 1820 13916 1876
rect 13972 1820 19404 1876
rect 19460 1820 19470 1876
rect 21522 1820 21532 1876
rect 21588 1820 25228 1876
rect 25284 1820 25294 1876
rect 26114 1820 26124 1876
rect 26180 1820 28700 1876
rect 28756 1820 28766 1876
rect 32722 1820 32732 1876
rect 32788 1820 44268 1876
rect 44324 1820 44334 1876
rect 49858 1820 49868 1876
rect 49924 1820 52752 1876
rect 0 1792 112 1820
rect 52640 1792 52752 1820
rect 8764 1708 9268 1764
rect 13346 1708 13356 1764
rect 13412 1708 30156 1764
rect 30212 1708 30222 1764
rect 32722 1708 32732 1764
rect 32788 1708 36932 1764
rect 8764 1652 8820 1708
rect 9212 1652 9268 1708
rect 36876 1652 36932 1708
rect 43652 1708 46172 1764
rect 46228 1708 46238 1764
rect 43652 1652 43708 1708
rect 6514 1596 6524 1652
rect 6580 1596 8820 1652
rect 8950 1596 8988 1652
rect 9044 1596 9054 1652
rect 9212 1596 11228 1652
rect 11284 1596 11294 1652
rect 11554 1596 11564 1652
rect 11620 1596 15148 1652
rect 16370 1596 16380 1652
rect 16436 1596 18620 1652
rect 18676 1596 18686 1652
rect 19394 1596 19404 1652
rect 19460 1596 21308 1652
rect 21364 1596 21374 1652
rect 21522 1596 21532 1652
rect 21588 1596 22204 1652
rect 22260 1596 22270 1652
rect 22530 1596 22540 1652
rect 22596 1596 23660 1652
rect 23716 1596 23726 1652
rect 24210 1596 24220 1652
rect 24276 1596 24780 1652
rect 24836 1596 24846 1652
rect 24994 1596 25004 1652
rect 25060 1596 35196 1652
rect 35252 1596 35262 1652
rect 36876 1596 43708 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 15092 1540 15148 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 6290 1484 6300 1540
rect 6356 1484 13356 1540
rect 13412 1484 13422 1540
rect 15092 1484 18676 1540
rect 18834 1484 18844 1540
rect 18900 1484 23100 1540
rect 23156 1484 23166 1540
rect 24210 1484 24220 1540
rect 24276 1484 24892 1540
rect 24948 1484 24958 1540
rect 25218 1484 25228 1540
rect 25284 1484 30828 1540
rect 30884 1484 30894 1540
rect 31042 1484 31052 1540
rect 31108 1484 40236 1540
rect 40292 1484 40302 1540
rect 0 1428 112 1456
rect 18620 1428 18676 1484
rect 52640 1428 52752 1456
rect 0 1372 5628 1428
rect 5684 1372 5694 1428
rect 13458 1372 13468 1428
rect 13524 1372 17948 1428
rect 18004 1372 18014 1428
rect 18620 1372 19180 1428
rect 19236 1372 19246 1428
rect 20178 1372 20188 1428
rect 20244 1372 21532 1428
rect 21588 1372 21598 1428
rect 21858 1372 21868 1428
rect 21924 1372 28588 1428
rect 28644 1372 28654 1428
rect 28802 1372 28812 1428
rect 28868 1372 35588 1428
rect 37874 1372 37884 1428
rect 37940 1372 45948 1428
rect 46004 1372 46014 1428
rect 49746 1372 49756 1428
rect 49812 1372 52752 1428
rect 0 1344 112 1372
rect 35532 1316 35588 1372
rect 52640 1344 52752 1372
rect 14466 1260 14476 1316
rect 14532 1260 35308 1316
rect 35364 1260 35374 1316
rect 35532 1260 38108 1316
rect 38164 1260 38174 1316
rect 5058 1148 5068 1204
rect 5124 1148 15372 1204
rect 15428 1148 15438 1204
rect 15586 1148 15596 1204
rect 15652 1148 20300 1204
rect 20356 1148 20366 1204
rect 20850 1148 20860 1204
rect 20916 1148 21084 1204
rect 21140 1148 25004 1204
rect 25060 1148 25070 1204
rect 26338 1148 26348 1204
rect 26404 1148 33740 1204
rect 33796 1148 33806 1204
rect 36642 1148 36652 1204
rect 36708 1148 47180 1204
rect 47236 1148 47246 1204
rect 2482 1036 2492 1092
rect 2548 1036 26796 1092
rect 26852 1036 26862 1092
rect 30146 1036 30156 1092
rect 30212 1036 48748 1092
rect 48804 1036 48814 1092
rect 0 980 112 1008
rect 52640 980 52752 1008
rect 0 924 3276 980
rect 3332 924 3342 980
rect 12562 924 12572 980
rect 12628 924 19964 980
rect 20020 924 20030 980
rect 20132 924 30212 980
rect 30370 924 30380 980
rect 30436 924 50428 980
rect 50484 924 50764 980
rect 50820 924 50830 980
rect 50988 924 52752 980
rect 0 896 112 924
rect 20132 868 20188 924
rect 30156 868 30212 924
rect 50988 868 51044 924
rect 52640 896 52752 924
rect 13458 812 13468 868
rect 13524 812 20188 868
rect 20626 812 20636 868
rect 20692 812 24332 868
rect 24388 812 24398 868
rect 24892 812 27692 868
rect 27748 812 27758 868
rect 30156 812 33516 868
rect 33572 812 33582 868
rect 33730 812 33740 868
rect 33796 812 43260 868
rect 43316 812 43326 868
rect 48178 812 48188 868
rect 48244 812 51044 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 8372 700 20412 756
rect 20468 700 20478 756
rect 21186 700 21196 756
rect 21252 700 22540 756
rect 22596 700 22606 756
rect 22754 700 22764 756
rect 22820 700 23996 756
rect 24052 700 24062 756
rect 0 532 112 560
rect 8372 532 8428 700
rect 24892 644 24948 812
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 15362 588 15372 644
rect 15428 588 16996 644
rect 17602 588 17612 644
rect 17668 588 24948 644
rect 25004 700 30044 756
rect 30100 700 30110 756
rect 16940 532 16996 588
rect 25004 532 25060 700
rect 25218 588 25228 644
rect 25284 588 47292 644
rect 47348 588 47358 644
rect 52640 532 52752 560
rect 0 476 4172 532
rect 4228 476 4238 532
rect 6738 476 6748 532
rect 6804 476 8428 532
rect 11890 476 11900 532
rect 11956 476 16716 532
rect 16772 476 16782 532
rect 16940 476 22876 532
rect 22932 476 22942 532
rect 23090 476 23100 532
rect 23156 476 25060 532
rect 25218 476 25228 532
rect 25284 476 36988 532
rect 37044 476 37054 532
rect 50530 476 50540 532
rect 50596 476 52752 532
rect 0 448 112 476
rect 52640 448 52752 476
rect 4050 364 4060 420
rect 4116 364 8316 420
rect 8372 364 8382 420
rect 12674 364 12684 420
rect 12740 364 22316 420
rect 22372 364 22382 420
rect 22530 364 22540 420
rect 22596 364 26628 420
rect 26786 364 26796 420
rect 26852 364 41804 420
rect 41860 364 41870 420
rect 26572 308 26628 364
rect 19842 252 19852 308
rect 19908 252 22316 308
rect 22372 252 22382 308
rect 22642 252 22652 308
rect 22708 252 26516 308
rect 26572 252 34188 308
rect 34244 252 34254 308
rect 37538 252 37548 308
rect 37604 252 50876 308
rect 50932 252 50942 308
rect 26460 196 26516 252
rect 7410 140 7420 196
rect 7476 140 23772 196
rect 23828 140 23838 196
rect 23986 140 23996 196
rect 24052 140 25228 196
rect 25284 140 25294 196
rect 26226 140 26236 196
rect 26292 140 26302 196
rect 26460 140 32732 196
rect 32788 140 32798 196
rect 37986 140 37996 196
rect 38052 140 38556 196
rect 38612 140 38622 196
rect 39778 140 39788 196
rect 39844 140 48412 196
rect 48468 140 48478 196
rect 0 84 112 112
rect 26236 84 26292 140
rect 52640 84 52752 112
rect 0 28 5180 84
rect 5236 28 5246 84
rect 9650 28 9660 84
rect 9716 28 26292 84
rect 26898 28 26908 84
rect 26964 28 31052 84
rect 31108 28 31118 84
rect 51538 28 51548 84
rect 51604 28 52752 84
rect 0 0 112 28
rect 52640 0 52752 28
<< via3 >>
rect 16156 14028 16212 14084
rect 16380 14028 16436 14084
rect 26684 14028 26740 14084
rect 32060 14028 32116 14084
rect 14924 13916 14980 13972
rect 21420 13916 21476 13972
rect 22876 13916 22932 13972
rect 29372 13804 29428 13860
rect 13580 13692 13636 13748
rect 24892 13580 24948 13636
rect 25116 13580 25172 13636
rect 16156 13468 16212 13524
rect 32732 13468 32788 13524
rect 18732 13356 18788 13412
rect 21868 13356 21924 13412
rect 22204 13356 22260 13412
rect 24220 13356 24276 13412
rect 26460 13356 26516 13412
rect 32060 13356 32116 13412
rect 33852 13356 33908 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 20748 13244 20804 13300
rect 24892 13244 24948 13300
rect 26908 13244 26964 13300
rect 30940 13244 30996 13300
rect 23660 13132 23716 13188
rect 24220 13132 24276 13188
rect 31164 13020 31220 13076
rect 33628 13020 33684 13076
rect 13244 12908 13300 12964
rect 28252 12908 28308 12964
rect 32732 12908 32788 12964
rect 39564 12908 39620 12964
rect 18732 12796 18788 12852
rect 25340 12796 25396 12852
rect 30940 12796 30996 12852
rect 15148 12684 15204 12740
rect 16492 12684 16548 12740
rect 30604 12684 30660 12740
rect 33852 12684 33908 12740
rect 19292 12572 19348 12628
rect 24220 12572 24276 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 19740 12348 19796 12404
rect 24892 12348 24948 12404
rect 31948 12348 32004 12404
rect 33964 12348 34020 12404
rect 39564 12348 39620 12404
rect 17724 12236 17780 12292
rect 19404 12236 19460 12292
rect 20748 12236 20804 12292
rect 23436 12236 23492 12292
rect 15148 12124 15204 12180
rect 17612 12124 17668 12180
rect 20524 12124 20580 12180
rect 26348 12012 26404 12068
rect 28252 12012 28308 12068
rect 28476 12012 28532 12068
rect 33964 12012 34020 12068
rect 39116 12012 39172 12068
rect 17948 11900 18004 11956
rect 18620 11900 18676 11956
rect 22316 11900 22372 11956
rect 24892 11900 24948 11956
rect 26796 11900 26852 11956
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 13468 11788 13524 11844
rect 14924 11788 14980 11844
rect 18060 11788 18116 11844
rect 18732 11788 18788 11844
rect 20188 11788 20244 11844
rect 25116 11788 25172 11844
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 18508 11676 18564 11732
rect 20300 11676 20356 11732
rect 22540 11676 22596 11732
rect 24220 11676 24276 11732
rect 24892 11676 24948 11732
rect 28476 11676 28532 11732
rect 13468 11564 13524 11620
rect 35532 11564 35588 11620
rect 41804 11564 41860 11620
rect 16492 11452 16548 11508
rect 20188 11452 20244 11508
rect 27356 11452 27412 11508
rect 16268 11340 16324 11396
rect 17724 11340 17780 11396
rect 21420 11340 21476 11396
rect 22988 11228 23044 11284
rect 26348 11228 26404 11284
rect 27356 11228 27412 11284
rect 16716 11116 16772 11172
rect 28252 11116 28308 11172
rect 29932 11116 29988 11172
rect 23100 11004 23156 11060
rect 24892 11004 24948 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 13580 10892 13636 10948
rect 16044 10892 16100 10948
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 16492 10892 16548 10948
rect 19068 10892 19124 10948
rect 26796 10892 26852 10948
rect 27020 10892 27076 10948
rect 31500 10892 31556 10948
rect 34188 10892 34244 10948
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 15932 10780 15988 10836
rect 21868 10780 21924 10836
rect 22428 10780 22484 10836
rect 24220 10780 24276 10836
rect 28252 10780 28308 10836
rect 8988 10668 9044 10724
rect 26684 10556 26740 10612
rect 26908 10556 26964 10612
rect 29932 10556 29988 10612
rect 21532 10444 21588 10500
rect 23100 10444 23156 10500
rect 33516 10444 33572 10500
rect 9548 10332 9604 10388
rect 14028 10332 14084 10388
rect 39228 10332 39284 10388
rect 23436 10220 23492 10276
rect 23660 10220 23716 10276
rect 26684 10220 26740 10276
rect 28476 10220 28532 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 17724 10108 17780 10164
rect 19068 10108 19124 10164
rect 20076 10108 20132 10164
rect 20300 10108 20356 10164
rect 28924 10108 28980 10164
rect 26572 9996 26628 10052
rect 19068 9884 19124 9940
rect 30940 9884 30996 9940
rect 20972 9772 21028 9828
rect 22652 9772 22708 9828
rect 31724 9772 31780 9828
rect 21868 9660 21924 9716
rect 16716 9548 16772 9604
rect 21532 9436 21588 9492
rect 22988 9436 23044 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 18508 9324 18564 9380
rect 25228 9324 25284 9380
rect 31500 9324 31556 9380
rect 17276 9212 17332 9268
rect 22092 9212 22148 9268
rect 37212 9212 37268 9268
rect 15148 9100 15204 9156
rect 17276 8988 17332 9044
rect 19292 8988 19348 9044
rect 28476 8988 28532 9044
rect 22428 8876 22484 8932
rect 23100 8876 23156 8932
rect 26908 8876 26964 8932
rect 37212 8876 37268 8932
rect 16828 8764 16884 8820
rect 19964 8764 20020 8820
rect 20188 8764 20244 8820
rect 21868 8764 21924 8820
rect 25564 8764 25620 8820
rect 30940 8764 30996 8820
rect 33292 8764 33348 8820
rect 11676 8652 11732 8708
rect 20076 8652 20132 8708
rect 20412 8652 20468 8708
rect 34860 8652 34916 8708
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 17500 8540 17556 8596
rect 23100 8540 23156 8596
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 33404 8540 33460 8596
rect 38444 8540 38500 8596
rect 11676 8316 11732 8372
rect 15820 8316 15876 8372
rect 16604 8316 16660 8372
rect 25676 8204 25732 8260
rect 14028 8092 14084 8148
rect 16604 8092 16660 8148
rect 16828 8092 16884 8148
rect 21868 7980 21924 8036
rect 25340 7868 25396 7924
rect 33516 7868 33572 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 9996 7756 10052 7812
rect 15148 7756 15204 7812
rect 20076 7756 20132 7812
rect 24220 7756 24276 7812
rect 31948 7644 32004 7700
rect 19404 7532 19460 7588
rect 22316 7532 22372 7588
rect 22876 7532 22932 7588
rect 26572 7532 26628 7588
rect 28924 7532 28980 7588
rect 13804 7420 13860 7476
rect 17612 7420 17668 7476
rect 20076 7420 20132 7476
rect 13356 7308 13412 7364
rect 28476 7308 28532 7364
rect 15932 7196 15988 7252
rect 16156 7196 16212 7252
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 15484 6972 15540 7028
rect 15708 6972 15764 7028
rect 27020 7196 27076 7252
rect 28140 7196 28196 7252
rect 31724 7196 31780 7252
rect 39228 7196 39284 7252
rect 22764 7084 22820 7140
rect 26684 7084 26740 7140
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 18508 6972 18564 7028
rect 19852 6972 19908 7028
rect 20076 6972 20132 7028
rect 28252 6972 28308 7028
rect 28476 6972 28532 7028
rect 38556 6972 38612 7028
rect 19404 6860 19460 6916
rect 23212 6748 23268 6804
rect 20972 6636 21028 6692
rect 22764 6636 22820 6692
rect 29708 6636 29764 6692
rect 14700 6524 14756 6580
rect 15708 6524 15764 6580
rect 15932 6524 15988 6580
rect 16940 6412 16996 6468
rect 25452 6412 25508 6468
rect 13804 6300 13860 6356
rect 16604 6300 16660 6356
rect 17052 6300 17108 6356
rect 29708 6300 29764 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 9548 6188 9604 6244
rect 24220 6188 24276 6244
rect 25004 6188 25060 6244
rect 25228 6188 25284 6244
rect 28140 6188 28196 6244
rect 29932 6188 29988 6244
rect 14700 6076 14756 6132
rect 15036 6076 15092 6132
rect 17500 6076 17556 6132
rect 24220 5964 24276 6020
rect 16268 5852 16324 5908
rect 27020 5852 27076 5908
rect 28252 5852 28308 5908
rect 35532 5852 35588 5908
rect 24892 5740 24948 5796
rect 20636 5628 20692 5684
rect 21756 5628 21812 5684
rect 15036 5516 15092 5572
rect 16716 5516 16772 5572
rect 21308 5516 21364 5572
rect 25004 5516 25060 5572
rect 26460 5516 26516 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 17836 5404 17892 5460
rect 23436 5404 23492 5460
rect 24892 5404 24948 5460
rect 11676 5292 11732 5348
rect 25116 5292 25172 5348
rect 27804 5180 27860 5236
rect 9996 5068 10052 5124
rect 17836 5068 17892 5124
rect 18732 5068 18788 5124
rect 18956 5068 19012 5124
rect 22988 5068 23044 5124
rect 25116 5068 25172 5124
rect 26572 5068 26628 5124
rect 11676 4956 11732 5012
rect 16492 4956 16548 5012
rect 25228 4956 25284 5012
rect 28588 5068 28644 5124
rect 33404 5068 33460 5124
rect 29596 4956 29652 5012
rect 26852 4844 26908 4900
rect 8316 4732 8372 4788
rect 18732 4732 18788 4788
rect 29148 4732 29204 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 25900 4620 25956 4676
rect 26908 4620 26964 4676
rect 13020 4508 13076 4564
rect 13244 4508 13300 4564
rect 14700 4396 14756 4452
rect 15260 4396 15316 4452
rect 24892 4396 24948 4452
rect 26796 4396 26852 4452
rect 16268 4284 16324 4340
rect 16492 4284 16548 4340
rect 20076 4284 20132 4340
rect 25564 4284 25620 4340
rect 25900 4284 25956 4340
rect 15148 4172 15204 4228
rect 23660 4172 23716 4228
rect 26460 4172 26516 4228
rect 21196 4060 21252 4116
rect 26348 4060 26404 4116
rect 27020 4060 27076 4116
rect 30380 4060 30436 4116
rect 13020 3948 13076 4004
rect 15260 3948 15316 4004
rect 16380 3948 16436 4004
rect 17612 3948 17668 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 21196 3836 21252 3892
rect 24220 3836 24276 3892
rect 25228 3836 25284 3892
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 16828 3724 16884 3780
rect 29372 3724 29428 3780
rect 25228 3612 25284 3668
rect 28700 3612 28756 3668
rect 17052 3500 17108 3556
rect 18844 3500 18900 3556
rect 26572 3500 26628 3556
rect 17612 3388 17668 3444
rect 19292 3388 19348 3444
rect 18620 3276 18676 3332
rect 22428 3276 22484 3332
rect 23548 3276 23604 3332
rect 25564 3276 25620 3332
rect 16940 3164 16996 3220
rect 19292 3164 19348 3220
rect 26796 3164 26852 3220
rect 27020 3164 27076 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 17164 3052 17220 3108
rect 23548 3052 23604 3108
rect 25788 3052 25844 3108
rect 14140 2828 14196 2884
rect 17052 2828 17108 2884
rect 22204 2828 22260 2884
rect 22428 2828 22484 2884
rect 26908 2828 26964 2884
rect 29932 2828 29988 2884
rect 18396 2716 18452 2772
rect 18732 2716 18788 2772
rect 26236 2716 26292 2772
rect 23436 2604 23492 2660
rect 16156 2492 16212 2548
rect 20300 2492 20356 2548
rect 14140 2380 14196 2436
rect 28588 2380 28644 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 23660 2268 23716 2324
rect 25676 2268 25732 2324
rect 16716 2156 16772 2212
rect 18620 2156 18676 2212
rect 26236 2156 26292 2212
rect 28588 2156 28644 2212
rect 29148 2156 29204 2212
rect 39116 2156 39172 2212
rect 32620 2044 32676 2100
rect 34860 2044 34916 2100
rect 18060 1932 18116 1988
rect 29596 1932 29652 1988
rect 19404 1820 19460 1876
rect 32732 1820 32788 1876
rect 8988 1596 9044 1652
rect 24220 1596 24276 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 24892 1484 24948 1540
rect 31052 1484 31108 1540
rect 17948 1372 18004 1428
rect 28588 1372 28644 1428
rect 15372 1148 15428 1204
rect 15596 1148 15652 1204
rect 20300 1148 20356 1204
rect 25004 1148 25060 1204
rect 33740 1148 33796 1204
rect 30380 924 30436 980
rect 13468 812 13524 868
rect 20636 812 20692 868
rect 33740 812 33796 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 20412 700 20468 756
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 15372 588 15428 644
rect 25228 588 25284 644
rect 23100 476 23156 532
rect 8316 364 8372 420
rect 22316 364 22372 420
rect 41804 364 41860 420
rect 22652 252 22708 308
rect 34188 252 34244 308
rect 25228 140 25284 196
rect 31052 28 31108 84
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14224
rect 16156 14084 16212 14094
rect 14924 13972 14980 13982
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 13580 13748 13636 13758
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 13244 12964 13300 12974
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 8988 10724 9044 10734
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 8316 4788 8372 4798
rect 8316 420 8372 4732
rect 8988 1652 9044 10668
rect 9548 10388 9604 10398
rect 9548 6244 9604 10332
rect 11676 8708 11732 8718
rect 11676 8372 11732 8652
rect 11676 8306 11732 8316
rect 9548 6178 9604 6188
rect 9996 7812 10052 7822
rect 9996 5124 10052 7756
rect 9996 5058 10052 5068
rect 11676 5348 11732 5358
rect 11676 5012 11732 5292
rect 11676 4946 11732 4956
rect 13020 4564 13076 4574
rect 13020 4004 13076 4508
rect 13244 4564 13300 12908
rect 13468 11844 13524 11854
rect 13468 11620 13524 11788
rect 13468 11554 13524 11564
rect 13580 10948 13636 13692
rect 14924 11844 14980 13916
rect 16156 13524 16212 14028
rect 16156 13458 16212 13468
rect 16380 14084 16436 14094
rect 15148 12740 15204 12750
rect 15148 12180 15204 12684
rect 15148 12114 15204 12124
rect 14924 11778 14980 11788
rect 16380 11638 16436 14028
rect 21420 13972 21476 13982
rect 18732 13412 18788 13422
rect 18732 12852 18788 13356
rect 18732 12786 18788 12796
rect 20748 13300 20804 13310
rect 13580 10882 13636 10892
rect 15820 11582 16436 11638
rect 16492 12740 16548 12750
rect 14028 10388 14084 10398
rect 14028 8148 14084 10332
rect 14028 8082 14084 8092
rect 15148 9156 15204 9166
rect 15148 7812 15204 9100
rect 15820 8372 15876 11582
rect 16492 11508 16548 12684
rect 19292 12628 19348 12638
rect 16492 11442 16548 11452
rect 16940 12302 17780 12358
rect 16268 11396 16324 11406
rect 16268 11098 16324 11340
rect 15932 11042 16324 11098
rect 16716 11172 16772 11182
rect 15932 10836 15988 11042
rect 15932 10770 15988 10780
rect 16044 10948 16100 10958
rect 16044 10558 16100 10892
rect 16492 10948 16548 10958
rect 16492 10558 16548 10892
rect 16044 10502 16548 10558
rect 16716 9604 16772 11116
rect 16716 9538 16772 9548
rect 16828 8820 16884 8830
rect 15820 8306 15876 8316
rect 16604 8372 16660 8382
rect 16604 8148 16660 8316
rect 16604 8082 16660 8092
rect 16828 8148 16884 8764
rect 16828 8082 16884 8092
rect 15148 7746 15204 7756
rect 13804 7476 13860 7486
rect 13356 7364 13412 7374
rect 13412 7308 13524 7318
rect 13356 7262 13524 7308
rect 13244 4498 13300 4508
rect 13020 3938 13076 3948
rect 8988 1586 9044 1596
rect 13468 868 13524 7262
rect 13804 6356 13860 7420
rect 15932 7252 15988 7262
rect 15484 7028 15540 7038
rect 15484 6778 15540 6972
rect 15708 7028 15764 7038
rect 15484 6722 15652 6778
rect 13804 6290 13860 6300
rect 14700 6580 14756 6590
rect 14700 6132 14756 6524
rect 14700 6066 14756 6076
rect 15036 6132 15092 6142
rect 15036 5572 15092 6076
rect 15036 5506 15092 5516
rect 14700 4452 14756 4462
rect 15260 4452 15316 4462
rect 14756 4396 15204 4438
rect 14700 4382 15204 4396
rect 15148 4228 15204 4382
rect 15148 4162 15204 4172
rect 15260 4004 15316 4396
rect 15260 3938 15316 3948
rect 14140 2884 14196 2894
rect 14140 2436 14196 2828
rect 14140 2370 14196 2380
rect 13468 802 13524 812
rect 15372 1204 15428 1214
rect 15372 644 15428 1148
rect 15596 1204 15652 6722
rect 15708 6580 15764 6972
rect 15708 6514 15764 6524
rect 15932 6580 15988 7196
rect 15932 6514 15988 6524
rect 16156 7252 16212 7262
rect 16156 2548 16212 7196
rect 16940 6778 16996 12302
rect 17724 12292 17780 12302
rect 17724 12226 17780 12236
rect 17612 12180 17668 12190
rect 17276 9268 17332 9278
rect 17276 9044 17332 9212
rect 17276 8978 17332 8988
rect 16380 6722 16996 6778
rect 17500 8596 17556 8606
rect 16268 5908 16324 5918
rect 16268 4340 16324 5852
rect 16268 4274 16324 4284
rect 16380 4004 16436 6722
rect 16940 6468 16996 6478
rect 16604 6412 16940 6418
rect 16604 6362 16996 6412
rect 16604 6356 16660 6362
rect 16604 6290 16660 6300
rect 17052 6356 17108 6366
rect 17052 5698 17108 6300
rect 17500 6132 17556 8540
rect 17612 7476 17668 12124
rect 17948 12122 18788 12178
rect 17948 11956 18004 12122
rect 17948 11890 18004 11900
rect 18060 11956 18676 11998
rect 18060 11942 18620 11956
rect 18060 11844 18116 11942
rect 18620 11890 18676 11900
rect 18060 11778 18116 11788
rect 18732 11844 18788 12122
rect 18732 11778 18788 11788
rect 18508 11732 18564 11742
rect 17724 11396 17780 11406
rect 17724 10164 17780 11340
rect 18508 11098 18564 11676
rect 18508 11042 19124 11098
rect 19068 10948 19124 11042
rect 19068 10882 19124 10892
rect 17724 10098 17780 10108
rect 19068 10164 19124 10174
rect 19068 9940 19124 10108
rect 19068 9874 19124 9884
rect 17612 7410 17668 7420
rect 18508 9380 18564 9390
rect 18508 7318 18564 9324
rect 19292 9044 19348 12572
rect 19740 12404 19796 12414
rect 19404 12348 19740 12358
rect 19404 12302 19796 12348
rect 19404 12292 19460 12302
rect 19404 12226 19460 12236
rect 20748 12292 20804 13244
rect 20748 12226 20804 12236
rect 20524 12180 20580 12190
rect 20524 11998 20580 12124
rect 20076 11942 20580 11998
rect 20076 10164 20132 11942
rect 20188 11844 20244 11854
rect 20188 11508 20244 11788
rect 20188 11442 20244 11452
rect 20300 11732 20356 11742
rect 20076 10098 20132 10108
rect 20300 10164 20356 11676
rect 21420 11396 21476 13916
rect 22876 13972 22932 13982
rect 21420 11330 21476 11340
rect 21868 13412 21924 13422
rect 21868 10836 21924 13356
rect 21868 10770 21924 10780
rect 22204 13412 22260 13422
rect 21532 10500 21588 10510
rect 21532 10198 21588 10444
rect 20300 10098 20356 10108
rect 20412 10142 21588 10198
rect 20412 9118 20468 10142
rect 19292 8978 19348 8988
rect 19964 9062 20468 9118
rect 20972 9828 21028 9838
rect 19964 8820 20020 9062
rect 19964 8754 20020 8764
rect 20188 8820 20244 8830
rect 20076 8708 20132 8718
rect 20076 7812 20132 8652
rect 20076 7746 20132 7756
rect 19404 7588 19460 7598
rect 19404 7498 19460 7532
rect 19404 7476 20132 7498
rect 19404 7442 20076 7476
rect 20076 7410 20132 7420
rect 20188 7318 20244 8764
rect 17500 6066 17556 6076
rect 18396 7262 18564 7318
rect 19852 7262 20244 7318
rect 20412 8708 20468 8718
rect 16716 5642 17108 5698
rect 16716 5572 16772 5642
rect 16716 5506 16772 5516
rect 17836 5460 17892 5470
rect 17836 5124 17892 5404
rect 17836 5058 17892 5068
rect 16492 5012 16548 5022
rect 16492 4340 16548 4956
rect 16492 4274 16548 4284
rect 16380 3938 16436 3948
rect 17612 4004 17668 4014
rect 16828 3780 16884 3790
rect 16828 3718 16884 3724
rect 16156 2482 16212 2492
rect 16716 3662 16884 3718
rect 16716 2212 16772 3662
rect 17052 3556 17108 3566
rect 17108 3500 17220 3538
rect 17052 3482 17220 3500
rect 16940 3220 16996 3230
rect 16996 3164 17108 3178
rect 16940 3122 17108 3164
rect 17052 2884 17108 3122
rect 17164 3108 17220 3482
rect 17612 3444 17668 3948
rect 17612 3378 17668 3388
rect 17164 3042 17220 3052
rect 17052 2818 17108 2828
rect 18396 2772 18452 7262
rect 18396 2706 18452 2716
rect 18508 7028 18564 7038
rect 18508 2278 18564 6972
rect 19852 7028 19908 7262
rect 19852 6962 19908 6972
rect 20076 7028 20132 7038
rect 19404 6916 19460 6926
rect 18732 5124 18788 5134
rect 18732 4788 18788 5068
rect 18732 4722 18788 4732
rect 18956 5124 19012 5134
rect 18956 3718 19012 5068
rect 18844 3662 19012 3718
rect 18844 3556 18900 3662
rect 18844 3490 18900 3500
rect 19292 3444 19348 3454
rect 16716 2146 16772 2156
rect 17948 2222 18564 2278
rect 18620 3332 18676 3342
rect 17948 1428 18004 2222
rect 18620 2212 18676 3276
rect 19292 3220 19348 3388
rect 19292 3154 19348 3164
rect 18620 2146 18676 2156
rect 18732 2772 18788 2782
rect 18060 1988 18116 1998
rect 18060 1918 18116 1932
rect 18732 1918 18788 2716
rect 18060 1862 18788 1918
rect 19404 1876 19460 6860
rect 20076 4340 20132 6972
rect 20076 4274 20132 4284
rect 19404 1810 19460 1820
rect 20300 2548 20356 2558
rect 17948 1362 18004 1372
rect 15596 1138 15652 1148
rect 20300 1204 20356 2492
rect 20300 1138 20356 1148
rect 20412 756 20468 8652
rect 20972 6692 21028 9772
rect 21868 9716 21924 9726
rect 21868 9658 21924 9660
rect 21868 9602 22148 9658
rect 21532 9492 21588 9502
rect 21532 8578 21588 9436
rect 22092 9268 22148 9602
rect 22092 9202 22148 9212
rect 22204 9118 22260 13356
rect 22316 11956 22372 11966
rect 22316 11818 22372 11900
rect 22316 11762 22596 11818
rect 22540 11732 22596 11762
rect 22540 11666 22596 11676
rect 22428 10836 22484 10846
rect 22428 10738 22484 10780
rect 22428 10682 22820 10738
rect 22652 9828 22708 9838
rect 22204 9062 22596 9118
rect 22428 8938 22484 8942
rect 21868 8932 22484 8938
rect 21868 8882 22428 8932
rect 21868 8820 21924 8882
rect 22428 8866 22484 8876
rect 21868 8754 21924 8764
rect 22540 8758 22596 9062
rect 22204 8702 22596 8758
rect 21532 8522 21924 8578
rect 21868 8036 21924 8522
rect 21868 7970 21924 7980
rect 20972 6626 21028 6636
rect 20636 5684 20692 5694
rect 20636 868 20692 5628
rect 21308 5684 21812 5698
rect 21308 5642 21756 5684
rect 21308 5572 21364 5642
rect 21756 5618 21812 5628
rect 21308 5506 21364 5516
rect 21196 4116 21252 4126
rect 21196 3892 21252 4060
rect 21196 3826 21252 3836
rect 22204 2884 22260 8702
rect 22204 2818 22260 2828
rect 22316 7588 22372 7598
rect 20636 802 20692 812
rect 20412 690 20468 700
rect 15372 578 15428 588
rect 8316 354 8372 364
rect 22316 420 22372 7532
rect 22428 3332 22484 3342
rect 22428 2884 22484 3276
rect 22428 2818 22484 2828
rect 22316 354 22372 364
rect 22652 308 22708 9772
rect 22764 7140 22820 10682
rect 22876 7588 22932 13916
rect 23660 13188 23716 13198
rect 23436 12292 23492 12302
rect 22988 11284 23044 11294
rect 22988 9492 23044 11228
rect 23100 11060 23156 11070
rect 23100 10500 23156 11004
rect 23100 10434 23156 10444
rect 23436 10276 23492 12236
rect 23436 10210 23492 10220
rect 23660 10276 23716 13132
rect 23660 10210 23716 10220
rect 23776 12572 24096 14224
rect 24220 13412 24276 13422
rect 24220 13188 24276 13356
rect 24220 13122 24276 13132
rect 24436 13356 24756 14224
rect 26684 14084 26740 14094
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 24220 12628 24276 12638
rect 24220 11732 24276 12572
rect 24220 11666 24276 11676
rect 24436 11788 24756 13300
rect 24892 13636 24948 13646
rect 24892 13300 24948 13580
rect 24892 13234 24948 13244
rect 25116 13636 25172 13646
rect 24892 12404 24948 12414
rect 24892 11956 24948 12348
rect 24892 11890 24948 11900
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 25116 11844 25172 13580
rect 26460 13412 26516 13422
rect 26460 12898 26516 13356
rect 26684 13258 26740 14028
rect 32060 14084 32116 14094
rect 29372 13860 29428 13870
rect 26908 13300 26964 13310
rect 26684 13244 26908 13258
rect 26684 13202 26964 13244
rect 28252 12964 28308 12974
rect 25116 11778 25172 11788
rect 25340 12852 25396 12862
rect 26460 12842 27076 12898
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 22988 9426 23044 9436
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23100 8932 23156 8942
rect 23100 8596 23156 8876
rect 23100 8530 23156 8540
rect 22876 7522 22932 7532
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 22764 7074 22820 7084
rect 23212 6804 23268 6814
rect 22764 6748 23212 6778
rect 22764 6722 23268 6748
rect 22764 6692 22820 6722
rect 22764 6626 22820 6636
rect 23776 6300 24096 7812
rect 24220 10836 24276 10846
rect 24220 7812 24276 10780
rect 24220 7746 24276 7756
rect 24436 10220 24756 11732
rect 24892 11732 24948 11742
rect 24892 11060 24948 11676
rect 24892 10994 24948 11004
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 24436 7084 24756 8596
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 23436 5460 23492 5470
rect 22988 5124 23044 5134
rect 22988 658 23044 5068
rect 23436 2660 23492 5404
rect 23776 4732 24096 6244
rect 24220 6244 24276 6254
rect 24220 6020 24276 6188
rect 24220 5954 24276 5964
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23660 4228 23716 4238
rect 23548 3332 23604 3342
rect 23548 3108 23604 3276
rect 23548 3042 23604 3052
rect 23436 2594 23492 2604
rect 23660 2324 23716 4172
rect 23660 2258 23716 2268
rect 23776 3164 24096 4676
rect 24436 5516 24756 7028
rect 25228 9380 25284 9390
rect 25228 6418 25284 9324
rect 25340 7924 25396 12796
rect 26348 12068 26404 12078
rect 26348 11818 26404 12012
rect 26796 11956 26852 11966
rect 26348 11762 26628 11818
rect 26348 11284 26404 11294
rect 25340 7858 25396 7868
rect 25564 8820 25620 8830
rect 25004 6362 25284 6418
rect 25452 6468 25508 6478
rect 25004 6244 25060 6362
rect 25004 6178 25060 6188
rect 25228 6244 25284 6254
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 24892 5796 24948 5806
rect 24892 5460 24948 5740
rect 24892 5394 24948 5404
rect 25004 5572 25060 5582
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 24220 3892 24276 3902
rect 24220 1652 24276 3836
rect 24220 1586 24276 1596
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 22988 602 23156 658
rect 23100 532 23156 602
rect 23100 466 23156 476
rect 22652 242 22708 252
rect 23776 0 24096 1540
rect 24436 812 24756 2324
rect 24892 4452 24948 4462
rect 24892 1540 24948 4396
rect 24892 1474 24948 1484
rect 25004 1204 25060 5516
rect 25116 5348 25172 5358
rect 25116 5124 25172 5292
rect 25116 5058 25172 5068
rect 25228 5012 25284 6188
rect 25228 4946 25284 4956
rect 25228 3892 25284 3902
rect 25228 3668 25284 3836
rect 25228 3602 25284 3612
rect 25452 3358 25508 6412
rect 25564 4340 25620 8764
rect 25564 4274 25620 4284
rect 25676 8260 25732 8270
rect 25452 3332 25620 3358
rect 25452 3302 25564 3332
rect 25564 3266 25620 3276
rect 25676 2324 25732 8204
rect 25900 4676 25956 4686
rect 25900 4340 25956 4620
rect 25900 4274 25956 4284
rect 26348 4116 26404 11228
rect 26572 10052 26628 11762
rect 26796 10948 26852 11900
rect 26796 10882 26852 10892
rect 27020 10948 27076 12842
rect 28252 12068 28308 12908
rect 28252 12002 28308 12012
rect 28476 12068 28532 12078
rect 28476 11732 28532 12012
rect 28476 11666 28532 11676
rect 27356 11508 27412 11518
rect 27356 11284 27412 11452
rect 27356 11218 27412 11228
rect 27020 10882 27076 10892
rect 28252 11172 28308 11182
rect 28252 10836 28308 11116
rect 28252 10770 28308 10780
rect 26684 10612 26740 10622
rect 26684 10276 26740 10556
rect 26684 10210 26740 10220
rect 26908 10612 26964 10622
rect 26572 9986 26628 9996
rect 26908 8932 26964 10556
rect 28476 10276 28532 10286
rect 28476 9044 28532 10220
rect 28476 8978 28532 8988
rect 28924 10164 28980 10174
rect 26908 8866 26964 8876
rect 26572 7588 26628 7598
rect 26460 5572 26516 5582
rect 26460 4228 26516 5516
rect 26572 5124 26628 7532
rect 28924 7588 28980 10108
rect 28924 7522 28980 7532
rect 28476 7364 28532 7374
rect 27020 7252 27076 7262
rect 26684 7140 26740 7150
rect 27020 7138 27076 7196
rect 26740 7084 27076 7138
rect 26684 7082 27076 7084
rect 28140 7252 28196 7262
rect 26684 7074 26740 7082
rect 28140 6244 28196 7196
rect 28140 6178 28196 6188
rect 28252 7028 28308 7038
rect 27020 5908 27076 5918
rect 28252 5908 28308 6972
rect 28476 7028 28532 7308
rect 28476 6962 28532 6972
rect 27076 5852 27860 5878
rect 27020 5822 27860 5852
rect 28252 5842 28308 5852
rect 27804 5236 27860 5822
rect 27804 5170 27860 5180
rect 26572 5058 26628 5068
rect 28588 5124 28644 5134
rect 28588 4978 28644 5068
rect 26852 4922 28644 4978
rect 26852 4900 26908 4922
rect 26852 4834 26908 4844
rect 29148 4788 29204 4798
rect 26908 4676 26964 4686
rect 26796 4452 26852 4462
rect 26908 4438 26964 4620
rect 26852 4396 26964 4438
rect 26796 4382 26964 4396
rect 26460 4162 26516 4172
rect 26348 4050 26404 4060
rect 27020 4116 27076 4126
rect 27020 3718 27076 4060
rect 26572 3662 27076 3718
rect 28700 3668 28756 3678
rect 26572 3556 26628 3662
rect 26572 3490 26628 3500
rect 26796 3220 26852 3230
rect 27020 3220 27076 3230
rect 26852 3164 27020 3178
rect 26796 3122 27076 3164
rect 25788 3108 25844 3118
rect 25788 2998 25844 3052
rect 25788 2942 26964 2998
rect 26908 2884 26964 2942
rect 26908 2818 26964 2828
rect 25676 2258 25732 2268
rect 26236 2772 26292 2782
rect 26236 2212 26292 2716
rect 26236 2146 26292 2156
rect 28588 2436 28644 2446
rect 28588 2212 28644 2380
rect 28588 2146 28644 2156
rect 28700 1558 28756 3612
rect 29148 2212 29204 4732
rect 29372 3780 29428 13804
rect 32060 13412 32116 14028
rect 32060 13346 32116 13356
rect 32732 13524 32788 13534
rect 30940 13300 30996 13310
rect 30940 12852 30996 13244
rect 31164 13076 31220 13086
rect 31164 12898 31220 13020
rect 32732 12964 32788 13468
rect 33852 13412 33908 13422
rect 32732 12898 32788 12908
rect 33628 13076 33684 13086
rect 30940 12786 30996 12796
rect 31052 12842 31220 12898
rect 30604 12740 30660 12750
rect 31052 12718 31108 12842
rect 30660 12684 31108 12718
rect 30604 12662 31108 12684
rect 31948 12404 32004 12414
rect 29932 11172 29988 11182
rect 29932 10612 29988 11116
rect 29932 10546 29988 10556
rect 31500 10948 31556 10958
rect 30940 9940 30996 9950
rect 30940 8820 30996 9884
rect 31500 9380 31556 10892
rect 31500 9314 31556 9324
rect 31724 9828 31780 9838
rect 30940 8754 30996 8764
rect 31724 7252 31780 9772
rect 31948 7700 32004 12348
rect 33516 10500 33572 10510
rect 33292 8820 33348 8830
rect 33292 8758 33348 8764
rect 33292 8702 33460 8758
rect 33404 8596 33460 8702
rect 33404 8530 33460 8540
rect 33516 7924 33572 10444
rect 33516 7858 33572 7868
rect 31948 7634 32004 7644
rect 31724 7186 31780 7196
rect 29708 6692 29764 6702
rect 29708 6356 29764 6636
rect 29708 6290 29764 6300
rect 29932 6244 29988 6254
rect 29372 3714 29428 3724
rect 29596 5012 29652 5022
rect 29148 2146 29204 2156
rect 29596 1988 29652 4956
rect 29932 2884 29988 6188
rect 33628 5158 33684 13020
rect 33852 12740 33908 13356
rect 33852 12674 33908 12684
rect 39564 12964 39620 12974
rect 33964 12404 34020 12414
rect 33964 12068 34020 12348
rect 39564 12404 39620 12908
rect 39564 12338 39620 12348
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 33964 12002 34020 12012
rect 39116 12068 39172 12078
rect 35532 11620 35588 11630
rect 33404 5124 33684 5158
rect 33460 5102 33684 5124
rect 34188 10948 34244 10958
rect 33404 5058 33460 5068
rect 29932 2818 29988 2828
rect 30380 4116 30436 4126
rect 29596 1922 29652 1932
rect 28588 1502 28756 1558
rect 28588 1428 28644 1502
rect 28588 1362 28644 1372
rect 25004 1138 25060 1148
rect 30380 980 30436 4060
rect 32620 2100 32676 2110
rect 32676 2044 32788 2098
rect 32620 2042 32788 2044
rect 32620 2034 32676 2042
rect 32732 1876 32788 2042
rect 32732 1810 32788 1820
rect 30380 914 30436 924
rect 31052 1540 31108 1550
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 25228 644 25284 654
rect 25228 196 25284 588
rect 25228 130 25284 140
rect 31052 84 31108 1484
rect 33740 1204 33796 1214
rect 33740 868 33796 1148
rect 33740 802 33796 812
rect 34188 308 34244 10892
rect 34860 8708 34916 8718
rect 34860 2100 34916 8652
rect 35532 5908 35588 11564
rect 37212 9268 37268 9278
rect 37212 8932 37268 9212
rect 37212 8866 37268 8876
rect 38444 8596 38500 8606
rect 38500 8540 38612 8578
rect 38444 8522 38612 8540
rect 38556 7028 38612 8522
rect 38556 6962 38612 6972
rect 35532 5842 35588 5852
rect 39116 2212 39172 12012
rect 41804 11620 41860 11630
rect 39228 10388 39284 10398
rect 39228 7252 39284 10332
rect 39228 7186 39284 7196
rect 39116 2146 39172 2156
rect 34860 2034 34916 2044
rect 41804 420 41860 11564
rect 41804 354 41860 364
rect 43776 11004 44096 12516
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 43776 9436 44096 10948
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 43776 6300 44096 7812
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 43776 4732 44096 6244
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 43776 3164 44096 4676
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 34188 242 34244 252
rect 31052 18 31108 28
rect 43776 0 44096 1540
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44436 3948 44756 5460
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 38528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 37632 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 5712 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 5712 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 45248 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 29232 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 47600 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 36064 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 46816 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 43792 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 27776 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 47600 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 32704 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 17024 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 44576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 34384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 50624 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 30464 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 26208 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 38976 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 1456 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 10528 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 13776 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 32816 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 26320 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 38752 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 24192 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 25088 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 45696 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 24752 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 50624 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 44688 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform 1 0 46256 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 48496 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 29232 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 29232 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform 1 0 24752 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 13552 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 6048 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 8400 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 19152 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 30128 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform 1 0 13104 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 3360 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 6720 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 2352 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 5712 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 25312 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 17808 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 25312 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 22960 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform -1 0 10304 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform 1 0 26544 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 29120 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform -1 0 22624 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform -1 0 21056 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform -1 0 19712 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 42448 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 47936 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 47600 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 49392 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform -1 0 19488 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform -1 0 17584 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 42112 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform -1 0 24080 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform -1 0 24528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform -1 0 28000 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 27104 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 38752 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 26992 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform 1 0 49168 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform 1 0 38416 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform 1 0 46592 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 6496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 44464 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 10080 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 41664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 7504 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform -1 0 2576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 21728 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 43680 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 11536 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 15008 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 9744 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 23296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 36960 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 37856 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 15568 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 20496 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 10864 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 20944 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 4592 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 9632 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform 1 0 12320 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 23520 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 9184 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 12432 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 25312 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 11200 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform 1 0 32480 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform 1 0 27216 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__000__I
timestamp 1486834041
transform 1 0 38304 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__001__I
timestamp 1486834041
transform -1 0 37632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I
timestamp 1486834041
transform 1 0 5488 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1486834041
transform 1 0 5488 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__I
timestamp 1486834041
transform -1 0 45248 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__I
timestamp 1486834041
transform 1 0 29008 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__006__I
timestamp 1486834041
transform 1 0 31808 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__007__I
timestamp 1486834041
transform -1 0 47600 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__008__I
timestamp 1486834041
transform 1 0 35840 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__009__I
timestamp 1486834041
transform -1 0 46816 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__010__I
timestamp 1486834041
transform 1 0 43568 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__011__I
timestamp 1486834041
transform 1 0 27552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__012__I
timestamp 1486834041
transform -1 0 47600 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__013__I
timestamp 1486834041
transform -1 0 32704 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__014__I
timestamp 1486834041
transform 1 0 16800 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__015__I
timestamp 1486834041
transform -1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__016__I
timestamp 1486834041
transform -1 0 44576 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__017__I
timestamp 1486834041
transform 1 0 34160 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__018__I
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__019__I
timestamp 1486834041
transform -1 0 30464 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__020__I
timestamp 1486834041
transform -1 0 26208 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__021__I
timestamp 1486834041
transform -1 0 38976 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__022__I
timestamp 1486834041
transform 1 0 1232 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__023__I
timestamp 1486834041
transform -1 0 10528 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__024__I
timestamp 1486834041
transform -1 0 13776 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__025__I
timestamp 1486834041
transform -1 0 32816 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__026__I
timestamp 1486834041
transform 1 0 26096 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__027__I
timestamp 1486834041
transform -1 0 38752 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__028__I
timestamp 1486834041
transform 1 0 23744 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__029__I
timestamp 1486834041
transform 1 0 23968 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I
timestamp 1486834041
transform -1 0 45696 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__I
timestamp 1486834041
transform -1 0 24752 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__032__I
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__I
timestamp 1486834041
transform 1 0 44464 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__I
timestamp 1486834041
transform -1 0 46256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__I
timestamp 1486834041
transform 1 0 48272 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__I
timestamp 1486834041
transform -1 0 29232 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__I
timestamp 1486834041
transform 1 0 29008 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__I
timestamp 1486834041
transform 1 0 24528 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__I
timestamp 1486834041
transform -1 0 13776 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__I
timestamp 1486834041
transform 1 0 6048 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__041__I
timestamp 1486834041
transform -1 0 8624 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I
timestamp 1486834041
transform -1 0 19376 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1486834041
transform 1 0 30128 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I
timestamp 1486834041
transform -1 0 13104 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1486834041
transform -1 0 3584 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1486834041
transform 1 0 6720 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1486834041
transform -1 0 2576 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I
timestamp 1486834041
transform -1 0 6832 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I
timestamp 1486834041
transform 1 0 25312 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1486834041
transform 1 0 17808 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1486834041
transform 1 0 22960 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1486834041
transform -1 0 10528 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1486834041
transform 1 0 26320 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1486834041
transform -1 0 29120 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1486834041
transform -1 0 22848 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1486834041
transform 1 0 21056 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1486834041
transform -1 0 19936 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1486834041
transform 1 0 42224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1486834041
transform 1 0 47712 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1486834041
transform 1 0 47376 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1486834041
transform -1 0 48272 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1486834041
transform -1 0 19712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1486834041
transform 1 0 17584 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1486834041
transform 1 0 41888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1486834041
transform 1 0 43568 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1486834041
transform 1 0 24528 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1486834041
transform 1 0 28000 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1486834041
transform 1 0 26880 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1486834041
transform 1 0 38528 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1486834041
transform -1 0 27216 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1486834041
transform 1 0 48944 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1486834041
transform 1 0 38192 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1486834041
transform -1 0 46592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1486834041
transform 1 0 6496 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1486834041
transform -1 0 44464 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1486834041
transform -1 0 10304 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1486834041
transform -1 0 41664 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1486834041
transform -1 0 7728 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1486834041
transform -1 0 2800 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1486834041
transform -1 0 21952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1486834041
transform -1 0 43680 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1486834041
transform -1 0 11760 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I
timestamp 1486834041
transform -1 0 15232 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1486834041
transform -1 0 9968 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I
timestamp 1486834041
transform -1 0 23520 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1486834041
transform 1 0 36736 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1486834041
transform -1 0 37856 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1486834041
transform 1 0 15568 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1486834041
transform -1 0 20720 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1486834041
transform 1 0 10864 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1486834041
transform -1 0 21168 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1486834041
transform -1 0 9856 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1486834041
transform -1 0 12320 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1486834041
transform -1 0 23744 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1486834041
transform 1 0 9184 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1486834041
transform -1 0 25536 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1486834041
transform 1 0 11200 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1486834041
transform -1 0 7168 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1486834041
transform 1 0 32256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1486834041
transform 1 0 26992 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_184
timestamp 1486834041
transform 1 0 21280 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_200
timestamp 1486834041
transform 1 0 23072 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_454
timestamp 1486834041
transform 1 0 51520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_456
timestamp 1486834041
transform 1 0 51744 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_88
timestamp 1486834041
transform 1 0 10528 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_96
timestamp 1486834041
transform 1 0 11424 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_99
timestamp 1486834041
transform 1 0 11760 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_125
timestamp 1486834041
transform 1 0 14672 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_133
timestamp 1486834041
transform 1 0 15568 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1486834041
transform 1 0 16016 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_158
timestamp 1486834041
transform 1 0 18368 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_172
timestamp 1486834041
transform 1 0 19936 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_183
timestamp 1486834041
transform 1 0 21168 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_199
timestamp 1486834041
transform 1 0 22960 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1486834041
transform 1 0 23856 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 24080 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_276
timestamp 1486834041
transform 1 0 31584 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_294
timestamp 1486834041
transform 1 0 33600 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_326
timestamp 1486834041
transform 1 0 37184 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_334
timestamp 1486834041
transform 1 0 38080 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_338
timestamp 1486834041
transform 1 0 38528 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_368
timestamp 1486834041
transform 1 0 41888 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_376
timestamp 1486834041
transform 1 0 42784 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_380
timestamp 1486834041
transform 1 0 43232 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_392
timestamp 1486834041
transform 1 0 44576 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_408
timestamp 1486834041
transform 1 0 46368 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_426
timestamp 1486834041
transform 1 0 48384 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1486834041
transform 1 0 48608 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_4
timestamp 1486834041
transform 1 0 1120 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_15
timestamp 1486834041
transform 1 0 2352 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_23
timestamp 1486834041
transform 1 0 3248 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_39
timestamp 1486834041
transform 1 0 5040 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_71
timestamp 1486834041
transform 1 0 8624 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_87
timestamp 1486834041
transform 1 0 10416 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_109
timestamp 1486834041
transform 1 0 12880 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_141
timestamp 1486834041
transform 1 0 16464 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_153
timestamp 1486834041
transform 1 0 17808 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_169
timestamp 1486834041
transform 1 0 19600 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_173
timestamp 1486834041
transform 1 0 20048 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 27664 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_247
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1486834041
transform 1 0 35504 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1486834041
transform 1 0 36624 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_332
timestamp 1486834041
transform 1 0 37856 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_336
timestamp 1486834041
transform 1 0 38304 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_348
timestamp 1486834041
transform 1 0 39648 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_380
timestamp 1486834041
transform 1 0 43232 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_384
timestamp 1486834041
transform 1 0 43680 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_395
timestamp 1486834041
transform 1 0 44912 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_406
timestamp 1486834041
transform 1 0 46144 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_410
timestamp 1486834041
transform 1 0 46592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_412
timestamp 1486834041
transform 1 0 46816 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_6
timestamp 1486834041
transform 1 0 1344 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_8
timestamp 1486834041
transform 1 0 1568 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_19
timestamp 1486834041
transform 1 0 2800 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_51
timestamp 1486834041
transform 1 0 6384 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_67
timestamp 1486834041
transform 1 0 8176 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_69
timestamp 1486834041
transform 1 0 8400 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_158
timestamp 1486834041
transform 1 0 18368 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_166
timestamp 1486834041
transform 1 0 19264 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_168
timestamp 1486834041
transform 1 0 19488 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_179
timestamp 1486834041
transform 1 0 20720 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_195
timestamp 1486834041
transform 1 0 22512 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_203
timestamp 1486834041
transform 1 0 23408 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_207
timestamp 1486834041
transform 1 0 23856 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_222
timestamp 1486834041
transform 1 0 25536 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_230
timestamp 1486834041
transform 1 0 26432 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_234
timestamp 1486834041
transform 1 0 26880 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_246
timestamp 1486834041
transform 1 0 28224 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_250
timestamp 1486834041
transform 1 0 28672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_262
timestamp 1486834041
transform 1 0 30016 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_278
timestamp 1486834041
transform 1 0 31808 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1486834041
transform 1 0 32256 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_284
timestamp 1486834041
transform 1 0 32480 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_295
timestamp 1486834041
transform 1 0 33712 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_327
timestamp 1486834041
transform 1 0 37296 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_343
timestamp 1486834041
transform 1 0 39088 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_347
timestamp 1486834041
transform 1 0 39536 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 39760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_384
timestamp 1486834041
transform 1 0 43680 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_388
timestamp 1486834041
transform 1 0 44128 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_418
timestamp 1486834041
transform 1 0 47488 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_426
timestamp 1486834041
transform 1 0 48384 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1486834041
transform 1 0 48608 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_77
timestamp 1486834041
transform 1 0 9296 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_81
timestamp 1486834041
transform 1 0 9744 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_93
timestamp 1486834041
transform 1 0 11088 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 11984 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_123
timestamp 1486834041
transform 1 0 14448 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_135
timestamp 1486834041
transform 1 0 15792 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_167
timestamp 1486834041
transform 1 0 19376 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_209
timestamp 1486834041
transform 1 0 24080 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_225
timestamp 1486834041
transform 1 0 25872 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_237
timestamp 1486834041
transform 1 0 27216 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_279
timestamp 1486834041
transform 1 0 31920 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_281
timestamp 1486834041
transform 1 0 32144 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_292
timestamp 1486834041
transform 1 0 33376 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_308
timestamp 1486834041
transform 1 0 35168 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_312
timestamp 1486834041
transform 1 0 35616 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_314
timestamp 1486834041
transform 1 0 35840 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_317
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_349
timestamp 1486834041
transform 1 0 39760 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_365
timestamp 1486834041
transform 1 0 41552 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_367
timestamp 1486834041
transform 1 0 41776 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_378
timestamp 1486834041
transform 1 0 43008 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_382
timestamp 1486834041
transform 1 0 43456 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_395
timestamp 1486834041
transform 1 0 44912 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_403
timestamp 1486834041
transform 1 0 45808 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_415
timestamp 1486834041
transform 1 0 47152 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_34
timestamp 1486834041
transform 1 0 4480 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_42
timestamp 1486834041
transform 1 0 5376 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_45
timestamp 1486834041
transform 1 0 5712 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_56
timestamp 1486834041
transform 1 0 6944 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_64
timestamp 1486834041
transform 1 0 7840 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1486834041
transform 1 0 8288 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_80
timestamp 1486834041
transform 1 0 9632 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_84
timestamp 1486834041
transform 1 0 10080 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_88
timestamp 1486834041
transform 1 0 10528 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_130
timestamp 1486834041
transform 1 0 15232 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_138
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1486834041
transform 1 0 16800 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_155
timestamp 1486834041
transform 1 0 18032 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_187
timestamp 1486834041
transform 1 0 21616 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_191
timestamp 1486834041
transform 1 0 22064 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_193
timestamp 1486834041
transform 1 0 22288 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_204
timestamp 1486834041
transform 1 0 23520 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_208
timestamp 1486834041
transform 1 0 23968 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_223
timestamp 1486834041
transform 1 0 25648 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_255
timestamp 1486834041
transform 1 0 29232 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_271
timestamp 1486834041
transform 1 0 31024 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 31920 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_314
timestamp 1486834041
transform 1 0 35840 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_330
timestamp 1486834041
transform 1 0 37632 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_334
timestamp 1486834041
transform 1 0 38080 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_348
timestamp 1486834041
transform 1 0 39648 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 47264 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_426
timestamp 1486834041
transform 1 0 48384 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1486834041
transform 1 0 48608 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_55
timestamp 1486834041
transform 1 0 6832 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_71
timestamp 1486834041
transform 1 0 8624 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_75
timestamp 1486834041
transform 1 0 9072 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_77
timestamp 1486834041
transform 1 0 9296 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_96
timestamp 1486834041
transform 1 0 11424 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_193
timestamp 1486834041
transform 1 0 22288 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_201
timestamp 1486834041
transform 1 0 23184 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_215
timestamp 1486834041
transform 1 0 24752 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_231
timestamp 1486834041
transform 1 0 26544 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_239
timestamp 1486834041
transform 1 0 27440 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_243
timestamp 1486834041
transform 1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_311
timestamp 1486834041
transform 1 0 35504 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_325
timestamp 1486834041
transform 1 0 37072 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_327
timestamp 1486834041
transform 1 0 37296 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_346
timestamp 1486834041
transform 1 0 39424 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_378
timestamp 1486834041
transform 1 0 43008 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_382
timestamp 1486834041
transform 1 0 43456 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 43680 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1486834041
transform 1 0 47600 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_430
timestamp 1486834041
transform 1 0 48832 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_34
timestamp 1486834041
transform 1 0 4480 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_42
timestamp 1486834041
transform 1 0 5376 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_53
timestamp 1486834041
transform 1 0 6608 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_69
timestamp 1486834041
transform 1 0 8400 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_83
timestamp 1486834041
transform 1 0 9968 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_115
timestamp 1486834041
transform 1 0 13552 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_131
timestamp 1486834041
transform 1 0 15344 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 16240 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_158
timestamp 1486834041
transform 1 0 18368 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_170
timestamp 1486834041
transform 1 0 19712 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_186
timestamp 1486834041
transform 1 0 21504 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_194
timestamp 1486834041
transform 1 0 22400 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_244
timestamp 1486834041
transform 1 0 28000 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_252
timestamp 1486834041
transform 1 0 28896 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_263
timestamp 1486834041
transform 1 0 30128 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_279
timestamp 1486834041
transform 1 0 31920 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_384
timestamp 1486834041
transform 1 0 43680 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_388
timestamp 1486834041
transform 1 0 44128 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_399
timestamp 1486834041
transform 1 0 45360 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_415
timestamp 1486834041
transform 1 0 47152 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1486834041
transform 1 0 47600 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_426
timestamp 1486834041
transform 1 0 48384 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1486834041
transform 1 0 48608 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 11984 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_135
timestamp 1486834041
transform 1 0 15792 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_151
timestamp 1486834041
transform 1 0 17584 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_167
timestamp 1486834041
transform 1 0 19376 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_185
timestamp 1486834041
transform 1 0 21392 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_187
timestamp 1486834041
transform 1 0 21616 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_190
timestamp 1486834041
transform 1 0 21952 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_198
timestamp 1486834041
transform 1 0 22848 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_200
timestamp 1486834041
transform 1 0 23072 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_211
timestamp 1486834041
transform 1 0 24304 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_243
timestamp 1486834041
transform 1 0 27888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_251
timestamp 1486834041
transform 1 0 28784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_263
timestamp 1486834041
transform 1 0 30128 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_295
timestamp 1486834041
transform 1 0 33712 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_311
timestamp 1486834041
transform 1 0 35504 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 8064 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_86
timestamp 1486834041
transform 1 0 10304 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_150
timestamp 1486834041
transform 1 0 17472 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_169
timestamp 1486834041
transform 1 0 19600 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_177
timestamp 1486834041
transform 1 0 20496 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_179
timestamp 1486834041
transform 1 0 20720 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_198
timestamp 1486834041
transform 1 0 22848 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 23744 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_223
timestamp 1486834041
transform 1 0 25648 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_265
timestamp 1486834041
transform 1 0 30352 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_273
timestamp 1486834041
transform 1 0 31248 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_277
timestamp 1486834041
transform 1 0 31696 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_290
timestamp 1486834041
transform 1 0 33152 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_322
timestamp 1486834041
transform 1 0 36736 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_338
timestamp 1486834041
transform 1 0 38528 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 39424 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 47264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_61
timestamp 1486834041
transform 1 0 7504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_65
timestamp 1486834041
transform 1 0 7952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_67
timestamp 1486834041
transform 1 0 8176 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_78
timestamp 1486834041
transform 1 0 9408 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_86
timestamp 1486834041
transform 1 0 10304 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_90
timestamp 1486834041
transform 1 0 10752 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_201
timestamp 1486834041
transform 1 0 23184 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_205
timestamp 1486834041
transform 1 0 23632 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_226
timestamp 1486834041
transform 1 0 25984 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_234
timestamp 1486834041
transform 1 0 26880 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_237
timestamp 1486834041
transform 1 0 27216 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_333
timestamp 1486834041
transform 1 0 37968 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_345
timestamp 1486834041
transform 1 0 39312 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_363
timestamp 1486834041
transform 1 0 41328 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_366
timestamp 1486834041
transform 1 0 41664 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_382
timestamp 1486834041
transform 1 0 43456 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_384
timestamp 1486834041
transform 1 0 43680 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_393
timestamp 1486834041
transform 1 0 44688 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_409
timestamp 1486834041
transform 1 0 46480 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 8064 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_82
timestamp 1486834041
transform 1 0 9856 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_96
timestamp 1486834041
transform 1 0 11424 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1486834041
transform 1 0 16800 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 24080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_222
timestamp 1486834041
transform 1 0 25536 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_226
timestamp 1486834041
transform 1 0 25984 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_243
timestamp 1486834041
transform 1 0 27888 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_275
timestamp 1486834041
transform 1 0 31472 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_298
timestamp 1486834041
transform 1 0 34048 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_309
timestamp 1486834041
transform 1 0 35280 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_313
timestamp 1486834041
transform 1 0 35728 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_324
timestamp 1486834041
transform 1 0 36960 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_332
timestamp 1486834041
transform 1 0 37856 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_334
timestamp 1486834041
transform 1 0 38080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_349
timestamp 1486834041
transform 1 0 39760 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_374
timestamp 1486834041
transform 1 0 42560 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_382
timestamp 1486834041
transform 1 0 43456 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_401
timestamp 1486834041
transform 1 0 45584 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_417
timestamp 1486834041
transform 1 0 47376 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_426
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1486834041
transform 1 0 48608 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_17
timestamp 1486834041
transform 1 0 2576 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1486834041
transform 1 0 4368 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_45
timestamp 1486834041
transform 1 0 5712 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_47
timestamp 1486834041
transform 1 0 5936 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_50
timestamp 1486834041
transform 1 0 6272 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_66
timestamp 1486834041
transform 1 0 8064 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_74
timestamp 1486834041
transform 1 0 8960 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_76
timestamp 1486834041
transform 1 0 9184 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_115
timestamp 1486834041
transform 1 0 13552 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_181
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_211
timestamp 1486834041
transform 1 0 24304 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_219
timestamp 1486834041
transform 1 0 25200 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_223
timestamp 1486834041
transform 1 0 25648 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_225
timestamp 1486834041
transform 1 0 25872 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_244
timestamp 1486834041
transform 1 0 28000 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 35504 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_381
timestamp 1486834041
transform 1 0 43344 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_403
timestamp 1486834041
transform 1 0 45808 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_411
timestamp 1486834041
transform 1 0 46704 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_415
timestamp 1486834041
transform 1 0 47152 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_34
timestamp 1486834041
transform 1 0 4480 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_38
timestamp 1486834041
transform 1 0 4928 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_58
timestamp 1486834041
transform 1 0 7168 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_60
timestamp 1486834041
transform 1 0 7392 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_63
timestamp 1486834041
transform 1 0 7728 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_67
timestamp 1486834041
transform 1 0 8176 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_69
timestamp 1486834041
transform 1 0 8400 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_222
timestamp 1486834041
transform 1 0 25536 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_230
timestamp 1486834041
transform 1 0 26432 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_236
timestamp 1486834041
transform 1 0 27104 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_250
timestamp 1486834041
transform 1 0 28672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_252
timestamp 1486834041
transform 1 0 28896 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_255
timestamp 1486834041
transform 1 0 29232 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_271
timestamp 1486834041
transform 1 0 31024 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 31920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_314
timestamp 1486834041
transform 1 0 35840 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_318
timestamp 1486834041
transform 1 0 36288 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_347
timestamp 1486834041
transform 1 0 39536 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_349
timestamp 1486834041
transform 1 0 39760 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_380
timestamp 1486834041
transform 1 0 43232 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_412
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_426
timestamp 1486834041
transform 1 0 48384 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1486834041
transform 1 0 48608 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_10
timestamp 1486834041
transform 1 0 1792 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_14
timestamp 1486834041
transform 1 0 2240 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_26
timestamp 1486834041
transform 1 0 3584 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 4480 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_41
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_43
timestamp 1486834041
transform 1 0 5488 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_52
timestamp 1486834041
transform 1 0 6496 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_71
timestamp 1486834041
transform 1 0 8624 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_75
timestamp 1486834041
transform 1 0 9072 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_117
timestamp 1486834041
transform 1 0 13776 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_219
timestamp 1486834041
transform 1 0 25200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_227
timestamp 1486834041
transform 1 0 26096 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_239
timestamp 1486834041
transform 1 0 27440 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_263
timestamp 1486834041
transform 1 0 30128 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_274
timestamp 1486834041
transform 1 0 31360 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_306
timestamp 1486834041
transform 1 0 34944 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_314
timestamp 1486834041
transform 1 0 35840 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_381
timestamp 1486834041
transform 1 0 43344 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_403
timestamp 1486834041
transform 1 0 45808 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_411
timestamp 1486834041
transform 1 0 46704 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_54
timestamp 1486834041
transform 1 0 6720 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_62
timestamp 1486834041
transform 1 0 7616 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_66
timestamp 1486834041
transform 1 0 8064 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_206
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_221
timestamp 1486834041
transform 1 0 25424 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_237
timestamp 1486834041
transform 1 0 27216 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_329
timestamp 1486834041
transform 1 0 37520 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_370
timestamp 1486834041
transform 1 0 42112 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_373
timestamp 1486834041
transform 1 0 42448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_404
timestamp 1486834041
transform 1 0 45920 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_454
timestamp 1486834041
transform 1 0 51520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_456
timestamp 1486834041
transform 1 0 51744 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 48496 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 48720 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 50064 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 50288 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 48720 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 50064 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 48496 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 50288 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 50288 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform -1 0 51632 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 46928 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 50288 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 50064 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 50288 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 50064 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 48720 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 48496 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 48608 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 47040 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 46928 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 47040 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 48720 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 48496 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 48608 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 48720 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 50288 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 48720 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 50064 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 48496 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 50288 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 37520 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 38192 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 40880 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 40208 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 41664 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 39760 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 41776 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 44352 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 37744 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 37968 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 39312 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 37072 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 37968 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 39312 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 40544 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 38640 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 12432 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 9296 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 14224 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 12432 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 14784 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 13216 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 15792 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 12432 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 16352 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 14784 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 15568 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 16352 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 15568 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 17136 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 14336 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 20272 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 20048 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 18704 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 17920 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 17136 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 16352 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 17136 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 19600 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 16912 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 17136 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 22064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 22736 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 22624 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 23632 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 23632 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 25424 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 21616 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 19488 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 21616 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 21168 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 21056 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform 1 0 35280 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 52080 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 52080 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 52080 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 52080 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 52080 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 52080 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 52080 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 52080 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 52080 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 52080 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 52080 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 52080 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 52080 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 52080 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 52080 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 52080 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_45
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_51
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_52
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_58
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_59
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_64
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_65
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_66
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_71
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_72
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_73
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_77
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_78
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_79
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_80
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_84
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_91
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_92
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_93
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_94
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_97
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_98
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_99
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_100
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_101
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_103
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_104
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_105
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_106
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_107
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_108
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_110
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_111
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_112
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_113
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_114
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_115
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_116
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_117
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_118
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_119
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_120
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_121
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_122
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_123
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_124
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_125
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_126
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_127
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_128
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_129
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_130
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_131
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_132
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_133
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_136
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_137
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_140
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_141
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_142
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_143
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 52640 0 52752 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 52640 4480 52752 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 52640 4928 52752 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 52640 5376 52752 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 52640 5824 52752 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 52640 6272 52752 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 52640 6720 52752 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 52640 7168 52752 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 52640 7616 52752 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 52640 8064 52752 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 52640 8512 52752 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 52640 448 52752 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 52640 8960 52752 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 52640 9408 52752 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 52640 9856 52752 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 52640 10304 52752 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 52640 10752 52752 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 52640 11200 52752 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 52640 11648 52752 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 52640 12096 52752 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 52640 12544 52752 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 52640 12992 52752 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 52640 896 52752 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 52640 13440 52752 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 52640 13888 52752 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 52640 1344 52752 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 52640 1792 52752 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 52640 2240 52752 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 52640 2688 52752 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 52640 3136 52752 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 52640 3584 52752 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 52640 4032 52752 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 4032 0 4144 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 28672 0 28784 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 31136 0 31248 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 33600 0 33712 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 36064 0 36176 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 38528 0 38640 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 40992 0 41104 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 43456 0 43568 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 45920 0 46032 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 48384 0 48496 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 50848 0 50960 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 6496 0 6608 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 8960 0 9072 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 13888 0 14000 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 16352 0 16464 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 18816 0 18928 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 21280 0 21392 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 23744 0 23856 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 35840 14112 35952 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 38080 14112 38192 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 38528 14112 38640 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 38976 14112 39088 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 39424 14112 39536 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 39872 14112 39984 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 36288 14112 36400 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 36736 14112 36848 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 37184 14112 37296 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 37632 14112 37744 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 12544 14112 12656 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 12992 14112 13104 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 13440 14112 13552 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 13888 14112 14000 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 14336 14112 14448 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 14784 14112 14896 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 15232 14112 15344 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 15680 14112 15792 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 16128 14112 16240 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 16576 14112 16688 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 19264 14112 19376 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 19712 14112 19824 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 20160 14112 20272 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 17024 14112 17136 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 17472 14112 17584 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 17920 14112 18032 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 18368 14112 18480 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 18816 14112 18928 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 22848 14112 22960 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 23296 14112 23408 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 23744 14112 23856 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 20608 14112 20720 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 21056 14112 21168 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 21504 14112 21616 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 21952 14112 22064 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 22400 14112 22512 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 24192 14112 24304 14224 0 FreeSans 448 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 24640 14112 24752 14224 0 FreeSans 448 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 26880 14112 26992 14224 0 FreeSans 448 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 27328 14112 27440 14224 0 FreeSans 448 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 27776 14112 27888 14224 0 FreeSans 448 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 28224 14112 28336 14224 0 FreeSans 448 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 25088 14112 25200 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 25536 14112 25648 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 25984 14112 26096 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 26432 14112 26544 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 30912 14112 31024 14224 0 FreeSans 448 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 31360 14112 31472 14224 0 FreeSans 448 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 31808 14112 31920 14224 0 FreeSans 448 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 28672 14112 28784 14224 0 FreeSans 448 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 29120 14112 29232 14224 0 FreeSans 448 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 29568 14112 29680 14224 0 FreeSans 448 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 30016 14112 30128 14224 0 FreeSans 448 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 30464 14112 30576 14224 0 FreeSans 448 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 34496 14112 34608 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 34944 14112 35056 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 35392 14112 35504 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 32256 14112 32368 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 32704 14112 32816 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 33152 14112 33264 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 33600 14112 33712 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 34048 14112 34160 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1568 0 1680 112 0 FreeSans 448 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 26376 12544 26376 12544 0 VDD
rlabel metal1 26376 13328 26376 13328 0 VSS
rlabel metal3 2646 56 2646 56 0 FrameData[0]
rlabel metal2 43960 9744 43960 9744 0 FrameData[10]
rlabel metal3 1638 4984 1638 4984 0 FrameData[11]
rlabel metal3 1694 5432 1694 5432 0 FrameData[12]
rlabel metal2 6552 9016 6552 9016 0 FrameData[13]
rlabel metal3 1694 6328 1694 6328 0 FrameData[14]
rlabel metal3 630 6776 630 6776 0 FrameData[15]
rlabel metal3 1414 7224 1414 7224 0 FrameData[16]
rlabel metal3 854 7672 854 7672 0 FrameData[17]
rlabel metal3 50624 952 50624 952 0 FrameData[18]
rlabel metal4 24248 6104 24248 6104 0 FrameData[19]
rlabel metal3 2142 504 2142 504 0 FrameData[1]
rlabel metal2 26152 10248 26152 10248 0 FrameData[20]
rlabel metal3 39032 2184 39032 2184 0 FrameData[21]
rlabel metal2 1624 2800 1624 2800 0 FrameData[22]
rlabel metal3 854 10360 854 10360 0 FrameData[23]
rlabel metal2 13832 2184 13832 2184 0 FrameData[24]
rlabel metal2 16744 1512 16744 1512 0 FrameData[25]
rlabel metal3 1694 11704 1694 11704 0 FrameData[26]
rlabel metal2 14168 2800 14168 2800 0 FrameData[27]
rlabel metal3 462 12600 462 12600 0 FrameData[28]
rlabel metal3 1190 13048 1190 13048 0 FrameData[29]
rlabel metal2 3304 3024 3304 3024 0 FrameData[2]
rlabel metal3 45752 3528 45752 3528 0 FrameData[30]
rlabel metal3 182 13944 182 13944 0 FrameData[31]
rlabel metal2 5600 6552 5600 6552 0 FrameData[3]
rlabel metal2 45416 2800 45416 2800 0 FrameData[4]
rlabel metal3 2142 2296 2142 2296 0 FrameData[5]
rlabel metal2 11592 2184 11592 2184 0 FrameData[6]
rlabel metal3 1862 3192 1862 3192 0 FrameData[7]
rlabel metal3 1134 3640 1134 3640 0 FrameData[8]
rlabel metal3 46872 2072 46872 2072 0 FrameData[9]
rlabel metal3 52122 56 52122 56 0 FrameData_O[0]
rlabel metal3 51898 4536 51898 4536 0 FrameData_O[10]
rlabel metal2 51240 4760 51240 4760 0 FrameData_O[11]
rlabel metal2 51240 5320 51240 5320 0 FrameData_O[12]
rlabel metal3 51226 5880 51226 5880 0 FrameData_O[13]
rlabel metal2 51240 6216 51240 6216 0 FrameData_O[14]
rlabel metal3 51170 6776 51170 6776 0 FrameData_O[15]
rlabel metal2 51464 6888 51464 6888 0 FrameData_O[16]
rlabel metal3 52066 7672 52066 7672 0 FrameData_O[17]
rlabel metal3 51786 8120 51786 8120 0 FrameData_O[18]
rlabel metal3 51842 8568 51842 8568 0 FrameData_O[19]
rlabel metal3 51618 504 51618 504 0 FrameData_O[1]
rlabel metal3 52066 9016 52066 9016 0 FrameData_O[20]
rlabel metal3 51842 9464 51842 9464 0 FrameData_O[21]
rlabel metal3 52066 9912 52066 9912 0 FrameData_O[22]
rlabel metal3 51170 10360 51170 10360 0 FrameData_O[23]
rlabel metal3 51954 10808 51954 10808 0 FrameData_O[24]
rlabel metal3 51282 11256 51282 11256 0 FrameData_O[25]
rlabel metal3 51842 11704 51842 11704 0 FrameData_O[26]
rlabel metal3 51226 12152 51226 12152 0 FrameData_O[27]
rlabel metal3 50442 12600 50442 12600 0 FrameData_O[28]
rlabel metal2 48104 12712 48104 12712 0 FrameData_O[29]
rlabel metal3 51842 952 51842 952 0 FrameData_O[2]
rlabel metal3 50400 9688 50400 9688 0 FrameData_O[30]
rlabel metal3 50400 9240 50400 9240 0 FrameData_O[31]
rlabel metal3 51226 1400 51226 1400 0 FrameData_O[3]
rlabel metal3 51282 1848 51282 1848 0 FrameData_O[4]
rlabel metal2 51464 2072 51464 2072 0 FrameData_O[5]
rlabel metal3 51898 2744 51898 2744 0 FrameData_O[6]
rlabel metal2 51240 3080 51240 3080 0 FrameData_O[7]
rlabel metal3 51058 3640 51058 3640 0 FrameData_O[8]
rlabel metal2 51464 3752 51464 3752 0 FrameData_O[9]
rlabel metal2 4088 238 4088 238 0 FrameStrobe[0]
rlabel metal2 19320 7168 19320 7168 0 FrameStrobe[10]
rlabel metal3 30688 8120 30688 8120 0 FrameStrobe[11]
rlabel metal2 33656 1134 33656 1134 0 FrameStrobe[12]
rlabel metal4 26376 11915 26376 11915 0 FrameStrobe[13]
rlabel metal3 26152 12824 26152 12824 0 FrameStrobe[14]
rlabel metal2 2352 10360 2352 10360 0 FrameStrobe[15]
rlabel metal2 43512 3486 43512 3486 0 FrameStrobe[16]
rlabel metal2 45976 742 45976 742 0 FrameStrobe[17]
rlabel metal2 48440 126 48440 126 0 FrameStrobe[18]
rlabel metal2 50904 182 50904 182 0 FrameStrobe[19]
rlabel metal2 6552 854 6552 854 0 FrameStrobe[1]
rlabel metal2 46200 2912 46200 2912 0 FrameStrobe[2]
rlabel metal2 48328 7784 48328 7784 0 FrameStrobe[3]
rlabel metal3 25256 6720 25256 6720 0 FrameStrobe[4]
rlabel metal2 16408 854 16408 854 0 FrameStrobe[5]
rlabel metal2 18872 798 18872 798 0 FrameStrobe[6]
rlabel metal2 21336 854 21336 854 0 FrameStrobe[7]
rlabel metal2 23800 126 23800 126 0 FrameStrobe[8]
rlabel metal2 9576 56 9576 56 0 FrameStrobe[9]
rlabel metal2 35896 13482 35896 13482 0 FrameStrobe_O[0]
rlabel metal2 38920 10864 38920 10864 0 FrameStrobe_O[10]
rlabel metal2 41608 12712 41608 12712 0 FrameStrobe_O[11]
rlabel metal2 40824 12096 40824 12096 0 FrameStrobe_O[12]
rlabel metal2 38808 13146 38808 13146 0 FrameStrobe_O[13]
rlabel metal2 43736 13272 43736 13272 0 FrameStrobe_O[14]
rlabel metal2 39256 13426 39256 13426 0 FrameStrobe_O[15]
rlabel metal2 39480 13314 39480 13314 0 FrameStrobe_O[16]
rlabel metal2 39704 12810 39704 12810 0 FrameStrobe_O[17]
rlabel metal2 39928 12474 39928 12474 0 FrameStrobe_O[18]
rlabel metal2 40152 13650 40152 13650 0 FrameStrobe_O[19]
rlabel metal2 36568 12712 36568 12712 0 FrameStrobe_O[1]
rlabel metal2 36344 13594 36344 13594 0 FrameStrobe_O[2]
rlabel metal2 38136 12824 38136 12824 0 FrameStrobe_O[3]
rlabel metal2 40040 13272 40040 13272 0 FrameStrobe_O[4]
rlabel metal2 37016 12474 37016 12474 0 FrameStrobe_O[5]
rlabel metal2 38696 12152 38696 12152 0 FrameStrobe_O[6]
rlabel metal2 40040 12432 40040 12432 0 FrameStrobe_O[7]
rlabel metal2 41272 13272 41272 13272 0 FrameStrobe_O[8]
rlabel metal2 39368 11592 39368 11592 0 FrameStrobe_O[9]
rlabel metal2 12376 14098 12376 14098 0 N1BEG[0]
rlabel metal3 11536 10808 11536 10808 0 N1BEG[1]
rlabel metal2 12992 7672 12992 7672 0 N1BEG[2]
rlabel metal2 10920 11704 10920 11704 0 N1BEG[3]
rlabel metal2 13272 13202 13272 13202 0 N2BEG[0]
rlabel metal2 13496 11130 13496 11130 0 N2BEG[1]
rlabel metal3 13048 10024 13048 10024 0 N2BEG[2]
rlabel metal2 13944 13874 13944 13874 0 N2BEG[3]
rlabel metal2 14560 7672 14560 7672 0 N2BEG[4]
rlabel metal2 9800 13272 9800 13272 0 N2BEG[5]
rlabel metal2 14616 13258 14616 13258 0 N2BEG[6]
rlabel metal2 12488 12096 12488 12096 0 N2BEG[7]
rlabel metal2 15176 9352 15176 9352 0 N2BEGb[0]
rlabel metal2 15288 12026 15288 12026 0 N2BEGb[1]
rlabel metal2 15512 13986 15512 13986 0 N2BEGb[2]
rlabel metal2 15736 13818 15736 13818 0 N2BEGb[3]
rlabel metal2 15960 13930 15960 13930 0 N2BEGb[4]
rlabel metal2 15624 11200 15624 11200 0 N2BEGb[5]
rlabel metal2 16408 13370 16408 13370 0 N2BEGb[6]
rlabel metal2 16632 11690 16632 11690 0 N2BEGb[7]
rlabel metal2 16856 13650 16856 13650 0 N4BEG[0]
rlabel metal2 19096 11690 19096 11690 0 N4BEG[10]
rlabel metal2 19320 12082 19320 12082 0 N4BEG[11]
rlabel metal3 18928 12376 18928 12376 0 N4BEG[12]
rlabel metal2 19880 11536 19880 11536 0 N4BEG[13]
rlabel metal3 19432 11480 19432 11480 0 N4BEG[14]
rlabel metal2 17416 13216 17416 13216 0 N4BEG[15]
rlabel metal2 17080 13258 17080 13258 0 N4BEG[1]
rlabel metal2 15512 12432 15512 12432 0 N4BEG[2]
rlabel metal2 17528 13202 17528 13202 0 N4BEG[3]
rlabel metal2 17752 12810 17752 12810 0 N4BEG[4]
rlabel metal2 17976 13650 17976 13650 0 N4BEG[5]
rlabel metal2 18144 9688 18144 9688 0 N4BEG[6]
rlabel metal2 18424 13930 18424 13930 0 N4BEG[7]
rlabel metal2 18312 11088 18312 11088 0 N4BEG[8]
rlabel metal2 16744 12432 16744 12432 0 N4BEG[9]
rlabel metal2 20832 9240 20832 9240 0 NN4BEG[0]
rlabel metal2 22680 12474 22680 12474 0 NN4BEG[10]
rlabel metal2 22904 13930 22904 13930 0 NN4BEG[11]
rlabel metal2 23128 13258 23128 13258 0 NN4BEG[12]
rlabel metal2 22904 13272 22904 13272 0 NN4BEG[13]
rlabel metal2 23576 13202 23576 13202 0 NN4BEG[14]
rlabel metal2 23800 13426 23800 13426 0 NN4BEG[15]
rlabel metal2 20664 13202 20664 13202 0 NN4BEG[1]
rlabel metal3 20216 12264 20216 12264 0 NN4BEG[2]
rlabel metal2 20216 11928 20216 11928 0 NN4BEG[3]
rlabel metal3 20272 12824 20272 12824 0 NN4BEG[4]
rlabel metal2 21560 12922 21560 12922 0 NN4BEG[5]
rlabel metal2 21784 13650 21784 13650 0 NN4BEG[6]
rlabel metal2 22008 12810 22008 12810 0 NN4BEG[7]
rlabel metal3 21952 12376 21952 12376 0 NN4BEG[8]
rlabel metal3 21840 13160 21840 13160 0 NN4BEG[9]
rlabel metal2 29064 3920 29064 3920 0 S1END[0]
rlabel metal2 26376 12712 26376 12712 0 S1END[1]
rlabel metal2 24472 13818 24472 13818 0 S1END[2]
rlabel metal2 23016 10528 23016 10528 0 S1END[3]
rlabel metal2 38920 2856 38920 2856 0 S2END[0]
rlabel metal2 26936 12866 26936 12866 0 S2END[1]
rlabel metal2 27328 12824 27328 12824 0 S2END[2]
rlabel metal3 25536 5992 25536 5992 0 S2END[3]
rlabel metal2 43624 4368 43624 4368 0 S2END[4]
rlabel metal3 24920 7560 24920 7560 0 S2END[5]
rlabel metal2 41944 4536 41944 4536 0 S2END[6]
rlabel metal2 17640 1568 17640 1568 0 S2END[7]
rlabel metal2 19656 7112 19656 7112 0 S2MID[0]
rlabel metal2 48216 7672 48216 7672 0 S2MID[1]
rlabel metal3 47600 4088 47600 4088 0 S2MID[2]
rlabel metal3 46760 5992 46760 5992 0 S2MID[3]
rlabel metal2 42616 12992 42616 12992 0 S2MID[4]
rlabel metal3 20776 2184 20776 2184 0 S2MID[5]
rlabel metal3 21000 1176 21000 1176 0 S2MID[6]
rlabel metal3 24472 12712 24472 12712 0 S2MID[7]
rlabel metal2 23464 6104 23464 6104 0 S4END[0]
rlabel metal2 44408 6496 44408 6496 0 S4END[10]
rlabel metal2 6328 12600 6328 12600 0 S4END[11]
rlabel metal2 46760 4424 46760 4424 0 S4END[12]
rlabel metal3 37296 9128 37296 9128 0 S4END[13]
rlabel metal2 49000 6048 49000 6048 0 S4END[14]
rlabel metal3 27664 9800 27664 9800 0 S4END[15]
rlabel metal3 21560 14056 21560 14056 0 S4END[1]
rlabel metal3 17808 2184 17808 2184 0 S4END[2]
rlabel metal2 15848 3752 15848 3752 0 S4END[3]
rlabel metal2 43624 2800 43624 2800 0 S4END[4]
rlabel metal3 21840 8232 21840 8232 0 S4END[5]
rlabel metal3 2576 3528 2576 3528 0 S4END[6]
rlabel metal3 11592 2408 11592 2408 0 S4END[7]
rlabel metal2 41776 10024 41776 10024 0 S4END[8]
rlabel metal3 21000 8176 21000 8176 0 S4END[9]
rlabel metal2 32312 5936 32312 5936 0 SS4END[0]
rlabel metal2 20944 2184 20944 2184 0 SS4END[10]
rlabel metal2 10920 4816 10920 4816 0 SS4END[11]
rlabel metal2 20664 5600 20664 5600 0 SS4END[12]
rlabel metal2 15624 4648 15624 4648 0 SS4END[13]
rlabel metal3 36512 13160 36512 13160 0 SS4END[14]
rlabel metal2 36848 2856 36848 2856 0 SS4END[15]
rlabel metal2 7112 12880 7112 12880 0 SS4END[1]
rlabel metal2 25816 2632 25816 2632 0 SS4END[2]
rlabel metal2 25144 9744 25144 9744 0 SS4END[3]
rlabel metal2 32984 14042 32984 14042 0 SS4END[4]
rlabel metal2 21224 8120 21224 8120 0 SS4END[5]
rlabel metal2 23688 6496 23688 6496 0 SS4END[6]
rlabel metal3 18312 7112 18312 7112 0 SS4END[7]
rlabel metal2 11928 8232 11928 8232 0 SS4END[8]
rlabel metal2 4424 2800 4424 2800 0 SS4END[9]
rlabel metal2 1624 1134 1624 1134 0 UserCLK
rlabel metal2 35728 13160 35728 13160 0 UserCLKo
rlabel metal2 48776 2464 48776 2464 0 net1
rlabel metal2 51352 4368 51352 4368 0 net10
rlabel metal3 21112 6552 21112 6552 0 net100
rlabel metal2 4088 2856 4088 2856 0 net101
rlabel metal2 18984 10528 18984 10528 0 net102
rlabel metal2 20160 9990 20160 9990 0 net103
rlabel metal2 22904 7560 22904 7560 0 net104
rlabel metal3 32872 3304 32872 3304 0 net105
rlabel metal3 49112 8680 49112 8680 0 net11
rlabel metal3 42672 2744 42672 2744 0 net12
rlabel metal2 42168 9632 42168 9632 0 net13
rlabel metal3 47992 10416 47992 10416 0 net14
rlabel metal3 4592 2856 4592 2856 0 net15
rlabel metal2 48776 10696 48776 10696 0 net16
rlabel metal2 14504 1568 14504 1568 0 net17
rlabel metal3 47264 11368 47264 11368 0 net18
rlabel metal2 41160 9184 41160 9184 0 net19
rlabel metal3 46816 9688 46816 9688 0 net2
rlabel metal2 49560 12936 49560 12936 0 net20
rlabel metal2 45192 11032 45192 11032 0 net21
rlabel metal2 47096 11032 47096 11032 0 net22
rlabel metal4 14168 2632 14168 2632 0 net23
rlabel metal2 48832 6888 48832 6888 0 net24
rlabel metal2 48776 8904 48776 8904 0 net25
rlabel metal2 13384 1624 13384 1624 0 net26
rlabel metal2 48888 2352 48888 2352 0 net27
rlabel metal3 49840 6888 49840 6888 0 net28
rlabel metal2 46200 6384 46200 6384 0 net29
rlabel metal2 50232 3976 50232 3976 0 net3
rlabel metal3 49336 8904 49336 8904 0 net30
rlabel metal3 47096 4312 47096 4312 0 net31
rlabel metal2 47544 2296 47544 2296 0 net32
rlabel metal2 37352 12880 37352 12880 0 net33
rlabel metal2 18536 7392 18536 7392 0 net34
rlabel metal2 38696 9856 38696 9856 0 net35
rlabel metal2 40600 9240 40600 9240 0 net36
rlabel metal3 3920 3304 3920 3304 0 net37
rlabel metal2 42952 12432 42952 12432 0 net38
rlabel metal2 1736 9968 1736 9968 0 net39
rlabel metal3 49448 10136 49448 10136 0 net4
rlabel metal2 25928 12768 25928 12768 0 net40
rlabel metal2 39928 7840 39928 7840 0 net41
rlabel metal2 17080 5992 17080 5992 0 net42
rlabel metal2 44296 12320 44296 12320 0 net43
rlabel metal2 45304 10416 45304 10416 0 net44
rlabel metal2 46872 4648 46872 4648 0 net45
rlabel metal3 45304 8344 45304 8344 0 net46
rlabel metal2 38808 7924 38808 7924 0 net47
rlabel metal3 30912 6664 30912 6664 0 net48
rlabel metal2 35336 5152 35336 5152 0 net49
rlabel metal2 49000 3472 49000 3472 0 net5
rlabel metal2 39480 12208 39480 12208 0 net50
rlabel metal2 40712 13328 40712 13328 0 net51
rlabel metal2 38808 10864 38808 10864 0 net52
rlabel metal3 17248 8904 17248 8904 0 net53
rlabel metal2 9576 6104 9576 6104 0 net54
rlabel metal3 17416 7504 17416 7504 0 net55
rlabel metal3 24304 2968 24304 2968 0 net56
rlabel metal4 21560 9007 21560 9007 0 net57
rlabel metal2 20440 1848 20440 1848 0 net58
rlabel metal3 17080 2968 17080 2968 0 net59
rlabel metal3 49168 6664 49168 6664 0 net6
rlabel metal2 40600 5712 40600 5712 0 net60
rlabel metal2 48552 6272 48552 6272 0 net61
rlabel metal2 48328 3920 48328 3920 0 net62
rlabel metal2 50008 7840 50008 7840 0 net63
rlabel metal2 13944 9016 13944 9016 0 net64
rlabel metal3 16520 2856 16520 2856 0 net65
rlabel metal2 42728 4704 42728 4704 0 net66
rlabel metal2 23352 7616 23352 7616 0 net67
rlabel metal2 18088 4144 18088 4144 0 net68
rlabel metal2 23744 5992 23744 5992 0 net69
rlabel metal2 48776 7392 48776 7392 0 net7
rlabel metal3 20384 3080 20384 3080 0 net70
rlabel metal2 15400 10416 15400 10416 0 net71
rlabel metal2 39480 2520 39480 2520 0 net72
rlabel metal2 26376 9744 26376 9744 0 net73
rlabel metal3 20552 8344 20552 8344 0 net74
rlabel metal3 24080 2184 24080 2184 0 net75
rlabel metal2 17304 12768 17304 12768 0 net76
rlabel metal2 14280 8064 14280 8064 0 net77
rlabel metal2 18088 11312 18088 11312 0 net78
rlabel metal3 19152 12152 19152 12152 0 net79
rlabel metal2 45304 3752 45304 3752 0 net8
rlabel metal2 49896 6104 49896 6104 0 net80
rlabel metal2 39144 7728 39144 7728 0 net81
rlabel metal2 47320 2016 47320 2016 0 net82
rlabel metal2 17304 8736 17304 8736 0 net83
rlabel metal2 45080 5936 45080 5936 0 net84
rlabel metal2 17080 9408 17080 9408 0 net85
rlabel metal2 38808 9856 38808 9856 0 net86
rlabel metal2 6888 11368 6888 11368 0 net87
rlabel metal2 1848 4704 1848 4704 0 net88
rlabel metal3 25032 616 25032 616 0 net89
rlabel metal2 35336 8960 35336 8960 0 net9
rlabel metal3 16520 11088 16520 11088 0 net90
rlabel metal2 11816 2968 11816 2968 0 net91
rlabel metal3 23912 9912 23912 9912 0 net92
rlabel metal2 10472 5600 10472 5600 0 net93
rlabel metal2 23800 11928 23800 11928 0 net94
rlabel metal3 26376 10192 26376 10192 0 net95
rlabel metal4 24920 5600 24920 5600 0 net96
rlabel metal2 17528 11088 17528 11088 0 net97
rlabel metal2 19768 7504 19768 7504 0 net98
rlabel metal2 16744 8960 16744 8960 0 net99
<< properties >>
string FIXED_BBOX 0 0 52752 14224
<< end >>
