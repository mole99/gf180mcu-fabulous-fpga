magic
tech gf180mcuD
magscale 1 10
timestamp 1764323338
<< metal1 >>
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 10670 13186 10722 13198
rect 2034 13134 2046 13186
rect 2098 13134 2110 13186
rect 10670 13122 10722 13134
rect 53118 13186 53170 13198
rect 53118 13122 53170 13134
rect 8082 13022 8094 13074
rect 8146 13022 8158 13074
rect 43362 13022 43374 13074
rect 43426 13022 43438 13074
rect 2382 12962 2434 12974
rect 6066 12910 6078 12962
rect 6130 12910 6142 12962
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 14018 12910 14030 12962
rect 14082 12910 14094 12962
rect 19394 12910 19406 12962
rect 19458 12910 19470 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 25106 12910 25118 12962
rect 25170 12910 25182 12962
rect 27122 12910 27134 12962
rect 27186 12910 27198 12962
rect 30034 12910 30046 12962
rect 30098 12910 30110 12962
rect 32834 12910 32846 12962
rect 32898 12910 32910 12962
rect 38210 12910 38222 12962
rect 38274 12910 38286 12962
rect 40898 12910 40910 12962
rect 40962 12910 40974 12962
rect 44146 12910 44158 12962
rect 44210 12910 44222 12962
rect 45938 12910 45950 12962
rect 46002 12910 46014 12962
rect 48962 12910 48974 12962
rect 49026 12910 49038 12962
rect 51762 12910 51774 12962
rect 51826 12910 51838 12962
rect 52546 12910 52558 12962
rect 52610 12910 52622 12962
rect 55122 12910 55134 12962
rect 55186 12910 55198 12962
rect 2382 12898 2434 12910
rect 5070 12850 5122 12862
rect 13022 12850 13074 12862
rect 7186 12798 7198 12850
rect 7250 12798 7262 12850
rect 5070 12786 5122 12798
rect 13022 12786 13074 12798
rect 18398 12850 18450 12862
rect 18398 12786 18450 12798
rect 21086 12850 21138 12862
rect 21086 12786 21138 12798
rect 24110 12850 24162 12862
rect 24110 12786 24162 12798
rect 26126 12850 26178 12862
rect 26126 12786 26178 12798
rect 29150 12850 29202 12862
rect 29150 12786 29202 12798
rect 31838 12850 31890 12862
rect 31838 12786 31890 12798
rect 37214 12850 37266 12862
rect 37214 12786 37266 12798
rect 39902 12850 39954 12862
rect 39902 12786 39954 12798
rect 45166 12850 45218 12862
rect 45166 12786 45218 12798
rect 47966 12850 48018 12862
rect 47966 12786 48018 12798
rect 50766 12850 50818 12862
rect 50766 12786 50818 12798
rect 56142 12738 56194 12750
rect 56142 12674 56194 12686
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 15710 12402 15762 12414
rect 15710 12338 15762 12350
rect 34526 12402 34578 12414
rect 34526 12338 34578 12350
rect 53006 12402 53058 12414
rect 53006 12338 53058 12350
rect 10446 12290 10498 12302
rect 20638 12290 20690 12302
rect 15026 12238 15038 12290
rect 15090 12238 15102 12290
rect 10446 12226 10498 12238
rect 20638 12226 20690 12238
rect 22318 12290 22370 12302
rect 22318 12226 22370 12238
rect 26462 12290 26514 12302
rect 39902 12290 39954 12302
rect 30594 12238 30606 12290
rect 30658 12238 30670 12290
rect 49970 12238 49982 12290
rect 50034 12238 50046 12290
rect 26462 12226 26514 12238
rect 39902 12226 39954 12238
rect 11006 12178 11058 12190
rect 11006 12114 11058 12126
rect 21198 12178 21250 12190
rect 21198 12114 21250 12126
rect 22878 12178 22930 12190
rect 29038 12178 29090 12190
rect 32398 12178 32450 12190
rect 23538 12126 23550 12178
rect 23602 12126 23614 12178
rect 28578 12126 28590 12178
rect 28642 12126 28654 12178
rect 30258 12126 30270 12178
rect 30322 12126 30334 12178
rect 22878 12114 22930 12126
rect 29038 12114 29090 12126
rect 32398 12114 32450 12126
rect 46846 12178 46898 12190
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 53554 12126 53566 12178
rect 53618 12126 53630 12178
rect 46846 12114 46898 12126
rect 23998 12066 24050 12078
rect 16706 12014 16718 12066
rect 16770 12014 16782 12066
rect 23998 12002 24050 12014
rect 26126 12066 26178 12078
rect 26126 12002 26178 12014
rect 32958 12066 33010 12078
rect 37102 12066 37154 12078
rect 35522 12014 35534 12066
rect 35586 12014 35598 12066
rect 32958 12002 33010 12014
rect 37102 12002 37154 12014
rect 47406 12066 47458 12078
rect 54338 12014 54350 12066
rect 54402 12014 54414 12066
rect 55122 12014 55134 12066
rect 55186 12014 55198 12066
rect 55906 12014 55918 12066
rect 55970 12014 55982 12066
rect 47406 12002 47458 12014
rect 14590 11954 14642 11966
rect 14590 11890 14642 11902
rect 25566 11954 25618 11966
rect 25566 11890 25618 11902
rect 27022 11954 27074 11966
rect 27022 11890 27074 11902
rect 37662 11954 37714 11966
rect 37662 11890 37714 11902
rect 40462 11954 40514 11966
rect 44942 11954 44994 11966
rect 44594 11902 44606 11954
rect 44658 11902 44670 11954
rect 40462 11890 40514 11902
rect 44942 11890 44994 11902
rect 49534 11954 49586 11966
rect 49534 11890 49586 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 14254 11506 14306 11518
rect 14254 11442 14306 11454
rect 18174 11506 18226 11518
rect 50978 11454 50990 11506
rect 51042 11454 51054 11506
rect 18174 11442 18226 11454
rect 14814 11394 14866 11406
rect 14814 11330 14866 11342
rect 18734 11394 18786 11406
rect 18734 11330 18786 11342
rect 24558 11394 24610 11406
rect 24558 11330 24610 11342
rect 35086 11394 35138 11406
rect 35086 11330 35138 11342
rect 47518 11394 47570 11406
rect 52546 11342 52558 11394
rect 52610 11342 52622 11394
rect 54114 11342 54126 11394
rect 54178 11342 54190 11394
rect 47518 11330 47570 11342
rect 25118 11282 25170 11294
rect 25118 11218 25170 11230
rect 35646 11282 35698 11294
rect 51998 11282 52050 11294
rect 47058 11230 47070 11282
rect 47122 11230 47134 11282
rect 35646 11218 35698 11230
rect 51998 11218 52050 11230
rect 53566 11170 53618 11182
rect 53566 11106 53618 11118
rect 55134 11170 55186 11182
rect 55134 11106 55186 11118
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 53006 10834 53058 10846
rect 53006 10770 53058 10782
rect 28702 10722 28754 10734
rect 28702 10658 28754 10670
rect 38558 10722 38610 10734
rect 38558 10658 38610 10670
rect 54574 10722 54626 10734
rect 54574 10658 54626 10670
rect 56142 10722 56194 10734
rect 56142 10658 56194 10670
rect 29262 10610 29314 10622
rect 29262 10546 29314 10558
rect 30830 10610 30882 10622
rect 30830 10546 30882 10558
rect 34526 10610 34578 10622
rect 34526 10546 34578 10558
rect 35086 10610 35138 10622
rect 52098 10558 52110 10610
rect 52162 10558 52174 10610
rect 35086 10546 35138 10558
rect 31390 10498 31442 10510
rect 53554 10446 53566 10498
rect 53618 10446 53630 10498
rect 55122 10446 55134 10498
rect 55186 10446 55198 10498
rect 31390 10434 31442 10446
rect 37998 10386 38050 10398
rect 37998 10322 38050 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 19406 10050 19458 10062
rect 19406 9986 19458 9998
rect 32622 9938 32674 9950
rect 32622 9874 32674 9886
rect 34638 9938 34690 9950
rect 34638 9874 34690 9886
rect 35198 9938 35250 9950
rect 35198 9874 35250 9886
rect 33182 9826 33234 9838
rect 52546 9774 52558 9826
rect 52610 9774 52622 9826
rect 54226 9774 54238 9826
rect 54290 9774 54302 9826
rect 33182 9762 33234 9774
rect 19966 9714 20018 9726
rect 19966 9650 20018 9662
rect 53566 9714 53618 9726
rect 53566 9650 53618 9662
rect 55134 9602 55186 9614
rect 55134 9538 55186 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 2942 9154 2994 9166
rect 28914 9102 28926 9154
rect 28978 9102 28990 9154
rect 2942 9090 2994 9102
rect 23214 9042 23266 9054
rect 23214 8978 23266 8990
rect 25566 9042 25618 9054
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 55234 8990 55246 9042
rect 55298 8990 55310 9042
rect 25566 8978 25618 8990
rect 22654 8930 22706 8942
rect 22654 8866 22706 8878
rect 26126 8930 26178 8942
rect 26126 8866 26178 8878
rect 41694 8930 41746 8942
rect 41694 8866 41746 8878
rect 44718 8930 44770 8942
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 55906 8878 55918 8930
rect 55970 8878 55982 8930
rect 44718 8866 44770 8878
rect 2382 8818 2434 8830
rect 2382 8754 2434 8766
rect 41134 8818 41186 8830
rect 41134 8754 41186 8766
rect 44158 8818 44210 8830
rect 44158 8754 44210 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 22430 8482 22482 8494
rect 22430 8418 22482 8430
rect 30718 8482 30770 8494
rect 30718 8418 30770 8430
rect 29262 8370 29314 8382
rect 29262 8306 29314 8318
rect 29822 8370 29874 8382
rect 54114 8318 54126 8370
rect 54178 8318 54190 8370
rect 54898 8318 54910 8370
rect 54962 8318 54974 8370
rect 29822 8306 29874 8318
rect 18286 8258 18338 8270
rect 18286 8194 18338 8206
rect 43598 8258 43650 8270
rect 43598 8194 43650 8206
rect 22990 8146 23042 8158
rect 44158 8146 44210 8158
rect 17826 8094 17838 8146
rect 17890 8094 17902 8146
rect 31154 8094 31166 8146
rect 31218 8094 31230 8146
rect 22990 8082 23042 8094
rect 44158 8082 44210 8094
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 56142 7698 56194 7710
rect 56142 7634 56194 7646
rect 35646 7586 35698 7598
rect 9202 7534 9214 7586
rect 9266 7534 9278 7586
rect 26338 7534 26350 7586
rect 26402 7534 26414 7586
rect 35646 7522 35698 7534
rect 54574 7586 54626 7598
rect 54574 7522 54626 7534
rect 20862 7474 20914 7486
rect 20862 7410 20914 7422
rect 25902 7474 25954 7486
rect 53554 7422 53566 7474
rect 53618 7422 53630 7474
rect 55122 7422 55134 7474
rect 55186 7422 55198 7474
rect 25902 7410 25954 7422
rect 5406 7362 5458 7374
rect 5406 7298 5458 7310
rect 21422 7362 21474 7374
rect 21422 7298 21474 7310
rect 5966 7250 6018 7262
rect 5966 7186 6018 7198
rect 9662 7250 9714 7262
rect 9662 7186 9714 7198
rect 35086 7250 35138 7262
rect 35086 7186 35138 7198
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 16158 6802 16210 6814
rect 16158 6738 16210 6750
rect 15598 6690 15650 6702
rect 15598 6626 15650 6638
rect 26462 6690 26514 6702
rect 26462 6626 26514 6638
rect 43262 6690 43314 6702
rect 43262 6626 43314 6638
rect 44830 6690 44882 6702
rect 54114 6638 54126 6690
rect 54178 6638 54190 6690
rect 44830 6626 44882 6638
rect 27022 6578 27074 6590
rect 43698 6526 43710 6578
rect 43762 6526 43774 6578
rect 45266 6526 45278 6578
rect 45330 6526 45342 6578
rect 27022 6514 27074 6526
rect 55134 6466 55186 6478
rect 55134 6402 55186 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 56142 6130 56194 6142
rect 56142 6066 56194 6078
rect 54574 6018 54626 6030
rect 40450 5966 40462 6018
rect 40514 5966 40526 6018
rect 54574 5954 54626 5966
rect 35758 5906 35810 5918
rect 46622 5906 46674 5918
rect 40114 5854 40126 5906
rect 40178 5854 40190 5906
rect 35758 5842 35810 5854
rect 46622 5842 46674 5854
rect 49422 5906 49474 5918
rect 53554 5854 53566 5906
rect 53618 5854 53630 5906
rect 55346 5854 55358 5906
rect 55410 5854 55422 5906
rect 49422 5842 49474 5854
rect 14254 5794 14306 5806
rect 14254 5730 14306 5742
rect 17166 5794 17218 5806
rect 17166 5730 17218 5742
rect 24446 5794 24498 5806
rect 24446 5730 24498 5742
rect 24782 5794 24834 5806
rect 24782 5730 24834 5742
rect 25342 5794 25394 5806
rect 25342 5730 25394 5742
rect 37886 5794 37938 5806
rect 37886 5730 37938 5742
rect 47182 5794 47234 5806
rect 47182 5730 47234 5742
rect 49982 5794 50034 5806
rect 49982 5730 50034 5742
rect 14814 5682 14866 5694
rect 14814 5618 14866 5630
rect 16606 5682 16658 5694
rect 16606 5618 16658 5630
rect 23886 5682 23938 5694
rect 23886 5618 23938 5630
rect 35198 5682 35250 5694
rect 35198 5618 35250 5630
rect 37326 5682 37378 5694
rect 37326 5618 37378 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 18622 5346 18674 5358
rect 18622 5282 18674 5294
rect 29822 5346 29874 5358
rect 29822 5282 29874 5294
rect 32398 5346 32450 5358
rect 32398 5282 32450 5294
rect 52894 5346 52946 5358
rect 52894 5282 52946 5294
rect 53230 5346 53282 5358
rect 53230 5282 53282 5294
rect 32958 5234 33010 5246
rect 32958 5170 33010 5182
rect 52334 5234 52386 5246
rect 52334 5170 52386 5182
rect 10894 5122 10946 5134
rect 10894 5058 10946 5070
rect 20078 5122 20130 5134
rect 20078 5058 20130 5070
rect 28926 5122 28978 5134
rect 28926 5058 28978 5070
rect 34638 5122 34690 5134
rect 34638 5058 34690 5070
rect 35198 5122 35250 5134
rect 39118 5122 39170 5134
rect 38658 5070 38670 5122
rect 38722 5070 38734 5122
rect 35198 5058 35250 5070
rect 39118 5058 39170 5070
rect 42590 5122 42642 5134
rect 42590 5058 42642 5070
rect 43150 5122 43202 5134
rect 47518 5122 47570 5134
rect 47058 5070 47070 5122
rect 47122 5070 47134 5122
rect 54226 5070 54238 5122
rect 54290 5070 54302 5122
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 43150 5058 43202 5070
rect 47518 5058 47570 5070
rect 19182 5010 19234 5022
rect 29486 5010 29538 5022
rect 10434 4958 10446 5010
rect 10498 4958 10510 5010
rect 19618 4958 19630 5010
rect 19682 4958 19694 5010
rect 19182 4946 19234 4958
rect 29486 4946 29538 4958
rect 30382 5010 30434 5022
rect 30382 4946 30434 4958
rect 53790 5010 53842 5022
rect 53790 4946 53842 4958
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 54574 4562 54626 4574
rect 54574 4498 54626 4510
rect 56142 4562 56194 4574
rect 56142 4498 56194 4510
rect 52670 4450 52722 4462
rect 11778 4398 11790 4450
rect 11842 4398 11854 4450
rect 18162 4398 18174 4450
rect 18226 4398 18238 4450
rect 24322 4398 24334 4450
rect 24386 4398 24398 4450
rect 35634 4398 35646 4450
rect 35698 4398 35710 4450
rect 36754 4398 36766 4450
rect 36818 4398 36830 4450
rect 45378 4398 45390 4450
rect 45442 4398 45454 4450
rect 52670 4386 52722 4398
rect 2606 4338 2658 4350
rect 39230 4338 39282 4350
rect 32610 4286 32622 4338
rect 32674 4286 32686 4338
rect 35298 4286 35310 4338
rect 35362 4286 35374 4338
rect 2606 4274 2658 4286
rect 39230 4274 39282 4286
rect 41470 4338 41522 4350
rect 41470 4274 41522 4286
rect 44942 4338 44994 4350
rect 53666 4286 53678 4338
rect 53730 4286 53742 4338
rect 55234 4286 55246 4338
rect 55298 4286 55310 4338
rect 44942 4274 44994 4286
rect 10110 4226 10162 4238
rect 10110 4162 10162 4174
rect 33070 4226 33122 4238
rect 33070 4162 33122 4174
rect 39790 4226 39842 4238
rect 39790 4162 39842 4174
rect 42030 4226 42082 4238
rect 46610 4174 46622 4226
rect 46674 4174 46686 4226
rect 42030 4162 42082 4174
rect 3166 4114 3218 4126
rect 3166 4050 3218 4062
rect 10670 4114 10722 4126
rect 10670 4050 10722 4062
rect 12238 4114 12290 4126
rect 12238 4050 12290 4062
rect 18622 4114 18674 4126
rect 18622 4050 18674 4062
rect 23886 4114 23938 4126
rect 23886 4050 23938 4062
rect 36318 4114 36370 4126
rect 36318 4050 36370 4062
rect 47182 4114 47234 4126
rect 47182 4050 47234 4062
rect 53230 4114 53282 4126
rect 53230 4050 53282 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 27582 3778 27634 3790
rect 27582 3714 27634 3726
rect 46510 3778 46562 3790
rect 46510 3714 46562 3726
rect 49758 3778 49810 3790
rect 49758 3714 49810 3726
rect 51326 3778 51378 3790
rect 51326 3714 51378 3726
rect 24558 3666 24610 3678
rect 49198 3666 49250 3678
rect 26002 3614 26014 3666
rect 26066 3614 26078 3666
rect 37538 3614 37550 3666
rect 37602 3614 37614 3666
rect 39106 3614 39118 3666
rect 39170 3614 39182 3666
rect 41794 3614 41806 3666
rect 41858 3614 41870 3666
rect 43362 3614 43374 3666
rect 43426 3614 43438 3666
rect 24558 3602 24610 3614
rect 49198 3602 49250 3614
rect 50766 3666 50818 3678
rect 50766 3602 50818 3614
rect 51662 3666 51714 3678
rect 52546 3614 52558 3666
rect 52610 3614 52622 3666
rect 54114 3614 54126 3666
rect 54178 3614 54190 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 51662 3602 51714 3614
rect 48302 3554 48354 3566
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 33394 3502 33406 3554
rect 33458 3502 33470 3554
rect 35746 3502 35758 3554
rect 35810 3502 35822 3554
rect 41346 3502 41358 3554
rect 41410 3502 41422 3554
rect 45042 3502 45054 3554
rect 45106 3502 45118 3554
rect 48302 3490 48354 3502
rect 48862 3554 48914 3566
rect 48862 3490 48914 3502
rect 52222 3554 52274 3566
rect 52222 3490 52274 3502
rect 23998 3442 24050 3454
rect 28142 3442 28194 3454
rect 43934 3442 43986 3454
rect 53566 3442 53618 3454
rect 24994 3390 25006 3442
rect 25058 3390 25070 3442
rect 38210 3390 38222 3442
rect 38274 3390 38286 3442
rect 40562 3390 40574 3442
rect 40626 3390 40638 3442
rect 46946 3390 46958 3442
rect 47010 3390 47022 3442
rect 23998 3378 24050 3390
rect 28142 3378 28194 3390
rect 43934 3378 43986 3390
rect 53566 3378 53618 3390
rect 26574 3330 26626 3342
rect 26574 3266 26626 3278
rect 32622 3330 32674 3342
rect 32622 3266 32674 3278
rect 34750 3330 34802 3342
rect 34750 3266 34802 3278
rect 36542 3330 36594 3342
rect 36542 3266 36594 3278
rect 42366 3330 42418 3342
rect 42366 3266 42418 3278
rect 45502 3330 45554 3342
rect 45502 3266 45554 3278
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 54574 2994 54626 3006
rect 54574 2930 54626 2942
rect 56142 2994 56194 3006
rect 56142 2930 56194 2942
rect 30158 2882 30210 2894
rect 30158 2818 30210 2830
rect 38110 2882 38162 2894
rect 38110 2818 38162 2830
rect 41246 2882 41298 2894
rect 53006 2882 53058 2894
rect 44818 2830 44830 2882
rect 44882 2830 44894 2882
rect 41246 2818 41298 2830
rect 53006 2818 53058 2830
rect 43038 2770 43090 2782
rect 50878 2770 50930 2782
rect 25218 2718 25230 2770
rect 25282 2718 25294 2770
rect 30482 2718 30494 2770
rect 30546 2718 30558 2770
rect 34850 2718 34862 2770
rect 34914 2718 34926 2770
rect 35298 2718 35310 2770
rect 35362 2718 35374 2770
rect 36306 2718 36318 2770
rect 36370 2718 36382 2770
rect 39106 2718 39118 2770
rect 39170 2718 39182 2770
rect 40674 2718 40686 2770
rect 40738 2718 40750 2770
rect 42242 2718 42254 2770
rect 42306 2718 42318 2770
rect 44258 2718 44270 2770
rect 44322 2718 44334 2770
rect 45714 2718 45726 2770
rect 45778 2718 45790 2770
rect 47282 2718 47294 2770
rect 47346 2718 47358 2770
rect 48962 2718 48974 2770
rect 49026 2718 49038 2770
rect 52098 2718 52110 2770
rect 52162 2718 52174 2770
rect 53554 2718 53566 2770
rect 53618 2718 53630 2770
rect 55122 2718 55134 2770
rect 55186 2718 55198 2770
rect 43038 2706 43090 2718
rect 50878 2706 50930 2718
rect 14366 2658 14418 2670
rect 14366 2594 14418 2606
rect 17838 2658 17890 2670
rect 29262 2658 29314 2670
rect 35758 2658 35810 2670
rect 43598 2658 43650 2670
rect 26674 2606 26686 2658
rect 26738 2606 26750 2658
rect 32050 2606 32062 2658
rect 32114 2606 32126 2658
rect 34066 2606 34078 2658
rect 34130 2606 34142 2658
rect 37090 2606 37102 2658
rect 37154 2606 37166 2658
rect 39890 2606 39902 2658
rect 39954 2606 39966 2658
rect 17838 2594 17890 2606
rect 29262 2594 29314 2606
rect 35758 2594 35810 2606
rect 43598 2594 43650 2606
rect 51438 2658 51490 2670
rect 51438 2594 51490 2606
rect 13806 2546 13858 2558
rect 13806 2482 13858 2494
rect 17278 2546 17330 2558
rect 17278 2482 17330 2494
rect 25678 2546 25730 2558
rect 25678 2482 25730 2494
rect 27246 2546 27298 2558
rect 27246 2482 27298 2494
rect 28702 2546 28754 2558
rect 28702 2482 28754 2494
rect 29598 2546 29650 2558
rect 29598 2482 29650 2494
rect 31054 2546 31106 2558
rect 31054 2482 31106 2494
rect 32622 2546 32674 2558
rect 32622 2482 32674 2494
rect 46286 2546 46338 2558
rect 46286 2482 46338 2494
rect 47854 2546 47906 2558
rect 47854 2482 47906 2494
rect 49422 2546 49474 2558
rect 49422 2482 49474 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 19182 2210 19234 2222
rect 19182 2146 19234 2158
rect 20862 2210 20914 2222
rect 20862 2146 20914 2158
rect 25118 2210 25170 2222
rect 25118 2146 25170 2158
rect 31278 2210 31330 2222
rect 31278 2146 31330 2158
rect 1710 2098 1762 2110
rect 1710 2034 1762 2046
rect 21422 2098 21474 2110
rect 21422 2034 21474 2046
rect 22430 2098 22482 2110
rect 31838 2098 31890 2110
rect 46510 2098 46562 2110
rect 51214 2098 51266 2110
rect 22754 2046 22766 2098
rect 22818 2046 22830 2098
rect 26002 2046 26014 2098
rect 26066 2046 26078 2098
rect 28802 2046 28814 2098
rect 28866 2046 28878 2098
rect 30370 2046 30382 2098
rect 30434 2046 30446 2098
rect 32386 2046 32398 2098
rect 32450 2046 32462 2098
rect 35186 2046 35198 2098
rect 35250 2046 35262 2098
rect 41458 2046 41470 2098
rect 41522 2046 41534 2098
rect 43362 2046 43374 2098
rect 43426 2046 43438 2098
rect 44930 2046 44942 2098
rect 44994 2046 45006 2098
rect 48066 2046 48078 2098
rect 48130 2046 48142 2098
rect 49634 2046 49646 2098
rect 49698 2046 49710 2098
rect 52546 2046 52558 2098
rect 52610 2046 52622 2098
rect 54114 2046 54126 2098
rect 54178 2046 54190 2098
rect 54898 2046 54910 2098
rect 54962 2046 54974 2098
rect 22430 2034 22482 2046
rect 31838 2034 31890 2046
rect 46510 2034 46562 2046
rect 51214 2034 51266 2046
rect 2270 1986 2322 1998
rect 2270 1922 2322 1934
rect 9550 1986 9602 1998
rect 9550 1922 9602 1934
rect 21870 1986 21922 1998
rect 38670 1986 38722 1998
rect 36754 1934 36766 1986
rect 36818 1934 36830 1986
rect 38098 1934 38110 1986
rect 38162 1934 38174 1986
rect 21870 1922 21922 1934
rect 38670 1922 38722 1934
rect 39230 1986 39282 1998
rect 47070 1986 47122 1998
rect 43026 1934 43038 1986
rect 43090 1934 43102 1986
rect 39230 1922 39282 1934
rect 47070 1922 47122 1934
rect 51774 1986 51826 1998
rect 51774 1922 51826 1934
rect 19742 1874 19794 1886
rect 9986 1822 9998 1874
rect 10050 1822 10062 1874
rect 19742 1810 19794 1822
rect 25678 1874 25730 1886
rect 32958 1874 33010 1886
rect 28018 1822 28030 1874
rect 28082 1822 28094 1874
rect 25678 1810 25730 1822
rect 32958 1810 33010 1822
rect 35758 1874 35810 1886
rect 53566 1874 53618 1886
rect 45714 1822 45726 1874
rect 45778 1822 45790 1874
rect 48738 1822 48750 1874
rect 48802 1822 48814 1874
rect 50530 1822 50542 1874
rect 50594 1822 50606 1874
rect 35758 1810 35810 1822
rect 53566 1810 53618 1822
rect 23774 1762 23826 1774
rect 23774 1698 23826 1710
rect 27022 1762 27074 1774
rect 27022 1698 27074 1710
rect 29374 1762 29426 1774
rect 29374 1698 29426 1710
rect 34190 1762 34242 1774
rect 34190 1698 34242 1710
rect 37326 1762 37378 1774
rect 37326 1698 37378 1710
rect 40462 1762 40514 1774
rect 40462 1698 40514 1710
rect 42030 1762 42082 1774
rect 42030 1698 42082 1710
rect 43934 1762 43986 1774
rect 43934 1698 43986 1710
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 53566 1426 53618 1438
rect 53566 1362 53618 1374
rect 56142 1426 56194 1438
rect 56142 1362 56194 1374
rect 26910 1314 26962 1326
rect 26910 1250 26962 1262
rect 40910 1314 40962 1326
rect 40910 1250 40962 1262
rect 51998 1314 52050 1326
rect 51998 1250 52050 1262
rect 22082 1150 22094 1202
rect 22146 1150 22158 1202
rect 24322 1150 24334 1202
rect 24386 1150 24398 1202
rect 26114 1150 26126 1202
rect 26178 1150 26190 1202
rect 29138 1150 29150 1202
rect 29202 1150 29214 1202
rect 29586 1150 29598 1202
rect 29650 1150 29662 1202
rect 31490 1150 31502 1202
rect 31554 1150 31566 1202
rect 33058 1150 33070 1202
rect 33122 1150 33134 1202
rect 35298 1150 35310 1202
rect 35362 1150 35374 1202
rect 37090 1150 37102 1202
rect 37154 1150 37166 1202
rect 40114 1150 40126 1202
rect 40178 1150 40190 1202
rect 41906 1150 41918 1202
rect 41970 1150 41982 1202
rect 44146 1150 44158 1202
rect 44210 1150 44222 1202
rect 44482 1150 44494 1202
rect 44546 1150 44558 1202
rect 46722 1150 46734 1202
rect 46786 1150 46798 1202
rect 48402 1150 48414 1202
rect 48466 1150 48478 1202
rect 50978 1150 50990 1202
rect 51042 1150 51054 1202
rect 52770 1150 52782 1202
rect 52834 1150 52846 1202
rect 55122 1150 55134 1202
rect 55186 1150 55198 1202
rect 22866 1038 22878 1090
rect 22930 1038 22942 1090
rect 25106 1038 25118 1090
rect 25170 1038 25182 1090
rect 28466 1038 28478 1090
rect 28530 1038 28542 1090
rect 39554 1038 39566 1090
rect 39618 1038 39630 1090
rect 43362 1038 43374 1090
rect 43426 1038 43438 1090
rect 30158 978 30210 990
rect 30158 914 30210 926
rect 32062 978 32114 990
rect 32062 914 32114 926
rect 33630 978 33682 990
rect 33630 914 33682 926
rect 35870 978 35922 990
rect 35870 914 35922 926
rect 37438 978 37490 990
rect 37438 914 37490 926
rect 45054 978 45106 990
rect 45054 914 45106 926
rect 47294 978 47346 990
rect 47294 914 47346 926
rect 48862 978 48914 990
rect 48862 914 48914 926
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 2046 13134 2098 13186
rect 10670 13134 10722 13186
rect 53118 13134 53170 13186
rect 8094 13022 8146 13074
rect 43374 13022 43426 13074
rect 2382 12910 2434 12962
rect 6078 12910 6130 12962
rect 10334 12910 10386 12962
rect 14030 12910 14082 12962
rect 19406 12910 19458 12962
rect 22094 12910 22146 12962
rect 25118 12910 25170 12962
rect 27134 12910 27186 12962
rect 30046 12910 30098 12962
rect 32846 12910 32898 12962
rect 38222 12910 38274 12962
rect 40910 12910 40962 12962
rect 44158 12910 44210 12962
rect 45950 12910 46002 12962
rect 48974 12910 49026 12962
rect 51774 12910 51826 12962
rect 52558 12910 52610 12962
rect 55134 12910 55186 12962
rect 5070 12798 5122 12850
rect 7198 12798 7250 12850
rect 13022 12798 13074 12850
rect 18398 12798 18450 12850
rect 21086 12798 21138 12850
rect 24110 12798 24162 12850
rect 26126 12798 26178 12850
rect 29150 12798 29202 12850
rect 31838 12798 31890 12850
rect 37214 12798 37266 12850
rect 39902 12798 39954 12850
rect 45166 12798 45218 12850
rect 47966 12798 48018 12850
rect 50766 12798 50818 12850
rect 56142 12686 56194 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 15710 12350 15762 12402
rect 34526 12350 34578 12402
rect 53006 12350 53058 12402
rect 10446 12238 10498 12290
rect 15038 12238 15090 12290
rect 20638 12238 20690 12290
rect 22318 12238 22370 12290
rect 26462 12238 26514 12290
rect 30606 12238 30658 12290
rect 39902 12238 39954 12290
rect 49982 12238 50034 12290
rect 11006 12126 11058 12178
rect 21198 12126 21250 12178
rect 22878 12126 22930 12178
rect 23550 12126 23602 12178
rect 28590 12126 28642 12178
rect 29038 12126 29090 12178
rect 30270 12126 30322 12178
rect 32398 12126 32450 12178
rect 46846 12126 46898 12178
rect 52222 12126 52274 12178
rect 53566 12126 53618 12178
rect 16718 12014 16770 12066
rect 23998 12014 24050 12066
rect 26126 12014 26178 12066
rect 32958 12014 33010 12066
rect 35534 12014 35586 12066
rect 37102 12014 37154 12066
rect 47406 12014 47458 12066
rect 54350 12014 54402 12066
rect 55134 12014 55186 12066
rect 55918 12014 55970 12066
rect 14590 11902 14642 11954
rect 25566 11902 25618 11954
rect 27022 11902 27074 11954
rect 37662 11902 37714 11954
rect 40462 11902 40514 11954
rect 44606 11902 44658 11954
rect 44942 11902 44994 11954
rect 49534 11902 49586 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 14254 11454 14306 11506
rect 18174 11454 18226 11506
rect 50990 11454 51042 11506
rect 14814 11342 14866 11394
rect 18734 11342 18786 11394
rect 24558 11342 24610 11394
rect 35086 11342 35138 11394
rect 47518 11342 47570 11394
rect 52558 11342 52610 11394
rect 54126 11342 54178 11394
rect 25118 11230 25170 11282
rect 35646 11230 35698 11282
rect 47070 11230 47122 11282
rect 51998 11230 52050 11282
rect 53566 11118 53618 11170
rect 55134 11118 55186 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 53006 10782 53058 10834
rect 28702 10670 28754 10722
rect 38558 10670 38610 10722
rect 54574 10670 54626 10722
rect 56142 10670 56194 10722
rect 29262 10558 29314 10610
rect 30830 10558 30882 10610
rect 34526 10558 34578 10610
rect 35086 10558 35138 10610
rect 52110 10558 52162 10610
rect 31390 10446 31442 10498
rect 53566 10446 53618 10498
rect 55134 10446 55186 10498
rect 37998 10334 38050 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 19406 9998 19458 10050
rect 32622 9886 32674 9938
rect 34638 9886 34690 9938
rect 35198 9886 35250 9938
rect 33182 9774 33234 9826
rect 52558 9774 52610 9826
rect 54238 9774 54290 9826
rect 19966 9662 20018 9714
rect 53566 9662 53618 9714
rect 55134 9550 55186 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 2942 9102 2994 9154
rect 28926 9102 28978 9154
rect 23214 8990 23266 9042
rect 25566 8990 25618 9042
rect 28590 8990 28642 9042
rect 55246 8990 55298 9042
rect 22654 8878 22706 8930
rect 26126 8878 26178 8930
rect 41694 8878 41746 8930
rect 44718 8878 44770 8930
rect 53566 8878 53618 8930
rect 54350 8878 54402 8930
rect 55918 8878 55970 8930
rect 2382 8766 2434 8818
rect 41134 8766 41186 8818
rect 44158 8766 44210 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 22430 8430 22482 8482
rect 30718 8430 30770 8482
rect 29262 8318 29314 8370
rect 29822 8318 29874 8370
rect 54126 8318 54178 8370
rect 54910 8318 54962 8370
rect 18286 8206 18338 8258
rect 43598 8206 43650 8258
rect 17838 8094 17890 8146
rect 22990 8094 23042 8146
rect 31166 8094 31218 8146
rect 44158 8094 44210 8146
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 56142 7646 56194 7698
rect 9214 7534 9266 7586
rect 26350 7534 26402 7586
rect 35646 7534 35698 7586
rect 54574 7534 54626 7586
rect 20862 7422 20914 7474
rect 25902 7422 25954 7474
rect 53566 7422 53618 7474
rect 55134 7422 55186 7474
rect 5406 7310 5458 7362
rect 21422 7310 21474 7362
rect 5966 7198 6018 7250
rect 9662 7198 9714 7250
rect 35086 7198 35138 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 16158 6750 16210 6802
rect 15598 6638 15650 6690
rect 26462 6638 26514 6690
rect 43262 6638 43314 6690
rect 44830 6638 44882 6690
rect 54126 6638 54178 6690
rect 27022 6526 27074 6578
rect 43710 6526 43762 6578
rect 45278 6526 45330 6578
rect 55134 6414 55186 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 56142 6078 56194 6130
rect 40462 5966 40514 6018
rect 54574 5966 54626 6018
rect 35758 5854 35810 5906
rect 40126 5854 40178 5906
rect 46622 5854 46674 5906
rect 49422 5854 49474 5906
rect 53566 5854 53618 5906
rect 55358 5854 55410 5906
rect 14254 5742 14306 5794
rect 17166 5742 17218 5794
rect 24446 5742 24498 5794
rect 24782 5742 24834 5794
rect 25342 5742 25394 5794
rect 37886 5742 37938 5794
rect 47182 5742 47234 5794
rect 49982 5742 50034 5794
rect 14814 5630 14866 5682
rect 16606 5630 16658 5682
rect 23886 5630 23938 5682
rect 35198 5630 35250 5682
rect 37326 5630 37378 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 18622 5294 18674 5346
rect 29822 5294 29874 5346
rect 32398 5294 32450 5346
rect 52894 5294 52946 5346
rect 53230 5294 53282 5346
rect 32958 5182 33010 5234
rect 52334 5182 52386 5234
rect 10894 5070 10946 5122
rect 20078 5070 20130 5122
rect 28926 5070 28978 5122
rect 34638 5070 34690 5122
rect 35198 5070 35250 5122
rect 38670 5070 38722 5122
rect 39118 5070 39170 5122
rect 42590 5070 42642 5122
rect 43150 5070 43202 5122
rect 47070 5070 47122 5122
rect 47518 5070 47570 5122
rect 54238 5070 54290 5122
rect 54910 5070 54962 5122
rect 10446 4958 10498 5010
rect 19182 4958 19234 5010
rect 19630 4958 19682 5010
rect 29486 4958 29538 5010
rect 30382 4958 30434 5010
rect 53790 4958 53842 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 54574 4510 54626 4562
rect 56142 4510 56194 4562
rect 11790 4398 11842 4450
rect 18174 4398 18226 4450
rect 24334 4398 24386 4450
rect 35646 4398 35698 4450
rect 36766 4398 36818 4450
rect 45390 4398 45442 4450
rect 52670 4398 52722 4450
rect 2606 4286 2658 4338
rect 32622 4286 32674 4338
rect 35310 4286 35362 4338
rect 39230 4286 39282 4338
rect 41470 4286 41522 4338
rect 44942 4286 44994 4338
rect 53678 4286 53730 4338
rect 55246 4286 55298 4338
rect 10110 4174 10162 4226
rect 33070 4174 33122 4226
rect 39790 4174 39842 4226
rect 42030 4174 42082 4226
rect 46622 4174 46674 4226
rect 3166 4062 3218 4114
rect 10670 4062 10722 4114
rect 12238 4062 12290 4114
rect 18622 4062 18674 4114
rect 23886 4062 23938 4114
rect 36318 4062 36370 4114
rect 47182 4062 47234 4114
rect 53230 4062 53282 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 27582 3726 27634 3778
rect 46510 3726 46562 3778
rect 49758 3726 49810 3778
rect 51326 3726 51378 3778
rect 24558 3614 24610 3666
rect 26014 3614 26066 3666
rect 37550 3614 37602 3666
rect 39118 3614 39170 3666
rect 41806 3614 41858 3666
rect 43374 3614 43426 3666
rect 49198 3614 49250 3666
rect 50766 3614 50818 3666
rect 51662 3614 51714 3666
rect 52558 3614 52610 3666
rect 54126 3614 54178 3666
rect 54910 3614 54962 3666
rect 23550 3502 23602 3554
rect 33406 3502 33458 3554
rect 35758 3502 35810 3554
rect 41358 3502 41410 3554
rect 45054 3502 45106 3554
rect 48302 3502 48354 3554
rect 48862 3502 48914 3554
rect 52222 3502 52274 3554
rect 23998 3390 24050 3442
rect 25006 3390 25058 3442
rect 28142 3390 28194 3442
rect 38222 3390 38274 3442
rect 40574 3390 40626 3442
rect 43934 3390 43986 3442
rect 46958 3390 47010 3442
rect 53566 3390 53618 3442
rect 26574 3278 26626 3330
rect 32622 3278 32674 3330
rect 34750 3278 34802 3330
rect 36542 3278 36594 3330
rect 42366 3278 42418 3330
rect 45502 3278 45554 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 54574 2942 54626 2994
rect 56142 2942 56194 2994
rect 30158 2830 30210 2882
rect 38110 2830 38162 2882
rect 41246 2830 41298 2882
rect 44830 2830 44882 2882
rect 53006 2830 53058 2882
rect 25230 2718 25282 2770
rect 30494 2718 30546 2770
rect 34862 2718 34914 2770
rect 35310 2718 35362 2770
rect 36318 2718 36370 2770
rect 39118 2718 39170 2770
rect 40686 2718 40738 2770
rect 42254 2718 42306 2770
rect 43038 2718 43090 2770
rect 44270 2718 44322 2770
rect 45726 2718 45778 2770
rect 47294 2718 47346 2770
rect 48974 2718 49026 2770
rect 50878 2718 50930 2770
rect 52110 2718 52162 2770
rect 53566 2718 53618 2770
rect 55134 2718 55186 2770
rect 14366 2606 14418 2658
rect 17838 2606 17890 2658
rect 26686 2606 26738 2658
rect 29262 2606 29314 2658
rect 32062 2606 32114 2658
rect 34078 2606 34130 2658
rect 35758 2606 35810 2658
rect 37102 2606 37154 2658
rect 39902 2606 39954 2658
rect 43598 2606 43650 2658
rect 51438 2606 51490 2658
rect 13806 2494 13858 2546
rect 17278 2494 17330 2546
rect 25678 2494 25730 2546
rect 27246 2494 27298 2546
rect 28702 2494 28754 2546
rect 29598 2494 29650 2546
rect 31054 2494 31106 2546
rect 32622 2494 32674 2546
rect 46286 2494 46338 2546
rect 47854 2494 47906 2546
rect 49422 2494 49474 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 19182 2158 19234 2210
rect 20862 2158 20914 2210
rect 25118 2158 25170 2210
rect 31278 2158 31330 2210
rect 1710 2046 1762 2098
rect 21422 2046 21474 2098
rect 22430 2046 22482 2098
rect 22766 2046 22818 2098
rect 26014 2046 26066 2098
rect 28814 2046 28866 2098
rect 30382 2046 30434 2098
rect 31838 2046 31890 2098
rect 32398 2046 32450 2098
rect 35198 2046 35250 2098
rect 41470 2046 41522 2098
rect 43374 2046 43426 2098
rect 44942 2046 44994 2098
rect 46510 2046 46562 2098
rect 48078 2046 48130 2098
rect 49646 2046 49698 2098
rect 51214 2046 51266 2098
rect 52558 2046 52610 2098
rect 54126 2046 54178 2098
rect 54910 2046 54962 2098
rect 2270 1934 2322 1986
rect 9550 1934 9602 1986
rect 21870 1934 21922 1986
rect 36766 1934 36818 1986
rect 38110 1934 38162 1986
rect 38670 1934 38722 1986
rect 39230 1934 39282 1986
rect 43038 1934 43090 1986
rect 47070 1934 47122 1986
rect 51774 1934 51826 1986
rect 9998 1822 10050 1874
rect 19742 1822 19794 1874
rect 25678 1822 25730 1874
rect 28030 1822 28082 1874
rect 32958 1822 33010 1874
rect 35758 1822 35810 1874
rect 45726 1822 45778 1874
rect 48750 1822 48802 1874
rect 50542 1822 50594 1874
rect 53566 1822 53618 1874
rect 23774 1710 23826 1762
rect 27022 1710 27074 1762
rect 29374 1710 29426 1762
rect 34190 1710 34242 1762
rect 37326 1710 37378 1762
rect 40462 1710 40514 1762
rect 42030 1710 42082 1762
rect 43934 1710 43986 1762
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 53566 1374 53618 1426
rect 56142 1374 56194 1426
rect 26910 1262 26962 1314
rect 40910 1262 40962 1314
rect 51998 1262 52050 1314
rect 22094 1150 22146 1202
rect 24334 1150 24386 1202
rect 26126 1150 26178 1202
rect 29150 1150 29202 1202
rect 29598 1150 29650 1202
rect 31502 1150 31554 1202
rect 33070 1150 33122 1202
rect 35310 1150 35362 1202
rect 37102 1150 37154 1202
rect 40126 1150 40178 1202
rect 41918 1150 41970 1202
rect 44158 1150 44210 1202
rect 44494 1150 44546 1202
rect 46734 1150 46786 1202
rect 48414 1150 48466 1202
rect 50990 1150 51042 1202
rect 52782 1150 52834 1202
rect 55134 1150 55186 1202
rect 22878 1038 22930 1090
rect 25118 1038 25170 1090
rect 28478 1038 28530 1090
rect 39566 1038 39618 1090
rect 43374 1038 43426 1090
rect 30158 926 30210 978
rect 32062 926 32114 978
rect 33630 926 33682 978
rect 35870 926 35922 978
rect 37438 926 37490 978
rect 45054 926 45106 978
rect 47294 926 47346 978
rect 48862 926 48914 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 1792 14112 1904 14224
rect 4480 14112 4592 14224
rect 7168 14112 7280 14224
rect 9856 14112 9968 14224
rect 12544 14112 12656 14224
rect 15232 14112 15344 14224
rect 17920 14112 18032 14224
rect 20608 14112 20720 14224
rect 23296 14112 23408 14224
rect 25984 14112 26096 14224
rect 28672 14112 28784 14224
rect 31360 14112 31472 14224
rect 34048 14112 34160 14224
rect 36736 14112 36848 14224
rect 39424 14112 39536 14224
rect 42112 14112 42224 14224
rect 44800 14112 44912 14224
rect 47488 14112 47600 14224
rect 50176 14112 50288 14224
rect 52864 14112 52976 14224
rect 55552 14112 55664 14224
rect 1820 13636 1876 14112
rect 4508 14084 4564 14112
rect 4508 14018 4564 14028
rect 5068 14084 5124 14094
rect 1820 13580 2100 13636
rect 2044 13186 2100 13580
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 2044 13134 2046 13186
rect 2098 13134 2100 13186
rect 2044 13122 2100 13134
rect 2380 12962 2436 12974
rect 2380 12910 2382 12962
rect 2434 12910 2436 12962
rect 1596 12628 1652 12638
rect 364 12180 420 12190
rect 364 10052 420 12124
rect 1596 11508 1652 12572
rect 1596 11442 1652 11452
rect 2380 10724 2436 12910
rect 5068 12850 5124 14028
rect 6860 13076 6916 13086
rect 5068 12798 5070 12850
rect 5122 12798 5124 12850
rect 5068 12786 5124 12798
rect 5292 12964 5348 12974
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 5292 11732 5348 12908
rect 6076 12962 6132 12974
rect 6076 12910 6078 12962
rect 6130 12910 6132 12962
rect 6076 12852 6132 12910
rect 6076 12786 6132 12796
rect 6860 11956 6916 13020
rect 7196 12850 7252 14112
rect 8092 14084 8148 14094
rect 7196 12798 7198 12850
rect 7250 12798 7252 12850
rect 7196 12786 7252 12798
rect 7308 13972 7364 13982
rect 6860 11890 6916 11900
rect 6972 12068 7028 12078
rect 5292 11666 5348 11676
rect 6636 11284 6692 11294
rect 6692 11228 6916 11284
rect 6636 11218 6692 11228
rect 2380 10658 2436 10668
rect 3052 11172 3108 11182
rect 364 9986 420 9996
rect 1596 9492 1652 9502
rect 1596 8372 1652 9436
rect 2940 9156 2996 9166
rect 2940 9062 2996 9100
rect 1596 8306 1652 8316
rect 2380 8818 2436 8830
rect 2380 8766 2382 8818
rect 2434 8766 2436 8818
rect 1148 5796 1204 5806
rect 700 2884 756 2894
rect 700 112 756 2828
rect 1148 112 1204 5740
rect 2044 5124 2100 5134
rect 1708 4452 1764 4462
rect 1708 2098 1764 4396
rect 1708 2046 1710 2098
rect 1762 2046 1764 2098
rect 1708 2034 1764 2046
rect 1820 2548 1876 2558
rect 1820 1316 1876 2492
rect 1596 1260 1876 1316
rect 1596 112 1652 1260
rect 2044 112 2100 5068
rect 2268 1986 2324 1998
rect 2268 1934 2270 1986
rect 2322 1934 2324 1986
rect 2268 1092 2324 1934
rect 2380 1876 2436 8766
rect 2828 5684 2884 5694
rect 2380 1810 2436 1820
rect 2492 5236 2548 5246
rect 2268 1026 2324 1036
rect 2492 112 2548 5180
rect 2604 4340 2660 4350
rect 2604 4246 2660 4284
rect 2828 2884 2884 5628
rect 2940 4116 2996 4126
rect 3052 4116 3108 11116
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 6748 10612 6804 10622
rect 3164 10388 3220 10398
rect 3164 8932 3220 10332
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 3164 8866 3220 8876
rect 3276 9940 3332 9950
rect 3276 8260 3332 9884
rect 6636 9492 6692 9502
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4956 9268 5012 9278
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3276 8194 3332 8204
rect 4284 7924 4340 7934
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3388 7588 3444 7598
rect 2996 4060 3108 4116
rect 3164 4116 3220 4126
rect 2940 4050 2996 4060
rect 3164 4022 3220 4060
rect 2828 2828 2996 2884
rect 2940 112 2996 2828
rect 3388 112 3444 7532
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 3836 1316 3892 1326
rect 3836 112 3892 1260
rect 4284 112 4340 7868
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4956 6804 5012 9212
rect 6412 8820 6468 8830
rect 5404 7364 5460 7374
rect 5404 7270 5460 7308
rect 4956 6738 5012 6748
rect 5964 7250 6020 7262
rect 5964 7198 5966 7250
rect 6018 7198 6020 7250
rect 5068 6580 5124 6590
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 5068 3668 5124 6524
rect 5964 6020 6020 7198
rect 5964 5954 6020 5964
rect 6076 4116 6132 4126
rect 5068 3602 5124 3612
rect 5628 3892 5684 3902
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 4844 2100 4900 2110
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 4844 644 4900 2044
rect 4732 588 4900 644
rect 5180 980 5236 990
rect 4732 112 4788 588
rect 5180 112 5236 924
rect 5628 112 5684 3836
rect 6076 2996 6132 4060
rect 6076 2930 6132 2940
rect 6188 4004 6244 4014
rect 6188 2772 6244 3948
rect 6076 2716 6244 2772
rect 6076 112 6132 2716
rect 6412 1316 6468 8764
rect 6636 8148 6692 9436
rect 6748 9156 6804 10556
rect 6860 9380 6916 11228
rect 6860 9314 6916 9324
rect 6748 9090 6804 9100
rect 6972 9044 7028 12012
rect 6972 8978 7028 8988
rect 7084 11172 7140 11182
rect 6860 8708 6916 8718
rect 6860 8428 6916 8652
rect 6748 8372 6916 8428
rect 6748 8306 6804 8316
rect 6636 8082 6692 8092
rect 6972 8148 7028 8158
rect 6748 7700 6804 7710
rect 6636 5348 6692 5358
rect 6636 4452 6692 5292
rect 6748 4676 6804 7644
rect 6748 4610 6804 4620
rect 6860 6132 6916 6142
rect 6636 4396 6804 4452
rect 6748 2212 6804 4396
rect 6860 2436 6916 6076
rect 6972 5684 7028 8092
rect 7084 5908 7140 11116
rect 7308 10948 7364 13916
rect 7308 10882 7364 10892
rect 7644 13188 7700 13198
rect 7084 5842 7140 5852
rect 7196 10724 7252 10734
rect 6972 5628 7140 5684
rect 6860 2370 6916 2380
rect 6972 5460 7028 5470
rect 6748 2146 6804 2156
rect 6972 2100 7028 5404
rect 6972 2034 7028 2044
rect 7084 1876 7140 5628
rect 7196 4228 7252 10668
rect 7420 7812 7476 7822
rect 7196 4162 7252 4172
rect 7308 6916 7364 6926
rect 7308 2660 7364 6860
rect 7420 4004 7476 7756
rect 7532 7476 7588 7486
rect 7532 5796 7588 7420
rect 7532 5730 7588 5740
rect 7532 5572 7588 5582
rect 7532 5124 7588 5516
rect 7532 5058 7588 5068
rect 7420 3938 7476 3948
rect 7644 3332 7700 13132
rect 8092 13074 8148 14028
rect 9884 13636 9940 14112
rect 9884 13570 9940 13580
rect 10668 13636 10724 13646
rect 10668 13186 10724 13580
rect 10668 13134 10670 13186
rect 10722 13134 10724 13186
rect 10668 13122 10724 13134
rect 8092 13022 8094 13074
rect 8146 13022 8148 13074
rect 8092 13010 8148 13022
rect 10332 12962 10388 12974
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 10332 12292 10388 12910
rect 12572 12852 12628 14112
rect 13356 13972 13412 13982
rect 13020 12852 13076 12862
rect 12572 12850 13076 12852
rect 12572 12798 13022 12850
rect 13074 12798 13076 12850
rect 12572 12796 13076 12798
rect 13020 12786 13076 12796
rect 10444 12292 10500 12302
rect 10332 12290 10500 12292
rect 10332 12238 10446 12290
rect 10498 12238 10500 12290
rect 10332 12236 10500 12238
rect 10444 12226 10500 12236
rect 11004 12292 11060 12302
rect 11004 12178 11060 12236
rect 11004 12126 11006 12178
rect 11058 12126 11060 12178
rect 11004 12114 11060 12126
rect 11228 11956 11284 11966
rect 8540 10276 8596 10286
rect 8428 10164 8484 10174
rect 8428 8260 8484 10108
rect 8428 8194 8484 8204
rect 8540 6580 8596 10220
rect 9212 10052 9268 10062
rect 9212 7586 9268 9996
rect 9212 7534 9214 7586
rect 9266 7534 9268 7586
rect 9212 7522 9268 7534
rect 10108 8484 10164 8494
rect 9660 7252 9716 7262
rect 9660 7158 9716 7196
rect 8540 6514 8596 6524
rect 7644 3266 7700 3276
rect 7756 5236 7812 5246
rect 10108 5236 10164 8428
rect 7308 2594 7364 2604
rect 7420 3108 7476 3118
rect 6412 1250 6468 1260
rect 6972 1820 7140 1876
rect 6524 1204 6580 1214
rect 6524 112 6580 1148
rect 6972 112 7028 1820
rect 7420 112 7476 3052
rect 7756 2884 7812 5180
rect 9996 5180 10164 5236
rect 10556 5348 10612 5358
rect 9996 4564 10052 5180
rect 9996 4498 10052 4508
rect 10444 5010 10500 5022
rect 10444 4958 10446 5010
rect 10498 4958 10500 5010
rect 10108 4228 10164 4238
rect 10108 4226 10388 4228
rect 10108 4174 10110 4226
rect 10162 4174 10388 4226
rect 10108 4172 10388 4174
rect 10108 4162 10164 4172
rect 9660 4116 9716 4126
rect 9212 3780 9268 3790
rect 7756 2818 7812 2828
rect 8316 2884 8372 2894
rect 7868 1652 7924 1662
rect 7868 112 7924 1596
rect 8316 112 8372 2828
rect 8764 1316 8820 1326
rect 8764 112 8820 1260
rect 9212 112 9268 3724
rect 9548 1986 9604 1998
rect 9548 1934 9550 1986
rect 9602 1934 9604 1986
rect 9548 868 9604 1934
rect 9548 802 9604 812
rect 9660 112 9716 4060
rect 10332 3332 10388 4172
rect 10444 3556 10500 4958
rect 10444 3490 10500 3500
rect 10332 3266 10388 3276
rect 10556 3108 10612 5292
rect 10892 5122 10948 5134
rect 10892 5070 10894 5122
rect 10946 5070 10948 5122
rect 10108 3052 10612 3108
rect 10668 4114 10724 4126
rect 10668 4062 10670 4114
rect 10722 4062 10724 4114
rect 9996 1876 10052 1886
rect 9996 1782 10052 1820
rect 10108 112 10164 3052
rect 10556 868 10612 878
rect 10556 112 10612 812
rect 10668 644 10724 4062
rect 10668 578 10724 588
rect 10892 420 10948 5070
rect 10892 354 10948 364
rect 11004 5012 11060 5022
rect 11004 112 11060 4956
rect 11228 4116 11284 11900
rect 13356 9940 13412 13916
rect 15036 13636 15092 13646
rect 14028 12964 14084 12974
rect 14028 12962 14308 12964
rect 14028 12910 14030 12962
rect 14082 12910 14308 12962
rect 14028 12908 14308 12910
rect 14028 12898 14084 12908
rect 13468 11620 13524 11630
rect 13468 10052 13524 11564
rect 14252 11506 14308 12908
rect 15036 12290 15092 13580
rect 15260 12404 15316 14112
rect 15820 13860 15876 13870
rect 15708 12404 15764 12414
rect 15260 12402 15764 12404
rect 15260 12350 15710 12402
rect 15762 12350 15764 12402
rect 15260 12348 15764 12350
rect 15708 12338 15764 12348
rect 15036 12238 15038 12290
rect 15090 12238 15092 12290
rect 15036 12226 15092 12238
rect 14252 11454 14254 11506
rect 14306 11454 14308 11506
rect 14252 11442 14308 11454
rect 14364 12180 14420 12190
rect 13468 9986 13524 9996
rect 13916 10164 13972 10174
rect 13356 9874 13412 9884
rect 13916 9268 13972 10108
rect 13916 9202 13972 9212
rect 14252 9716 14308 9726
rect 13468 9156 13524 9166
rect 13356 7700 13412 7710
rect 12796 7028 12852 7038
rect 11788 4452 11844 4462
rect 11788 4358 11844 4396
rect 11228 4050 11284 4060
rect 12236 4116 12292 4126
rect 12236 4022 12292 4060
rect 12348 3668 12404 3678
rect 11676 3444 11732 3454
rect 11452 1652 11508 1662
rect 11452 112 11508 1596
rect 11564 1204 11620 1214
rect 11564 980 11620 1148
rect 11564 914 11620 924
rect 11676 756 11732 3388
rect 11676 690 11732 700
rect 11900 1204 11956 1214
rect 11900 112 11956 1148
rect 12348 112 12404 3612
rect 12796 868 12852 6972
rect 13356 3780 13412 7644
rect 13468 4452 13524 9100
rect 13916 8148 13972 8158
rect 13692 6244 13748 6254
rect 13468 4386 13524 4396
rect 13580 5796 13636 5806
rect 13356 3714 13412 3724
rect 13580 3332 13636 5740
rect 13692 3668 13748 6188
rect 13916 4788 13972 8092
rect 14252 6020 14308 9660
rect 14364 8428 14420 12124
rect 14588 11954 14644 11966
rect 14588 11902 14590 11954
rect 14642 11902 14644 11954
rect 14588 11284 14644 11902
rect 14588 11218 14644 11228
rect 14812 11394 14868 11406
rect 14812 11342 14814 11394
rect 14866 11342 14868 11394
rect 14700 11060 14756 11070
rect 14476 10948 14532 10958
rect 14476 9716 14532 10892
rect 14476 9650 14532 9660
rect 14588 10612 14644 10622
rect 14364 8372 14532 8428
rect 14252 5954 14308 5964
rect 13916 4722 13972 4732
rect 14140 5908 14196 5918
rect 14140 3780 14196 5852
rect 14252 5794 14308 5806
rect 14252 5742 14254 5794
rect 14306 5742 14308 5794
rect 14252 4452 14308 5742
rect 14476 5348 14532 8372
rect 14588 7588 14644 10556
rect 14588 7522 14644 7532
rect 14476 5282 14532 5292
rect 14588 6804 14644 6814
rect 14252 4386 14308 4396
rect 14140 3714 14196 3724
rect 14252 4004 14308 4014
rect 13692 3602 13748 3612
rect 13580 3266 13636 3276
rect 14140 3332 14196 3342
rect 13916 2660 13972 2670
rect 13804 2546 13860 2558
rect 13804 2494 13806 2546
rect 13858 2494 13860 2546
rect 13804 1316 13860 2494
rect 13804 1250 13860 1260
rect 12796 802 12852 812
rect 13692 1204 13748 1214
rect 13244 756 13300 766
rect 12796 196 12852 206
rect 12796 112 12852 140
rect 13244 112 13300 700
rect 13692 112 13748 1148
rect 672 0 784 112
rect 1120 0 1232 112
rect 1568 0 1680 112
rect 2016 0 2128 112
rect 2464 0 2576 112
rect 2912 0 3024 112
rect 3360 0 3472 112
rect 3808 0 3920 112
rect 4256 0 4368 112
rect 4704 0 4816 112
rect 5152 0 5264 112
rect 5600 0 5712 112
rect 6048 0 6160 112
rect 6496 0 6608 112
rect 6944 0 7056 112
rect 7392 0 7504 112
rect 7840 0 7952 112
rect 8288 0 8400 112
rect 8736 0 8848 112
rect 9184 0 9296 112
rect 9632 0 9744 112
rect 10080 0 10192 112
rect 10528 0 10640 112
rect 10976 0 11088 112
rect 11424 0 11536 112
rect 11872 0 11984 112
rect 12320 0 12432 112
rect 12768 0 12880 112
rect 13216 0 13328 112
rect 13664 0 13776 112
rect 13916 84 13972 2604
rect 14140 2212 14196 3276
rect 14252 3108 14308 3948
rect 14252 3042 14308 3052
rect 14364 2658 14420 2670
rect 14364 2606 14366 2658
rect 14418 2606 14420 2658
rect 14364 2324 14420 2606
rect 14364 2258 14420 2268
rect 14140 2146 14196 2156
rect 14476 2212 14532 2222
rect 14140 1988 14196 1998
rect 14140 112 14196 1932
rect 14476 532 14532 2156
rect 14476 466 14532 476
rect 14588 112 14644 6748
rect 14700 5124 14756 11004
rect 14812 9604 14868 11342
rect 14924 10948 14980 10958
rect 14924 10276 14980 10892
rect 14924 10210 14980 10220
rect 15148 10388 15204 10398
rect 14812 9538 14868 9548
rect 14924 9492 14980 9502
rect 14924 8372 14980 9436
rect 15148 8428 15204 10332
rect 14924 8306 14980 8316
rect 15036 8372 15204 8428
rect 15036 7812 15092 8372
rect 15036 7746 15092 7756
rect 15036 7140 15092 7150
rect 14700 5058 14756 5068
rect 14812 5682 14868 5694
rect 14812 5630 14814 5682
rect 14866 5630 14868 5682
rect 14700 2996 14756 3006
rect 14700 1652 14756 2940
rect 14700 1586 14756 1596
rect 14812 1316 14868 5630
rect 14812 1250 14868 1260
rect 15036 112 15092 7084
rect 15260 6916 15316 6926
rect 15260 5012 15316 6860
rect 15260 4946 15316 4956
rect 15596 6690 15652 6702
rect 15596 6638 15598 6690
rect 15650 6638 15652 6690
rect 15596 2436 15652 6638
rect 15820 3388 15876 13804
rect 17948 13412 18004 14112
rect 17948 13356 18452 13412
rect 18396 12850 18452 13356
rect 18396 12798 18398 12850
rect 18450 12798 18452 12850
rect 18396 12786 18452 12798
rect 19404 12962 19460 12974
rect 19404 12910 19406 12962
rect 19458 12910 19460 12962
rect 18284 12740 18340 12750
rect 16492 12068 16548 12078
rect 16492 10724 16548 12012
rect 16716 12068 16772 12078
rect 16716 11974 16772 12012
rect 18172 12068 18228 12078
rect 17052 11844 17108 11854
rect 16828 11620 16884 11630
rect 17052 11620 17108 11788
rect 16884 11564 17108 11620
rect 17276 11620 17332 11630
rect 16828 11554 16884 11564
rect 16492 10658 16548 10668
rect 16716 11172 16772 11182
rect 15932 10276 15988 10286
rect 15932 6804 15988 10220
rect 16716 10052 16772 11116
rect 17276 10836 17332 11564
rect 18172 11506 18228 12012
rect 18172 11454 18174 11506
rect 18226 11454 18228 11506
rect 18172 11442 18228 11454
rect 18284 11396 18340 12684
rect 18396 12292 18452 12302
rect 18396 11732 18452 12236
rect 19404 12292 19460 12910
rect 20636 12852 20692 14112
rect 21196 13748 21252 13758
rect 21084 12852 21140 12862
rect 20636 12850 21140 12852
rect 20636 12798 21086 12850
rect 21138 12798 21140 12850
rect 20636 12796 21140 12798
rect 21084 12786 21140 12796
rect 19404 12226 19460 12236
rect 20636 12292 20692 12302
rect 20636 12198 20692 12236
rect 20972 12180 21028 12190
rect 18396 11666 18452 11676
rect 18620 11956 18676 11966
rect 18508 11396 18564 11406
rect 18284 11330 18340 11340
rect 18396 11340 18508 11396
rect 18172 11172 18228 11182
rect 17276 10770 17332 10780
rect 18060 10836 18116 10846
rect 16716 9986 16772 9996
rect 15932 6738 15988 6748
rect 16044 8260 16100 8270
rect 15820 3332 15988 3388
rect 15932 2884 15988 3332
rect 15932 2818 15988 2828
rect 15596 2370 15652 2380
rect 16044 2100 16100 8204
rect 17836 8146 17892 8158
rect 17836 8094 17838 8146
rect 17890 8094 17892 8146
rect 17836 8036 17892 8094
rect 17836 7970 17892 7980
rect 16380 7476 16436 7486
rect 16156 6804 16212 6814
rect 16156 6710 16212 6748
rect 16380 5348 16436 7420
rect 17724 7252 17780 7262
rect 16716 6132 16772 6142
rect 16604 5682 16660 5694
rect 16604 5630 16606 5682
rect 16658 5630 16660 5682
rect 16604 5572 16660 5630
rect 16604 5506 16660 5516
rect 16380 5282 16436 5292
rect 16044 2034 16100 2044
rect 16492 4900 16548 4910
rect 16492 1988 16548 4844
rect 16492 1922 16548 1932
rect 15260 1428 15316 1438
rect 15260 532 15316 1372
rect 16380 1092 16436 1102
rect 15260 466 15316 476
rect 15932 868 15988 878
rect 15484 252 15764 308
rect 15484 112 15540 252
rect 13916 18 13972 28
rect 14112 0 14224 112
rect 14560 0 14672 112
rect 15008 0 15120 112
rect 15456 0 15568 112
rect 15708 84 15764 252
rect 15932 112 15988 812
rect 16380 112 16436 1036
rect 16716 1092 16772 6076
rect 17164 5794 17220 5806
rect 17164 5742 17166 5794
rect 17218 5742 17220 5794
rect 16828 4116 16884 4126
rect 16828 2100 16884 4060
rect 16828 2034 16884 2044
rect 16940 2996 16996 3006
rect 16716 1026 16772 1036
rect 16828 1652 16884 1662
rect 16828 112 16884 1596
rect 16940 1204 16996 2940
rect 17164 1988 17220 5742
rect 17276 2548 17332 2558
rect 17276 2454 17332 2492
rect 17164 1922 17220 1932
rect 16940 1138 16996 1148
rect 17276 1092 17332 1102
rect 17276 112 17332 1036
rect 17724 112 17780 7196
rect 18060 5124 18116 10780
rect 18172 5796 18228 11116
rect 18396 10836 18452 11340
rect 18508 11330 18564 11340
rect 18396 10770 18452 10780
rect 18284 10724 18340 10734
rect 18284 9716 18340 10668
rect 18620 10724 18676 11900
rect 20076 11844 20132 11854
rect 20076 11508 20132 11788
rect 20076 11442 20132 11452
rect 18732 11394 18788 11406
rect 18732 11342 18734 11394
rect 18786 11342 18788 11394
rect 18732 10836 18788 11342
rect 18732 10770 18788 10780
rect 19852 11284 19908 11294
rect 18620 10658 18676 10668
rect 18284 9650 18340 9660
rect 18396 10500 18452 10510
rect 18396 9044 18452 10444
rect 19404 10164 19460 10174
rect 19404 10050 19460 10108
rect 19404 9998 19406 10050
rect 19458 9998 19460 10050
rect 19404 9986 19460 9998
rect 18396 8978 18452 8988
rect 18172 5730 18228 5740
rect 18284 8258 18340 8270
rect 18284 8206 18286 8258
rect 18338 8206 18340 8258
rect 18060 5058 18116 5068
rect 18172 5572 18228 5582
rect 18172 4450 18228 5516
rect 18172 4398 18174 4450
rect 18226 4398 18228 4450
rect 18172 4386 18228 4398
rect 17836 4116 17892 4126
rect 17836 3444 17892 4060
rect 17836 3378 17892 3388
rect 17836 2658 17892 2670
rect 17836 2606 17838 2658
rect 17890 2606 17892 2658
rect 17836 1204 17892 2606
rect 18284 1652 18340 8206
rect 18508 6692 18564 6702
rect 18396 4228 18452 4238
rect 18508 4228 18564 6636
rect 19852 6356 19908 11228
rect 20748 11060 20804 11070
rect 19964 9714 20020 9726
rect 19964 9662 19966 9714
rect 20018 9662 20020 9714
rect 19964 8372 20020 9662
rect 20748 8596 20804 11004
rect 20972 9044 21028 12124
rect 21196 12178 21252 13692
rect 23324 13412 23380 14112
rect 23324 13346 23380 13356
rect 23548 13524 23604 13534
rect 22092 12964 22148 12974
rect 22092 12962 22372 12964
rect 22092 12910 22094 12962
rect 22146 12910 22372 12962
rect 22092 12908 22372 12910
rect 22092 12898 22148 12908
rect 21980 12852 22036 12862
rect 21196 12126 21198 12178
rect 21250 12126 21252 12178
rect 21196 12114 21252 12126
rect 21868 12404 21924 12414
rect 21868 11732 21924 12348
rect 21868 11666 21924 11676
rect 21980 11396 22036 12796
rect 22316 12290 22372 12908
rect 22316 12238 22318 12290
rect 22370 12238 22372 12290
rect 22316 12226 22372 12238
rect 22428 12852 22484 12862
rect 21980 11330 22036 11340
rect 22092 11844 22148 11854
rect 20972 8978 21028 8988
rect 21196 10724 21252 10734
rect 20748 8530 20804 8540
rect 19964 8306 20020 8316
rect 20860 8484 20916 8494
rect 20860 7474 20916 8428
rect 20860 7422 20862 7474
rect 20914 7422 20916 7474
rect 20860 7410 20916 7422
rect 20636 7140 20692 7150
rect 19852 6290 19908 6300
rect 19964 6916 20020 6926
rect 19964 6244 20020 6860
rect 20076 6804 20132 6814
rect 20076 6468 20132 6748
rect 20076 6402 20132 6412
rect 19964 6178 20020 6188
rect 19964 6020 20020 6030
rect 18620 5348 18676 5358
rect 18620 5254 18676 5292
rect 19180 5010 19236 5022
rect 19180 4958 19182 5010
rect 19234 4958 19236 5010
rect 18452 4172 18564 4228
rect 18732 4564 18788 4574
rect 18396 4162 18452 4172
rect 18620 4114 18676 4126
rect 18620 4062 18622 4114
rect 18674 4062 18676 4114
rect 18620 1764 18676 4062
rect 18732 3108 18788 4508
rect 18732 3042 18788 3052
rect 19180 2660 19236 4958
rect 19180 2594 19236 2604
rect 19628 5010 19684 5022
rect 19628 4958 19630 5010
rect 19682 4958 19684 5010
rect 19180 2436 19236 2446
rect 19180 2210 19236 2380
rect 19180 2158 19182 2210
rect 19234 2158 19236 2210
rect 19180 2146 19236 2158
rect 18620 1698 18676 1708
rect 19068 2100 19124 2110
rect 18284 1586 18340 1596
rect 17836 1138 17892 1148
rect 18172 644 18228 654
rect 18172 112 18228 588
rect 18620 420 18676 430
rect 18620 112 18676 364
rect 19068 112 19124 2044
rect 19516 1316 19572 1326
rect 19516 112 19572 1260
rect 19628 308 19684 4958
rect 19964 3668 20020 5964
rect 20636 6020 20692 7084
rect 20636 5954 20692 5964
rect 20972 5908 21028 5918
rect 20860 5236 20916 5246
rect 20076 5124 20132 5134
rect 20076 5030 20132 5068
rect 20636 5124 20692 5134
rect 19964 3602 20020 3612
rect 20188 3556 20244 3566
rect 19852 3444 19908 3454
rect 19852 2884 19908 3388
rect 19852 2818 19908 2828
rect 20188 2884 20244 3500
rect 20188 2818 20244 2828
rect 20636 1988 20692 5068
rect 20860 2210 20916 5180
rect 20972 4116 21028 5852
rect 21196 5348 21252 10668
rect 21868 10724 21924 10734
rect 21644 10164 21700 10174
rect 21420 7364 21476 7374
rect 21420 7270 21476 7308
rect 21196 5282 21252 5292
rect 21532 6804 21588 6814
rect 20972 4050 21028 4060
rect 21420 4116 21476 4126
rect 20860 2158 20862 2210
rect 20914 2158 20916 2210
rect 20860 2146 20916 2158
rect 21420 2098 21476 4060
rect 21532 3332 21588 6748
rect 21644 5572 21700 10108
rect 21868 8428 21924 10668
rect 21756 8372 21924 8428
rect 21756 6580 21812 8372
rect 22092 7588 22148 11788
rect 22204 11284 22260 11294
rect 22204 9604 22260 11228
rect 22428 9828 22484 12796
rect 22876 12180 22932 12190
rect 22876 12086 22932 12124
rect 23548 12178 23604 13468
rect 24108 13412 24164 13422
rect 24108 12850 24164 13356
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24108 12798 24110 12850
rect 24162 12798 24164 12850
rect 24108 12786 24164 12798
rect 25116 12962 25172 12974
rect 25116 12910 25118 12962
rect 25170 12910 25172 12962
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 23548 12126 23550 12178
rect 23602 12126 23604 12178
rect 23548 12114 23604 12126
rect 24332 12292 24388 12302
rect 23996 12068 24052 12078
rect 23996 12066 24276 12068
rect 23996 12014 23998 12066
rect 24050 12014 24276 12066
rect 23996 12012 24276 12014
rect 23996 12002 24052 12012
rect 23548 11956 23604 11966
rect 23548 10164 23604 11900
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23548 10098 23604 10108
rect 22428 9762 22484 9772
rect 24220 9828 24276 12012
rect 24332 11060 24388 12236
rect 25116 12292 25172 12910
rect 26012 12852 26068 14112
rect 28588 13076 28644 13086
rect 27132 12962 27188 12974
rect 27132 12910 27134 12962
rect 27186 12910 27188 12962
rect 26124 12852 26180 12862
rect 26012 12850 26180 12852
rect 26012 12798 26126 12850
rect 26178 12798 26180 12850
rect 26012 12796 26180 12798
rect 26124 12786 26180 12796
rect 25116 12226 25172 12236
rect 26460 12292 26516 12302
rect 26460 12198 26516 12236
rect 26124 12068 26180 12078
rect 26124 12066 26292 12068
rect 26124 12014 26126 12066
rect 26178 12014 26292 12066
rect 26124 12012 26292 12014
rect 26124 12002 26180 12012
rect 25564 11954 25620 11966
rect 25564 11902 25566 11954
rect 25618 11902 25620 11954
rect 24892 11844 24948 11854
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24892 11508 24948 11788
rect 24892 11442 24948 11452
rect 24332 10994 24388 11004
rect 24556 11394 24612 11406
rect 24556 11342 24558 11394
rect 24610 11342 24612 11394
rect 24556 10724 24612 11342
rect 25116 11284 25172 11294
rect 25116 11282 25284 11284
rect 25116 11230 25118 11282
rect 25170 11230 25284 11282
rect 25116 11228 25284 11230
rect 25116 11218 25172 11228
rect 24556 10658 24612 10668
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 25116 10164 25172 10174
rect 24220 9762 24276 9772
rect 25116 9716 25172 10108
rect 25116 9650 25172 9660
rect 22204 9538 22260 9548
rect 24220 9492 24276 9502
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 22092 7522 22148 7532
rect 22204 9044 22260 9054
rect 21756 6514 21812 6524
rect 21980 6580 22036 6590
rect 21980 6356 22036 6524
rect 21980 6290 22036 6300
rect 21644 5506 21700 5516
rect 22204 5572 22260 8988
rect 23212 9044 23268 9054
rect 23212 8950 23268 8988
rect 22652 8932 22708 8942
rect 22652 8838 22708 8876
rect 22428 8708 22484 8718
rect 22428 8482 22484 8652
rect 22428 8430 22430 8482
rect 22482 8430 22484 8482
rect 22428 8418 22484 8430
rect 24220 8372 24276 9436
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24220 8306 24276 8316
rect 22988 8146 23044 8158
rect 22988 8094 22990 8146
rect 23042 8094 23044 8146
rect 22988 7476 23044 8094
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 24108 7700 24164 7710
rect 24668 7700 24724 7710
rect 24164 7644 24668 7700
rect 24108 7634 24164 7644
rect 24668 7634 24724 7644
rect 25228 7588 25284 11228
rect 25564 10052 25620 11902
rect 25564 9986 25620 9996
rect 25564 9156 25620 9166
rect 25564 9042 25620 9100
rect 25564 8990 25566 9042
rect 25618 8990 25620 9042
rect 25564 8978 25620 8990
rect 26124 8932 26180 8942
rect 26124 8838 26180 8876
rect 25228 7522 25284 7532
rect 25900 8148 25956 8158
rect 22988 7410 23044 7420
rect 25900 7474 25956 8092
rect 26236 7924 26292 12012
rect 27020 11954 27076 11966
rect 27020 11902 27022 11954
rect 27074 11902 27076 11954
rect 27020 11508 27076 11902
rect 27020 11442 27076 11452
rect 27132 10724 27188 12910
rect 28588 12178 28644 13020
rect 28700 12852 28756 14112
rect 29708 13860 29764 13870
rect 29148 12852 29204 12862
rect 28700 12850 29204 12852
rect 28700 12798 29150 12850
rect 29202 12798 29204 12850
rect 28700 12796 29204 12798
rect 29148 12786 29204 12796
rect 28588 12126 28590 12178
rect 28642 12126 28644 12178
rect 28588 12114 28644 12126
rect 29036 12180 29092 12190
rect 29036 12086 29092 12124
rect 29484 11956 29540 11966
rect 27132 10658 27188 10668
rect 28140 11844 28196 11854
rect 26796 9940 26852 9950
rect 26796 8428 26852 9884
rect 26796 8372 26964 8428
rect 26908 8306 26964 8316
rect 26236 7858 26292 7868
rect 26796 8260 26852 8270
rect 26348 7588 26404 7598
rect 25900 7422 25902 7474
rect 25954 7422 25956 7474
rect 25900 7410 25956 7422
rect 26124 7586 26404 7588
rect 26124 7534 26350 7586
rect 26402 7534 26404 7586
rect 26124 7532 26404 7534
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 24892 7028 24948 7038
rect 24220 6804 24276 6814
rect 24220 6356 24276 6748
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24220 6290 24276 6300
rect 23804 6234 24068 6244
rect 23772 6020 23828 6030
rect 22204 5506 22260 5516
rect 22652 5796 22708 5806
rect 21532 3266 21588 3276
rect 21644 5236 21700 5246
rect 21420 2046 21422 2098
rect 21474 2046 21476 2098
rect 21420 2034 21476 2046
rect 21532 3108 21588 3118
rect 21308 1988 21364 1998
rect 20636 1932 20916 1988
rect 19740 1874 19796 1886
rect 19740 1822 19742 1874
rect 19794 1822 19796 1874
rect 19740 1316 19796 1822
rect 19740 1250 19796 1260
rect 19964 1652 20020 1662
rect 19628 242 19684 252
rect 19964 112 20020 1596
rect 20412 1652 20468 1662
rect 20412 112 20468 1596
rect 20860 112 20916 1932
rect 21308 112 21364 1932
rect 21532 420 21588 3052
rect 21644 2996 21700 5180
rect 22428 4564 22484 4574
rect 22204 3668 22260 3678
rect 21644 2930 21700 2940
rect 21756 3556 21812 3566
rect 21644 2436 21700 2446
rect 21644 868 21700 2380
rect 21644 802 21700 812
rect 21532 354 21588 364
rect 21756 112 21812 3500
rect 21868 1988 21924 1998
rect 21868 1894 21924 1932
rect 22092 1204 22148 1214
rect 22092 1110 22148 1148
rect 22204 112 22260 3612
rect 22428 2098 22484 4508
rect 22428 2046 22430 2098
rect 22482 2046 22484 2098
rect 22428 2034 22484 2046
rect 22652 112 22708 5740
rect 23772 5572 23828 5964
rect 24892 5908 24948 6972
rect 25452 6916 25508 6926
rect 25452 6692 25508 6860
rect 25452 6626 25508 6636
rect 24892 5842 24948 5852
rect 24444 5794 24500 5806
rect 24444 5742 24446 5794
rect 24498 5742 24500 5794
rect 23772 5506 23828 5516
rect 23884 5682 23940 5694
rect 23884 5630 23886 5682
rect 23938 5630 23940 5682
rect 23884 5460 23940 5630
rect 24444 5684 24500 5742
rect 24780 5796 24836 5806
rect 24780 5702 24836 5740
rect 25340 5796 25396 5806
rect 25340 5702 25396 5740
rect 24444 5618 24500 5628
rect 25900 5684 25956 5694
rect 25228 5572 25284 5582
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24892 5460 24948 5470
rect 23884 5394 23940 5404
rect 23772 5348 23828 5358
rect 24892 5348 24948 5404
rect 23772 5236 23828 5292
rect 23996 5292 24948 5348
rect 23996 5236 24052 5292
rect 23772 5180 24052 5236
rect 23100 5124 23156 5134
rect 22764 2100 22820 2110
rect 22764 2006 22820 2044
rect 22876 1092 22932 1102
rect 22876 998 22932 1036
rect 23100 112 23156 5068
rect 23324 5012 23380 5022
rect 23380 4956 23492 5012
rect 23324 4946 23380 4956
rect 23324 4788 23380 4798
rect 23324 1428 23380 4732
rect 23436 2996 23492 4956
rect 25116 4900 25172 4910
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24892 4564 24948 4574
rect 24332 4450 24388 4462
rect 24332 4398 24334 4450
rect 24386 4398 24388 4450
rect 23884 4114 23940 4126
rect 23884 4062 23886 4114
rect 23938 4062 23940 4114
rect 23884 3892 23940 4062
rect 23884 3826 23940 3836
rect 23548 3556 23604 3566
rect 23548 3462 23604 3500
rect 23996 3444 24052 3482
rect 23996 3378 24052 3388
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24220 3108 24276 3118
rect 23436 2930 23492 2940
rect 23996 2772 24052 2782
rect 23996 2100 24052 2716
rect 24220 2436 24276 3052
rect 24220 2370 24276 2380
rect 23996 2034 24052 2044
rect 23324 1362 23380 1372
rect 23548 1988 23604 1998
rect 23548 112 23604 1932
rect 23772 1764 23828 1774
rect 23772 1762 24276 1764
rect 23772 1710 23774 1762
rect 23826 1710 24276 1762
rect 23772 1708 24276 1710
rect 23772 1698 23828 1708
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 24220 644 24276 1708
rect 24332 1202 24388 4398
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 24556 3668 24612 3678
rect 24556 3574 24612 3612
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24892 1988 24948 4508
rect 25116 4116 25172 4844
rect 25228 4340 25284 5516
rect 25340 5236 25396 5246
rect 25340 4900 25396 5180
rect 25340 4834 25396 4844
rect 25228 4274 25284 4284
rect 25676 4676 25732 4686
rect 25676 4228 25732 4620
rect 25676 4162 25732 4172
rect 25116 4060 25396 4116
rect 25228 3556 25284 3566
rect 24892 1922 24948 1932
rect 25004 3442 25060 3454
rect 25004 3390 25006 3442
rect 25058 3390 25060 3442
rect 24332 1150 24334 1202
rect 24386 1150 24388 1202
rect 24332 1138 24388 1150
rect 24892 1092 24948 1102
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24220 588 24500 644
rect 24444 112 24500 588
rect 24892 112 24948 1036
rect 25004 644 25060 3390
rect 25228 2996 25284 3500
rect 25340 3220 25396 4060
rect 25340 3154 25396 3164
rect 25116 2940 25284 2996
rect 25116 2210 25172 2940
rect 25228 2770 25284 2782
rect 25228 2718 25230 2770
rect 25282 2718 25284 2770
rect 25228 2660 25284 2718
rect 25228 2594 25284 2604
rect 25676 2548 25732 2558
rect 25116 2158 25118 2210
rect 25170 2158 25172 2210
rect 25116 2146 25172 2158
rect 25340 2546 25732 2548
rect 25340 2494 25678 2546
rect 25730 2494 25732 2546
rect 25340 2492 25732 2494
rect 25116 1092 25172 1102
rect 25116 998 25172 1036
rect 25004 578 25060 588
rect 25340 112 25396 2492
rect 25676 2482 25732 2492
rect 25900 2100 25956 5628
rect 26012 4116 26068 4126
rect 26012 3666 26068 4060
rect 26012 3614 26014 3666
rect 26066 3614 26068 3666
rect 26012 3602 26068 3614
rect 26012 2100 26068 2110
rect 25900 2098 26068 2100
rect 25900 2046 26014 2098
rect 26066 2046 26068 2098
rect 25900 2044 26068 2046
rect 26012 2034 26068 2044
rect 25676 1874 25732 1886
rect 25676 1822 25678 1874
rect 25730 1822 25732 1874
rect 25676 1428 25732 1822
rect 25676 1362 25732 1372
rect 25788 1652 25844 1662
rect 25788 112 25844 1596
rect 26124 1202 26180 7532
rect 26348 7522 26404 7532
rect 26460 6690 26516 6702
rect 26460 6638 26462 6690
rect 26514 6638 26516 6690
rect 26236 5684 26292 5694
rect 26236 4564 26292 5628
rect 26460 5124 26516 6638
rect 26460 5058 26516 5068
rect 26684 5124 26740 5134
rect 26684 4788 26740 5068
rect 26684 4722 26740 4732
rect 26236 4498 26292 4508
rect 26236 3556 26292 3566
rect 26236 1764 26292 3500
rect 26236 1698 26292 1708
rect 26572 3330 26628 3342
rect 26572 3278 26574 3330
rect 26626 3278 26628 3330
rect 26572 1652 26628 3278
rect 26684 2658 26740 2670
rect 26684 2606 26686 2658
rect 26738 2606 26740 2658
rect 26684 1876 26740 2606
rect 26684 1810 26740 1820
rect 26796 1764 26852 8204
rect 27692 8148 27748 8158
rect 27580 7700 27636 7710
rect 27020 6578 27076 6590
rect 27020 6526 27022 6578
rect 27074 6526 27076 6578
rect 27020 2324 27076 6526
rect 27580 3778 27636 7644
rect 27692 4228 27748 8092
rect 28140 8036 28196 11788
rect 28700 10724 28756 10734
rect 28700 10630 28756 10668
rect 29260 10724 29316 10734
rect 29260 10610 29316 10668
rect 29260 10558 29262 10610
rect 29314 10558 29316 10610
rect 29260 10546 29316 10558
rect 28140 7970 28196 7980
rect 28476 10500 28532 10510
rect 27692 4162 27748 4172
rect 27916 7028 27972 7038
rect 27580 3726 27582 3778
rect 27634 3726 27636 3778
rect 27580 3714 27636 3726
rect 27020 2258 27076 2268
rect 27244 2546 27300 2558
rect 27244 2494 27246 2546
rect 27298 2494 27300 2546
rect 26796 1698 26852 1708
rect 27020 1764 27076 1774
rect 27020 1762 27188 1764
rect 27020 1710 27022 1762
rect 27074 1710 27188 1762
rect 27020 1708 27188 1710
rect 27020 1698 27076 1708
rect 26572 1586 26628 1596
rect 26908 1316 26964 1326
rect 26908 1222 26964 1260
rect 26124 1150 26126 1202
rect 26178 1150 26180 1202
rect 26124 1138 26180 1150
rect 26236 1092 26292 1102
rect 26236 112 26292 1036
rect 26684 1092 26740 1102
rect 26684 112 26740 1036
rect 27132 112 27188 1708
rect 27244 1092 27300 2494
rect 27916 2100 27972 6972
rect 28476 5908 28532 10444
rect 28924 9156 28980 9166
rect 28812 9154 28980 9156
rect 28812 9102 28926 9154
rect 28978 9102 28980 9154
rect 28812 9100 28980 9102
rect 28588 9042 28644 9054
rect 28588 8990 28590 9042
rect 28642 8990 28644 9042
rect 28588 8820 28644 8990
rect 28588 8754 28644 8764
rect 28476 5842 28532 5852
rect 28588 3668 28644 3678
rect 27916 2034 27972 2044
rect 28140 3442 28196 3454
rect 28140 3390 28142 3442
rect 28194 3390 28196 3442
rect 28028 1874 28084 1886
rect 28028 1822 28030 1874
rect 28082 1822 28084 1874
rect 27244 1026 27300 1036
rect 27580 1316 27636 1326
rect 27580 112 27636 1260
rect 28028 112 28084 1822
rect 28140 1204 28196 3390
rect 28588 2996 28644 3612
rect 28588 2930 28644 2940
rect 28700 2548 28756 2558
rect 28700 2454 28756 2492
rect 28812 2098 28868 9100
rect 28924 9090 28980 9100
rect 29484 9156 29540 11900
rect 29708 11732 29764 13804
rect 30044 12962 30100 12974
rect 30044 12910 30046 12962
rect 30098 12910 30100 12962
rect 29708 11666 29764 11676
rect 29820 12740 29876 12750
rect 29484 9090 29540 9100
rect 29596 11060 29652 11070
rect 29260 8372 29316 8382
rect 29260 8278 29316 8316
rect 29596 8148 29652 11004
rect 29820 11060 29876 12684
rect 29820 10994 29876 11004
rect 29932 11844 29988 11854
rect 29820 10500 29876 10510
rect 29708 10388 29764 10398
rect 29708 8596 29764 10332
rect 29708 8530 29764 8540
rect 29820 8370 29876 10444
rect 29932 9492 29988 11788
rect 30044 9940 30100 12910
rect 31388 12852 31444 14112
rect 33068 13972 33124 13982
rect 32396 13188 32452 13198
rect 31836 12852 31892 12862
rect 31388 12850 31892 12852
rect 31388 12798 31838 12850
rect 31890 12798 31892 12850
rect 31388 12796 31892 12798
rect 31836 12786 31892 12796
rect 30604 12290 30660 12302
rect 30604 12238 30606 12290
rect 30658 12238 30660 12290
rect 30268 12180 30324 12190
rect 30268 12178 30436 12180
rect 30268 12126 30270 12178
rect 30322 12126 30436 12178
rect 30268 12124 30436 12126
rect 30268 12114 30324 12124
rect 30268 11620 30324 11630
rect 30044 9874 30100 9884
rect 30156 10948 30212 10958
rect 29932 9426 29988 9436
rect 29820 8318 29822 8370
rect 29874 8318 29876 8370
rect 29820 8306 29876 8318
rect 30044 9268 30100 9278
rect 29596 8082 29652 8092
rect 29820 5348 29876 5358
rect 29820 5254 29876 5292
rect 28924 5122 28980 5134
rect 28924 5070 28926 5122
rect 28978 5070 28980 5122
rect 28924 3780 28980 5070
rect 28924 3714 28980 3724
rect 29484 5010 29540 5022
rect 29484 4958 29486 5010
rect 29538 4958 29540 5010
rect 28812 2046 28814 2098
rect 28866 2046 28868 2098
rect 28812 2034 28868 2046
rect 29148 2996 29204 3006
rect 28140 1138 28196 1148
rect 29148 1202 29204 2940
rect 29260 2658 29316 2670
rect 29260 2606 29262 2658
rect 29314 2606 29316 2658
rect 29260 2548 29316 2606
rect 29260 2482 29316 2492
rect 29372 1762 29428 1774
rect 29372 1710 29374 1762
rect 29426 1710 29428 1762
rect 29372 1204 29428 1710
rect 29148 1150 29150 1202
rect 29202 1150 29204 1202
rect 29148 1138 29204 1150
rect 29260 1148 29428 1204
rect 29484 1204 29540 4958
rect 30044 4900 30100 9212
rect 30156 5348 30212 10892
rect 30268 10052 30324 11564
rect 30268 9986 30324 9996
rect 30156 5282 30212 5292
rect 30380 5236 30436 12124
rect 30604 9268 30660 12238
rect 32396 12178 32452 13132
rect 32844 12964 32900 12974
rect 32844 12870 32900 12908
rect 32396 12126 32398 12178
rect 32450 12126 32452 12178
rect 32396 12114 32452 12126
rect 30828 12068 30884 12078
rect 30604 9202 30660 9212
rect 30716 10612 30772 10622
rect 30268 5180 30436 5236
rect 30492 8708 30548 8718
rect 30156 5124 30212 5134
rect 30268 5124 30324 5180
rect 30212 5068 30324 5124
rect 30156 5058 30212 5068
rect 30044 4834 30100 4844
rect 30380 5010 30436 5022
rect 30380 4958 30382 5010
rect 30434 4958 30436 5010
rect 30156 3780 30212 3790
rect 30156 2882 30212 3724
rect 30156 2830 30158 2882
rect 30210 2830 30212 2882
rect 30156 2818 30212 2830
rect 29596 2546 29652 2558
rect 29596 2494 29598 2546
rect 29650 2494 29652 2546
rect 29596 2212 29652 2494
rect 29596 2146 29652 2156
rect 30380 2098 30436 4958
rect 30492 4340 30548 8652
rect 30716 8482 30772 10556
rect 30828 10610 30884 12012
rect 32956 12066 33012 12078
rect 32956 12014 32958 12066
rect 33010 12014 33012 12066
rect 32956 10836 33012 12014
rect 32956 10770 33012 10780
rect 30828 10558 30830 10610
rect 30882 10558 30884 10610
rect 30828 10546 30884 10558
rect 30716 8430 30718 8482
rect 30770 8430 30772 8482
rect 30716 8418 30772 8430
rect 31388 10498 31444 10510
rect 31388 10446 31390 10498
rect 31442 10446 31444 10498
rect 31388 8372 31444 10446
rect 32956 10388 33012 10398
rect 32396 10164 32452 10174
rect 31388 8306 31444 8316
rect 31612 8596 31668 8606
rect 30492 4274 30548 4284
rect 31164 8146 31220 8158
rect 31164 8094 31166 8146
rect 31218 8094 31220 8146
rect 30940 3220 30996 3230
rect 30940 2884 30996 3164
rect 31164 2996 31220 8094
rect 31500 8036 31556 8046
rect 31164 2930 31220 2940
rect 31276 7140 31332 7150
rect 30940 2818 30996 2828
rect 30492 2772 30548 2782
rect 30492 2678 30548 2716
rect 31052 2548 31108 2558
rect 30380 2046 30382 2098
rect 30434 2046 30436 2098
rect 30380 2034 30436 2046
rect 30604 2546 31108 2548
rect 30604 2494 31054 2546
rect 31106 2494 31108 2546
rect 30604 2492 31108 2494
rect 30156 1988 30212 1998
rect 30156 1652 30212 1932
rect 30156 1586 30212 1596
rect 30604 1316 30660 2492
rect 31052 2482 31108 2492
rect 30268 1260 30660 1316
rect 30716 2324 30772 2334
rect 29596 1204 29652 1214
rect 29484 1202 29652 1204
rect 29484 1150 29598 1202
rect 29650 1150 29652 1202
rect 29484 1148 29652 1150
rect 28476 1090 28532 1102
rect 28476 1038 28478 1090
rect 28530 1038 28532 1090
rect 28476 112 28532 1038
rect 29260 868 29316 1148
rect 29596 1138 29652 1148
rect 28924 812 29316 868
rect 29372 980 29428 990
rect 28924 112 28980 812
rect 29372 112 29428 924
rect 30156 980 30212 990
rect 30156 886 30212 924
rect 29820 868 29876 878
rect 29820 112 29876 812
rect 30268 112 30324 1260
rect 30716 756 30772 2268
rect 31276 2210 31332 7084
rect 31500 4564 31556 7980
rect 31612 4676 31668 8540
rect 31836 8484 31892 8494
rect 31836 6244 31892 8428
rect 31836 6178 31892 6188
rect 32060 6692 32116 6702
rect 31836 5908 31892 5918
rect 32060 5908 32116 6636
rect 31892 5852 32004 5908
rect 31836 5842 31892 5852
rect 31612 4610 31668 4620
rect 31724 5572 31780 5582
rect 31500 4498 31556 4508
rect 31276 2158 31278 2210
rect 31330 2158 31332 2210
rect 31276 2146 31332 2158
rect 31388 2772 31444 2782
rect 31388 1988 31444 2716
rect 31388 1922 31444 1932
rect 31612 2548 31668 2558
rect 30716 690 30772 700
rect 31164 1876 31220 1886
rect 30716 532 30772 542
rect 30716 112 30772 476
rect 31164 112 31220 1820
rect 31500 1204 31556 1214
rect 31500 1110 31556 1148
rect 31612 112 31668 2492
rect 31724 1316 31780 5516
rect 31948 5572 32004 5852
rect 32060 5842 32116 5852
rect 31948 5506 32004 5516
rect 32396 5346 32452 10108
rect 32620 9940 32676 9950
rect 32620 9846 32676 9884
rect 32844 9604 32900 9614
rect 32396 5294 32398 5346
rect 32450 5294 32452 5346
rect 32396 5282 32452 5294
rect 32732 5572 32788 5582
rect 32732 4900 32788 5516
rect 32844 5012 32900 9548
rect 32956 5234 33012 10332
rect 33068 9940 33124 13916
rect 34076 13076 34132 14112
rect 34076 13020 34580 13076
rect 34524 12402 34580 13020
rect 34524 12350 34526 12402
rect 34578 12350 34580 12402
rect 34524 12338 34580 12350
rect 34748 12964 34804 12974
rect 34524 11060 34580 11070
rect 34524 10610 34580 11004
rect 34524 10558 34526 10610
rect 34578 10558 34580 10610
rect 34524 10546 34580 10558
rect 33068 9874 33124 9884
rect 34636 9940 34692 9950
rect 34636 9846 34692 9884
rect 33180 9826 33236 9838
rect 33180 9774 33182 9826
rect 33234 9774 33236 9826
rect 33180 9716 33236 9774
rect 33180 9650 33236 9660
rect 33740 8148 33796 8158
rect 33740 6804 33796 8092
rect 33740 6738 33796 6748
rect 32956 5182 32958 5234
rect 33010 5182 33012 5234
rect 32956 5170 33012 5182
rect 33628 6132 33684 6142
rect 32844 4956 33012 5012
rect 32732 4844 32900 4900
rect 32620 4340 32676 4350
rect 32620 4338 32788 4340
rect 32620 4286 32622 4338
rect 32674 4286 32788 4338
rect 32620 4284 32788 4286
rect 32620 4274 32676 4284
rect 32620 3332 32676 3342
rect 32172 3330 32676 3332
rect 32172 3278 32622 3330
rect 32674 3278 32676 3330
rect 32172 3276 32676 3278
rect 32060 2660 32116 2670
rect 31836 2658 32116 2660
rect 31836 2606 32062 2658
rect 32114 2606 32116 2658
rect 31836 2604 32116 2606
rect 31836 2098 31892 2604
rect 32060 2594 32116 2604
rect 31836 2046 31838 2098
rect 31890 2046 31892 2098
rect 31836 2034 31892 2046
rect 31724 1250 31780 1260
rect 32060 978 32116 990
rect 32060 926 32062 978
rect 32114 926 32116 978
rect 32060 868 32116 926
rect 32060 802 32116 812
rect 32172 644 32228 3276
rect 32620 3266 32676 3276
rect 32732 2772 32788 4284
rect 32844 3332 32900 4844
rect 32844 3266 32900 3276
rect 32732 2706 32788 2716
rect 32956 2772 33012 4956
rect 33628 4340 33684 6076
rect 33852 6132 33908 6142
rect 33740 5572 33796 5582
rect 33740 4900 33796 5516
rect 33852 5124 33908 6076
rect 33852 5058 33908 5068
rect 33964 5348 34020 5358
rect 33740 4834 33796 4844
rect 33628 4274 33684 4284
rect 33068 4228 33124 4238
rect 33068 4226 33460 4228
rect 33068 4174 33070 4226
rect 33122 4174 33460 4226
rect 33068 4172 33460 4174
rect 33068 4162 33124 4172
rect 33404 3554 33460 4172
rect 33404 3502 33406 3554
rect 33458 3502 33460 3554
rect 33404 3490 33460 3502
rect 32956 2706 33012 2716
rect 33628 3108 33684 3118
rect 32396 2660 32452 2670
rect 32396 2098 32452 2604
rect 33068 2660 33124 2670
rect 32620 2548 32676 2558
rect 32620 2454 32676 2492
rect 32396 2046 32398 2098
rect 32450 2046 32452 2098
rect 32396 2034 32452 2046
rect 32956 1876 33012 1886
rect 32956 1782 33012 1820
rect 32060 588 32228 644
rect 32508 1764 32564 1774
rect 32060 112 32116 588
rect 32508 112 32564 1708
rect 33068 1652 33124 2604
rect 32956 1596 33124 1652
rect 33516 2324 33572 2334
rect 32956 112 33012 1596
rect 33068 1428 33124 1438
rect 33068 1202 33124 1372
rect 33068 1150 33070 1202
rect 33122 1150 33124 1202
rect 33068 1138 33124 1150
rect 33516 1092 33572 2268
rect 33628 1652 33684 3052
rect 33964 2884 34020 5292
rect 34636 5122 34692 5134
rect 34636 5070 34638 5122
rect 34690 5070 34692 5122
rect 34636 5012 34692 5070
rect 34636 4946 34692 4956
rect 34748 3668 34804 12908
rect 36764 12852 36820 14112
rect 38220 12962 38276 12974
rect 38220 12910 38222 12962
rect 38274 12910 38276 12962
rect 37212 12852 37268 12862
rect 36764 12850 37268 12852
rect 36764 12798 37214 12850
rect 37266 12798 37268 12850
rect 36764 12796 37268 12798
rect 37212 12786 37268 12796
rect 36876 12404 36932 12414
rect 35532 12068 35588 12078
rect 35532 11974 35588 12012
rect 35308 11844 35364 11854
rect 35084 11394 35140 11406
rect 35084 11342 35086 11394
rect 35138 11342 35140 11394
rect 35084 11172 35140 11342
rect 35084 11106 35140 11116
rect 35196 11396 35252 11406
rect 34972 10836 35028 10846
rect 34972 8820 35028 10780
rect 35084 10612 35140 10622
rect 35084 10518 35140 10556
rect 35196 9938 35252 11340
rect 35196 9886 35198 9938
rect 35250 9886 35252 9938
rect 35196 9874 35252 9886
rect 35308 9940 35364 11788
rect 35980 11732 36036 11742
rect 35644 11282 35700 11294
rect 35644 11230 35646 11282
rect 35698 11230 35700 11282
rect 35644 11172 35700 11230
rect 35644 11106 35700 11116
rect 35308 9874 35364 9884
rect 34972 8764 35476 8820
rect 35308 8596 35364 8606
rect 35084 7250 35140 7262
rect 35084 7198 35086 7250
rect 35138 7198 35140 7250
rect 34748 3602 34804 3612
rect 34860 7140 34916 7150
rect 34748 3332 34804 3342
rect 33964 2818 34020 2828
rect 34412 3330 34804 3332
rect 34412 3278 34750 3330
rect 34802 3278 34804 3330
rect 34412 3276 34804 3278
rect 34076 2660 34132 2670
rect 34076 2566 34132 2604
rect 33628 1586 33684 1596
rect 33852 1876 33908 1886
rect 33516 1026 33572 1036
rect 33404 980 33460 990
rect 33404 112 33460 924
rect 33628 978 33684 990
rect 33628 926 33630 978
rect 33682 926 33684 978
rect 33628 532 33684 926
rect 33628 466 33684 476
rect 33852 112 33908 1820
rect 34188 1764 34244 1774
rect 34188 1670 34244 1708
rect 34412 1652 34468 3276
rect 34748 3266 34804 3276
rect 34860 3220 34916 7084
rect 35084 7028 35140 7198
rect 35084 6962 35140 6972
rect 35308 6580 35364 8540
rect 35308 6514 35364 6524
rect 35196 5908 35252 5918
rect 35252 5852 35364 5908
rect 35196 5842 35252 5852
rect 35196 5682 35252 5694
rect 35196 5630 35198 5682
rect 35250 5630 35252 5682
rect 35196 5460 35252 5630
rect 35196 5394 35252 5404
rect 35196 5124 35252 5134
rect 35196 5030 35252 5068
rect 35196 4676 35252 4686
rect 35196 4340 35252 4620
rect 35308 4564 35364 5852
rect 35420 4900 35476 8764
rect 35644 7700 35700 7710
rect 35644 7586 35700 7644
rect 35644 7534 35646 7586
rect 35698 7534 35700 7586
rect 35644 7522 35700 7534
rect 35756 5908 35812 5918
rect 35756 5814 35812 5852
rect 35420 4834 35476 4844
rect 35644 5012 35700 5022
rect 35644 4676 35700 4956
rect 35980 5012 36036 11676
rect 35980 4946 36036 4956
rect 36092 8708 36148 8718
rect 35308 4498 35364 4508
rect 35420 4620 35700 4676
rect 35308 4340 35364 4350
rect 35196 4338 35364 4340
rect 35196 4286 35310 4338
rect 35362 4286 35364 4338
rect 35196 4284 35364 4286
rect 35308 4274 35364 4284
rect 35420 3388 35476 4620
rect 35644 4450 35700 4462
rect 35644 4398 35646 4450
rect 35698 4398 35700 4450
rect 35420 3332 35588 3388
rect 34860 3154 34916 3164
rect 35532 3108 35588 3332
rect 35532 3042 35588 3052
rect 34860 2772 34916 2782
rect 34860 2678 34916 2716
rect 35308 2770 35364 2782
rect 35308 2718 35310 2770
rect 35362 2718 35364 2770
rect 34300 1596 34468 1652
rect 35084 2660 35140 2670
rect 34300 112 34356 1596
rect 35084 1316 35140 2604
rect 35308 2212 35364 2718
rect 35644 2772 35700 4398
rect 36092 4116 36148 8652
rect 36092 4050 36148 4060
rect 36204 5908 36260 5918
rect 35756 3554 35812 3566
rect 35756 3502 35758 3554
rect 35810 3502 35812 3554
rect 35756 3332 35812 3502
rect 35756 3266 35812 3276
rect 36204 2772 36260 5852
rect 36764 4450 36820 4462
rect 36764 4398 36766 4450
rect 36818 4398 36820 4450
rect 36316 4114 36372 4126
rect 36316 4062 36318 4114
rect 36370 4062 36372 4114
rect 36316 3892 36372 4062
rect 36764 4116 36820 4398
rect 36764 4050 36820 4060
rect 36316 3826 36372 3836
rect 36876 3388 36932 12348
rect 38220 12292 38276 12910
rect 39452 12852 39508 14112
rect 42140 13076 42196 14112
rect 44828 13972 44884 14112
rect 44828 13916 45220 13972
rect 45052 13748 45108 13758
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 42140 13010 42196 13020
rect 43372 13076 43428 13086
rect 43372 12982 43428 13020
rect 40908 12962 40964 12974
rect 40908 12910 40910 12962
rect 40962 12910 40964 12962
rect 39900 12852 39956 12862
rect 39452 12850 39956 12852
rect 39452 12798 39902 12850
rect 39954 12798 39956 12850
rect 39452 12796 39956 12798
rect 39900 12786 39956 12796
rect 40124 12516 40180 12526
rect 38220 12226 38276 12236
rect 39900 12292 39956 12302
rect 39900 12198 39956 12236
rect 37100 12068 37156 12078
rect 37100 11974 37156 12012
rect 36988 11956 37044 11966
rect 36988 6692 37044 11900
rect 37660 11954 37716 11966
rect 37660 11902 37662 11954
rect 37714 11902 37716 11954
rect 36988 6626 37044 6636
rect 37100 8820 37156 8830
rect 37100 6356 37156 8764
rect 37660 7588 37716 11902
rect 38556 10836 38612 10846
rect 38556 10722 38612 10780
rect 38556 10670 38558 10722
rect 38610 10670 38612 10722
rect 38556 10658 38612 10670
rect 37996 10386 38052 10398
rect 37996 10334 37998 10386
rect 38050 10334 38052 10386
rect 37996 10052 38052 10334
rect 40124 10164 40180 12460
rect 40236 12068 40292 12078
rect 40236 10948 40292 12012
rect 40460 11954 40516 11966
rect 40460 11902 40462 11954
rect 40514 11902 40516 11954
rect 40460 11844 40516 11902
rect 40460 11778 40516 11788
rect 40236 10882 40292 10892
rect 40124 10108 40404 10164
rect 37996 9986 38052 9996
rect 40348 8148 40404 10108
rect 40348 8082 40404 8092
rect 37660 7522 37716 7532
rect 37100 6290 37156 6300
rect 40684 6580 40740 6590
rect 40460 6018 40516 6030
rect 40460 5966 40462 6018
rect 40514 5966 40516 6018
rect 40124 5906 40180 5918
rect 40124 5854 40126 5906
rect 40178 5854 40180 5906
rect 37884 5794 37940 5806
rect 37884 5742 37886 5794
rect 37938 5742 37940 5794
rect 37324 5682 37380 5694
rect 37324 5630 37326 5682
rect 37378 5630 37380 5682
rect 37324 5348 37380 5630
rect 37324 5282 37380 5292
rect 36540 3332 36596 3342
rect 36428 3330 36596 3332
rect 36428 3278 36542 3330
rect 36594 3278 36596 3330
rect 36428 3276 36596 3278
rect 36316 2772 36372 2782
rect 36204 2770 36372 2772
rect 36204 2718 36318 2770
rect 36370 2718 36372 2770
rect 36204 2716 36372 2718
rect 35644 2706 35700 2716
rect 36316 2706 36372 2716
rect 35308 2146 35364 2156
rect 35756 2658 35812 2670
rect 35756 2606 35758 2658
rect 35810 2606 35812 2658
rect 35196 2100 35252 2110
rect 35196 2006 35252 2044
rect 35756 2100 35812 2606
rect 35756 2034 35812 2044
rect 35756 1876 35812 1886
rect 35756 1782 35812 1820
rect 35644 1764 35700 1774
rect 36428 1764 36484 3276
rect 36540 3266 36596 3276
rect 36652 3332 36932 3388
rect 37212 5124 37268 5134
rect 35084 1260 35252 1316
rect 34748 868 34804 878
rect 34748 112 34804 812
rect 35196 112 35252 1260
rect 35308 1204 35364 1214
rect 35308 1110 35364 1148
rect 35644 112 35700 1708
rect 36092 1708 36484 1764
rect 36652 1764 36708 3332
rect 36988 2884 37044 2894
rect 36876 2548 36932 2558
rect 36764 1988 36820 1998
rect 36764 1894 36820 1932
rect 36652 1708 36820 1764
rect 35868 980 35924 990
rect 35868 886 35924 924
rect 36092 112 36148 1708
rect 36540 1092 36596 1102
rect 36540 112 36596 1036
rect 15708 18 15764 28
rect 15904 0 16016 112
rect 16352 0 16464 112
rect 16800 0 16912 112
rect 17248 0 17360 112
rect 17696 0 17808 112
rect 18144 0 18256 112
rect 18592 0 18704 112
rect 19040 0 19152 112
rect 19488 0 19600 112
rect 19936 0 20048 112
rect 20384 0 20496 112
rect 20832 0 20944 112
rect 21280 0 21392 112
rect 21728 0 21840 112
rect 22176 0 22288 112
rect 22624 0 22736 112
rect 23072 0 23184 112
rect 23520 0 23632 112
rect 23968 0 24080 112
rect 24416 0 24528 112
rect 24864 0 24976 112
rect 25312 0 25424 112
rect 25760 0 25872 112
rect 26208 0 26320 112
rect 26656 0 26768 112
rect 27104 0 27216 112
rect 27552 0 27664 112
rect 28000 0 28112 112
rect 28448 0 28560 112
rect 28896 0 29008 112
rect 29344 0 29456 112
rect 29792 0 29904 112
rect 30240 0 30352 112
rect 30688 0 30800 112
rect 31136 0 31248 112
rect 31584 0 31696 112
rect 32032 0 32144 112
rect 32480 0 32592 112
rect 32928 0 33040 112
rect 33376 0 33488 112
rect 33824 0 33936 112
rect 34272 0 34384 112
rect 34720 0 34832 112
rect 35168 0 35280 112
rect 35616 0 35728 112
rect 36064 0 36176 112
rect 36512 0 36624 112
rect 36764 84 36820 1708
rect 36876 1316 36932 2492
rect 36876 1250 36932 1260
rect 36988 112 37044 2828
rect 37100 2660 37156 2670
rect 37100 2566 37156 2604
rect 37100 1204 37156 1214
rect 37212 1204 37268 5068
rect 37548 5124 37604 5134
rect 37548 3666 37604 5068
rect 37548 3614 37550 3666
rect 37602 3614 37604 3666
rect 37548 3602 37604 3614
rect 37884 3388 37940 5742
rect 38668 5122 38724 5134
rect 38668 5070 38670 5122
rect 38722 5070 38724 5122
rect 38668 4788 38724 5070
rect 39116 5124 39172 5134
rect 39116 5030 39172 5068
rect 38668 4722 38724 4732
rect 39228 4340 39284 4350
rect 39228 4246 39284 4284
rect 39788 4226 39844 4238
rect 39788 4174 39790 4226
rect 39842 4174 39844 4226
rect 39116 4116 39172 4126
rect 39116 3666 39172 4060
rect 39116 3614 39118 3666
rect 39170 3614 39172 3666
rect 39116 3602 39172 3614
rect 38220 3442 38276 3454
rect 38220 3390 38222 3442
rect 38274 3390 38276 3442
rect 37884 3332 38052 3388
rect 37996 1988 38052 3332
rect 38108 2884 38164 2894
rect 38108 2790 38164 2828
rect 38108 1988 38164 1998
rect 37996 1986 38164 1988
rect 37996 1934 38110 1986
rect 38162 1934 38164 1986
rect 37996 1932 38164 1934
rect 38108 1922 38164 1932
rect 37324 1764 37380 1774
rect 37324 1670 37380 1708
rect 38220 1316 38276 3390
rect 39788 3388 39844 4174
rect 40124 3388 40180 5854
rect 40348 3556 40404 3566
rect 39788 3332 40068 3388
rect 40124 3332 40292 3388
rect 39116 2772 39172 2782
rect 39116 2678 39172 2716
rect 37100 1202 37268 1204
rect 37100 1150 37102 1202
rect 37154 1150 37268 1202
rect 37100 1148 37268 1150
rect 37548 1260 38276 1316
rect 38332 2660 38388 2670
rect 37100 1138 37156 1148
rect 37436 980 37492 990
rect 37436 886 37492 924
rect 37548 756 37604 1260
rect 37436 700 37604 756
rect 37436 112 37492 700
rect 37884 532 37940 542
rect 37884 112 37940 476
rect 38332 112 38388 2604
rect 39900 2660 39956 2670
rect 39900 2566 39956 2604
rect 38668 1986 38724 1998
rect 38668 1934 38670 1986
rect 38722 1934 38724 1986
rect 38668 1652 38724 1934
rect 39228 1988 39284 1998
rect 39228 1894 39284 1932
rect 38668 1586 38724 1596
rect 39676 1652 39732 1662
rect 39564 1092 39620 1102
rect 39564 998 39620 1036
rect 38780 868 38836 878
rect 38780 112 38836 812
rect 39228 756 39284 766
rect 39228 112 39284 700
rect 39676 112 39732 1596
rect 40012 1204 40068 3332
rect 40124 1204 40180 1214
rect 40012 1202 40180 1204
rect 40012 1150 40126 1202
rect 40178 1150 40180 1202
rect 40012 1148 40180 1150
rect 40124 1138 40180 1148
rect 40124 980 40180 990
rect 40124 112 40180 924
rect 40236 308 40292 3332
rect 40348 2660 40404 3500
rect 40460 2772 40516 5966
rect 40460 2706 40516 2716
rect 40572 3442 40628 3454
rect 40572 3390 40574 3442
rect 40626 3390 40628 3442
rect 40348 2594 40404 2604
rect 40460 1762 40516 1774
rect 40460 1710 40462 1762
rect 40514 1710 40516 1762
rect 40460 868 40516 1710
rect 40572 1652 40628 3390
rect 40684 2770 40740 6524
rect 40908 5348 40964 12910
rect 44156 12964 44212 12974
rect 44156 12962 44324 12964
rect 44156 12910 44158 12962
rect 44210 12910 44324 12962
rect 44156 12908 44324 12910
rect 44156 12898 44212 12908
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 43372 11844 43428 11854
rect 41692 8930 41748 8942
rect 41692 8878 41694 8930
rect 41746 8878 41748 8930
rect 41132 8820 41188 8830
rect 41132 8726 41188 8764
rect 41692 8820 41748 8878
rect 41692 8754 41748 8764
rect 43148 7588 43204 7598
rect 43148 6468 43204 7532
rect 43372 6804 43428 11788
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 44156 8818 44212 8830
rect 44156 8766 44158 8818
rect 44210 8766 44212 8818
rect 44156 8708 44212 8766
rect 44156 8642 44212 8652
rect 43372 6738 43428 6748
rect 43484 8484 43540 8494
rect 43260 6692 43316 6702
rect 43260 6598 43316 6636
rect 43148 6412 43316 6468
rect 40908 5282 40964 5292
rect 41692 6244 41748 6254
rect 41356 5012 41412 5022
rect 41132 4676 41188 4686
rect 41132 3892 41188 4620
rect 41132 3826 41188 3836
rect 41356 3554 41412 4956
rect 41468 4564 41524 4574
rect 41468 4338 41524 4508
rect 41468 4286 41470 4338
rect 41522 4286 41524 4338
rect 41468 4274 41524 4286
rect 41692 4340 41748 6188
rect 41692 4274 41748 4284
rect 41804 5796 41860 5806
rect 41804 3666 41860 5740
rect 41804 3614 41806 3666
rect 41858 3614 41860 3666
rect 41804 3602 41860 3614
rect 41916 5124 41972 5134
rect 41356 3502 41358 3554
rect 41410 3502 41412 3554
rect 41356 3490 41412 3502
rect 40684 2718 40686 2770
rect 40738 2718 40740 2770
rect 40684 2706 40740 2718
rect 41244 2882 41300 2894
rect 41244 2830 41246 2882
rect 41298 2830 41300 2882
rect 40572 1586 40628 1596
rect 41020 1540 41076 1550
rect 40908 1314 40964 1326
rect 40908 1262 40910 1314
rect 40962 1262 40964 1314
rect 40460 802 40516 812
rect 40572 1092 40628 1102
rect 40236 242 40292 252
rect 40572 112 40628 1036
rect 40908 532 40964 1262
rect 40908 466 40964 476
rect 41020 112 41076 1484
rect 41244 980 41300 2830
rect 41468 2884 41524 2894
rect 41468 2098 41524 2828
rect 41468 2046 41470 2098
rect 41522 2046 41524 2098
rect 41468 2034 41524 2046
rect 41244 914 41300 924
rect 41468 1652 41524 1662
rect 41468 112 41524 1596
rect 41916 1202 41972 5068
rect 42588 5122 42644 5134
rect 42588 5070 42590 5122
rect 42642 5070 42644 5122
rect 42028 4226 42084 4238
rect 42028 4174 42030 4226
rect 42082 4174 42084 4226
rect 42028 4116 42084 4174
rect 42028 4050 42084 4060
rect 42252 4116 42308 4126
rect 42252 2770 42308 4060
rect 42252 2718 42254 2770
rect 42306 2718 42308 2770
rect 42252 2706 42308 2718
rect 42364 3330 42420 3342
rect 42364 3278 42366 3330
rect 42418 3278 42420 3330
rect 41916 1150 41918 1202
rect 41970 1150 41972 1202
rect 41916 1138 41972 1150
rect 42028 1762 42084 1774
rect 42028 1710 42030 1762
rect 42082 1710 42084 1762
rect 41916 980 41972 990
rect 41916 112 41972 924
rect 42028 756 42084 1710
rect 42364 1652 42420 3278
rect 42588 1764 42644 5070
rect 43148 5124 43204 5134
rect 43148 5030 43204 5068
rect 42588 1698 42644 1708
rect 42812 3556 42868 3566
rect 42364 1586 42420 1596
rect 42028 690 42084 700
rect 42364 196 42420 206
rect 42364 112 42420 140
rect 42812 112 42868 3500
rect 43260 3388 43316 6412
rect 43484 5908 43540 8428
rect 43484 5842 43540 5852
rect 43596 8258 43652 8270
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 43372 4004 43428 4014
rect 43372 3666 43428 3948
rect 43596 3892 43652 8206
rect 44156 8146 44212 8158
rect 44156 8094 44158 8146
rect 44210 8094 44212 8146
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 43820 7588 43876 7598
rect 43820 7140 43876 7532
rect 43820 7074 43876 7084
rect 44156 6804 44212 8094
rect 44156 6738 44212 6748
rect 43708 6580 43764 6590
rect 43708 6486 43764 6524
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 44268 5012 44324 12908
rect 44604 11956 44660 11994
rect 44604 11890 44660 11900
rect 44940 11956 44996 11966
rect 44940 11862 44996 11900
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44940 11172 44996 11182
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44716 8932 44772 8942
rect 44716 8838 44772 8876
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44828 6690 44884 6702
rect 44828 6638 44830 6690
rect 44882 6638 44884 6690
rect 44828 6020 44884 6638
rect 44828 5954 44884 5964
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 44268 4946 44324 4956
rect 44156 4900 44212 4910
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 44156 4564 44212 4844
rect 44940 4676 44996 11116
rect 45052 6356 45108 13692
rect 45164 12850 45220 13916
rect 45948 12964 46004 12974
rect 45164 12798 45166 12850
rect 45218 12798 45220 12850
rect 45164 12786 45220 12798
rect 45612 12962 46004 12964
rect 45612 12910 45950 12962
rect 46002 12910 46004 12962
rect 45612 12908 46004 12910
rect 45388 11844 45444 11854
rect 45388 9044 45444 11788
rect 45388 8978 45444 8988
rect 45052 6290 45108 6300
rect 45164 8260 45220 8270
rect 45052 4676 45108 4686
rect 44940 4620 45052 4676
rect 45052 4610 45108 4620
rect 44380 4564 44436 4574
rect 44156 4508 44380 4564
rect 44380 4498 44436 4508
rect 45052 4452 45108 4462
rect 44940 4340 44996 4350
rect 44940 4246 44996 4284
rect 44268 4060 44884 4116
rect 44268 4004 44324 4060
rect 44828 4004 44884 4060
rect 44268 3938 44324 3948
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44828 3938 44884 3948
rect 44464 3882 44728 3892
rect 43596 3826 43652 3836
rect 43372 3614 43374 3666
rect 43426 3614 43428 3666
rect 43372 3602 43428 3614
rect 43932 3556 43988 3566
rect 43932 3442 43988 3500
rect 45052 3554 45108 4396
rect 45052 3502 45054 3554
rect 45106 3502 45108 3554
rect 45052 3490 45108 3502
rect 43932 3390 43934 3442
rect 43986 3390 43988 3442
rect 43260 3332 43540 3388
rect 43932 3378 43988 3390
rect 45164 3388 45220 8204
rect 45276 6578 45332 6590
rect 45276 6526 45278 6578
rect 45330 6526 45332 6578
rect 45276 5124 45332 6526
rect 45276 5058 45332 5068
rect 45500 5124 45556 5134
rect 45388 4450 45444 4462
rect 45388 4398 45390 4450
rect 45442 4398 45444 4450
rect 45388 3444 45444 4398
rect 45500 4116 45556 5068
rect 45500 4050 45556 4060
rect 43036 3108 43092 3118
rect 43036 2770 43092 3052
rect 43036 2718 43038 2770
rect 43090 2718 43092 2770
rect 43036 2706 43092 2718
rect 43372 2100 43428 2110
rect 43372 2006 43428 2044
rect 43036 1988 43092 1998
rect 43036 1894 43092 1932
rect 43260 1316 43316 1326
rect 43260 112 43316 1260
rect 43372 1092 43428 1102
rect 43484 1092 43540 3332
rect 45052 3332 45220 3388
rect 45276 3388 45444 3444
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 45052 3108 45108 3332
rect 45052 3042 45108 3052
rect 44828 2882 44884 2894
rect 44828 2830 44830 2882
rect 44882 2830 44884 2882
rect 44268 2770 44324 2782
rect 44268 2718 44270 2770
rect 44322 2718 44324 2770
rect 43596 2658 43652 2670
rect 43596 2606 43598 2658
rect 43650 2606 43652 2658
rect 43596 2100 43652 2606
rect 43596 2034 43652 2044
rect 43932 1764 43988 1802
rect 43932 1698 43988 1708
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 44156 1540 44212 1550
rect 44156 1202 44212 1484
rect 44156 1150 44158 1202
rect 44210 1150 44212 1202
rect 44156 1138 44212 1150
rect 43596 1092 43652 1102
rect 43484 1036 43596 1092
rect 43372 998 43428 1036
rect 43596 1026 43652 1036
rect 43708 532 43764 542
rect 43708 112 43764 476
rect 44268 420 44324 2718
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 44828 1316 44884 2830
rect 45276 2884 45332 3388
rect 45500 3332 45556 3342
rect 45276 2818 45332 2828
rect 45388 3330 45556 3332
rect 45388 3278 45502 3330
rect 45554 3278 45556 3330
rect 45388 3276 45556 3278
rect 44940 2660 44996 2670
rect 44940 2098 44996 2604
rect 44940 2046 44942 2098
rect 44994 2046 44996 2098
rect 44940 2034 44996 2046
rect 44828 1250 44884 1260
rect 44492 1204 44548 1214
rect 44492 1110 44548 1148
rect 45052 980 45108 990
rect 45052 886 45108 924
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 44268 354 44324 364
rect 44604 644 44660 654
rect 44156 308 44212 318
rect 44156 112 44212 252
rect 44604 112 44660 588
rect 45388 644 45444 3276
rect 45500 3266 45556 3276
rect 45612 3220 45668 12908
rect 45948 12898 46004 12908
rect 47516 12852 47572 14112
rect 49980 14084 50036 14094
rect 48972 12964 49028 12974
rect 48972 12962 49252 12964
rect 48972 12910 48974 12962
rect 49026 12910 49252 12962
rect 48972 12908 49252 12910
rect 48972 12898 49028 12908
rect 47964 12852 48020 12862
rect 47516 12850 48020 12852
rect 47516 12798 47966 12850
rect 48018 12798 48020 12850
rect 47516 12796 48020 12798
rect 47964 12786 48020 12796
rect 46844 12740 46900 12750
rect 46844 12178 46900 12684
rect 46844 12126 46846 12178
rect 46898 12126 46900 12178
rect 46844 12114 46900 12126
rect 47180 12068 47236 12078
rect 47404 12068 47460 12078
rect 47236 12012 47348 12068
rect 47180 12002 47236 12012
rect 47068 11284 47124 11294
rect 47068 11190 47124 11228
rect 46172 9716 46228 9726
rect 45724 3444 45780 3454
rect 45724 3332 45780 3388
rect 45724 3266 45780 3276
rect 45612 3154 45668 3164
rect 45724 3108 45780 3118
rect 45724 2770 45780 3052
rect 45724 2718 45726 2770
rect 45778 2718 45780 2770
rect 45724 2706 45780 2718
rect 45724 1874 45780 1886
rect 45724 1822 45726 1874
rect 45778 1822 45780 1874
rect 45388 578 45444 588
rect 45500 868 45556 878
rect 45052 420 45108 430
rect 45052 112 45108 364
rect 45500 112 45556 812
rect 45724 196 45780 1822
rect 45724 130 45780 140
rect 45948 1764 46004 1774
rect 45948 112 46004 1708
rect 46172 1204 46228 9660
rect 46508 7252 46564 7262
rect 46508 3778 46564 7196
rect 46620 5908 46676 5918
rect 46620 5814 46676 5852
rect 47180 5794 47236 5806
rect 47180 5742 47182 5794
rect 47234 5742 47236 5794
rect 47180 5460 47236 5742
rect 47180 5394 47236 5404
rect 46732 5348 46788 5358
rect 46620 4228 46676 4238
rect 46620 4134 46676 4172
rect 46508 3726 46510 3778
rect 46562 3726 46564 3778
rect 46508 3714 46564 3726
rect 46620 3668 46676 3678
rect 46508 3220 46564 3230
rect 46172 1138 46228 1148
rect 46284 2546 46340 2558
rect 46284 2494 46286 2546
rect 46338 2494 46340 2546
rect 46284 308 46340 2494
rect 46508 2098 46564 3164
rect 46508 2046 46510 2098
rect 46562 2046 46564 2098
rect 46508 2034 46564 2046
rect 46620 1316 46676 3612
rect 46732 3332 46788 5292
rect 47068 5236 47124 5246
rect 47068 5122 47124 5180
rect 47068 5070 47070 5122
rect 47122 5070 47124 5122
rect 47068 5058 47124 5070
rect 47292 4900 47348 12012
rect 47404 11974 47460 12012
rect 47740 11956 47796 11966
rect 47516 11394 47572 11406
rect 47516 11342 47518 11394
rect 47570 11342 47572 11394
rect 47516 7252 47572 11342
rect 47516 7186 47572 7196
rect 47516 5124 47572 5134
rect 47516 5030 47572 5068
rect 47292 4834 47348 4844
rect 47180 4114 47236 4126
rect 47180 4062 47182 4114
rect 47234 4062 47236 4114
rect 47180 3668 47236 4062
rect 47180 3602 47236 3612
rect 46732 3266 46788 3276
rect 46956 3442 47012 3454
rect 46956 3390 46958 3442
rect 47010 3390 47012 3442
rect 46956 1988 47012 3390
rect 47292 2772 47348 2782
rect 47292 2678 47348 2716
rect 46956 1922 47012 1932
rect 47068 1986 47124 1998
rect 47068 1934 47070 1986
rect 47122 1934 47124 1986
rect 47068 1876 47124 1934
rect 47068 1810 47124 1820
rect 46284 242 46340 252
rect 46396 1260 46676 1316
rect 46732 1428 46788 1438
rect 46396 112 46452 1260
rect 46732 1202 46788 1372
rect 46732 1150 46734 1202
rect 46786 1150 46788 1202
rect 46732 1138 46788 1150
rect 46844 1316 46900 1326
rect 46844 112 46900 1260
rect 47292 978 47348 990
rect 47292 926 47294 978
rect 47346 926 47348 978
rect 47292 532 47348 926
rect 47292 466 47348 476
rect 47292 308 47348 318
rect 47292 112 47348 252
rect 47740 112 47796 11900
rect 49084 11508 49140 11518
rect 48860 9268 48916 9278
rect 48748 8036 48804 8046
rect 48188 7252 48244 7262
rect 48076 3444 48132 3454
rect 47852 2546 47908 2558
rect 47852 2494 47854 2546
rect 47906 2494 47908 2546
rect 47852 1764 47908 2494
rect 48076 2098 48132 3388
rect 48076 2046 48078 2098
rect 48130 2046 48132 2098
rect 48076 2034 48132 2046
rect 47852 1698 47908 1708
rect 48188 112 48244 7196
rect 48748 5908 48804 7980
rect 48860 6804 48916 9212
rect 48860 6738 48916 6748
rect 48972 7588 49028 7598
rect 48748 5842 48804 5852
rect 48748 4788 48804 4798
rect 48412 4004 48468 4014
rect 48300 3556 48356 3566
rect 48300 3462 48356 3500
rect 48412 1202 48468 3948
rect 48636 2660 48692 2670
rect 48636 1540 48692 2604
rect 48748 2324 48804 4732
rect 48860 3556 48916 3566
rect 48860 3462 48916 3500
rect 48972 2770 49028 7532
rect 48972 2718 48974 2770
rect 49026 2718 49028 2770
rect 48972 2706 49028 2718
rect 48748 2258 48804 2268
rect 48636 1474 48692 1484
rect 48748 1874 48804 1886
rect 48748 1822 48750 1874
rect 48802 1822 48804 1874
rect 48412 1150 48414 1202
rect 48466 1150 48468 1202
rect 48412 1138 48468 1150
rect 48748 868 48804 1822
rect 49084 1652 49140 11452
rect 49196 3666 49252 12908
rect 49980 12290 50036 14028
rect 50204 14084 50260 14112
rect 50204 14018 50260 14028
rect 50764 14084 50820 14094
rect 50764 12850 50820 14028
rect 52892 13188 52948 14112
rect 54908 13636 54964 13646
rect 53116 13188 53172 13198
rect 52892 13186 53172 13188
rect 52892 13134 53118 13186
rect 53170 13134 53172 13186
rect 52892 13132 53172 13134
rect 53116 13122 53172 13132
rect 51772 12964 51828 12974
rect 52556 12964 52612 12974
rect 51772 12870 51828 12908
rect 52332 12962 52612 12964
rect 52332 12910 52558 12962
rect 52610 12910 52612 12962
rect 52332 12908 52612 12910
rect 50764 12798 50766 12850
rect 50818 12798 50820 12850
rect 50764 12786 50820 12798
rect 49980 12238 49982 12290
rect 50034 12238 50036 12290
rect 49980 12226 50036 12238
rect 52220 12178 52276 12190
rect 52220 12126 52222 12178
rect 52274 12126 52276 12178
rect 50988 12068 51044 12078
rect 49532 11956 49588 11966
rect 49196 3614 49198 3666
rect 49250 3614 49252 3666
rect 49196 3602 49252 3614
rect 49308 11954 49588 11956
rect 49308 11902 49534 11954
rect 49586 11902 49588 11954
rect 49308 11900 49588 11902
rect 49084 1586 49140 1596
rect 48748 802 48804 812
rect 48860 978 48916 990
rect 48860 926 48862 978
rect 48914 926 48916 978
rect 48636 756 48692 766
rect 48636 112 48692 700
rect 48860 420 48916 926
rect 49308 756 49364 11900
rect 49532 11890 49588 11900
rect 50988 11506 51044 12012
rect 50988 11454 50990 11506
rect 51042 11454 51044 11506
rect 50988 11442 51044 11454
rect 51996 11284 52052 11294
rect 51996 11190 52052 11228
rect 51884 10724 51940 10734
rect 50204 6356 50260 6366
rect 49420 6132 49476 6142
rect 49420 5906 49476 6076
rect 49420 5854 49422 5906
rect 49474 5854 49476 5906
rect 49420 5842 49476 5854
rect 49532 5796 49588 5806
rect 49420 2546 49476 2558
rect 49420 2494 49422 2546
rect 49474 2494 49476 2546
rect 49420 1316 49476 2494
rect 49420 1250 49476 1260
rect 49308 690 49364 700
rect 48860 354 48916 364
rect 49084 196 49140 206
rect 49084 112 49140 140
rect 49532 112 49588 5740
rect 49980 5796 50036 5806
rect 49980 5702 50036 5740
rect 49980 4900 50036 4910
rect 49756 3892 49812 3902
rect 49756 3778 49812 3836
rect 49756 3726 49758 3778
rect 49810 3726 49812 3778
rect 49756 3714 49812 3726
rect 49644 2548 49700 2558
rect 49644 2098 49700 2492
rect 49644 2046 49646 2098
rect 49698 2046 49700 2098
rect 49644 2034 49700 2046
rect 49980 112 50036 4844
rect 50204 196 50260 6300
rect 50988 5460 51044 5470
rect 50428 4564 50484 4574
rect 50428 2772 50484 4508
rect 50764 3668 50820 3678
rect 50764 3574 50820 3612
rect 50428 2706 50484 2716
rect 50876 2996 50932 3006
rect 50876 2770 50932 2940
rect 50876 2718 50878 2770
rect 50930 2718 50932 2770
rect 50876 2706 50932 2718
rect 50876 2324 50932 2334
rect 50540 1874 50596 1886
rect 50540 1822 50542 1874
rect 50594 1822 50596 1874
rect 50540 308 50596 1822
rect 50540 242 50596 252
rect 50204 130 50260 140
rect 50428 196 50484 206
rect 50428 112 50484 140
rect 50876 112 50932 2268
rect 50988 1202 51044 5404
rect 51660 4788 51716 4798
rect 51324 4004 51380 4014
rect 51324 3778 51380 3948
rect 51324 3726 51326 3778
rect 51378 3726 51380 3778
rect 51324 3714 51380 3726
rect 51660 3666 51716 4732
rect 51660 3614 51662 3666
rect 51714 3614 51716 3666
rect 51660 3602 51716 3614
rect 51212 3332 51268 3342
rect 51212 2098 51268 3276
rect 51212 2046 51214 2098
rect 51266 2046 51268 2098
rect 51212 2034 51268 2046
rect 51436 2658 51492 2670
rect 51436 2606 51438 2658
rect 51490 2606 51492 2658
rect 51436 2100 51492 2606
rect 51436 2034 51492 2044
rect 51772 1988 51828 1998
rect 51772 1894 51828 1932
rect 51884 1764 51940 10668
rect 52108 10612 52164 10622
rect 52108 10518 52164 10556
rect 52220 10276 52276 12126
rect 52220 10210 52276 10220
rect 52108 8820 52164 8830
rect 52108 6916 52164 8764
rect 52108 6850 52164 6860
rect 52332 5234 52388 12908
rect 52556 12898 52612 12908
rect 52668 12964 52724 12974
rect 52556 11396 52612 11406
rect 52556 11302 52612 11340
rect 52556 9828 52612 9838
rect 52556 9734 52612 9772
rect 52332 5182 52334 5234
rect 52386 5182 52388 5234
rect 52332 5170 52388 5182
rect 52444 8596 52500 8606
rect 52220 3554 52276 3566
rect 52220 3502 52222 3554
rect 52274 3502 52276 3554
rect 52220 3444 52276 3502
rect 52220 3378 52276 3388
rect 52108 2770 52164 2782
rect 52108 2718 52110 2770
rect 52162 2718 52164 2770
rect 52108 2212 52164 2718
rect 52108 2146 52164 2156
rect 52444 2100 52500 8540
rect 52668 4450 52724 12908
rect 53004 12404 53060 12414
rect 53004 12310 53060 12348
rect 53564 12180 53620 12190
rect 53564 12086 53620 12124
rect 54348 12068 54404 12078
rect 54348 11974 54404 12012
rect 54124 11394 54180 11406
rect 54124 11342 54126 11394
rect 54178 11342 54180 11394
rect 53564 11172 53620 11182
rect 53564 11078 53620 11116
rect 53004 11060 53060 11070
rect 53004 10834 53060 11004
rect 53004 10782 53006 10834
rect 53058 10782 53060 10834
rect 53004 10770 53060 10782
rect 54124 10836 54180 11342
rect 54124 10770 54180 10780
rect 54572 10722 54628 10734
rect 54572 10670 54574 10722
rect 54626 10670 54628 10722
rect 53564 10500 53620 10510
rect 53564 10406 53620 10444
rect 53116 10276 53172 10286
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 52780 5796 52836 5806
rect 52556 3780 52612 3790
rect 52556 3666 52612 3724
rect 52556 3614 52558 3666
rect 52610 3614 52612 3666
rect 52556 3602 52612 3614
rect 52668 3556 52724 3566
rect 52556 2100 52612 2110
rect 52444 2098 52612 2100
rect 52444 2046 52558 2098
rect 52610 2046 52612 2098
rect 52444 2044 52612 2046
rect 52556 2034 52612 2044
rect 51772 1708 51940 1764
rect 50988 1150 50990 1202
rect 51042 1150 51044 1202
rect 50988 1138 51044 1150
rect 51324 1652 51380 1662
rect 51324 112 51380 1596
rect 51772 112 51828 1708
rect 51996 1314 52052 1326
rect 51996 1262 51998 1314
rect 52050 1262 52052 1314
rect 51996 980 52052 1262
rect 51996 914 52052 924
rect 52220 1204 52276 1214
rect 52220 112 52276 1148
rect 52668 112 52724 3500
rect 52780 1202 52836 5740
rect 52892 5348 52948 5358
rect 52892 5254 52948 5292
rect 53116 3668 53172 10220
rect 54572 10164 54628 10670
rect 54572 10098 54628 10108
rect 54236 9826 54292 9838
rect 54236 9774 54238 9826
rect 54290 9774 54292 9826
rect 53564 9716 53620 9726
rect 53564 9622 53620 9660
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 7700 53620 8878
rect 54124 8372 54180 8382
rect 54124 8278 54180 8316
rect 53564 7634 53620 7644
rect 53564 7476 53620 7486
rect 53564 7382 53620 7420
rect 54236 7028 54292 9774
rect 54348 8930 54404 8942
rect 54348 8878 54350 8930
rect 54402 8878 54404 8930
rect 54348 8596 54404 8878
rect 54908 8932 54964 13580
rect 55132 12964 55188 12974
rect 55020 12962 55188 12964
rect 55020 12910 55134 12962
rect 55186 12910 55188 12962
rect 55020 12908 55188 12910
rect 55020 9156 55076 12908
rect 55132 12898 55188 12908
rect 55580 12404 55636 14112
rect 55580 12338 55636 12348
rect 55804 13972 55860 13982
rect 55132 12066 55188 12078
rect 55132 12014 55134 12066
rect 55186 12014 55188 12066
rect 55132 11844 55188 12014
rect 55132 11778 55188 11788
rect 55804 11284 55860 13916
rect 56476 13524 56532 13534
rect 56140 12738 56196 12750
rect 56140 12686 56142 12738
rect 56194 12686 56196 12738
rect 55804 11218 55860 11228
rect 55916 12066 55972 12078
rect 55916 12014 55918 12066
rect 55970 12014 55972 12066
rect 55132 11170 55188 11182
rect 55132 11118 55134 11170
rect 55186 11118 55188 11170
rect 55132 10836 55188 11118
rect 55132 10770 55188 10780
rect 55132 10498 55188 10510
rect 55132 10446 55134 10498
rect 55186 10446 55188 10498
rect 55132 10388 55188 10446
rect 55132 10322 55188 10332
rect 55916 10388 55972 12014
rect 56140 11284 56196 12686
rect 56140 11218 56196 11228
rect 56364 12180 56420 12190
rect 56364 11172 56420 12124
rect 56364 11106 56420 11116
rect 55916 10322 55972 10332
rect 56140 10722 56196 10734
rect 56140 10670 56142 10722
rect 56194 10670 56196 10722
rect 55356 9940 55412 9950
rect 55132 9602 55188 9614
rect 55132 9550 55134 9602
rect 55186 9550 55188 9602
rect 55132 9492 55188 9550
rect 55132 9426 55188 9436
rect 55020 9090 55076 9100
rect 55244 9042 55300 9054
rect 55244 8990 55246 9042
rect 55298 8990 55300 9042
rect 55132 8932 55188 8942
rect 54908 8876 55076 8932
rect 54348 8530 54404 8540
rect 54908 8372 54964 8382
rect 54908 8278 54964 8316
rect 54572 7586 54628 7598
rect 54572 7534 54574 7586
rect 54626 7534 54628 7586
rect 54572 7252 54628 7534
rect 54572 7186 54628 7196
rect 54236 6962 54292 6972
rect 53676 6804 53732 6814
rect 53452 6580 53508 6590
rect 53228 5684 53284 5694
rect 53228 5346 53284 5628
rect 53228 5294 53230 5346
rect 53282 5294 53284 5346
rect 53228 5282 53284 5294
rect 53228 4116 53284 4126
rect 53228 4022 53284 4060
rect 53116 3602 53172 3612
rect 53004 2884 53060 2894
rect 53004 2790 53060 2828
rect 52780 1150 52782 1202
rect 52834 1150 52836 1202
rect 52780 1138 52836 1150
rect 53116 1092 53172 1102
rect 53116 112 53172 1036
rect 53452 644 53508 6524
rect 53564 5908 53620 5918
rect 53564 5814 53620 5852
rect 53676 4338 53732 6748
rect 54124 6690 54180 6702
rect 54124 6638 54126 6690
rect 54178 6638 54180 6690
rect 54124 6468 54180 6638
rect 54124 6402 54180 6412
rect 54236 6692 54292 6702
rect 54236 5122 54292 6636
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 5908 54628 5966
rect 54572 5842 54628 5852
rect 54236 5070 54238 5122
rect 54290 5070 54292 5122
rect 54236 5058 54292 5070
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 53676 4286 53678 4338
rect 53730 4286 53732 4338
rect 53676 4274 53732 4286
rect 53788 5010 53844 5022
rect 53788 4958 53790 5010
rect 53842 4958 53844 5010
rect 53788 4116 53844 4958
rect 53676 4060 53844 4116
rect 54124 4676 54180 4686
rect 53564 3556 53620 3566
rect 53564 3442 53620 3500
rect 53564 3390 53566 3442
rect 53618 3390 53620 3442
rect 53564 3378 53620 3390
rect 53564 2772 53620 2782
rect 53564 2678 53620 2716
rect 53676 2660 53732 4060
rect 54124 3666 54180 4620
rect 54572 4564 54628 4574
rect 54572 4470 54628 4508
rect 54124 3614 54126 3666
rect 54178 3614 54180 3666
rect 54124 3602 54180 3614
rect 54908 3668 54964 3678
rect 54908 3574 54964 3612
rect 53676 2594 53732 2604
rect 54460 3444 54516 3454
rect 54124 2100 54180 2110
rect 54124 2006 54180 2044
rect 54012 1988 54068 1998
rect 53564 1876 53620 1886
rect 53564 1782 53620 1820
rect 53564 1428 53620 1438
rect 53564 1334 53620 1372
rect 53452 588 53620 644
rect 53564 112 53620 588
rect 54012 112 54068 1932
rect 54460 112 54516 3388
rect 54572 3220 54628 3230
rect 54572 2994 54628 3164
rect 54572 2942 54574 2994
rect 54626 2942 54628 2994
rect 54572 2930 54628 2942
rect 55020 2772 55076 8876
rect 55132 7474 55188 8876
rect 55132 7422 55134 7474
rect 55186 7422 55188 7474
rect 55132 7410 55188 7422
rect 55244 7364 55300 8990
rect 55244 7298 55300 7308
rect 55244 6916 55300 6926
rect 55132 6466 55188 6478
rect 55132 6414 55134 6466
rect 55186 6414 55188 6466
rect 55132 6356 55188 6414
rect 55132 6290 55188 6300
rect 55244 4338 55300 6860
rect 55356 5906 55412 9884
rect 56140 9044 56196 10670
rect 56476 9716 56532 13468
rect 57036 13076 57092 13086
rect 56700 12628 56756 12638
rect 56700 11060 56756 12572
rect 56700 10994 56756 11004
rect 56476 9650 56532 9660
rect 56140 8978 56196 8988
rect 55916 8930 55972 8942
rect 55916 8878 55918 8930
rect 55970 8878 55972 8930
rect 55916 8148 55972 8878
rect 57036 8372 57092 13020
rect 57260 10164 57316 10174
rect 57260 9940 57316 10108
rect 57260 9874 57316 9884
rect 57036 8306 57092 8316
rect 55916 8082 55972 8092
rect 56140 7700 56196 7710
rect 56140 7606 56196 7644
rect 56140 6804 56196 6814
rect 56140 6130 56196 6748
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 55356 5854 55358 5906
rect 55410 5854 55412 5906
rect 55356 5842 55412 5854
rect 56140 5460 56196 5470
rect 56140 4562 56196 5404
rect 56140 4510 56142 4562
rect 56194 4510 56196 4562
rect 56140 4498 56196 4510
rect 56252 5348 56308 5358
rect 55244 4286 55246 4338
rect 55298 4286 55300 4338
rect 55244 4274 55300 4286
rect 55804 4116 55860 4126
rect 55356 3892 55412 3902
rect 55132 2772 55188 2782
rect 55020 2770 55188 2772
rect 55020 2718 55134 2770
rect 55186 2718 55188 2770
rect 55020 2716 55188 2718
rect 55132 2706 55188 2716
rect 54908 2324 54964 2334
rect 54908 2098 54964 2268
rect 54908 2046 54910 2098
rect 54962 2046 54964 2098
rect 54908 2034 54964 2046
rect 55132 1764 55188 1774
rect 54908 1540 54964 1550
rect 54908 112 54964 1484
rect 55132 1202 55188 1708
rect 55132 1150 55134 1202
rect 55186 1150 55188 1202
rect 55132 1138 55188 1150
rect 55356 112 55412 3836
rect 55804 112 55860 4060
rect 56140 4116 56196 4126
rect 56140 2994 56196 4060
rect 56140 2942 56142 2994
rect 56194 2942 56196 2994
rect 56140 2930 56196 2942
rect 56140 2772 56196 2782
rect 56140 1426 56196 2716
rect 56140 1374 56142 1426
rect 56194 1374 56196 1426
rect 56140 1362 56196 1374
rect 56252 112 56308 5292
rect 56700 4004 56756 4014
rect 56700 112 56756 3948
rect 56812 3556 56868 3566
rect 56812 532 56868 3500
rect 56812 466 56868 476
rect 56924 2884 56980 2894
rect 36764 18 36820 28
rect 36960 0 37072 112
rect 37408 0 37520 112
rect 37856 0 37968 112
rect 38304 0 38416 112
rect 38752 0 38864 112
rect 39200 0 39312 112
rect 39648 0 39760 112
rect 40096 0 40208 112
rect 40544 0 40656 112
rect 40992 0 41104 112
rect 41440 0 41552 112
rect 41888 0 42000 112
rect 42336 0 42448 112
rect 42784 0 42896 112
rect 43232 0 43344 112
rect 43680 0 43792 112
rect 44128 0 44240 112
rect 44576 0 44688 112
rect 45024 0 45136 112
rect 45472 0 45584 112
rect 45920 0 46032 112
rect 46368 0 46480 112
rect 46816 0 46928 112
rect 47264 0 47376 112
rect 47712 0 47824 112
rect 48160 0 48272 112
rect 48608 0 48720 112
rect 49056 0 49168 112
rect 49504 0 49616 112
rect 49952 0 50064 112
rect 50400 0 50512 112
rect 50848 0 50960 112
rect 51296 0 51408 112
rect 51744 0 51856 112
rect 52192 0 52304 112
rect 52640 0 52752 112
rect 53088 0 53200 112
rect 53536 0 53648 112
rect 53984 0 54096 112
rect 54432 0 54544 112
rect 54880 0 54992 112
rect 55328 0 55440 112
rect 55776 0 55888 112
rect 56224 0 56336 112
rect 56672 0 56784 112
rect 56924 84 56980 2828
rect 56924 18 56980 28
<< via2 >>
rect 4508 14028 4564 14084
rect 5068 14028 5124 14084
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 1596 12572 1652 12628
rect 364 12124 420 12180
rect 1596 11452 1652 11508
rect 6860 13020 6916 13076
rect 5292 12908 5348 12964
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 6076 12796 6132 12852
rect 8092 14028 8148 14084
rect 7308 13916 7364 13972
rect 6860 11900 6916 11956
rect 6972 12012 7028 12068
rect 5292 11676 5348 11732
rect 6636 11228 6692 11284
rect 2380 10668 2436 10724
rect 3052 11116 3108 11172
rect 364 9996 420 10052
rect 1596 9436 1652 9492
rect 2940 9154 2996 9156
rect 2940 9102 2942 9154
rect 2942 9102 2994 9154
rect 2994 9102 2996 9154
rect 2940 9100 2996 9102
rect 1596 8316 1652 8372
rect 1148 5740 1204 5796
rect 700 2828 756 2884
rect 2044 5068 2100 5124
rect 1708 4396 1764 4452
rect 1820 2492 1876 2548
rect 2828 5628 2884 5684
rect 2380 1820 2436 1876
rect 2492 5180 2548 5236
rect 2268 1036 2324 1092
rect 2604 4338 2660 4340
rect 2604 4286 2606 4338
rect 2606 4286 2658 4338
rect 2658 4286 2660 4338
rect 2604 4284 2660 4286
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 6748 10556 6804 10612
rect 3164 10332 3220 10388
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 3164 8876 3220 8932
rect 3276 9884 3332 9940
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 6636 9436 6692 9492
rect 4956 9212 5012 9268
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3276 8204 3332 8260
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4284 7868 4340 7924
rect 3388 7532 3444 7588
rect 2940 4060 2996 4116
rect 3164 4114 3220 4116
rect 3164 4062 3166 4114
rect 3166 4062 3218 4114
rect 3218 4062 3220 4114
rect 3164 4060 3220 4062
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 3836 1260 3892 1316
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 6412 8764 6468 8820
rect 5404 7362 5460 7364
rect 5404 7310 5406 7362
rect 5406 7310 5458 7362
rect 5458 7310 5460 7362
rect 5404 7308 5460 7310
rect 4956 6748 5012 6804
rect 5068 6524 5124 6580
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 5964 5964 6020 6020
rect 6076 4060 6132 4116
rect 5068 3612 5124 3668
rect 5628 3836 5684 3892
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 4844 2044 4900 2100
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 5180 924 5236 980
rect 6076 2940 6132 2996
rect 6188 3948 6244 4004
rect 6860 9324 6916 9380
rect 6748 9100 6804 9156
rect 6972 8988 7028 9044
rect 7084 11116 7140 11172
rect 6860 8652 6916 8708
rect 6748 8316 6804 8372
rect 6636 8092 6692 8148
rect 6972 8092 7028 8148
rect 6748 7644 6804 7700
rect 6636 5292 6692 5348
rect 6748 4620 6804 4676
rect 6860 6076 6916 6132
rect 7308 10892 7364 10948
rect 7644 13132 7700 13188
rect 7084 5852 7140 5908
rect 7196 10668 7252 10724
rect 6860 2380 6916 2436
rect 6972 5404 7028 5460
rect 6748 2156 6804 2212
rect 6972 2044 7028 2100
rect 7420 7756 7476 7812
rect 7196 4172 7252 4228
rect 7308 6860 7364 6916
rect 7532 7420 7588 7476
rect 7532 5740 7588 5796
rect 7532 5516 7588 5572
rect 7532 5068 7588 5124
rect 7420 3948 7476 4004
rect 9884 13580 9940 13636
rect 10668 13580 10724 13636
rect 13356 13916 13412 13972
rect 11004 12236 11060 12292
rect 11228 11900 11284 11956
rect 8540 10220 8596 10276
rect 8428 10108 8484 10164
rect 8428 8204 8484 8260
rect 9212 9996 9268 10052
rect 10108 8428 10164 8484
rect 9660 7250 9716 7252
rect 9660 7198 9662 7250
rect 9662 7198 9714 7250
rect 9714 7198 9716 7250
rect 9660 7196 9716 7198
rect 8540 6524 8596 6580
rect 7644 3276 7700 3332
rect 7756 5180 7812 5236
rect 7308 2604 7364 2660
rect 7420 3052 7476 3108
rect 6412 1260 6468 1316
rect 6524 1148 6580 1204
rect 10556 5292 10612 5348
rect 9996 4508 10052 4564
rect 9660 4060 9716 4116
rect 9212 3724 9268 3780
rect 7756 2828 7812 2884
rect 8316 2828 8372 2884
rect 7868 1596 7924 1652
rect 8764 1260 8820 1316
rect 9548 812 9604 868
rect 10444 3500 10500 3556
rect 10332 3276 10388 3332
rect 9996 1874 10052 1876
rect 9996 1822 9998 1874
rect 9998 1822 10050 1874
rect 10050 1822 10052 1874
rect 9996 1820 10052 1822
rect 10556 812 10612 868
rect 10668 588 10724 644
rect 10892 364 10948 420
rect 11004 4956 11060 5012
rect 15036 13580 15092 13636
rect 13468 11564 13524 11620
rect 15820 13804 15876 13860
rect 14364 12124 14420 12180
rect 13468 9996 13524 10052
rect 13916 10108 13972 10164
rect 13356 9884 13412 9940
rect 13916 9212 13972 9268
rect 14252 9660 14308 9716
rect 13468 9100 13524 9156
rect 13356 7644 13412 7700
rect 12796 6972 12852 7028
rect 11788 4450 11844 4452
rect 11788 4398 11790 4450
rect 11790 4398 11842 4450
rect 11842 4398 11844 4450
rect 11788 4396 11844 4398
rect 11228 4060 11284 4116
rect 12236 4114 12292 4116
rect 12236 4062 12238 4114
rect 12238 4062 12290 4114
rect 12290 4062 12292 4114
rect 12236 4060 12292 4062
rect 12348 3612 12404 3668
rect 11676 3388 11732 3444
rect 11452 1596 11508 1652
rect 11564 1148 11620 1204
rect 11564 924 11620 980
rect 11676 700 11732 756
rect 11900 1148 11956 1204
rect 13916 8092 13972 8148
rect 13692 6188 13748 6244
rect 13468 4396 13524 4452
rect 13580 5740 13636 5796
rect 13356 3724 13412 3780
rect 14588 11228 14644 11284
rect 14700 11004 14756 11060
rect 14476 10892 14532 10948
rect 14476 9660 14532 9716
rect 14588 10556 14644 10612
rect 14252 5964 14308 6020
rect 13916 4732 13972 4788
rect 14140 5852 14196 5908
rect 14588 7532 14644 7588
rect 14476 5292 14532 5348
rect 14588 6748 14644 6804
rect 14252 4396 14308 4452
rect 14140 3724 14196 3780
rect 14252 3948 14308 4004
rect 13692 3612 13748 3668
rect 13580 3276 13636 3332
rect 14140 3276 14196 3332
rect 13916 2604 13972 2660
rect 13804 1260 13860 1316
rect 12796 812 12852 868
rect 13692 1148 13748 1204
rect 13244 700 13300 756
rect 12796 140 12852 196
rect 14252 3052 14308 3108
rect 14364 2268 14420 2324
rect 14140 2156 14196 2212
rect 14476 2156 14532 2212
rect 14140 1932 14196 1988
rect 14476 476 14532 532
rect 14924 10892 14980 10948
rect 14924 10220 14980 10276
rect 15148 10332 15204 10388
rect 14812 9548 14868 9604
rect 14924 9436 14980 9492
rect 14924 8316 14980 8372
rect 15036 7756 15092 7812
rect 15036 7084 15092 7140
rect 14700 5068 14756 5124
rect 14700 2940 14756 2996
rect 14700 1596 14756 1652
rect 14812 1260 14868 1316
rect 15260 6860 15316 6916
rect 15260 4956 15316 5012
rect 18284 12684 18340 12740
rect 16492 12012 16548 12068
rect 16716 12066 16772 12068
rect 16716 12014 16718 12066
rect 16718 12014 16770 12066
rect 16770 12014 16772 12066
rect 16716 12012 16772 12014
rect 18172 12012 18228 12068
rect 17052 11788 17108 11844
rect 16828 11564 16884 11620
rect 17276 11564 17332 11620
rect 16492 10668 16548 10724
rect 16716 11116 16772 11172
rect 15932 10220 15988 10276
rect 18396 12236 18452 12292
rect 21196 13692 21252 13748
rect 19404 12236 19460 12292
rect 20636 12290 20692 12292
rect 20636 12238 20638 12290
rect 20638 12238 20690 12290
rect 20690 12238 20692 12290
rect 20636 12236 20692 12238
rect 20972 12124 21028 12180
rect 18396 11676 18452 11732
rect 18620 11900 18676 11956
rect 18284 11340 18340 11396
rect 18508 11340 18564 11396
rect 18172 11116 18228 11172
rect 17276 10780 17332 10836
rect 18060 10780 18116 10836
rect 16716 9996 16772 10052
rect 15932 6748 15988 6804
rect 16044 8204 16100 8260
rect 15932 2828 15988 2884
rect 15596 2380 15652 2436
rect 17836 7980 17892 8036
rect 16380 7420 16436 7476
rect 16156 6802 16212 6804
rect 16156 6750 16158 6802
rect 16158 6750 16210 6802
rect 16210 6750 16212 6802
rect 16156 6748 16212 6750
rect 17724 7196 17780 7252
rect 16716 6076 16772 6132
rect 16604 5516 16660 5572
rect 16380 5292 16436 5348
rect 16044 2044 16100 2100
rect 16492 4844 16548 4900
rect 16492 1932 16548 1988
rect 15260 1372 15316 1428
rect 16380 1036 16436 1092
rect 15260 476 15316 532
rect 15932 812 15988 868
rect 13916 28 13972 84
rect 16828 4060 16884 4116
rect 16828 2044 16884 2100
rect 16940 2940 16996 2996
rect 16716 1036 16772 1092
rect 16828 1596 16884 1652
rect 17276 2546 17332 2548
rect 17276 2494 17278 2546
rect 17278 2494 17330 2546
rect 17330 2494 17332 2546
rect 17276 2492 17332 2494
rect 17164 1932 17220 1988
rect 16940 1148 16996 1204
rect 17276 1036 17332 1092
rect 18396 10780 18452 10836
rect 18284 10668 18340 10724
rect 20076 11788 20132 11844
rect 20076 11452 20132 11508
rect 18732 10780 18788 10836
rect 19852 11228 19908 11284
rect 18620 10668 18676 10724
rect 18284 9660 18340 9716
rect 18396 10444 18452 10500
rect 19404 10108 19460 10164
rect 18396 8988 18452 9044
rect 18172 5740 18228 5796
rect 18060 5068 18116 5124
rect 18172 5516 18228 5572
rect 17836 4060 17892 4116
rect 17836 3388 17892 3444
rect 18508 6636 18564 6692
rect 20748 11004 20804 11060
rect 23324 13356 23380 13412
rect 23548 13468 23604 13524
rect 21980 12796 22036 12852
rect 21868 12348 21924 12404
rect 21868 11676 21924 11732
rect 22428 12796 22484 12852
rect 21980 11340 22036 11396
rect 22092 11788 22148 11844
rect 20972 8988 21028 9044
rect 21196 10668 21252 10724
rect 20748 8540 20804 8596
rect 19964 8316 20020 8372
rect 20860 8428 20916 8484
rect 20636 7084 20692 7140
rect 19852 6300 19908 6356
rect 19964 6860 20020 6916
rect 20076 6748 20132 6804
rect 20076 6412 20132 6468
rect 19964 6188 20020 6244
rect 19964 5964 20020 6020
rect 18620 5346 18676 5348
rect 18620 5294 18622 5346
rect 18622 5294 18674 5346
rect 18674 5294 18676 5346
rect 18620 5292 18676 5294
rect 18396 4172 18452 4228
rect 18732 4508 18788 4564
rect 18732 3052 18788 3108
rect 19180 2604 19236 2660
rect 19180 2380 19236 2436
rect 18620 1708 18676 1764
rect 19068 2044 19124 2100
rect 18284 1596 18340 1652
rect 17836 1148 17892 1204
rect 18172 588 18228 644
rect 18620 364 18676 420
rect 19516 1260 19572 1316
rect 20636 5964 20692 6020
rect 20972 5852 21028 5908
rect 20860 5180 20916 5236
rect 20076 5122 20132 5124
rect 20076 5070 20078 5122
rect 20078 5070 20130 5122
rect 20130 5070 20132 5122
rect 20076 5068 20132 5070
rect 20636 5068 20692 5124
rect 19964 3612 20020 3668
rect 20188 3500 20244 3556
rect 19852 3388 19908 3444
rect 19852 2828 19908 2884
rect 20188 2828 20244 2884
rect 21868 10668 21924 10724
rect 21644 10108 21700 10164
rect 21420 7362 21476 7364
rect 21420 7310 21422 7362
rect 21422 7310 21474 7362
rect 21474 7310 21476 7362
rect 21420 7308 21476 7310
rect 21196 5292 21252 5348
rect 21532 6748 21588 6804
rect 20972 4060 21028 4116
rect 21420 4060 21476 4116
rect 22204 11228 22260 11284
rect 22876 12178 22932 12180
rect 22876 12126 22878 12178
rect 22878 12126 22930 12178
rect 22930 12126 22932 12178
rect 22876 12124 22932 12126
rect 24108 13356 24164 13412
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 24332 12236 24388 12292
rect 23548 11900 23604 11956
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23548 10108 23604 10164
rect 22428 9772 22484 9828
rect 28588 13020 28644 13076
rect 25116 12236 25172 12292
rect 26460 12290 26516 12292
rect 26460 12238 26462 12290
rect 26462 12238 26514 12290
rect 26514 12238 26516 12290
rect 26460 12236 26516 12238
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 24892 11788 24948 11844
rect 24892 11452 24948 11508
rect 24332 11004 24388 11060
rect 24556 10668 24612 10724
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24220 9772 24276 9828
rect 25116 10108 25172 10164
rect 25116 9660 25172 9716
rect 22204 9548 22260 9604
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24220 9436 24276 9492
rect 22092 7532 22148 7588
rect 22204 8988 22260 9044
rect 21756 6524 21812 6580
rect 21980 6524 22036 6580
rect 21980 6300 22036 6356
rect 21644 5516 21700 5572
rect 23212 9042 23268 9044
rect 23212 8990 23214 9042
rect 23214 8990 23266 9042
rect 23266 8990 23268 9042
rect 23212 8988 23268 8990
rect 22652 8930 22708 8932
rect 22652 8878 22654 8930
rect 22654 8878 22706 8930
rect 22706 8878 22708 8930
rect 22652 8876 22708 8878
rect 22428 8652 22484 8708
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24220 8316 24276 8372
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24108 7644 24164 7700
rect 24668 7644 24724 7700
rect 25564 9996 25620 10052
rect 25564 9100 25620 9156
rect 26124 8930 26180 8932
rect 26124 8878 26126 8930
rect 26126 8878 26178 8930
rect 26178 8878 26180 8930
rect 26124 8876 26180 8878
rect 25228 7532 25284 7588
rect 25900 8092 25956 8148
rect 22988 7420 23044 7476
rect 27020 11452 27076 11508
rect 29708 13804 29764 13860
rect 29036 12178 29092 12180
rect 29036 12126 29038 12178
rect 29038 12126 29090 12178
rect 29090 12126 29092 12178
rect 29036 12124 29092 12126
rect 29484 11900 29540 11956
rect 27132 10668 27188 10724
rect 28140 11788 28196 11844
rect 26796 9884 26852 9940
rect 26908 8316 26964 8372
rect 26236 7868 26292 7924
rect 26796 8204 26852 8260
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 24892 6972 24948 7028
rect 24220 6748 24276 6804
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24220 6300 24276 6356
rect 24012 6244 24068 6246
rect 23772 5964 23828 6020
rect 22204 5516 22260 5572
rect 22652 5740 22708 5796
rect 21532 3276 21588 3332
rect 21644 5180 21700 5236
rect 21532 3052 21588 3108
rect 19740 1260 19796 1316
rect 19964 1596 20020 1652
rect 19628 252 19684 308
rect 20412 1596 20468 1652
rect 21308 1932 21364 1988
rect 22428 4508 22484 4564
rect 22204 3612 22260 3668
rect 21644 2940 21700 2996
rect 21756 3500 21812 3556
rect 21644 2380 21700 2436
rect 21644 812 21700 868
rect 21532 364 21588 420
rect 21868 1986 21924 1988
rect 21868 1934 21870 1986
rect 21870 1934 21922 1986
rect 21922 1934 21924 1986
rect 21868 1932 21924 1934
rect 22092 1202 22148 1204
rect 22092 1150 22094 1202
rect 22094 1150 22146 1202
rect 22146 1150 22148 1202
rect 22092 1148 22148 1150
rect 25452 6860 25508 6916
rect 25452 6636 25508 6692
rect 24892 5852 24948 5908
rect 23772 5516 23828 5572
rect 24780 5794 24836 5796
rect 24780 5742 24782 5794
rect 24782 5742 24834 5794
rect 24834 5742 24836 5794
rect 24780 5740 24836 5742
rect 25340 5794 25396 5796
rect 25340 5742 25342 5794
rect 25342 5742 25394 5794
rect 25394 5742 25396 5794
rect 25340 5740 25396 5742
rect 24444 5628 24500 5684
rect 25900 5628 25956 5684
rect 23884 5404 23940 5460
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 25228 5516 25284 5572
rect 24672 5460 24728 5462
rect 24892 5404 24948 5460
rect 23772 5292 23828 5348
rect 23100 5068 23156 5124
rect 22764 2098 22820 2100
rect 22764 2046 22766 2098
rect 22766 2046 22818 2098
rect 22818 2046 22820 2098
rect 22764 2044 22820 2046
rect 22876 1090 22932 1092
rect 22876 1038 22878 1090
rect 22878 1038 22930 1090
rect 22930 1038 22932 1090
rect 22876 1036 22932 1038
rect 23324 4956 23380 5012
rect 23324 4732 23380 4788
rect 25116 4844 25172 4900
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24892 4508 24948 4564
rect 23884 3836 23940 3892
rect 23548 3554 23604 3556
rect 23548 3502 23550 3554
rect 23550 3502 23602 3554
rect 23602 3502 23604 3554
rect 23548 3500 23604 3502
rect 23996 3442 24052 3444
rect 23996 3390 23998 3442
rect 23998 3390 24050 3442
rect 24050 3390 24052 3442
rect 23996 3388 24052 3390
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 23436 2940 23492 2996
rect 24220 3052 24276 3108
rect 23996 2716 24052 2772
rect 24220 2380 24276 2436
rect 23996 2044 24052 2100
rect 23324 1372 23380 1428
rect 23548 1932 23604 1988
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 24556 3666 24612 3668
rect 24556 3614 24558 3666
rect 24558 3614 24610 3666
rect 24610 3614 24612 3666
rect 24556 3612 24612 3614
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 25340 5180 25396 5236
rect 25340 4844 25396 4900
rect 25228 4284 25284 4340
rect 25676 4620 25732 4676
rect 25676 4172 25732 4228
rect 25228 3500 25284 3556
rect 24892 1932 24948 1988
rect 24892 1036 24948 1092
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 25340 3164 25396 3220
rect 25228 2604 25284 2660
rect 25116 1090 25172 1092
rect 25116 1038 25118 1090
rect 25118 1038 25170 1090
rect 25170 1038 25172 1090
rect 25116 1036 25172 1038
rect 25004 588 25060 644
rect 26012 4060 26068 4116
rect 25676 1372 25732 1428
rect 25788 1596 25844 1652
rect 26236 5628 26292 5684
rect 26460 5068 26516 5124
rect 26684 5068 26740 5124
rect 26684 4732 26740 4788
rect 26236 4508 26292 4564
rect 26236 3500 26292 3556
rect 26236 1708 26292 1764
rect 26684 1820 26740 1876
rect 27692 8092 27748 8148
rect 27580 7644 27636 7700
rect 28700 10722 28756 10724
rect 28700 10670 28702 10722
rect 28702 10670 28754 10722
rect 28754 10670 28756 10722
rect 28700 10668 28756 10670
rect 29260 10668 29316 10724
rect 28140 7980 28196 8036
rect 28476 10444 28532 10500
rect 27692 4172 27748 4228
rect 27916 6972 27972 7028
rect 27020 2268 27076 2324
rect 26796 1708 26852 1764
rect 26572 1596 26628 1652
rect 26908 1314 26964 1316
rect 26908 1262 26910 1314
rect 26910 1262 26962 1314
rect 26962 1262 26964 1314
rect 26908 1260 26964 1262
rect 26236 1036 26292 1092
rect 26684 1036 26740 1092
rect 28588 8764 28644 8820
rect 28476 5852 28532 5908
rect 28588 3612 28644 3668
rect 27916 2044 27972 2100
rect 27244 1036 27300 1092
rect 27580 1260 27636 1316
rect 28588 2940 28644 2996
rect 28700 2546 28756 2548
rect 28700 2494 28702 2546
rect 28702 2494 28754 2546
rect 28754 2494 28756 2546
rect 28700 2492 28756 2494
rect 29708 11676 29764 11732
rect 29820 12684 29876 12740
rect 29484 9100 29540 9156
rect 29596 11004 29652 11060
rect 29260 8370 29316 8372
rect 29260 8318 29262 8370
rect 29262 8318 29314 8370
rect 29314 8318 29316 8370
rect 29260 8316 29316 8318
rect 29820 11004 29876 11060
rect 29932 11788 29988 11844
rect 29820 10444 29876 10500
rect 29708 10332 29764 10388
rect 29708 8540 29764 8596
rect 33068 13916 33124 13972
rect 32396 13132 32452 13188
rect 30268 11564 30324 11620
rect 30044 9884 30100 9940
rect 30156 10892 30212 10948
rect 29932 9436 29988 9492
rect 30044 9212 30100 9268
rect 29596 8092 29652 8148
rect 29820 5346 29876 5348
rect 29820 5294 29822 5346
rect 29822 5294 29874 5346
rect 29874 5294 29876 5346
rect 29820 5292 29876 5294
rect 28924 3724 28980 3780
rect 29148 2940 29204 2996
rect 28140 1148 28196 1204
rect 29260 2492 29316 2548
rect 30268 9996 30324 10052
rect 30156 5292 30212 5348
rect 32844 12962 32900 12964
rect 32844 12910 32846 12962
rect 32846 12910 32898 12962
rect 32898 12910 32900 12962
rect 32844 12908 32900 12910
rect 30828 12012 30884 12068
rect 30604 9212 30660 9268
rect 30716 10556 30772 10612
rect 30492 8652 30548 8708
rect 30156 5068 30212 5124
rect 30044 4844 30100 4900
rect 30156 3724 30212 3780
rect 29596 2156 29652 2212
rect 32956 10780 33012 10836
rect 32956 10332 33012 10388
rect 32396 10108 32452 10164
rect 31388 8316 31444 8372
rect 31612 8540 31668 8596
rect 30492 4284 30548 4340
rect 30940 3164 30996 3220
rect 31500 7980 31556 8036
rect 31164 2940 31220 2996
rect 31276 7084 31332 7140
rect 30940 2828 30996 2884
rect 30492 2770 30548 2772
rect 30492 2718 30494 2770
rect 30494 2718 30546 2770
rect 30546 2718 30548 2770
rect 30492 2716 30548 2718
rect 30156 1932 30212 1988
rect 30156 1596 30212 1652
rect 30716 2268 30772 2324
rect 29372 924 29428 980
rect 30156 978 30212 980
rect 30156 926 30158 978
rect 30158 926 30210 978
rect 30210 926 30212 978
rect 30156 924 30212 926
rect 29820 812 29876 868
rect 31836 8428 31892 8484
rect 31836 6188 31892 6244
rect 32060 6636 32116 6692
rect 31836 5852 31892 5908
rect 31612 4620 31668 4676
rect 31724 5516 31780 5572
rect 31500 4508 31556 4564
rect 31388 2716 31444 2772
rect 31388 1932 31444 1988
rect 31612 2492 31668 2548
rect 30716 700 30772 756
rect 31164 1820 31220 1876
rect 30716 476 30772 532
rect 31500 1202 31556 1204
rect 31500 1150 31502 1202
rect 31502 1150 31554 1202
rect 31554 1150 31556 1202
rect 31500 1148 31556 1150
rect 32060 5852 32116 5908
rect 31948 5516 32004 5572
rect 32620 9938 32676 9940
rect 32620 9886 32622 9938
rect 32622 9886 32674 9938
rect 32674 9886 32676 9938
rect 32620 9884 32676 9886
rect 32844 9548 32900 9604
rect 32732 5516 32788 5572
rect 34748 12908 34804 12964
rect 34524 11004 34580 11060
rect 33068 9884 33124 9940
rect 34636 9938 34692 9940
rect 34636 9886 34638 9938
rect 34638 9886 34690 9938
rect 34690 9886 34692 9938
rect 34636 9884 34692 9886
rect 33180 9660 33236 9716
rect 33740 8092 33796 8148
rect 33740 6748 33796 6804
rect 33628 6076 33684 6132
rect 31724 1260 31780 1316
rect 32060 812 32116 868
rect 32844 3276 32900 3332
rect 32732 2716 32788 2772
rect 33852 6076 33908 6132
rect 33740 5516 33796 5572
rect 33852 5068 33908 5124
rect 33964 5292 34020 5348
rect 33740 4844 33796 4900
rect 33628 4284 33684 4340
rect 32956 2716 33012 2772
rect 33628 3052 33684 3108
rect 32396 2604 32452 2660
rect 33068 2604 33124 2660
rect 32620 2546 32676 2548
rect 32620 2494 32622 2546
rect 32622 2494 32674 2546
rect 32674 2494 32676 2546
rect 32620 2492 32676 2494
rect 32956 1874 33012 1876
rect 32956 1822 32958 1874
rect 32958 1822 33010 1874
rect 33010 1822 33012 1874
rect 32956 1820 33012 1822
rect 32508 1708 32564 1764
rect 33516 2268 33572 2324
rect 33068 1372 33124 1428
rect 34636 4956 34692 5012
rect 36876 12348 36932 12404
rect 35532 12066 35588 12068
rect 35532 12014 35534 12066
rect 35534 12014 35586 12066
rect 35586 12014 35588 12066
rect 35532 12012 35588 12014
rect 35308 11788 35364 11844
rect 35084 11116 35140 11172
rect 35196 11340 35252 11396
rect 34972 10780 35028 10836
rect 35084 10610 35140 10612
rect 35084 10558 35086 10610
rect 35086 10558 35138 10610
rect 35138 10558 35140 10610
rect 35084 10556 35140 10558
rect 35980 11676 36036 11732
rect 35644 11116 35700 11172
rect 35308 9884 35364 9940
rect 35308 8540 35364 8596
rect 34748 3612 34804 3668
rect 34860 7084 34916 7140
rect 33964 2828 34020 2884
rect 34076 2658 34132 2660
rect 34076 2606 34078 2658
rect 34078 2606 34130 2658
rect 34130 2606 34132 2658
rect 34076 2604 34132 2606
rect 33628 1596 33684 1652
rect 33852 1820 33908 1876
rect 33516 1036 33572 1092
rect 33404 924 33460 980
rect 33628 476 33684 532
rect 34188 1762 34244 1764
rect 34188 1710 34190 1762
rect 34190 1710 34242 1762
rect 34242 1710 34244 1762
rect 34188 1708 34244 1710
rect 35084 6972 35140 7028
rect 35308 6524 35364 6580
rect 35196 5852 35252 5908
rect 35196 5404 35252 5460
rect 35196 5122 35252 5124
rect 35196 5070 35198 5122
rect 35198 5070 35250 5122
rect 35250 5070 35252 5122
rect 35196 5068 35252 5070
rect 35196 4620 35252 4676
rect 35644 7644 35700 7700
rect 35756 5906 35812 5908
rect 35756 5854 35758 5906
rect 35758 5854 35810 5906
rect 35810 5854 35812 5906
rect 35756 5852 35812 5854
rect 35420 4844 35476 4900
rect 35644 4956 35700 5012
rect 35980 4956 36036 5012
rect 36092 8652 36148 8708
rect 35308 4508 35364 4564
rect 34860 3164 34916 3220
rect 35532 3052 35588 3108
rect 34860 2770 34916 2772
rect 34860 2718 34862 2770
rect 34862 2718 34914 2770
rect 34914 2718 34916 2770
rect 34860 2716 34916 2718
rect 35084 2604 35140 2660
rect 36092 4060 36148 4116
rect 36204 5852 36260 5908
rect 35756 3276 35812 3332
rect 35644 2716 35700 2772
rect 36764 4060 36820 4116
rect 36316 3836 36372 3892
rect 45052 13692 45108 13748
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 42140 13020 42196 13076
rect 43372 13074 43428 13076
rect 43372 13022 43374 13074
rect 43374 13022 43426 13074
rect 43426 13022 43428 13074
rect 43372 13020 43428 13022
rect 40124 12460 40180 12516
rect 38220 12236 38276 12292
rect 39900 12290 39956 12292
rect 39900 12238 39902 12290
rect 39902 12238 39954 12290
rect 39954 12238 39956 12290
rect 39900 12236 39956 12238
rect 37100 12066 37156 12068
rect 37100 12014 37102 12066
rect 37102 12014 37154 12066
rect 37154 12014 37156 12066
rect 37100 12012 37156 12014
rect 36988 11900 37044 11956
rect 36988 6636 37044 6692
rect 37100 8764 37156 8820
rect 38556 10780 38612 10836
rect 40236 12012 40292 12068
rect 40460 11788 40516 11844
rect 40236 10892 40292 10948
rect 37996 9996 38052 10052
rect 40348 8092 40404 8148
rect 37660 7532 37716 7588
rect 37100 6300 37156 6356
rect 40684 6524 40740 6580
rect 37324 5292 37380 5348
rect 35308 2156 35364 2212
rect 35196 2098 35252 2100
rect 35196 2046 35198 2098
rect 35198 2046 35250 2098
rect 35250 2046 35252 2098
rect 35196 2044 35252 2046
rect 35756 2044 35812 2100
rect 35756 1874 35812 1876
rect 35756 1822 35758 1874
rect 35758 1822 35810 1874
rect 35810 1822 35812 1874
rect 35756 1820 35812 1822
rect 37212 5068 37268 5124
rect 35644 1708 35700 1764
rect 34748 812 34804 868
rect 35308 1202 35364 1204
rect 35308 1150 35310 1202
rect 35310 1150 35362 1202
rect 35362 1150 35364 1202
rect 35308 1148 35364 1150
rect 36988 2828 37044 2884
rect 36876 2492 36932 2548
rect 36764 1986 36820 1988
rect 36764 1934 36766 1986
rect 36766 1934 36818 1986
rect 36818 1934 36820 1986
rect 36764 1932 36820 1934
rect 35868 978 35924 980
rect 35868 926 35870 978
rect 35870 926 35922 978
rect 35922 926 35924 978
rect 35868 924 35924 926
rect 36540 1036 36596 1092
rect 15708 28 15764 84
rect 36876 1260 36932 1316
rect 37100 2658 37156 2660
rect 37100 2606 37102 2658
rect 37102 2606 37154 2658
rect 37154 2606 37156 2658
rect 37100 2604 37156 2606
rect 37548 5068 37604 5124
rect 39116 5122 39172 5124
rect 39116 5070 39118 5122
rect 39118 5070 39170 5122
rect 39170 5070 39172 5122
rect 39116 5068 39172 5070
rect 38668 4732 38724 4788
rect 39228 4338 39284 4340
rect 39228 4286 39230 4338
rect 39230 4286 39282 4338
rect 39282 4286 39284 4338
rect 39228 4284 39284 4286
rect 39116 4060 39172 4116
rect 38108 2882 38164 2884
rect 38108 2830 38110 2882
rect 38110 2830 38162 2882
rect 38162 2830 38164 2882
rect 38108 2828 38164 2830
rect 37324 1762 37380 1764
rect 37324 1710 37326 1762
rect 37326 1710 37378 1762
rect 37378 1710 37380 1762
rect 37324 1708 37380 1710
rect 40348 3500 40404 3556
rect 39116 2770 39172 2772
rect 39116 2718 39118 2770
rect 39118 2718 39170 2770
rect 39170 2718 39172 2770
rect 39116 2716 39172 2718
rect 38332 2604 38388 2660
rect 37436 978 37492 980
rect 37436 926 37438 978
rect 37438 926 37490 978
rect 37490 926 37492 978
rect 37436 924 37492 926
rect 37884 476 37940 532
rect 39900 2658 39956 2660
rect 39900 2606 39902 2658
rect 39902 2606 39954 2658
rect 39954 2606 39956 2658
rect 39900 2604 39956 2606
rect 39228 1986 39284 1988
rect 39228 1934 39230 1986
rect 39230 1934 39282 1986
rect 39282 1934 39284 1986
rect 39228 1932 39284 1934
rect 38668 1596 38724 1652
rect 39676 1596 39732 1652
rect 39564 1090 39620 1092
rect 39564 1038 39566 1090
rect 39566 1038 39618 1090
rect 39618 1038 39620 1090
rect 39564 1036 39620 1038
rect 38780 812 38836 868
rect 39228 700 39284 756
rect 40124 924 40180 980
rect 40460 2716 40516 2772
rect 40348 2604 40404 2660
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 43372 11788 43428 11844
rect 41132 8818 41188 8820
rect 41132 8766 41134 8818
rect 41134 8766 41186 8818
rect 41186 8766 41188 8818
rect 41132 8764 41188 8766
rect 41692 8764 41748 8820
rect 43148 7532 43204 7588
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 44156 8652 44212 8708
rect 43372 6748 43428 6804
rect 43484 8428 43540 8484
rect 43260 6690 43316 6692
rect 43260 6638 43262 6690
rect 43262 6638 43314 6690
rect 43314 6638 43316 6690
rect 43260 6636 43316 6638
rect 40908 5292 40964 5348
rect 41692 6188 41748 6244
rect 41356 4956 41412 5012
rect 41132 4620 41188 4676
rect 41132 3836 41188 3892
rect 41468 4508 41524 4564
rect 41692 4284 41748 4340
rect 41804 5740 41860 5796
rect 41916 5068 41972 5124
rect 40572 1596 40628 1652
rect 41020 1484 41076 1540
rect 40460 812 40516 868
rect 40572 1036 40628 1092
rect 40236 252 40292 308
rect 40908 476 40964 532
rect 41468 2828 41524 2884
rect 41244 924 41300 980
rect 41468 1596 41524 1652
rect 42028 4060 42084 4116
rect 42252 4060 42308 4116
rect 41916 924 41972 980
rect 43148 5122 43204 5124
rect 43148 5070 43150 5122
rect 43150 5070 43202 5122
rect 43202 5070 43204 5122
rect 43148 5068 43204 5070
rect 42588 1708 42644 1764
rect 42812 3500 42868 3556
rect 42364 1596 42420 1652
rect 42028 700 42084 756
rect 42364 140 42420 196
rect 43484 5852 43540 5908
rect 43372 3948 43428 4004
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 43820 7532 43876 7588
rect 43820 7084 43876 7140
rect 44156 6748 44212 6804
rect 43708 6578 43764 6580
rect 43708 6526 43710 6578
rect 43710 6526 43762 6578
rect 43762 6526 43764 6578
rect 43708 6524 43764 6526
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 44604 11954 44660 11956
rect 44604 11902 44606 11954
rect 44606 11902 44658 11954
rect 44658 11902 44660 11954
rect 44604 11900 44660 11902
rect 44940 11954 44996 11956
rect 44940 11902 44942 11954
rect 44942 11902 44994 11954
rect 44994 11902 44996 11954
rect 44940 11900 44996 11902
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44940 11116 44996 11172
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 44716 8930 44772 8932
rect 44716 8878 44718 8930
rect 44718 8878 44770 8930
rect 44770 8878 44772 8930
rect 44716 8876 44772 8878
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44828 5964 44884 6020
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 44268 4956 44324 5012
rect 44156 4844 44212 4900
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 45388 11788 45444 11844
rect 45388 8988 45444 9044
rect 45052 6300 45108 6356
rect 45164 8204 45220 8260
rect 45052 4620 45108 4676
rect 44380 4508 44436 4564
rect 45052 4396 45108 4452
rect 44940 4338 44996 4340
rect 44940 4286 44942 4338
rect 44942 4286 44994 4338
rect 44994 4286 44996 4338
rect 44940 4284 44996 4286
rect 44268 3948 44324 4004
rect 44464 3946 44520 3948
rect 43596 3836 43652 3892
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44828 3948 44884 4004
rect 44672 3892 44728 3894
rect 43932 3500 43988 3556
rect 45276 5068 45332 5124
rect 45500 5068 45556 5124
rect 45500 4060 45556 4116
rect 43036 3052 43092 3108
rect 43372 2098 43428 2100
rect 43372 2046 43374 2098
rect 43374 2046 43426 2098
rect 43426 2046 43428 2098
rect 43372 2044 43428 2046
rect 43036 1986 43092 1988
rect 43036 1934 43038 1986
rect 43038 1934 43090 1986
rect 43090 1934 43092 1986
rect 43036 1932 43092 1934
rect 43260 1260 43316 1316
rect 43372 1090 43428 1092
rect 43372 1038 43374 1090
rect 43374 1038 43426 1090
rect 43426 1038 43428 1090
rect 43372 1036 43428 1038
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 45052 3052 45108 3108
rect 43596 2044 43652 2100
rect 43932 1762 43988 1764
rect 43932 1710 43934 1762
rect 43934 1710 43986 1762
rect 43986 1710 43988 1762
rect 43932 1708 43988 1710
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 44156 1484 44212 1540
rect 43596 1036 43652 1092
rect 43708 476 43764 532
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 45276 2828 45332 2884
rect 44940 2604 44996 2660
rect 44828 1260 44884 1316
rect 44492 1202 44548 1204
rect 44492 1150 44494 1202
rect 44494 1150 44546 1202
rect 44546 1150 44548 1202
rect 44492 1148 44548 1150
rect 45052 978 45108 980
rect 45052 926 45054 978
rect 45054 926 45106 978
rect 45106 926 45108 978
rect 45052 924 45108 926
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 44268 364 44324 420
rect 44604 588 44660 644
rect 44156 252 44212 308
rect 49980 14028 50036 14084
rect 46844 12684 46900 12740
rect 47180 12012 47236 12068
rect 47068 11282 47124 11284
rect 47068 11230 47070 11282
rect 47070 11230 47122 11282
rect 47122 11230 47124 11282
rect 47068 11228 47124 11230
rect 46172 9660 46228 9716
rect 45724 3388 45780 3444
rect 45724 3276 45780 3332
rect 45612 3164 45668 3220
rect 45724 3052 45780 3108
rect 45388 588 45444 644
rect 45500 812 45556 868
rect 45052 364 45108 420
rect 45724 140 45780 196
rect 45948 1708 46004 1764
rect 46508 7196 46564 7252
rect 46620 5906 46676 5908
rect 46620 5854 46622 5906
rect 46622 5854 46674 5906
rect 46674 5854 46676 5906
rect 46620 5852 46676 5854
rect 47180 5404 47236 5460
rect 46732 5292 46788 5348
rect 46620 4226 46676 4228
rect 46620 4174 46622 4226
rect 46622 4174 46674 4226
rect 46674 4174 46676 4226
rect 46620 4172 46676 4174
rect 46620 3612 46676 3668
rect 46508 3164 46564 3220
rect 46172 1148 46228 1204
rect 47068 5180 47124 5236
rect 47404 12066 47460 12068
rect 47404 12014 47406 12066
rect 47406 12014 47458 12066
rect 47458 12014 47460 12066
rect 47404 12012 47460 12014
rect 47740 11900 47796 11956
rect 47516 7196 47572 7252
rect 47516 5122 47572 5124
rect 47516 5070 47518 5122
rect 47518 5070 47570 5122
rect 47570 5070 47572 5122
rect 47516 5068 47572 5070
rect 47292 4844 47348 4900
rect 47180 3612 47236 3668
rect 46732 3276 46788 3332
rect 47292 2770 47348 2772
rect 47292 2718 47294 2770
rect 47294 2718 47346 2770
rect 47346 2718 47348 2770
rect 47292 2716 47348 2718
rect 46956 1932 47012 1988
rect 47068 1820 47124 1876
rect 46284 252 46340 308
rect 46732 1372 46788 1428
rect 46844 1260 46900 1316
rect 47292 476 47348 532
rect 47292 252 47348 308
rect 49084 11452 49140 11508
rect 48860 9212 48916 9268
rect 48748 7980 48804 8036
rect 48188 7196 48244 7252
rect 48076 3388 48132 3444
rect 47852 1708 47908 1764
rect 48860 6748 48916 6804
rect 48972 7532 49028 7588
rect 48748 5852 48804 5908
rect 48748 4732 48804 4788
rect 48412 3948 48468 4004
rect 48300 3554 48356 3556
rect 48300 3502 48302 3554
rect 48302 3502 48354 3554
rect 48354 3502 48356 3554
rect 48300 3500 48356 3502
rect 48636 2604 48692 2660
rect 48860 3554 48916 3556
rect 48860 3502 48862 3554
rect 48862 3502 48914 3554
rect 48914 3502 48916 3554
rect 48860 3500 48916 3502
rect 48748 2268 48804 2324
rect 48636 1484 48692 1540
rect 50204 14028 50260 14084
rect 50764 14028 50820 14084
rect 54908 13580 54964 13636
rect 51772 12962 51828 12964
rect 51772 12910 51774 12962
rect 51774 12910 51826 12962
rect 51826 12910 51828 12962
rect 51772 12908 51828 12910
rect 50988 12012 51044 12068
rect 49084 1596 49140 1652
rect 48748 812 48804 868
rect 48636 700 48692 756
rect 51996 11282 52052 11284
rect 51996 11230 51998 11282
rect 51998 11230 52050 11282
rect 52050 11230 52052 11282
rect 51996 11228 52052 11230
rect 51884 10668 51940 10724
rect 50204 6300 50260 6356
rect 49420 6076 49476 6132
rect 49532 5740 49588 5796
rect 49420 1260 49476 1316
rect 49308 700 49364 756
rect 48860 364 48916 420
rect 49084 140 49140 196
rect 49980 5794 50036 5796
rect 49980 5742 49982 5794
rect 49982 5742 50034 5794
rect 50034 5742 50036 5794
rect 49980 5740 50036 5742
rect 49980 4844 50036 4900
rect 49756 3836 49812 3892
rect 49644 2492 49700 2548
rect 50988 5404 51044 5460
rect 50428 4508 50484 4564
rect 50764 3666 50820 3668
rect 50764 3614 50766 3666
rect 50766 3614 50818 3666
rect 50818 3614 50820 3666
rect 50764 3612 50820 3614
rect 50428 2716 50484 2772
rect 50876 2940 50932 2996
rect 50876 2268 50932 2324
rect 50540 252 50596 308
rect 50204 140 50260 196
rect 50428 140 50484 196
rect 51660 4732 51716 4788
rect 51324 3948 51380 4004
rect 51212 3276 51268 3332
rect 51436 2044 51492 2100
rect 51772 1986 51828 1988
rect 51772 1934 51774 1986
rect 51774 1934 51826 1986
rect 51826 1934 51828 1986
rect 51772 1932 51828 1934
rect 52108 10610 52164 10612
rect 52108 10558 52110 10610
rect 52110 10558 52162 10610
rect 52162 10558 52164 10610
rect 52108 10556 52164 10558
rect 52220 10220 52276 10276
rect 52108 8764 52164 8820
rect 52108 6860 52164 6916
rect 52668 12908 52724 12964
rect 52556 11394 52612 11396
rect 52556 11342 52558 11394
rect 52558 11342 52610 11394
rect 52610 11342 52612 11394
rect 52556 11340 52612 11342
rect 52556 9826 52612 9828
rect 52556 9774 52558 9826
rect 52558 9774 52610 9826
rect 52610 9774 52612 9826
rect 52556 9772 52612 9774
rect 52444 8540 52500 8596
rect 52220 3388 52276 3444
rect 52108 2156 52164 2212
rect 53004 12402 53060 12404
rect 53004 12350 53006 12402
rect 53006 12350 53058 12402
rect 53058 12350 53060 12402
rect 53004 12348 53060 12350
rect 53564 12178 53620 12180
rect 53564 12126 53566 12178
rect 53566 12126 53618 12178
rect 53618 12126 53620 12178
rect 53564 12124 53620 12126
rect 54348 12066 54404 12068
rect 54348 12014 54350 12066
rect 54350 12014 54402 12066
rect 54402 12014 54404 12066
rect 54348 12012 54404 12014
rect 53564 11170 53620 11172
rect 53564 11118 53566 11170
rect 53566 11118 53618 11170
rect 53618 11118 53620 11170
rect 53564 11116 53620 11118
rect 53004 11004 53060 11060
rect 54124 10780 54180 10836
rect 53564 10498 53620 10500
rect 53564 10446 53566 10498
rect 53566 10446 53618 10498
rect 53618 10446 53620 10498
rect 53564 10444 53620 10446
rect 53116 10220 53172 10276
rect 52780 5740 52836 5796
rect 52556 3724 52612 3780
rect 52668 3500 52724 3556
rect 51324 1596 51380 1652
rect 51996 924 52052 980
rect 52220 1148 52276 1204
rect 52892 5346 52948 5348
rect 52892 5294 52894 5346
rect 52894 5294 52946 5346
rect 52946 5294 52948 5346
rect 52892 5292 52948 5294
rect 54572 10108 54628 10164
rect 53564 9714 53620 9716
rect 53564 9662 53566 9714
rect 53566 9662 53618 9714
rect 53618 9662 53620 9714
rect 53564 9660 53620 9662
rect 54124 8370 54180 8372
rect 54124 8318 54126 8370
rect 54126 8318 54178 8370
rect 54178 8318 54180 8370
rect 54124 8316 54180 8318
rect 53564 7644 53620 7700
rect 53564 7474 53620 7476
rect 53564 7422 53566 7474
rect 53566 7422 53618 7474
rect 53618 7422 53620 7474
rect 53564 7420 53620 7422
rect 55580 12348 55636 12404
rect 55804 13916 55860 13972
rect 55132 11788 55188 11844
rect 56476 13468 56532 13524
rect 55804 11228 55860 11284
rect 55132 10780 55188 10836
rect 55132 10332 55188 10388
rect 56140 11228 56196 11284
rect 56364 12124 56420 12180
rect 56364 11116 56420 11172
rect 55916 10332 55972 10388
rect 55356 9884 55412 9940
rect 55132 9436 55188 9492
rect 55020 9100 55076 9156
rect 54348 8540 54404 8596
rect 54908 8370 54964 8372
rect 54908 8318 54910 8370
rect 54910 8318 54962 8370
rect 54962 8318 54964 8370
rect 54908 8316 54964 8318
rect 54572 7196 54628 7252
rect 54236 6972 54292 7028
rect 53676 6748 53732 6804
rect 53452 6524 53508 6580
rect 53228 5628 53284 5684
rect 53228 4114 53284 4116
rect 53228 4062 53230 4114
rect 53230 4062 53282 4114
rect 53282 4062 53284 4114
rect 53228 4060 53284 4062
rect 53116 3612 53172 3668
rect 53004 2882 53060 2884
rect 53004 2830 53006 2882
rect 53006 2830 53058 2882
rect 53058 2830 53060 2882
rect 53004 2828 53060 2830
rect 53116 1036 53172 1092
rect 53564 5906 53620 5908
rect 53564 5854 53566 5906
rect 53566 5854 53618 5906
rect 53618 5854 53620 5906
rect 53564 5852 53620 5854
rect 54124 6412 54180 6468
rect 54236 6636 54292 6692
rect 54572 5852 54628 5908
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 54124 4620 54180 4676
rect 53564 3500 53620 3556
rect 53564 2770 53620 2772
rect 53564 2718 53566 2770
rect 53566 2718 53618 2770
rect 53618 2718 53620 2770
rect 53564 2716 53620 2718
rect 54572 4562 54628 4564
rect 54572 4510 54574 4562
rect 54574 4510 54626 4562
rect 54626 4510 54628 4562
rect 54572 4508 54628 4510
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 53676 2604 53732 2660
rect 54460 3388 54516 3444
rect 54124 2098 54180 2100
rect 54124 2046 54126 2098
rect 54126 2046 54178 2098
rect 54178 2046 54180 2098
rect 54124 2044 54180 2046
rect 54012 1932 54068 1988
rect 53564 1874 53620 1876
rect 53564 1822 53566 1874
rect 53566 1822 53618 1874
rect 53618 1822 53620 1874
rect 53564 1820 53620 1822
rect 53564 1426 53620 1428
rect 53564 1374 53566 1426
rect 53566 1374 53618 1426
rect 53618 1374 53620 1426
rect 53564 1372 53620 1374
rect 54572 3164 54628 3220
rect 55132 8876 55188 8932
rect 55244 7308 55300 7364
rect 55244 6860 55300 6916
rect 55132 6300 55188 6356
rect 57036 13020 57092 13076
rect 56700 12572 56756 12628
rect 56700 11004 56756 11060
rect 56476 9660 56532 9716
rect 56140 8988 56196 9044
rect 57260 10108 57316 10164
rect 57260 9884 57316 9940
rect 57036 8316 57092 8372
rect 55916 8092 55972 8148
rect 56140 7698 56196 7700
rect 56140 7646 56142 7698
rect 56142 7646 56194 7698
rect 56194 7646 56196 7698
rect 56140 7644 56196 7646
rect 56140 6748 56196 6804
rect 56140 5404 56196 5460
rect 56252 5292 56308 5348
rect 55804 4060 55860 4116
rect 55356 3836 55412 3892
rect 54908 2268 54964 2324
rect 55132 1708 55188 1764
rect 54908 1484 54964 1540
rect 56140 4060 56196 4116
rect 56140 2716 56196 2772
rect 56700 3948 56756 4004
rect 56812 3500 56868 3556
rect 56812 476 56868 532
rect 56924 2828 56980 2884
rect 36764 28 36820 84
rect 56924 28 56980 84
<< metal3 >>
rect 4498 14028 4508 14084
rect 4564 14028 5068 14084
rect 5124 14028 5134 14084
rect 8082 14028 8092 14084
rect 8148 14028 49980 14084
rect 50036 14028 50046 14084
rect 50194 14028 50204 14084
rect 50260 14028 50764 14084
rect 50820 14028 50830 14084
rect 0 13972 112 14000
rect 57344 13972 57456 14000
rect 0 13916 7308 13972
rect 7364 13916 7374 13972
rect 13346 13916 13356 13972
rect 13412 13916 33068 13972
rect 33124 13916 33134 13972
rect 55794 13916 55804 13972
rect 55860 13916 57456 13972
rect 0 13888 112 13916
rect 57344 13888 57456 13916
rect 15810 13804 15820 13860
rect 15876 13804 29708 13860
rect 29764 13804 29774 13860
rect 21186 13692 21196 13748
rect 21252 13692 45052 13748
rect 45108 13692 45118 13748
rect 9874 13580 9884 13636
rect 9940 13580 10668 13636
rect 10724 13580 10734 13636
rect 15026 13580 15036 13636
rect 15092 13580 54908 13636
rect 54964 13580 54974 13636
rect 0 13524 112 13552
rect 57344 13524 57456 13552
rect 0 13468 23548 13524
rect 23604 13468 23614 13524
rect 56466 13468 56476 13524
rect 56532 13468 57456 13524
rect 0 13440 112 13468
rect 57344 13440 57456 13468
rect 23314 13356 23324 13412
rect 23380 13356 24108 13412
rect 24164 13356 24174 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 7634 13132 7644 13188
rect 7700 13132 32396 13188
rect 32452 13132 32462 13188
rect 0 13076 112 13104
rect 57344 13076 57456 13104
rect 0 13020 4228 13076
rect 6850 13020 6860 13076
rect 6916 13020 28588 13076
rect 28644 13020 28654 13076
rect 42130 13020 42140 13076
rect 42196 13020 43372 13076
rect 43428 13020 43438 13076
rect 57026 13020 57036 13076
rect 57092 13020 57456 13076
rect 0 12992 112 13020
rect 4172 12964 4228 13020
rect 57344 12992 57456 13020
rect 4172 12908 5292 12964
rect 5348 12908 5358 12964
rect 32834 12908 32844 12964
rect 32900 12908 34748 12964
rect 34804 12908 34814 12964
rect 51762 12908 51772 12964
rect 51828 12908 52668 12964
rect 52724 12908 52734 12964
rect 6066 12796 6076 12852
rect 6132 12796 21980 12852
rect 22036 12796 22046 12852
rect 22418 12796 22428 12852
rect 22484 12796 38668 12852
rect 38612 12740 38668 12796
rect 18274 12684 18284 12740
rect 18340 12684 29820 12740
rect 29876 12684 29886 12740
rect 38612 12684 46844 12740
rect 46900 12684 46910 12740
rect 0 12628 112 12656
rect 57344 12628 57456 12656
rect 0 12572 1596 12628
rect 1652 12572 1662 12628
rect 56690 12572 56700 12628
rect 56756 12572 57456 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 57344 12544 57456 12572
rect 14242 12460 14252 12516
rect 14308 12460 21028 12516
rect 20972 12292 21028 12460
rect 37100 12460 40124 12516
rect 40180 12460 40190 12516
rect 21858 12348 21868 12404
rect 21924 12348 36876 12404
rect 36932 12348 36942 12404
rect 37100 12292 37156 12460
rect 52994 12348 53004 12404
rect 53060 12348 55580 12404
rect 55636 12348 55646 12404
rect 10994 12236 11004 12292
rect 11060 12236 18396 12292
rect 18452 12236 18462 12292
rect 19394 12236 19404 12292
rect 19460 12236 20636 12292
rect 20692 12236 20702 12292
rect 20972 12236 24332 12292
rect 24388 12236 24398 12292
rect 25106 12236 25116 12292
rect 25172 12236 26460 12292
rect 26516 12236 26526 12292
rect 26852 12236 37156 12292
rect 38210 12236 38220 12292
rect 38276 12236 39900 12292
rect 39956 12236 39966 12292
rect 0 12180 112 12208
rect 26852 12180 26908 12236
rect 57344 12180 57456 12208
rect 0 12124 364 12180
rect 420 12124 430 12180
rect 14354 12124 14364 12180
rect 14420 12124 20972 12180
rect 21028 12124 21038 12180
rect 22866 12124 22876 12180
rect 22932 12124 26908 12180
rect 29026 12124 29036 12180
rect 29092 12124 53564 12180
rect 53620 12124 53630 12180
rect 56354 12124 56364 12180
rect 56420 12124 57456 12180
rect 0 12096 112 12124
rect 57344 12096 57456 12124
rect 6962 12012 6972 12068
rect 7028 12012 16492 12068
rect 16548 12012 16558 12068
rect 16706 12012 16716 12068
rect 16772 12012 18172 12068
rect 18228 12012 18238 12068
rect 18844 12012 30828 12068
rect 30884 12012 30894 12068
rect 35522 12012 35532 12068
rect 35588 12012 37100 12068
rect 37156 12012 37166 12068
rect 40226 12012 40236 12068
rect 40292 12012 47180 12068
rect 47236 12012 47246 12068
rect 47394 12012 47404 12068
rect 47460 12012 50988 12068
rect 51044 12012 51054 12068
rect 54338 12012 54348 12068
rect 54404 12012 55468 12068
rect 1820 11900 6860 11956
rect 6916 11900 6926 11956
rect 11218 11900 11228 11956
rect 11284 11900 18620 11956
rect 18676 11900 18686 11956
rect 0 11732 112 11760
rect 1820 11732 1876 11900
rect 18844 11844 18900 12012
rect 23538 11900 23548 11956
rect 23604 11900 29484 11956
rect 29540 11900 29550 11956
rect 36978 11900 36988 11956
rect 37044 11900 44604 11956
rect 44660 11900 44670 11956
rect 44930 11900 44940 11956
rect 44996 11900 47740 11956
rect 47796 11900 47806 11956
rect 17042 11788 17052 11844
rect 17108 11788 18900 11844
rect 20066 11788 20076 11844
rect 20132 11788 22092 11844
rect 22148 11788 22158 11844
rect 24882 11788 24892 11844
rect 24948 11788 28140 11844
rect 28196 11788 28206 11844
rect 29922 11788 29932 11844
rect 29988 11788 35308 11844
rect 35364 11788 35374 11844
rect 40450 11788 40460 11844
rect 40516 11788 43372 11844
rect 43428 11788 43438 11844
rect 45378 11788 45388 11844
rect 45444 11788 55132 11844
rect 55188 11788 55198 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 55412 11732 55468 12012
rect 57344 11732 57456 11760
rect 0 11676 1876 11732
rect 5282 11676 5292 11732
rect 5348 11676 16828 11732
rect 18386 11676 18396 11732
rect 18452 11676 21868 11732
rect 21924 11676 21934 11732
rect 29698 11676 29708 11732
rect 29764 11676 35980 11732
rect 36036 11676 36046 11732
rect 55412 11676 57456 11732
rect 0 11648 112 11676
rect 13458 11564 13468 11620
rect 13524 11564 16660 11620
rect 16772 11564 16828 11676
rect 57344 11648 57456 11676
rect 16884 11564 16894 11620
rect 17266 11564 17276 11620
rect 17332 11564 30268 11620
rect 30324 11564 30334 11620
rect 16604 11508 16660 11564
rect 1586 11452 1596 11508
rect 1652 11452 8428 11508
rect 16604 11452 20076 11508
rect 20132 11452 20142 11508
rect 20300 11452 24892 11508
rect 24948 11452 24958 11508
rect 27010 11452 27020 11508
rect 27076 11452 49084 11508
rect 49140 11452 49150 11508
rect 8372 11396 8428 11452
rect 20300 11396 20356 11452
rect 8372 11340 18284 11396
rect 18340 11340 18350 11396
rect 18498 11340 18508 11396
rect 18564 11340 20356 11396
rect 21970 11340 21980 11396
rect 22036 11340 26908 11396
rect 35186 11340 35196 11396
rect 35252 11340 52556 11396
rect 52612 11340 52622 11396
rect 0 11284 112 11312
rect 26852 11284 26908 11340
rect 57344 11284 57456 11312
rect 0 11228 6636 11284
rect 6692 11228 6702 11284
rect 6860 11228 14588 11284
rect 14644 11228 14654 11284
rect 16258 11228 16268 11284
rect 16324 11228 19852 11284
rect 19908 11228 19918 11284
rect 20076 11228 22204 11284
rect 22260 11228 22270 11284
rect 26852 11228 47068 11284
rect 47124 11228 47134 11284
rect 51986 11228 51996 11284
rect 52052 11228 55804 11284
rect 55860 11228 55870 11284
rect 56130 11228 56140 11284
rect 56196 11228 57456 11284
rect 0 11200 112 11228
rect 6860 11172 6916 11228
rect 20076 11172 20132 11228
rect 57344 11200 57456 11228
rect 3042 11116 3052 11172
rect 3108 11116 6916 11172
rect 7074 11116 7084 11172
rect 7140 11116 16716 11172
rect 16772 11116 16782 11172
rect 18162 11116 18172 11172
rect 18228 11116 20132 11172
rect 20972 11116 35084 11172
rect 35140 11116 35150 11172
rect 35634 11116 35644 11172
rect 35700 11116 44940 11172
rect 44996 11116 45006 11172
rect 53554 11116 53564 11172
rect 53620 11116 56364 11172
rect 56420 11116 56430 11172
rect 14690 11004 14700 11060
rect 14756 11004 20748 11060
rect 20804 11004 20814 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 20972 10948 21028 11116
rect 24322 11004 24332 11060
rect 24388 11004 29596 11060
rect 29652 11004 29662 11060
rect 29810 11004 29820 11060
rect 29876 11004 34524 11060
rect 34580 11004 34590 11060
rect 52994 11004 53004 11060
rect 53060 11004 56700 11060
rect 56756 11004 56766 11060
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 7298 10892 7308 10948
rect 7364 10892 14476 10948
rect 14532 10892 14542 10948
rect 14914 10892 14924 10948
rect 14980 10892 21028 10948
rect 24210 10892 24220 10948
rect 24276 10892 30156 10948
rect 30212 10892 30222 10948
rect 31836 10892 40236 10948
rect 40292 10892 40302 10948
rect 0 10836 112 10864
rect 31836 10836 31892 10892
rect 57344 10836 57456 10864
rect 0 10780 17276 10836
rect 17332 10780 17342 10836
rect 18050 10780 18060 10836
rect 18116 10780 18396 10836
rect 18452 10780 18462 10836
rect 18722 10780 18732 10836
rect 18788 10780 31892 10836
rect 32946 10780 32956 10836
rect 33012 10780 34972 10836
rect 35028 10780 35038 10836
rect 38546 10780 38556 10836
rect 38612 10780 54124 10836
rect 54180 10780 54190 10836
rect 55122 10780 55132 10836
rect 55188 10780 57456 10836
rect 0 10752 112 10780
rect 57344 10752 57456 10780
rect 2370 10668 2380 10724
rect 2436 10668 7196 10724
rect 7252 10668 7262 10724
rect 8372 10668 16268 10724
rect 16324 10668 16334 10724
rect 16482 10668 16492 10724
rect 16548 10668 18284 10724
rect 18340 10668 18350 10724
rect 18610 10668 18620 10724
rect 18676 10668 21196 10724
rect 21252 10668 21262 10724
rect 21858 10668 21868 10724
rect 21924 10668 24556 10724
rect 24612 10668 24622 10724
rect 27122 10668 27132 10724
rect 27188 10668 28700 10724
rect 28756 10668 28766 10724
rect 29250 10668 29260 10724
rect 29316 10668 51884 10724
rect 51940 10668 51950 10724
rect 8372 10612 8428 10668
rect 6738 10556 6748 10612
rect 6804 10556 8428 10612
rect 14578 10556 14588 10612
rect 14644 10556 30716 10612
rect 30772 10556 30782 10612
rect 35074 10556 35084 10612
rect 35140 10556 52108 10612
rect 52164 10556 52174 10612
rect 18386 10444 18396 10500
rect 18452 10444 28476 10500
rect 28532 10444 28542 10500
rect 29810 10444 29820 10500
rect 29876 10444 53564 10500
rect 53620 10444 53630 10500
rect 0 10388 112 10416
rect 57344 10388 57456 10416
rect 0 10332 3164 10388
rect 3220 10332 3230 10388
rect 15138 10332 15148 10388
rect 15204 10332 29708 10388
rect 29764 10332 29774 10388
rect 32946 10332 32956 10388
rect 33012 10332 55132 10388
rect 55188 10332 55198 10388
rect 55906 10332 55916 10388
rect 55972 10332 57456 10388
rect 0 10304 112 10332
rect 57344 10304 57456 10332
rect 8530 10220 8540 10276
rect 8596 10220 14924 10276
rect 14980 10220 14990 10276
rect 15922 10220 15932 10276
rect 15988 10220 24220 10276
rect 24276 10220 24286 10276
rect 52210 10220 52220 10276
rect 52276 10220 53116 10276
rect 53172 10220 53182 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 8418 10108 8428 10164
rect 8484 10108 13748 10164
rect 13906 10108 13916 10164
rect 13972 10108 19404 10164
rect 19460 10108 19470 10164
rect 21634 10108 21644 10164
rect 21700 10108 23548 10164
rect 23604 10108 23614 10164
rect 25106 10108 25116 10164
rect 25172 10108 32396 10164
rect 32452 10108 32462 10164
rect 54562 10108 54572 10164
rect 54628 10108 57260 10164
rect 57316 10108 57326 10164
rect 354 9996 364 10052
rect 420 9996 8428 10052
rect 9202 9996 9212 10052
rect 9268 9996 13468 10052
rect 13524 9996 13534 10052
rect 0 9940 112 9968
rect 8372 9940 8428 9996
rect 0 9884 3276 9940
rect 3332 9884 3342 9940
rect 8372 9884 13356 9940
rect 13412 9884 13422 9940
rect 0 9856 112 9884
rect 13692 9828 13748 10108
rect 16706 9996 16716 10052
rect 16772 9996 25564 10052
rect 25620 9996 25630 10052
rect 30258 9996 30268 10052
rect 30324 9996 37996 10052
rect 38052 9996 38062 10052
rect 57344 9940 57456 9968
rect 15092 9884 26796 9940
rect 26852 9884 26862 9940
rect 30034 9884 30044 9940
rect 30100 9884 32620 9940
rect 32676 9884 32686 9940
rect 33058 9884 33068 9940
rect 33124 9884 34636 9940
rect 34692 9884 34702 9940
rect 35298 9884 35308 9940
rect 35364 9884 55356 9940
rect 55412 9884 55422 9940
rect 57250 9884 57260 9940
rect 57316 9884 57456 9940
rect 15092 9828 15148 9884
rect 57344 9856 57456 9884
rect 13692 9772 15148 9828
rect 18060 9772 22428 9828
rect 22484 9772 22494 9828
rect 24210 9772 24220 9828
rect 24276 9772 52556 9828
rect 52612 9772 52622 9828
rect 18060 9716 18116 9772
rect 4162 9660 4172 9716
rect 4228 9660 14252 9716
rect 14308 9660 14318 9716
rect 14466 9660 14476 9716
rect 14532 9660 18116 9716
rect 18274 9660 18284 9716
rect 18340 9660 25116 9716
rect 25172 9660 25182 9716
rect 33170 9660 33180 9716
rect 33236 9660 46172 9716
rect 46228 9660 46238 9716
rect 53554 9660 53564 9716
rect 53620 9660 56476 9716
rect 56532 9660 56542 9716
rect 14802 9548 14812 9604
rect 14868 9548 21140 9604
rect 22194 9548 22204 9604
rect 22260 9548 32844 9604
rect 32900 9548 32910 9604
rect 0 9492 112 9520
rect 0 9436 1596 9492
rect 1652 9436 1662 9492
rect 6626 9436 6636 9492
rect 6692 9436 14924 9492
rect 14980 9436 14990 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 6850 9324 6860 9380
rect 6916 9324 15148 9380
rect 15092 9268 15148 9324
rect 21084 9268 21140 9548
rect 57344 9492 57456 9520
rect 24210 9436 24220 9492
rect 24276 9436 29932 9492
rect 29988 9436 29998 9492
rect 55122 9436 55132 9492
rect 55188 9436 57456 9492
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 57344 9408 57456 9436
rect 4946 9212 4956 9268
rect 5012 9212 13916 9268
rect 13972 9212 13982 9268
rect 15092 9212 16772 9268
rect 21084 9212 30044 9268
rect 30100 9212 30110 9268
rect 30594 9212 30604 9268
rect 30660 9212 48860 9268
rect 48916 9212 48926 9268
rect 16716 9156 16772 9212
rect 2930 9100 2940 9156
rect 2996 9100 6748 9156
rect 6804 9100 6814 9156
rect 13458 9100 13468 9156
rect 13524 9100 15148 9156
rect 16716 9100 25564 9156
rect 25620 9100 25630 9156
rect 29474 9100 29484 9156
rect 29540 9100 33516 9156
rect 33572 9100 33582 9156
rect 43026 9100 43036 9156
rect 43092 9100 55020 9156
rect 55076 9100 55086 9156
rect 0 9044 112 9072
rect 15092 9044 15148 9100
rect 57344 9044 57456 9072
rect 0 8988 6972 9044
rect 7028 8988 7038 9044
rect 15092 8988 18396 9044
rect 18452 8988 18462 9044
rect 20962 8988 20972 9044
rect 21028 8988 22204 9044
rect 22260 8988 22270 9044
rect 23202 8988 23212 9044
rect 23268 8988 45388 9044
rect 45444 8988 45454 9044
rect 56130 8988 56140 9044
rect 56196 8988 57456 9044
rect 0 8960 112 8988
rect 57344 8960 57456 8988
rect 3154 8876 3164 8932
rect 3220 8876 22652 8932
rect 22708 8876 22718 8932
rect 26114 8876 26124 8932
rect 26180 8876 43036 8932
rect 43092 8876 43102 8932
rect 44706 8876 44716 8932
rect 44772 8876 55132 8932
rect 55188 8876 55198 8932
rect 6402 8764 6412 8820
rect 6468 8764 28588 8820
rect 28644 8764 28654 8820
rect 37090 8764 37100 8820
rect 37156 8764 41132 8820
rect 41188 8764 41198 8820
rect 41682 8764 41692 8820
rect 41748 8764 52108 8820
rect 52164 8764 52174 8820
rect 6850 8652 6860 8708
rect 6916 8652 22428 8708
rect 22484 8652 22494 8708
rect 30482 8652 30492 8708
rect 30548 8652 32564 8708
rect 36082 8652 36092 8708
rect 36148 8652 44156 8708
rect 44212 8652 44222 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 0 8540 4172 8596
rect 4228 8540 4238 8596
rect 20738 8540 20748 8596
rect 20804 8540 21140 8596
rect 29698 8540 29708 8596
rect 29764 8540 31612 8596
rect 31668 8540 31678 8596
rect 0 8512 112 8540
rect 21084 8484 21140 8540
rect 32508 8484 32564 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 57344 8596 57456 8624
rect 35298 8540 35308 8596
rect 35364 8540 44324 8596
rect 44268 8484 44324 8540
rect 50372 8540 52444 8596
rect 52500 8540 52510 8596
rect 54338 8540 54348 8596
rect 54404 8540 57456 8596
rect 50372 8484 50428 8540
rect 57344 8512 57456 8540
rect 10098 8428 10108 8484
rect 10164 8428 13300 8484
rect 13244 8372 13300 8428
rect 19516 8428 20860 8484
rect 20916 8428 20926 8484
rect 21084 8428 31836 8484
rect 31892 8428 31902 8484
rect 32508 8428 43484 8484
rect 43540 8428 43550 8484
rect 44268 8428 50428 8484
rect 19516 8372 19572 8428
rect 1586 8316 1596 8372
rect 1652 8316 6748 8372
rect 6804 8316 6814 8372
rect 13244 8316 14700 8372
rect 14756 8316 14766 8372
rect 14914 8316 14924 8372
rect 14980 8316 19572 8372
rect 19954 8316 19964 8372
rect 20020 8316 24220 8372
rect 24276 8316 24286 8372
rect 26898 8316 26908 8372
rect 26964 8316 29260 8372
rect 29316 8316 29326 8372
rect 31378 8316 31388 8372
rect 31444 8316 54124 8372
rect 54180 8316 54190 8372
rect 54898 8316 54908 8372
rect 54964 8316 57036 8372
rect 57092 8316 57102 8372
rect 3266 8204 3276 8260
rect 3332 8204 8428 8260
rect 8484 8204 8494 8260
rect 16034 8204 16044 8260
rect 16100 8204 26796 8260
rect 26852 8204 26862 8260
rect 27916 8204 45164 8260
rect 45220 8204 45230 8260
rect 0 8148 112 8176
rect 0 8092 6636 8148
rect 6692 8092 6702 8148
rect 6962 8092 6972 8148
rect 7028 8092 13916 8148
rect 13972 8092 13982 8148
rect 15092 8092 25900 8148
rect 25956 8092 25966 8148
rect 26114 8092 26124 8148
rect 26180 8092 27692 8148
rect 27748 8092 27758 8148
rect 0 8064 112 8092
rect 15092 7924 15148 8092
rect 27916 8036 27972 8204
rect 57344 8148 57456 8176
rect 29586 8092 29596 8148
rect 29652 8092 33740 8148
rect 33796 8092 33806 8148
rect 40338 8092 40348 8148
rect 40404 8092 44828 8148
rect 44884 8092 44894 8148
rect 55906 8092 55916 8148
rect 55972 8092 57456 8148
rect 57344 8064 57456 8092
rect 17826 7980 17836 8036
rect 17892 7980 27972 8036
rect 28130 7980 28140 8036
rect 28196 7980 31500 8036
rect 31556 7980 31566 8036
rect 38612 7980 48748 8036
rect 48804 7980 48814 8036
rect 38612 7924 38668 7980
rect 4274 7868 4284 7924
rect 4340 7868 15148 7924
rect 26226 7868 26236 7924
rect 26292 7868 38668 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 7410 7756 7420 7812
rect 7476 7756 15036 7812
rect 15092 7756 15102 7812
rect 24332 7756 26124 7812
rect 26180 7756 26190 7812
rect 0 7700 112 7728
rect 0 7644 6748 7700
rect 6804 7644 6814 7700
rect 13346 7644 13356 7700
rect 13412 7644 24108 7700
rect 24164 7644 24174 7700
rect 0 7616 112 7644
rect 24332 7588 24388 7756
rect 57344 7700 57456 7728
rect 24658 7644 24668 7700
rect 24724 7644 27580 7700
rect 27636 7644 27646 7700
rect 35634 7644 35644 7700
rect 35700 7644 53564 7700
rect 53620 7644 53630 7700
rect 56130 7644 56140 7700
rect 56196 7644 57456 7700
rect 57344 7616 57456 7644
rect 3378 7532 3388 7588
rect 3444 7532 14588 7588
rect 14644 7532 14654 7588
rect 22082 7532 22092 7588
rect 22148 7532 24388 7588
rect 25218 7532 25228 7588
rect 25284 7532 26068 7588
rect 37650 7532 37660 7588
rect 37716 7532 43148 7588
rect 43204 7532 43214 7588
rect 43810 7532 43820 7588
rect 43876 7532 48972 7588
rect 49028 7532 49038 7588
rect 26012 7476 26068 7532
rect 7522 7420 7532 7476
rect 7588 7420 16380 7476
rect 16436 7420 16446 7476
rect 22978 7420 22988 7476
rect 23044 7420 25676 7476
rect 25732 7420 25742 7476
rect 26012 7420 53564 7476
rect 53620 7420 53630 7476
rect 5394 7308 5404 7364
rect 5460 7308 14364 7364
rect 14420 7308 14430 7364
rect 14690 7308 14700 7364
rect 14756 7308 21196 7364
rect 21252 7308 21262 7364
rect 21410 7308 21420 7364
rect 21476 7308 55244 7364
rect 55300 7308 55310 7364
rect 0 7252 112 7280
rect 57344 7252 57456 7280
rect 0 7196 1652 7252
rect 9650 7196 9660 7252
rect 9716 7196 17724 7252
rect 17780 7196 17790 7252
rect 20972 7196 46508 7252
rect 46564 7196 46574 7252
rect 47506 7196 47516 7252
rect 47572 7196 48188 7252
rect 48244 7196 48254 7252
rect 54562 7196 54572 7252
rect 54628 7196 57456 7252
rect 0 7168 112 7196
rect 1596 6916 1652 7196
rect 15026 7084 15036 7140
rect 15092 7084 20636 7140
rect 20692 7084 20702 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 20972 7028 21028 7196
rect 57344 7168 57456 7196
rect 21186 7084 21196 7140
rect 21252 7084 24220 7140
rect 24276 7084 24286 7140
rect 26852 7084 31276 7140
rect 31332 7084 31342 7140
rect 34850 7084 34860 7140
rect 34916 7084 43820 7140
rect 43876 7084 43886 7140
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 26852 7028 26908 7084
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 12786 6972 12796 7028
rect 12852 6972 21028 7028
rect 24882 6972 24892 7028
rect 24948 6972 26908 7028
rect 27906 6972 27916 7028
rect 27972 6972 35084 7028
rect 35140 6972 35150 7028
rect 50372 6972 54236 7028
rect 54292 6972 54302 7028
rect 50372 6916 50428 6972
rect 1596 6860 5684 6916
rect 7298 6860 7308 6916
rect 7364 6860 15260 6916
rect 15316 6860 15326 6916
rect 19954 6860 19964 6916
rect 20020 6860 25452 6916
rect 25508 6860 25518 6916
rect 25666 6860 25676 6916
rect 25732 6860 50428 6916
rect 52098 6860 52108 6916
rect 52164 6860 55244 6916
rect 55300 6860 55310 6916
rect 0 6804 112 6832
rect 0 6748 4956 6804
rect 5012 6748 5022 6804
rect 0 6720 112 6748
rect 5628 6692 5684 6860
rect 57344 6804 57456 6832
rect 14578 6748 14588 6804
rect 14644 6748 15932 6804
rect 15988 6748 15998 6804
rect 16146 6748 16156 6804
rect 16212 6748 20076 6804
rect 20132 6748 20142 6804
rect 21522 6748 21532 6804
rect 21588 6748 24220 6804
rect 24276 6748 24286 6804
rect 25228 6748 33572 6804
rect 33730 6748 33740 6804
rect 33796 6748 38668 6804
rect 43362 6748 43372 6804
rect 43428 6748 43540 6804
rect 44146 6748 44156 6804
rect 44212 6748 47348 6804
rect 48850 6748 48860 6804
rect 48916 6748 53676 6804
rect 53732 6748 53742 6804
rect 56130 6748 56140 6804
rect 56196 6748 57456 6804
rect 25228 6692 25284 6748
rect 33516 6692 33572 6748
rect 38612 6692 38668 6748
rect 43484 6692 43540 6748
rect 47292 6692 47348 6748
rect 57344 6720 57456 6748
rect 5628 6636 15148 6692
rect 18498 6636 18508 6692
rect 18564 6636 25284 6692
rect 25442 6636 25452 6692
rect 25508 6636 32060 6692
rect 32116 6636 32126 6692
rect 33516 6636 36988 6692
rect 37044 6636 37054 6692
rect 38612 6636 43260 6692
rect 43316 6636 43326 6692
rect 43484 6636 45444 6692
rect 47292 6636 54236 6692
rect 54292 6636 54302 6692
rect 15092 6580 15148 6636
rect 45388 6580 45444 6636
rect 5058 6524 5068 6580
rect 5124 6524 8540 6580
rect 8596 6524 8606 6580
rect 15092 6524 21756 6580
rect 21812 6524 21822 6580
rect 21970 6524 21980 6580
rect 22036 6524 35308 6580
rect 35364 6524 35374 6580
rect 40674 6524 40684 6580
rect 40740 6524 43708 6580
rect 43764 6524 43774 6580
rect 45388 6524 53452 6580
rect 53508 6524 53518 6580
rect 20066 6412 20076 6468
rect 20132 6412 54124 6468
rect 54180 6412 54190 6468
rect 0 6356 112 6384
rect 57344 6356 57456 6384
rect 0 6300 3668 6356
rect 19842 6300 19852 6356
rect 19908 6300 21980 6356
rect 22036 6300 22046 6356
rect 24210 6300 24220 6356
rect 24276 6300 37100 6356
rect 37156 6300 37166 6356
rect 45042 6300 45052 6356
rect 45108 6300 50204 6356
rect 50260 6300 50270 6356
rect 55122 6300 55132 6356
rect 55188 6300 57456 6356
rect 0 6272 112 6300
rect 3612 6132 3668 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 57344 6272 57456 6300
rect 13682 6188 13692 6244
rect 13748 6188 19964 6244
rect 20020 6188 20030 6244
rect 31826 6188 31836 6244
rect 31892 6188 41692 6244
rect 41748 6188 41758 6244
rect 3612 6076 6860 6132
rect 6916 6076 6926 6132
rect 8372 6076 16716 6132
rect 16772 6076 16782 6132
rect 19282 6076 19292 6132
rect 19348 6076 33628 6132
rect 33684 6076 33694 6132
rect 33842 6076 33852 6132
rect 33908 6076 49420 6132
rect 49476 6076 49486 6132
rect 8372 6020 8428 6076
rect 5954 5964 5964 6020
rect 6020 5964 8428 6020
rect 14242 5964 14252 6020
rect 14308 5964 19964 6020
rect 20020 5964 20030 6020
rect 20626 5964 20636 6020
rect 20692 5964 23548 6020
rect 23604 5964 23614 6020
rect 23762 5964 23772 6020
rect 23828 5964 44828 6020
rect 44884 5964 44894 6020
rect 0 5908 112 5936
rect 57344 5908 57456 5936
rect 0 5852 7084 5908
rect 7140 5852 7150 5908
rect 9986 5852 9996 5908
rect 10052 5852 14140 5908
rect 14196 5852 14206 5908
rect 20962 5852 20972 5908
rect 21028 5852 24892 5908
rect 24948 5852 24958 5908
rect 28466 5852 28476 5908
rect 28532 5852 31836 5908
rect 31892 5852 31902 5908
rect 32050 5852 32060 5908
rect 32116 5852 35196 5908
rect 35252 5852 35262 5908
rect 35746 5852 35756 5908
rect 35812 5852 36204 5908
rect 36260 5852 36270 5908
rect 40674 5852 40684 5908
rect 40740 5852 42084 5908
rect 43474 5852 43484 5908
rect 43540 5852 46620 5908
rect 46676 5852 46686 5908
rect 48738 5852 48748 5908
rect 48804 5852 53564 5908
rect 53620 5852 53630 5908
rect 54562 5852 54572 5908
rect 54628 5852 57456 5908
rect 0 5824 112 5852
rect 42028 5796 42084 5852
rect 57344 5824 57456 5852
rect 1138 5740 1148 5796
rect 1204 5740 7532 5796
rect 7588 5740 7598 5796
rect 13570 5740 13580 5796
rect 13636 5740 18172 5796
rect 18228 5740 18238 5796
rect 22642 5740 22652 5796
rect 22708 5740 24780 5796
rect 24836 5740 24846 5796
rect 25330 5740 25340 5796
rect 25396 5740 41804 5796
rect 41860 5740 41870 5796
rect 42028 5740 49532 5796
rect 49588 5740 49598 5796
rect 49970 5740 49980 5796
rect 50036 5740 52780 5796
rect 52836 5740 52846 5796
rect 2818 5628 2828 5684
rect 2884 5628 24164 5684
rect 24434 5628 24444 5684
rect 24500 5628 25900 5684
rect 25956 5628 25966 5684
rect 26226 5628 26236 5684
rect 26292 5628 41860 5684
rect 7522 5516 7532 5572
rect 7588 5516 16604 5572
rect 16660 5516 16670 5572
rect 18162 5516 18172 5572
rect 18228 5516 21644 5572
rect 21700 5516 21710 5572
rect 22194 5516 22204 5572
rect 22260 5516 23772 5572
rect 23828 5516 23838 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 0 5404 4228 5460
rect 6962 5404 6972 5460
rect 7028 5404 23884 5460
rect 23940 5404 23950 5460
rect 0 5376 112 5404
rect 4172 5348 4228 5404
rect 24108 5348 24164 5628
rect 25218 5516 25228 5572
rect 25284 5516 31724 5572
rect 31780 5516 31790 5572
rect 31938 5516 31948 5572
rect 32004 5516 32732 5572
rect 32788 5516 32798 5572
rect 33730 5516 33740 5572
rect 33796 5516 38668 5572
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 24882 5404 24892 5460
rect 24948 5404 32396 5460
rect 32452 5404 32462 5460
rect 33740 5404 35196 5460
rect 35252 5404 35262 5460
rect 33740 5348 33796 5404
rect 38612 5348 38668 5516
rect 41804 5460 41860 5628
rect 42588 5628 53228 5684
rect 53284 5628 53294 5684
rect 42588 5460 42644 5628
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 57344 5460 57456 5488
rect 41804 5404 42644 5460
rect 47170 5404 47180 5460
rect 47236 5404 50988 5460
rect 51044 5404 51054 5460
rect 56130 5404 56140 5460
rect 56196 5404 57456 5460
rect 57344 5376 57456 5404
rect 4172 5292 6636 5348
rect 6692 5292 6702 5348
rect 6860 5292 9996 5348
rect 10052 5292 10062 5348
rect 10546 5292 10556 5348
rect 10612 5292 14476 5348
rect 14532 5292 14542 5348
rect 16370 5292 16380 5348
rect 16436 5292 18620 5348
rect 18676 5292 18686 5348
rect 21186 5292 21196 5348
rect 21252 5292 23772 5348
rect 23828 5292 23838 5348
rect 24108 5292 29820 5348
rect 29876 5292 29886 5348
rect 30146 5292 30156 5348
rect 30212 5292 33796 5348
rect 33954 5292 33964 5348
rect 34020 5292 37324 5348
rect 37380 5292 37390 5348
rect 38612 5292 40684 5348
rect 40740 5292 40750 5348
rect 40898 5292 40908 5348
rect 40964 5292 46732 5348
rect 46788 5292 46798 5348
rect 52882 5292 52892 5348
rect 52948 5292 56252 5348
rect 56308 5292 56318 5348
rect 6860 5236 6916 5292
rect 2482 5180 2492 5236
rect 2548 5180 6916 5236
rect 7746 5180 7756 5236
rect 7812 5180 20860 5236
rect 20916 5180 20926 5236
rect 21634 5180 21644 5236
rect 21700 5180 25340 5236
rect 25396 5180 25406 5236
rect 29362 5180 29372 5236
rect 29428 5180 31220 5236
rect 32834 5180 32844 5236
rect 32900 5180 47068 5236
rect 47124 5180 47134 5236
rect 31164 5124 31220 5180
rect 2034 5068 2044 5124
rect 2100 5068 7532 5124
rect 7588 5068 7598 5124
rect 11788 5068 14700 5124
rect 14756 5068 14766 5124
rect 14924 5068 18060 5124
rect 18116 5068 18126 5124
rect 20066 5068 20076 5124
rect 20132 5068 20636 5124
rect 20692 5068 20702 5124
rect 23090 5068 23100 5124
rect 23156 5068 26460 5124
rect 26516 5068 26526 5124
rect 26674 5068 26684 5124
rect 26740 5068 30156 5124
rect 30212 5068 30222 5124
rect 31164 5068 33852 5124
rect 33908 5068 33918 5124
rect 35186 5068 35196 5124
rect 35252 5068 37212 5124
rect 37268 5068 37278 5124
rect 37538 5068 37548 5124
rect 37604 5068 39116 5124
rect 39172 5068 39182 5124
rect 41906 5068 41916 5124
rect 41972 5068 43148 5124
rect 43204 5068 43214 5124
rect 43596 5068 45276 5124
rect 45332 5068 45342 5124
rect 45490 5068 45500 5124
rect 45556 5068 47516 5124
rect 47572 5068 47582 5124
rect 54898 5068 54908 5124
rect 54964 5068 55468 5124
rect 0 5012 112 5040
rect 11788 5012 11844 5068
rect 0 4956 8428 5012
rect 10994 4956 11004 5012
rect 11060 4956 11844 5012
rect 0 4928 112 4956
rect 8372 4900 8428 4956
rect 14924 4900 14980 5068
rect 43596 5012 43652 5068
rect 55412 5012 55468 5068
rect 57344 5012 57456 5040
rect 15250 4956 15260 5012
rect 15316 4956 23324 5012
rect 23380 4956 23390 5012
rect 23538 4956 23548 5012
rect 23604 4956 34636 5012
rect 34692 4956 34702 5012
rect 35634 4956 35644 5012
rect 35700 4956 35980 5012
rect 36036 4956 36046 5012
rect 41346 4956 41356 5012
rect 41412 4956 43652 5012
rect 44258 4956 44268 5012
rect 44324 4956 50428 5012
rect 55412 4956 57456 5012
rect 8372 4844 14980 4900
rect 16482 4844 16492 4900
rect 16548 4844 25116 4900
rect 25172 4844 25182 4900
rect 25330 4844 25340 4900
rect 25396 4844 26908 4900
rect 30034 4844 30044 4900
rect 30100 4844 33740 4900
rect 33796 4844 33806 4900
rect 35410 4844 35420 4900
rect 35476 4844 44156 4900
rect 44212 4844 44222 4900
rect 47282 4844 47292 4900
rect 47348 4844 49980 4900
rect 50036 4844 50046 4900
rect 26852 4788 26908 4844
rect 50372 4788 50428 4956
rect 57344 4928 57456 4956
rect 13906 4732 13916 4788
rect 13972 4732 23324 4788
rect 23380 4732 23390 4788
rect 24210 4732 24220 4788
rect 24276 4732 26684 4788
rect 26740 4732 26750 4788
rect 26852 4732 38668 4788
rect 38724 4732 38734 4788
rect 44818 4732 44828 4788
rect 44884 4732 48748 4788
rect 48804 4732 48814 4788
rect 50372 4732 51660 4788
rect 51716 4732 51726 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 6738 4620 6748 4676
rect 6804 4620 15036 4676
rect 15092 4620 15102 4676
rect 24220 4620 25676 4676
rect 25732 4620 25742 4676
rect 31602 4620 31612 4676
rect 31668 4620 35196 4676
rect 35252 4620 35262 4676
rect 35410 4620 35420 4676
rect 35476 4620 41132 4676
rect 41188 4620 41198 4676
rect 45042 4620 45052 4676
rect 45108 4620 54124 4676
rect 54180 4620 54190 4676
rect 0 4564 112 4592
rect 24220 4564 24276 4620
rect 57344 4564 57456 4592
rect 0 4508 9996 4564
rect 10052 4508 10062 4564
rect 11564 4508 18732 4564
rect 18788 4508 18798 4564
rect 22418 4508 22428 4564
rect 22484 4508 24276 4564
rect 24882 4508 24892 4564
rect 24948 4508 26236 4564
rect 26292 4508 26302 4564
rect 31490 4508 31500 4564
rect 31556 4508 35084 4564
rect 35140 4508 35150 4564
rect 35298 4508 35308 4564
rect 35364 4508 41468 4564
rect 41524 4508 41534 4564
rect 44370 4508 44380 4564
rect 44436 4508 50428 4564
rect 50484 4508 50494 4564
rect 54562 4508 54572 4564
rect 54628 4508 57456 4564
rect 0 4480 112 4508
rect 11564 4452 11620 4508
rect 57344 4480 57456 4508
rect 1698 4396 1708 4452
rect 1764 4396 11620 4452
rect 11778 4396 11788 4452
rect 11844 4396 13468 4452
rect 13524 4396 13534 4452
rect 14242 4396 14252 4452
rect 14308 4396 45052 4452
rect 45108 4396 45118 4452
rect 2594 4284 2604 4340
rect 2660 4284 25228 4340
rect 25284 4284 25294 4340
rect 25452 4284 30492 4340
rect 30548 4284 30558 4340
rect 33618 4284 33628 4340
rect 33684 4284 39228 4340
rect 39284 4284 39294 4340
rect 41682 4284 41692 4340
rect 41748 4284 44940 4340
rect 44996 4284 45006 4340
rect 25452 4228 25508 4284
rect 7186 4172 7196 4228
rect 7252 4172 18396 4228
rect 18452 4172 18462 4228
rect 18620 4172 25508 4228
rect 25666 4172 25676 4228
rect 25732 4172 26908 4228
rect 27682 4172 27692 4228
rect 27748 4172 46620 4228
rect 46676 4172 46686 4228
rect 0 4116 112 4144
rect 18620 4116 18676 4172
rect 0 4060 2940 4116
rect 2996 4060 3006 4116
rect 3154 4060 3164 4116
rect 3220 4060 6076 4116
rect 6132 4060 6142 4116
rect 9650 4060 9660 4116
rect 9716 4060 11228 4116
rect 11284 4060 11294 4116
rect 12226 4060 12236 4116
rect 12292 4060 16828 4116
rect 16884 4060 16894 4116
rect 17826 4060 17836 4116
rect 17892 4060 18676 4116
rect 18732 4060 20972 4116
rect 21028 4060 21038 4116
rect 21410 4060 21420 4116
rect 21476 4060 26012 4116
rect 26068 4060 26078 4116
rect 0 4032 112 4060
rect 18732 4004 18788 4060
rect 6178 3948 6188 4004
rect 6244 3948 7420 4004
rect 7476 3948 7486 4004
rect 14242 3948 14252 4004
rect 14308 3948 18788 4004
rect 26852 4004 26908 4172
rect 57344 4116 57456 4144
rect 28802 4060 28812 4116
rect 28868 4060 36092 4116
rect 36148 4060 36158 4116
rect 36726 4060 36764 4116
rect 36820 4060 36830 4116
rect 39106 4060 39116 4116
rect 39172 4060 42028 4116
rect 42084 4060 42094 4116
rect 42242 4060 42252 4116
rect 42308 4060 45500 4116
rect 45556 4060 45566 4116
rect 53218 4060 53228 4116
rect 53284 4060 55804 4116
rect 55860 4060 55870 4116
rect 56130 4060 56140 4116
rect 56196 4060 57456 4116
rect 57344 4032 57456 4060
rect 26852 3948 43372 4004
rect 43428 3948 43438 4004
rect 43586 3948 43596 4004
rect 43652 3948 44268 4004
rect 44324 3948 44334 4004
rect 44818 3948 44828 4004
rect 44884 3948 48412 4004
rect 48468 3948 48478 4004
rect 51314 3948 51324 4004
rect 51380 3948 56700 4004
rect 56756 3948 56766 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 5618 3836 5628 3892
rect 5684 3836 23884 3892
rect 23940 3836 23950 3892
rect 24882 3836 24892 3892
rect 24948 3836 36316 3892
rect 36372 3836 36382 3892
rect 41122 3836 41132 3892
rect 41188 3836 43596 3892
rect 43652 3836 43662 3892
rect 49746 3836 49756 3892
rect 49812 3836 55356 3892
rect 55412 3836 55422 3892
rect 9202 3724 9212 3780
rect 9268 3724 13356 3780
rect 13412 3724 13422 3780
rect 14130 3724 14140 3780
rect 14196 3724 28924 3780
rect 28980 3724 28990 3780
rect 30146 3724 30156 3780
rect 30212 3724 52556 3780
rect 52612 3724 52622 3780
rect 0 3668 112 3696
rect 57344 3668 57456 3696
rect 0 3612 5068 3668
rect 5124 3612 5134 3668
rect 12338 3612 12348 3668
rect 12404 3612 13692 3668
rect 13748 3612 13758 3668
rect 19954 3612 19964 3668
rect 20020 3612 20188 3668
rect 20244 3612 20254 3668
rect 22194 3612 22204 3668
rect 22260 3612 24556 3668
rect 24612 3612 24622 3668
rect 28578 3612 28588 3668
rect 28644 3612 33628 3668
rect 33684 3612 33694 3668
rect 34738 3612 34748 3668
rect 34804 3612 44212 3668
rect 46610 3612 46620 3668
rect 46676 3612 47180 3668
rect 47236 3612 47246 3668
rect 50754 3612 50764 3668
rect 50820 3612 53116 3668
rect 53172 3612 53182 3668
rect 54898 3612 54908 3668
rect 54964 3612 57456 3668
rect 0 3584 112 3612
rect 44156 3556 44212 3612
rect 57344 3584 57456 3612
rect 10434 3500 10444 3556
rect 10500 3500 20188 3556
rect 20244 3500 20254 3556
rect 21746 3500 21756 3556
rect 21812 3500 23548 3556
rect 23604 3500 23614 3556
rect 23772 3500 25228 3556
rect 25284 3500 25294 3556
rect 26226 3500 26236 3556
rect 26292 3500 28812 3556
rect 28868 3500 28878 3556
rect 29036 3500 40348 3556
rect 40404 3500 40414 3556
rect 42802 3500 42812 3556
rect 42868 3500 43932 3556
rect 43988 3500 43998 3556
rect 44156 3500 48300 3556
rect 48356 3500 48366 3556
rect 48850 3500 48860 3556
rect 48916 3500 52668 3556
rect 52724 3500 52734 3556
rect 53554 3500 53564 3556
rect 53620 3500 56812 3556
rect 56868 3500 56878 3556
rect 23772 3444 23828 3500
rect 29036 3444 29092 3500
rect 11666 3388 11676 3444
rect 11732 3388 17836 3444
rect 17892 3388 17902 3444
rect 19842 3388 19852 3444
rect 19908 3388 23828 3444
rect 23986 3388 23996 3444
rect 24052 3388 29092 3444
rect 35196 3388 43372 3444
rect 43428 3388 43438 3444
rect 43586 3388 43596 3444
rect 43652 3388 43764 3444
rect 45714 3388 45724 3444
rect 45780 3388 48076 3444
rect 48132 3388 48142 3444
rect 52210 3388 52220 3444
rect 52276 3388 54460 3444
rect 54516 3388 54526 3444
rect 35196 3332 35252 3388
rect 43708 3332 43764 3388
rect 3612 3276 7644 3332
rect 7700 3276 7710 3332
rect 10322 3276 10332 3332
rect 10388 3276 13580 3332
rect 13636 3276 13646 3332
rect 14130 3276 14140 3332
rect 14196 3276 21532 3332
rect 21588 3276 21598 3332
rect 23660 3276 31948 3332
rect 32834 3276 32844 3332
rect 32900 3276 35252 3332
rect 35746 3276 35756 3332
rect 35812 3276 36764 3332
rect 36820 3276 36830 3332
rect 43708 3276 45724 3332
rect 45780 3276 45790 3332
rect 46722 3276 46732 3332
rect 46788 3276 51212 3332
rect 51268 3276 51278 3332
rect 0 3220 112 3248
rect 3612 3220 3668 3276
rect 23660 3220 23716 3276
rect 31892 3220 31948 3276
rect 57344 3220 57456 3248
rect 0 3164 3668 3220
rect 14354 3164 14364 3220
rect 14420 3164 23716 3220
rect 25330 3164 25340 3220
rect 25396 3164 30940 3220
rect 30996 3164 31006 3220
rect 31892 3164 34860 3220
rect 34916 3164 34926 3220
rect 45602 3164 45612 3220
rect 45668 3164 46508 3220
rect 46564 3164 46574 3220
rect 54562 3164 54572 3220
rect 54628 3164 57456 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 57344 3136 57456 3164
rect 7410 3052 7420 3108
rect 7476 3052 14252 3108
rect 14308 3052 14318 3108
rect 18722 3052 18732 3108
rect 18788 3052 21532 3108
rect 21588 3052 21598 3108
rect 24210 3052 24220 3108
rect 24276 3052 33628 3108
rect 33684 3052 33694 3108
rect 35522 3052 35532 3108
rect 35588 3052 43036 3108
rect 43092 3052 43102 3108
rect 45042 3052 45052 3108
rect 45108 3052 45724 3108
rect 45780 3052 45790 3108
rect 6066 2940 6076 2996
rect 6132 2940 14700 2996
rect 14756 2940 14766 2996
rect 14914 2940 14924 2996
rect 14980 2940 16212 2996
rect 16930 2940 16940 2996
rect 16996 2940 21644 2996
rect 21700 2940 21710 2996
rect 23426 2940 23436 2996
rect 23492 2940 28588 2996
rect 28644 2940 28654 2996
rect 29138 2940 29148 2996
rect 29204 2940 31164 2996
rect 31220 2940 31230 2996
rect 33618 2940 33628 2996
rect 33684 2940 50876 2996
rect 50932 2940 50942 2996
rect 16156 2884 16212 2940
rect 690 2828 700 2884
rect 756 2828 7756 2884
rect 7812 2828 7822 2884
rect 8306 2828 8316 2884
rect 8372 2828 9044 2884
rect 0 2772 112 2800
rect 8988 2772 9044 2828
rect 9548 2828 15932 2884
rect 15988 2828 15998 2884
rect 16156 2828 19852 2884
rect 19908 2828 19918 2884
rect 20178 2828 20188 2884
rect 20244 2828 26012 2884
rect 26068 2828 26078 2884
rect 30930 2828 30940 2884
rect 30996 2828 33964 2884
rect 34020 2828 34030 2884
rect 34188 2828 35924 2884
rect 36978 2828 36988 2884
rect 37044 2828 38108 2884
rect 38164 2828 38174 2884
rect 38332 2828 40740 2884
rect 41458 2828 41468 2884
rect 41524 2828 45276 2884
rect 45332 2828 45342 2884
rect 52994 2828 53004 2884
rect 53060 2828 56924 2884
rect 56980 2828 56990 2884
rect 0 2716 8428 2772
rect 8988 2716 9324 2772
rect 9380 2716 9390 2772
rect 0 2688 112 2716
rect 8372 2660 8428 2716
rect 9548 2660 9604 2828
rect 34188 2772 34244 2828
rect 35868 2772 35924 2828
rect 38332 2772 38388 2828
rect 40684 2772 40740 2828
rect 57344 2772 57456 2800
rect 9762 2716 9772 2772
rect 9828 2716 14924 2772
rect 14980 2716 14990 2772
rect 20178 2716 20188 2772
rect 20244 2716 23996 2772
rect 24052 2716 24062 2772
rect 24210 2716 24220 2772
rect 24276 2716 30492 2772
rect 30548 2716 30558 2772
rect 31378 2716 31388 2772
rect 31444 2716 32732 2772
rect 32788 2716 32798 2772
rect 32946 2716 32956 2772
rect 33012 2716 34244 2772
rect 34850 2716 34860 2772
rect 34916 2716 35644 2772
rect 35700 2716 35710 2772
rect 35868 2716 38388 2772
rect 39106 2716 39116 2772
rect 39172 2716 40460 2772
rect 40516 2716 40526 2772
rect 40684 2716 47292 2772
rect 47348 2716 47358 2772
rect 50418 2716 50428 2772
rect 50484 2716 53564 2772
rect 53620 2716 53630 2772
rect 56130 2716 56140 2772
rect 56196 2716 57456 2772
rect 57344 2688 57456 2716
rect 1596 2604 7308 2660
rect 7364 2604 7374 2660
rect 8372 2604 9604 2660
rect 13906 2604 13916 2660
rect 13972 2604 17556 2660
rect 19170 2604 19180 2660
rect 19236 2604 25228 2660
rect 25284 2604 25294 2660
rect 30940 2604 32396 2660
rect 32452 2604 32462 2660
rect 33058 2604 33068 2660
rect 33124 2604 34076 2660
rect 34132 2604 34142 2660
rect 35074 2604 35084 2660
rect 35140 2604 37100 2660
rect 37156 2604 37166 2660
rect 38322 2604 38332 2660
rect 38388 2604 39900 2660
rect 39956 2604 39966 2660
rect 40338 2604 40348 2660
rect 40404 2604 44940 2660
rect 44996 2604 45006 2660
rect 48626 2604 48636 2660
rect 48692 2604 53676 2660
rect 53732 2604 53742 2660
rect 0 2324 112 2352
rect 1596 2324 1652 2604
rect 1810 2492 1820 2548
rect 1876 2492 17276 2548
rect 17332 2492 17342 2548
rect 17500 2436 17556 2604
rect 30940 2548 30996 2604
rect 20066 2492 20076 2548
rect 20132 2492 28700 2548
rect 28756 2492 28766 2548
rect 29250 2492 29260 2548
rect 29316 2492 30996 2548
rect 31602 2492 31612 2548
rect 31668 2492 32620 2548
rect 32676 2492 32686 2548
rect 36866 2492 36876 2548
rect 36932 2492 49644 2548
rect 49700 2492 49710 2548
rect 6850 2380 6860 2436
rect 6916 2380 15596 2436
rect 15652 2380 15662 2436
rect 17500 2380 19180 2436
rect 19236 2380 19246 2436
rect 21634 2380 21644 2436
rect 21700 2380 24220 2436
rect 24276 2380 24286 2436
rect 26002 2380 26012 2436
rect 26068 2380 43596 2436
rect 43652 2380 43662 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 57344 2324 57456 2352
rect 0 2268 1652 2324
rect 14354 2268 14364 2324
rect 14420 2268 24220 2324
rect 24276 2268 24286 2324
rect 27010 2268 27020 2324
rect 27076 2268 30548 2324
rect 30706 2268 30716 2324
rect 30772 2268 31780 2324
rect 33506 2268 33516 2324
rect 33572 2268 43708 2324
rect 48738 2268 48748 2324
rect 48804 2268 50876 2324
rect 50932 2268 50942 2324
rect 54898 2268 54908 2324
rect 54964 2268 57456 2324
rect 0 2240 112 2268
rect 6738 2156 6748 2212
rect 6804 2156 14140 2212
rect 14196 2156 14206 2212
rect 14466 2156 14476 2212
rect 14532 2156 29596 2212
rect 29652 2156 29662 2212
rect 30492 2100 30548 2268
rect 31724 2100 31780 2268
rect 43652 2212 43708 2268
rect 57344 2240 57456 2268
rect 31892 2156 35308 2212
rect 35364 2156 35374 2212
rect 43652 2156 52108 2212
rect 52164 2156 52174 2212
rect 31892 2100 31948 2156
rect 4834 2044 4844 2100
rect 4900 2044 6972 2100
rect 7028 2044 7038 2100
rect 13458 2044 13468 2100
rect 13524 2044 16044 2100
rect 16100 2044 16110 2100
rect 16818 2044 16828 2100
rect 16884 2044 19068 2100
rect 19124 2044 19134 2100
rect 20132 2044 22764 2100
rect 22820 2044 22830 2100
rect 23986 2044 23996 2100
rect 24052 2044 27916 2100
rect 27972 2044 27982 2100
rect 30492 2044 31668 2100
rect 31724 2044 31948 2100
rect 35186 2044 35196 2100
rect 35252 2044 35756 2100
rect 35812 2044 35822 2100
rect 36540 2044 43372 2100
rect 43428 2044 43438 2100
rect 43586 2044 43596 2100
rect 43652 2044 49476 2100
rect 51426 2044 51436 2100
rect 51492 2044 54124 2100
rect 54180 2044 54190 2100
rect 20132 1988 20188 2044
rect 31612 1988 31668 2044
rect 36540 1988 36596 2044
rect 14130 1932 14140 1988
rect 14196 1932 16492 1988
rect 16548 1932 16558 1988
rect 17154 1932 17164 1988
rect 17220 1932 20188 1988
rect 21298 1932 21308 1988
rect 21364 1932 21868 1988
rect 21924 1932 21934 1988
rect 23538 1932 23548 1988
rect 23604 1932 24892 1988
rect 24948 1932 24958 1988
rect 30146 1932 30156 1988
rect 30212 1932 31388 1988
rect 31444 1932 31454 1988
rect 31612 1932 36596 1988
rect 36754 1932 36764 1988
rect 36820 1932 39228 1988
rect 39284 1932 39294 1988
rect 43026 1932 43036 1988
rect 43092 1932 46956 1988
rect 47012 1932 47022 1988
rect 0 1876 112 1904
rect 0 1820 2380 1876
rect 2436 1820 2446 1876
rect 9986 1820 9996 1876
rect 10052 1820 22764 1876
rect 22820 1820 22830 1876
rect 23202 1820 23212 1876
rect 23268 1820 26684 1876
rect 26740 1820 26750 1876
rect 31154 1820 31164 1876
rect 31220 1820 32956 1876
rect 33012 1820 33022 1876
rect 33842 1820 33852 1876
rect 33908 1820 35756 1876
rect 35812 1820 35822 1876
rect 47058 1820 47068 1876
rect 47124 1820 48916 1876
rect 0 1792 112 1820
rect 18610 1708 18620 1764
rect 18676 1708 20188 1764
rect 20132 1652 20188 1708
rect 23100 1708 26236 1764
rect 26292 1708 26302 1764
rect 26786 1708 26796 1764
rect 26852 1708 31948 1764
rect 32498 1708 32508 1764
rect 32564 1708 34188 1764
rect 34244 1708 34254 1764
rect 35634 1708 35644 1764
rect 35700 1708 37324 1764
rect 37380 1708 37390 1764
rect 38892 1708 42588 1764
rect 42644 1708 42654 1764
rect 43652 1708 43932 1764
rect 43988 1708 43998 1764
rect 45938 1708 45948 1764
rect 46004 1708 47852 1764
rect 47908 1708 47918 1764
rect 7858 1596 7868 1652
rect 7924 1596 8428 1652
rect 11442 1596 11452 1652
rect 11508 1596 14252 1652
rect 14308 1596 14318 1652
rect 14690 1596 14700 1652
rect 14756 1596 16828 1652
rect 16884 1596 16894 1652
rect 18274 1596 18284 1652
rect 18340 1596 19964 1652
rect 20020 1596 20030 1652
rect 20132 1596 20412 1652
rect 20468 1596 20478 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 8372 1540 8428 1596
rect 8372 1484 20076 1540
rect 20132 1484 20142 1540
rect 0 1428 112 1456
rect 23100 1428 23156 1708
rect 25778 1596 25788 1652
rect 25844 1596 26572 1652
rect 26628 1596 26638 1652
rect 26796 1596 30156 1652
rect 30212 1596 30222 1652
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 26796 1540 26852 1596
rect 24220 1484 26852 1540
rect 31892 1540 31948 1708
rect 33618 1596 33628 1652
rect 33684 1596 38668 1652
rect 38724 1596 38734 1652
rect 38892 1540 38948 1708
rect 39666 1596 39676 1652
rect 39732 1596 40572 1652
rect 40628 1596 40638 1652
rect 41458 1596 41468 1652
rect 41524 1596 42364 1652
rect 42420 1596 42430 1652
rect 43652 1540 43708 1708
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 48860 1540 48916 1820
rect 49420 1764 49476 2044
rect 51762 1932 51772 1988
rect 51828 1932 54012 1988
rect 54068 1932 54078 1988
rect 57344 1876 57456 1904
rect 53554 1820 53564 1876
rect 53620 1820 57456 1876
rect 57344 1792 57456 1820
rect 49420 1708 55132 1764
rect 55188 1708 55198 1764
rect 49074 1596 49084 1652
rect 49140 1596 51324 1652
rect 51380 1596 51390 1652
rect 31892 1484 38948 1540
rect 41010 1484 41020 1540
rect 41076 1484 43708 1540
rect 44146 1484 44156 1540
rect 44212 1484 48636 1540
rect 48692 1484 48702 1540
rect 48860 1484 54908 1540
rect 54964 1484 54974 1540
rect 24220 1428 24276 1484
rect 57344 1428 57456 1456
rect 0 1372 15260 1428
rect 15316 1372 15326 1428
rect 15474 1372 15484 1428
rect 15540 1372 23156 1428
rect 23314 1372 23324 1428
rect 23380 1372 24276 1428
rect 25666 1372 25676 1428
rect 25732 1372 33068 1428
rect 33124 1372 33134 1428
rect 33506 1372 33516 1428
rect 33572 1372 46732 1428
rect 46788 1372 46798 1428
rect 53554 1372 53564 1428
rect 53620 1372 57456 1428
rect 0 1344 112 1372
rect 57344 1344 57456 1372
rect 3826 1260 3836 1316
rect 3892 1260 6412 1316
rect 6468 1260 6478 1316
rect 8754 1260 8764 1316
rect 8820 1260 13804 1316
rect 13860 1260 13870 1316
rect 14802 1260 14812 1316
rect 14868 1260 19516 1316
rect 19572 1260 19582 1316
rect 19730 1260 19740 1316
rect 19796 1260 26068 1316
rect 26898 1260 26908 1316
rect 26964 1260 27580 1316
rect 27636 1260 27646 1316
rect 31714 1260 31724 1316
rect 31780 1260 36876 1316
rect 36932 1260 36942 1316
rect 43250 1260 43260 1316
rect 43316 1260 44828 1316
rect 44884 1260 44894 1316
rect 46834 1260 46844 1316
rect 46900 1260 49420 1316
rect 49476 1260 49486 1316
rect 26012 1204 26068 1260
rect 6514 1148 6524 1204
rect 6580 1148 11564 1204
rect 11620 1148 11630 1204
rect 11890 1148 11900 1204
rect 11956 1148 13468 1204
rect 13524 1148 13534 1204
rect 13682 1148 13692 1204
rect 13748 1148 16940 1204
rect 16996 1148 17006 1204
rect 17826 1148 17836 1204
rect 17892 1148 22092 1204
rect 22148 1148 22158 1204
rect 26012 1148 27524 1204
rect 28130 1148 28140 1204
rect 28196 1148 31500 1204
rect 31556 1148 31566 1204
rect 31714 1148 31724 1204
rect 31780 1148 35308 1204
rect 35364 1148 35374 1204
rect 39788 1148 44492 1204
rect 44548 1148 44558 1204
rect 46162 1148 46172 1204
rect 46228 1148 52220 1204
rect 52276 1148 52286 1204
rect 27468 1092 27524 1148
rect 2258 1036 2268 1092
rect 2324 1036 16380 1092
rect 16436 1036 16446 1092
rect 16706 1036 16716 1092
rect 16772 1036 17276 1092
rect 17332 1036 17342 1092
rect 22866 1036 22876 1092
rect 22932 1036 24892 1092
rect 24948 1036 24958 1092
rect 25106 1036 25116 1092
rect 25172 1036 26236 1092
rect 26292 1036 26302 1092
rect 26674 1036 26684 1092
rect 26740 1036 27244 1092
rect 27300 1036 27310 1092
rect 27468 1036 33516 1092
rect 33572 1036 33582 1092
rect 36530 1036 36540 1092
rect 36596 1036 39564 1092
rect 39620 1036 39630 1092
rect 0 980 112 1008
rect 39788 980 39844 1148
rect 40562 1036 40572 1092
rect 40628 1036 43372 1092
rect 43428 1036 43438 1092
rect 43586 1036 43596 1092
rect 43652 1036 53116 1092
rect 53172 1036 53182 1092
rect 57344 980 57456 1008
rect 0 924 4900 980
rect 5170 924 5180 980
rect 5236 924 8596 980
rect 11554 924 11564 980
rect 11620 924 26068 980
rect 29362 924 29372 980
rect 29428 924 30156 980
rect 30212 924 30222 980
rect 33394 924 33404 980
rect 33460 924 35868 980
rect 35924 924 35934 980
rect 37426 924 37436 980
rect 37492 924 37502 980
rect 37772 924 39844 980
rect 40114 924 40124 980
rect 40180 924 41244 980
rect 41300 924 41310 980
rect 41906 924 41916 980
rect 41972 924 45052 980
rect 45108 924 45118 980
rect 51986 924 51996 980
rect 52052 924 57456 980
rect 0 896 112 924
rect 4844 868 4900 924
rect 8540 868 8596 924
rect 4844 812 8428 868
rect 8540 812 9548 868
rect 9604 812 9614 868
rect 10546 812 10556 868
rect 10612 812 12796 868
rect 12852 812 12862 868
rect 15922 812 15932 868
rect 15988 812 21644 868
rect 21700 812 21710 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 8372 756 8428 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 26012 756 26068 924
rect 37436 868 37492 924
rect 29810 812 29820 868
rect 29876 812 32060 868
rect 32116 812 32126 868
rect 34738 812 34748 868
rect 34804 812 37492 868
rect 8372 700 11676 756
rect 11732 700 11742 756
rect 13234 700 13244 756
rect 13300 700 19292 756
rect 19348 700 19358 756
rect 26012 700 30716 756
rect 30772 700 30782 756
rect 37772 644 37828 924
rect 57344 896 57456 924
rect 38770 812 38780 868
rect 38836 812 40460 868
rect 40516 812 40526 868
rect 45490 812 45500 868
rect 45556 812 48748 868
rect 48804 812 48814 868
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 39218 700 39228 756
rect 39284 700 42028 756
rect 42084 700 42094 756
rect 48626 700 48636 756
rect 48692 700 49308 756
rect 49364 700 49374 756
rect 10658 588 10668 644
rect 10724 588 18172 644
rect 18228 588 18238 644
rect 24994 588 25004 644
rect 25060 588 37828 644
rect 44594 588 44604 644
rect 44660 588 45388 644
rect 45444 588 45454 644
rect 0 532 112 560
rect 57344 532 57456 560
rect 0 476 14476 532
rect 14532 476 14542 532
rect 15250 476 15260 532
rect 15316 476 29372 532
rect 29428 476 29438 532
rect 30706 476 30716 532
rect 30772 476 33628 532
rect 33684 476 33694 532
rect 37874 476 37884 532
rect 37940 476 40908 532
rect 40964 476 40974 532
rect 43698 476 43708 532
rect 43764 476 47292 532
rect 47348 476 47358 532
rect 56802 476 56812 532
rect 56868 476 57456 532
rect 0 448 112 476
rect 57344 448 57456 476
rect 10882 364 10892 420
rect 10948 364 18620 420
rect 18676 364 18686 420
rect 21522 364 21532 420
rect 21588 364 31724 420
rect 31780 364 31790 420
rect 31892 364 44268 420
rect 44324 364 44334 420
rect 45042 364 45052 420
rect 45108 364 48860 420
rect 48916 364 48926 420
rect 31892 308 31948 364
rect 19618 252 19628 308
rect 19684 252 31948 308
rect 40226 252 40236 308
rect 40292 252 40302 308
rect 44146 252 44156 308
rect 44212 252 46284 308
rect 46340 252 46350 308
rect 47282 252 47292 308
rect 47348 252 50540 308
rect 50596 252 50606 308
rect 40236 196 40292 252
rect 12786 140 12796 196
rect 12852 140 40292 196
rect 42354 140 42364 196
rect 42420 140 45724 196
rect 45780 140 45790 196
rect 49074 140 49084 196
rect 49140 140 49150 196
rect 50194 140 50204 196
rect 50260 140 50428 196
rect 50484 140 50494 196
rect 0 84 112 112
rect 49084 84 49140 140
rect 57344 84 57456 112
rect 0 28 13916 84
rect 13972 28 13982 84
rect 15698 28 15708 84
rect 15764 28 24892 84
rect 24948 28 24958 84
rect 36754 28 36764 84
rect 36820 28 49140 84
rect 56914 28 56924 84
rect 56980 28 57456 84
rect 0 0 112 28
rect 57344 0 57456 28
<< via3 >>
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 14252 12460 14308 12516
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 16268 11228 16324 11284
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 24220 10892 24276 10948
rect 16268 10668 16324 10724
rect 24220 10220 24276 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 4172 9660 4228 9716
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 33516 9100 33572 9156
rect 43036 9100 43092 9156
rect 43036 8876 43092 8932
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 4172 8540 4228 8596
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 14700 8316 14756 8372
rect 26124 8092 26180 8148
rect 44828 8092 44884 8148
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 26124 7756 26180 7812
rect 25676 7420 25732 7476
rect 14364 7308 14420 7364
rect 14700 7308 14756 7364
rect 21196 7308 21252 7364
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 21196 7084 21252 7140
rect 24220 7084 24276 7140
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 25676 6860 25732 6916
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 19292 6076 19348 6132
rect 23548 5964 23604 6020
rect 9996 5852 10052 5908
rect 40684 5852 40740 5908
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 32396 5404 32452 5460
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 9996 5292 10052 5348
rect 40684 5292 40740 5348
rect 29372 5180 29428 5236
rect 32844 5180 32900 5236
rect 23548 4956 23604 5012
rect 24220 4732 24276 4788
rect 44828 4732 44884 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 15036 4620 15092 4676
rect 35420 4620 35476 4676
rect 35084 4508 35140 4564
rect 28812 4060 28868 4116
rect 36764 4060 36820 4116
rect 43596 3948 43652 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 24892 3836 24948 3892
rect 20188 3612 20244 3668
rect 33628 3612 33684 3668
rect 28812 3500 28868 3556
rect 43372 3388 43428 3444
rect 43596 3388 43652 3444
rect 36764 3276 36820 3332
rect 14364 3164 14420 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 14924 2940 14980 2996
rect 33628 2940 33684 2996
rect 26012 2828 26068 2884
rect 9324 2716 9380 2772
rect 9772 2716 9828 2772
rect 14924 2716 14980 2772
rect 20188 2716 20244 2772
rect 24220 2716 24276 2772
rect 20076 2492 20132 2548
rect 26012 2380 26068 2436
rect 43596 2380 43652 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 24220 2268 24276 2324
rect 13468 2044 13524 2100
rect 22764 1820 22820 1876
rect 23212 1820 23268 1876
rect 14252 1596 14308 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 20076 1484 20132 1540
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 15484 1372 15540 1428
rect 33516 1372 33572 1428
rect 13468 1148 13524 1204
rect 31724 1148 31780 1204
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 19292 700 19348 756
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 29372 476 29428 532
rect 31724 364 31780 420
rect 24892 28 24948 84
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 4436 13356 4756 14224
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 23776 12572 24096 14224
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 4172 9716 4228 9726
rect 4172 8596 4228 9660
rect 4172 8530 4228 8540
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 14252 12516 14308 12526
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 9996 5908 10052 5918
rect 9996 5348 10052 5852
rect 9996 5282 10052 5292
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 9324 2772 9828 2818
rect 9380 2762 9772 2772
rect 9324 2706 9380 2716
rect 9772 2706 9828 2716
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 13468 2100 13524 2110
rect 13468 1204 13524 2044
rect 14252 1652 14308 12460
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 16268 11284 16324 11294
rect 16268 10724 16324 11228
rect 16268 10658 16324 10668
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 24436 13356 24756 14224
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23776 9436 24096 10948
rect 24220 10948 24276 10958
rect 24220 10276 24276 10892
rect 24220 10210 24276 10220
rect 24436 10220 24756 11732
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 14700 8372 14756 8382
rect 14364 7364 14420 7374
rect 14364 3220 14420 7308
rect 14700 7364 14756 8316
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 14700 7298 14756 7308
rect 21196 7364 21252 7374
rect 21196 7140 21252 7308
rect 21196 7074 21252 7084
rect 23776 6300 24096 7812
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 43776 11004 44096 12516
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 43776 9436 44096 10948
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 19292 6132 19348 6142
rect 14364 3154 14420 3164
rect 15036 4676 15092 4686
rect 14924 2996 14980 3006
rect 14924 2772 14980 2940
rect 14924 2706 14980 2716
rect 14252 1586 14308 1596
rect 15036 1558 15092 4620
rect 15036 1502 15540 1558
rect 15484 1428 15540 1502
rect 15484 1362 15540 1372
rect 13468 1138 13524 1148
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 19292 756 19348 6076
rect 23548 6020 23604 6030
rect 23548 5012 23604 5964
rect 23548 4946 23604 4956
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 24220 7140 24276 7150
rect 24220 4788 24276 7084
rect 24220 4722 24276 4732
rect 24436 7084 24756 8596
rect 33516 9156 33572 9166
rect 26124 8148 26180 8158
rect 26124 7812 26180 8092
rect 26124 7746 26180 7756
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 25676 7476 25732 7486
rect 25676 6916 25732 7420
rect 25676 6850 25732 6860
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 20188 3668 20244 3678
rect 20188 2772 20244 3612
rect 20188 2706 20244 2716
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 20076 2548 20132 2558
rect 20076 1540 20132 2492
rect 22764 1876 22820 1886
rect 22764 1738 22820 1820
rect 23212 1876 23268 1886
rect 23212 1738 23268 1820
rect 22764 1682 23268 1738
rect 20076 1474 20132 1484
rect 23776 1596 24096 3108
rect 24436 3948 24756 5460
rect 32396 5460 32452 5470
rect 32396 5338 32452 5404
rect 32396 5282 32900 5338
rect 29372 5236 29428 5246
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 28812 4116 28868 4126
rect 24220 2772 24276 2782
rect 24220 2324 24276 2716
rect 24220 2258 24276 2268
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 19292 690 19348 700
rect 23776 0 24096 1540
rect 24436 812 24756 2324
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 24892 3892 24948 3902
rect 24892 84 24948 3836
rect 28812 3556 28868 4060
rect 28812 3490 28868 3500
rect 26012 2884 26068 2894
rect 26012 2436 26068 2828
rect 26012 2370 26068 2380
rect 29372 532 29428 5180
rect 32844 5236 32900 5282
rect 32844 5170 32900 5180
rect 33516 1428 33572 9100
rect 43036 9156 43092 9166
rect 43036 8932 43092 9100
rect 43036 8866 43092 8876
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 43776 6300 44096 7812
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 40684 5908 40740 5918
rect 40684 5348 40740 5852
rect 40684 5282 40740 5292
rect 43776 4732 44096 6244
rect 35420 4676 35476 4686
rect 35420 4618 35476 4620
rect 35084 4564 35476 4618
rect 35140 4562 35476 4564
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 35084 4498 35140 4508
rect 36764 4116 36820 4126
rect 33628 3668 33684 3678
rect 33628 2996 33684 3612
rect 36764 3332 36820 4060
rect 43596 4004 43652 4014
rect 43596 3898 43652 3948
rect 43372 3842 43652 3898
rect 43372 3444 43428 3842
rect 43372 3378 43428 3388
rect 43596 3444 43652 3454
rect 36764 3266 36820 3276
rect 33628 2930 33684 2940
rect 43596 2436 43652 3388
rect 43596 2370 43652 2380
rect 43776 3164 44096 4676
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 33516 1362 33572 1372
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 29372 466 29428 476
rect 31724 1204 31780 1214
rect 31724 420 31780 1148
rect 31724 354 31780 364
rect 24892 18 24948 28
rect 43776 0 44096 1540
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44436 3948 44756 5460
rect 44828 8148 44884 8158
rect 44828 4788 44884 8092
rect 44828 4722 44884 4732
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 19040 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 29456 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 46480 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 49280 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 2240 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 50736 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 42896 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 32256 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 34944 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 14448 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 30016 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 43456 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 40992 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 25424 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 15456 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 19264 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 20720 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 34944 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 22288 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 29120 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 22512 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 37856 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 25424 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 34496 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 34384 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 30688 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 23296 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 46704 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform -1 0 47712 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 49392 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 11200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform -1 0 15008 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform -1 0 18928 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform -1 0 21392 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 23072 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 27216 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 29456 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 33376 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 49056 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 37856 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 40656 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 51968 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 52416 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 47264 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 49952 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 53424 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 51520 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform 1 0 16464 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform 1 0 17136 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform 1 0 18480 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 20720 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 23744 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform 1 0 9408 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform 1 0 23744 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 25760 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 30576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 29680 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform 1 0 28784 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 27440 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 13664 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 24976 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 28560 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 31136 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 32368 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 35056 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 35056 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 2464 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform 1 0 38528 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform 1 0 34496 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform 1 0 35056 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 37184 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform 1 0 38416 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 39088 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform 1 0 39872 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 41328 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform 1 0 42448 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 43120 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform 1 0 44800 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform 1 0 46368 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform 1 0 44688 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform 1 0 46816 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 26320 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform 1 0 24640 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform 1 0 23296 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform 1 0 21728 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 20272 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 18816 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 18480 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 12432 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 11088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 10864 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 9856 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 6160 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 3360 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform -1 0 45136 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_188
timestamp 1486834041
transform 1 0 21728 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_242
timestamp 1486834041
transform 1 0 27776 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_271
timestamp 1486834041
transform 1 0 31024 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_302
timestamp 1486834041
transform 1 0 34496 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_336
timestamp 1486834041
transform 1 0 38304 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_370
timestamp 1486834041
transform 1 0 42112 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_404
timestamp 1486834041
transform 1 0 45920 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_438
timestamp 1486834041
transform 1 0 49728 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_444
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 54656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 54880 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1486834041
transform 1 0 1344 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_16
timestamp 1486834041
transform 1 0 2464 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_48
timestamp 1486834041
transform 1 0 6048 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_64
timestamp 1486834041
transform 1 0 7840 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1486834041
transform 1 0 8288 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_76
timestamp 1486834041
transform 1 0 9184 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_86
timestamp 1486834041
transform 1 0 10304 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_118
timestamp 1486834041
transform 1 0 13888 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_134
timestamp 1486834041
transform 1 0 15680 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_138
timestamp 1486834041
transform 1 0 16128 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_158
timestamp 1486834041
transform 1 0 18368 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_162
timestamp 1486834041
transform 1 0 18816 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_172
timestamp 1486834041
transform 1 0 19936 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1486834041
transform 1 0 20384 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_178
timestamp 1486834041
transform 1 0 20608 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_187
timestamp 1486834041
transform 1 0 21616 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_216
timestamp 1486834041
transform 1 0 24864 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_267
timestamp 1486834041
transform 1 0 30576 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_271
timestamp 1486834041
transform 1 0 31024 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_346
timestamp 1486834041
transform 1 0 39424 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_416
timestamp 1486834041
transform 1 0 47264 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_458
timestamp 1486834041
transform 1 0 51968 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 55776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 56224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_115
timestamp 1486834041
transform 1 0 13552 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_124
timestamp 1486834041
transform 1 0 14560 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_140
timestamp 1486834041
transform 1 0 16352 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_144
timestamp 1486834041
transform 1 0 16800 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_146
timestamp 1486834041
transform 1 0 17024 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_155
timestamp 1486834041
transform 1 0 18032 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_247
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_373
timestamp 1486834041
transform 1 0 42448 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_443
timestamp 1486834041
transform 1 0 50288 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_174
timestamp 1486834041
transform 1 0 20160 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_190
timestamp 1486834041
transform 1 0 21952 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_198
timestamp 1486834041
transform 1 0 22848 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_220
timestamp 1486834041
transform 1 0 25312 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_224
timestamp 1486834041
transform 1 0 25760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_247
timestamp 1486834041
transform 1 0 28336 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1486834041
transform 1 0 31920 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_296
timestamp 1486834041
transform 1 0 33824 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_300
timestamp 1486834041
transform 1 0 34272 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_315
timestamp 1486834041
transform 1 0 35952 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_345
timestamp 1486834041
transform 1 0 39312 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 39760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 47264 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_440
timestamp 1486834041
transform 1 0 49952 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_444
timestamp 1486834041
transform 1 0 50400 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 56224 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 56448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_10
timestamp 1486834041
transform 1 0 1792 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1486834041
transform 1 0 2240 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_24
timestamp 1486834041
transform 1 0 3360 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_32
timestamp 1486834041
transform 1 0 4256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_77
timestamp 1486834041
transform 1 0 9296 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_81
timestamp 1486834041
transform 1 0 9744 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_91
timestamp 1486834041
transform 1 0 10864 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_95
timestamp 1486834041
transform 1 0 11312 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_139
timestamp 1486834041
transform 1 0 16240 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_147
timestamp 1486834041
transform 1 0 17136 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_151
timestamp 1486834041
transform 1 0 17584 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_153
timestamp 1486834041
transform 1 0 17808 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_162
timestamp 1486834041
transform 1 0 18816 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_170
timestamp 1486834041
transform 1 0 19712 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_174
timestamp 1486834041
transform 1 0 20160 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_193
timestamp 1486834041
transform 1 0 22288 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_201
timestamp 1486834041
transform 1 0 23184 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_205
timestamp 1486834041
transform 1 0 23632 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_214
timestamp 1486834041
transform 1 0 24640 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_230
timestamp 1486834041
transform 1 0 26432 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_238
timestamp 1486834041
transform 1 0 27328 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_242
timestamp 1486834041
transform 1 0 27776 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_244
timestamp 1486834041
transform 1 0 28000 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_279
timestamp 1486834041
transform 1 0 31920 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_291
timestamp 1486834041
transform 1 0 33264 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_325
timestamp 1486834041
transform 1 0 37072 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_341
timestamp 1486834041
transform 1 0 38864 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_351
timestamp 1486834041
transform 1 0 39984 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_359
timestamp 1486834041
transform 1 0 40880 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_371
timestamp 1486834041
transform 1 0 42224 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_379
timestamp 1486834041
transform 1 0 43120 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_383
timestamp 1486834041
transform 1 0 43568 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_387
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_391
timestamp 1486834041
transform 1 0 44464 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_393
timestamp 1486834041
transform 1 0 44688 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_402
timestamp 1486834041
transform 1 0 45696 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_406
timestamp 1486834041
transform 1 0 46144 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_408
timestamp 1486834041
transform 1 0 46368 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_423
timestamp 1486834041
transform 1 0 48048 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_457
timestamp 1486834041
transform 1 0 51856 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_461
timestamp 1486834041
transform 1 0 52304 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 8064 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_80
timestamp 1486834041
transform 1 0 9632 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_84
timestamp 1486834041
transform 1 0 10080 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_93
timestamp 1486834041
transform 1 0 11088 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_125
timestamp 1486834041
transform 1 0 14672 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_133
timestamp 1486834041
transform 1 0 15568 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_137
timestamp 1486834041
transform 1 0 16016 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_139
timestamp 1486834041
transform 1 0 16240 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_158
timestamp 1486834041
transform 1 0 18368 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_175
timestamp 1486834041
transform 1 0 20272 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_207
timestamp 1486834041
transform 1 0 23856 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 24080 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_244
timestamp 1486834041
transform 1 0 28000 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_248
timestamp 1486834041
transform 1 0 28448 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_250
timestamp 1486834041
transform 1 0 28672 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_267
timestamp 1486834041
transform 1 0 30576 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_275
timestamp 1486834041
transform 1 0 31472 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 31920 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_290
timestamp 1486834041
transform 1 0 33152 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_298
timestamp 1486834041
transform 1 0 34048 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_310
timestamp 1486834041
transform 1 0 35392 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_326
timestamp 1486834041
transform 1 0 37184 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_334
timestamp 1486834041
transform 1 0 38080 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_336
timestamp 1486834041
transform 1 0 38304 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_345
timestamp 1486834041
transform 1 0 39312 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_349
timestamp 1486834041
transform 1 0 39760 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_368
timestamp 1486834041
transform 1 0 41888 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_372
timestamp 1486834041
transform 1 0 42336 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_381
timestamp 1486834041
transform 1 0 43344 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_397
timestamp 1486834041
transform 1 0 45136 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_405
timestamp 1486834041
transform 1 0 46032 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_409
timestamp 1486834041
transform 1 0 46480 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_411
timestamp 1486834041
transform 1 0 46704 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_454
timestamp 1486834041
transform 1 0 51520 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_458
timestamp 1486834041
transform 1 0 51968 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 55776 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 56224 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 11984 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1486834041
transform 1 0 13552 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_119
timestamp 1486834041
transform 1 0 14000 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_128
timestamp 1486834041
transform 1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_136
timestamp 1486834041
transform 1 0 15904 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_140
timestamp 1486834041
transform 1 0 16352 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_149
timestamp 1486834041
transform 1 0 17360 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_165
timestamp 1486834041
transform 1 0 19152 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_173
timestamp 1486834041
transform 1 0 20048 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_193
timestamp 1486834041
transform 1 0 22288 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_201
timestamp 1486834041
transform 1 0 23184 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_205
timestamp 1486834041
transform 1 0 23632 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_222
timestamp 1486834041
transform 1 0 25536 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_238
timestamp 1486834041
transform 1 0 27328 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1486834041
transform 1 0 27776 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1486834041
transform 1 0 28000 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_279
timestamp 1486834041
transform 1 0 31920 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_295
timestamp 1486834041
transform 1 0 33712 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_303
timestamp 1486834041
transform 1 0 34608 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_325
timestamp 1486834041
transform 1 0 37072 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_334
timestamp 1486834041
transform 1 0 38080 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_358
timestamp 1486834041
transform 1 0 40768 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_374
timestamp 1486834041
transform 1 0 42560 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_382
timestamp 1486834041
transform 1 0 43456 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 43680 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_403
timestamp 1486834041
transform 1 0 45808 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_407
timestamp 1486834041
transform 1 0 46256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_417
timestamp 1486834041
transform 1 0 47376 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_433
timestamp 1486834041
transform 1 0 49168 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_442
timestamp 1486834041
transform 1 0 50176 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_450
timestamp 1486834041
transform 1 0 51072 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1486834041
transform 1 0 51520 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_457
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_465
timestamp 1486834041
transform 1 0 52752 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_469
timestamp 1486834041
transform 1 0 53200 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 8064 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_104
timestamp 1486834041
transform 1 0 12320 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_120
timestamp 1486834041
transform 1 0 14112 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_128
timestamp 1486834041
transform 1 0 15008 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_228
timestamp 1486834041
transform 1 0 26208 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_237
timestamp 1486834041
transform 1 0 27216 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_269
timestamp 1486834041
transform 1 0 30800 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_277
timestamp 1486834041
transform 1 0 31696 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_279
timestamp 1486834041
transform 1 0 31920 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_368
timestamp 1486834041
transform 1 0 41888 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_376
timestamp 1486834041
transform 1 0 42784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_378
timestamp 1486834041
transform 1 0 43008 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_387
timestamp 1486834041
transform 1 0 44016 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_391
timestamp 1486834041
transform 1 0 44464 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_401
timestamp 1486834041
transform 1 0 45584 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1486834041
transform 1 0 47376 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1486834041
transform 1 0 47600 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_454
timestamp 1486834041
transform 1 0 51520 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_470
timestamp 1486834041
transform 1 0 53312 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_474
timestamp 1486834041
transform 1 0 53760 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 55776 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 56224 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_49
timestamp 1486834041
transform 1 0 6160 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_65
timestamp 1486834041
transform 1 0 7952 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_73
timestamp 1486834041
transform 1 0 8848 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_82
timestamp 1486834041
transform 1 0 9856 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_98
timestamp 1486834041
transform 1 0 11648 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_102
timestamp 1486834041
transform 1 0 12096 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_104
timestamp 1486834041
transform 1 0 12320 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_171
timestamp 1486834041
transform 1 0 19824 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_187
timestamp 1486834041
transform 1 0 21616 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_219
timestamp 1486834041
transform 1 0 25200 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_223
timestamp 1486834041
transform 1 0 25648 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_232
timestamp 1486834041
transform 1 0 26656 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_240
timestamp 1486834041
transform 1 0 27552 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_244
timestamp 1486834041
transform 1 0 28000 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_279
timestamp 1486834041
transform 1 0 31920 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_295
timestamp 1486834041
transform 1 0 33712 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_303
timestamp 1486834041
transform 1 0 34608 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_305
timestamp 1486834041
transform 1 0 34832 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 35840 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_451
timestamp 1486834041
transform 1 0 51184 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_457
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_465
timestamp 1486834041
transform 1 0 52752 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_469
timestamp 1486834041
transform 1 0 53200 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 8064 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 15904 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_150
timestamp 1486834041
transform 1 0 17472 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_159
timestamp 1486834041
transform 1 0 18480 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_191
timestamp 1486834041
transform 1 0 22064 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_201
timestamp 1486834041
transform 1 0 23184 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_244
timestamp 1486834041
transform 1 0 28000 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_252
timestamp 1486834041
transform 1 0 28896 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_262
timestamp 1486834041
transform 1 0 30016 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_266
timestamp 1486834041
transform 1 0 30464 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_275
timestamp 1486834041
transform 1 0 31472 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 31920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_282
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 39424 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_368
timestamp 1486834041
transform 1 0 41888 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_376
timestamp 1486834041
transform 1 0 42784 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_380
timestamp 1486834041
transform 1 0 43232 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_390
timestamp 1486834041
transform 1 0 44352 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_406
timestamp 1486834041
transform 1 0 46144 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_414
timestamp 1486834041
transform 1 0 47040 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_418
timestamp 1486834041
transform 1 0 47488 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_454
timestamp 1486834041
transform 1 0 51520 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_470
timestamp 1486834041
transform 1 0 53312 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_474
timestamp 1486834041
transform 1 0 53760 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 56224 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 56448 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_10
timestamp 1486834041
transform 1 0 1792 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_22
timestamp 1486834041
transform 1 0 3136 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_30
timestamp 1486834041
transform 1 0 4032 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 11984 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 19824 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_193
timestamp 1486834041
transform 1 0 22288 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_203
timestamp 1486834041
transform 1 0 23408 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_219
timestamp 1486834041
transform 1 0 25200 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_229
timestamp 1486834041
transform 1 0 26320 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_255
timestamp 1486834041
transform 1 0 29232 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_287
timestamp 1486834041
transform 1 0 32816 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_303
timestamp 1486834041
transform 1 0 34608 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_349
timestamp 1486834041
transform 1 0 39760 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_357
timestamp 1486834041
transform 1 0 40656 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_359
timestamp 1486834041
transform 1 0 40880 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_368
timestamp 1486834041
transform 1 0 41888 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_384
timestamp 1486834041
transform 1 0 43680 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_395
timestamp 1486834041
transform 1 0 44912 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_427
timestamp 1486834041
transform 1 0 48496 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_443
timestamp 1486834041
transform 1 0 50288 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_451
timestamp 1486834041
transform 1 0 51184 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_457
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_465
timestamp 1486834041
transform 1 0 52752 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_469
timestamp 1486834041
transform 1 0 53200 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 8064 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_136
timestamp 1486834041
transform 1 0 15904 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_158
timestamp 1486834041
transform 1 0 18368 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_174
timestamp 1486834041
transform 1 0 20160 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 23744 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 31584 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_292
timestamp 1486834041
transform 1 0 33376 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_300
timestamp 1486834041
transform 1 0 34272 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_310
timestamp 1486834041
transform 1 0 35392 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_342
timestamp 1486834041
transform 1 0 38976 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1486834041
transform 1 0 47264 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_454
timestamp 1486834041
transform 1 0 51520 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 56224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 56448 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 4480 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1486834041
transform 1 0 11984 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_171
timestamp 1486834041
transform 1 0 19824 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_241
timestamp 1486834041
transform 1 0 27664 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_257
timestamp 1486834041
transform 1 0 29456 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_265
timestamp 1486834041
transform 1 0 30352 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_267
timestamp 1486834041
transform 1 0 30576 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_276
timestamp 1486834041
transform 1 0 31584 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_292
timestamp 1486834041
transform 1 0 33376 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_300
timestamp 1486834041
transform 1 0 34272 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_309
timestamp 1486834041
transform 1 0 35280 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_313
timestamp 1486834041
transform 1 0 35728 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_325
timestamp 1486834041
transform 1 0 37072 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_329
timestamp 1486834041
transform 1 0 37520 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_331
timestamp 1486834041
transform 1 0 37744 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_340
timestamp 1486834041
transform 1 0 38752 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_372
timestamp 1486834041
transform 1 0 42336 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_380
timestamp 1486834041
transform 1 0 43232 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 43680 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_451
timestamp 1486834041
transform 1 0 51184 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1486834041
transform 1 0 8064 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_104
timestamp 1486834041
transform 1 0 12320 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_128
timestamp 1486834041
transform 1 0 15008 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_136
timestamp 1486834041
transform 1 0 15904 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_150
timestamp 1486834041
transform 1 0 17472 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_154
timestamp 1486834041
transform 1 0 17920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_163
timestamp 1486834041
transform 1 0 18928 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_195
timestamp 1486834041
transform 1 0 22512 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_203
timestamp 1486834041
transform 1 0 23408 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_207
timestamp 1486834041
transform 1 0 23856 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_209
timestamp 1486834041
transform 1 0 24080 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_252
timestamp 1486834041
transform 1 0 28896 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_268
timestamp 1486834041
transform 1 0 30688 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_276
timestamp 1486834041
transform 1 0 31584 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_298
timestamp 1486834041
transform 1 0 34048 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_314
timestamp 1486834041
transform 1 0 35840 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_346
timestamp 1486834041
transform 1 0 39424 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_384
timestamp 1486834041
transform 1 0 43680 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_400
timestamp 1486834041
transform 1 0 45472 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_408
timestamp 1486834041
transform 1 0 46368 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_438
timestamp 1486834041
transform 1 0 49728 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_446
timestamp 1486834041
transform 1 0 50624 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 56224 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 56448 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 4480 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_69
timestamp 1486834041
transform 1 0 8400 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_85
timestamp 1486834041
transform 1 0 10192 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_94
timestamp 1486834041
transform 1 0 11200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_102
timestamp 1486834041
transform 1 0 12096 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_104
timestamp 1486834041
transform 1 0 12320 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_107
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_145
timestamp 1486834041
transform 1 0 16912 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_161
timestamp 1486834041
transform 1 0 18704 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_169
timestamp 1486834041
transform 1 0 19600 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_173
timestamp 1486834041
transform 1 0 20048 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_185
timestamp 1486834041
transform 1 0 21392 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_189
timestamp 1486834041
transform 1 0 21840 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_191
timestamp 1486834041
transform 1 0 22064 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_200
timestamp 1486834041
transform 1 0 23072 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_210
timestamp 1486834041
transform 1 0 24192 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_218
timestamp 1486834041
transform 1 0 25088 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_220
timestamp 1486834041
transform 1 0 25312 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_237
timestamp 1486834041
transform 1 0 27216 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_255
timestamp 1486834041
transform 1 0 29232 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_259
timestamp 1486834041
transform 1 0 29680 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_261
timestamp 1486834041
transform 1 0 29904 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_270
timestamp 1486834041
transform 1 0 30912 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_278
timestamp 1486834041
transform 1 0 31808 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_290
timestamp 1486834041
transform 1 0 33152 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_298
timestamp 1486834041
transform 1 0 34048 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 35728 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_317
timestamp 1486834041
transform 1 0 36176 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_321
timestamp 1486834041
transform 1 0 36624 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_323
timestamp 1486834041
transform 1 0 36848 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_332
timestamp 1486834041
transform 1 0 37856 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_348
timestamp 1486834041
transform 1 0 39648 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_357
timestamp 1486834041
transform 1 0 40656 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_373
timestamp 1486834041
transform 1 0 42448 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_381
timestamp 1486834041
transform 1 0 43344 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_397
timestamp 1486834041
transform 1 0 45136 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_405
timestamp 1486834041
transform 1 0 46032 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_409
timestamp 1486834041
transform 1 0 46480 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_419
timestamp 1486834041
transform 1 0 47600 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_443
timestamp 1486834041
transform 1 0 50288 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 51184 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_10
timestamp 1486834041
transform 1 0 1792 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_17
timestamp 1486834041
transform 1 0 2576 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_33
timestamp 1486834041
transform 1 0 4368 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_50
timestamp 1486834041
transform 1 0 6272 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_78
timestamp 1486834041
transform 1 0 9408 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_82
timestamp 1486834041
transform 1 0 9856 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_97
timestamp 1486834041
transform 1 0 11536 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_101
timestamp 1486834041
transform 1 0 11984 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_106
timestamp 1486834041
transform 1 0 12544 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_121
timestamp 1486834041
transform 1 0 14224 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_129
timestamp 1486834041
transform 1 0 15120 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_133
timestamp 1486834041
transform 1 0 15568 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_135
timestamp 1486834041
transform 1 0 15792 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_154
timestamp 1486834041
transform 1 0 17920 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_169
timestamp 1486834041
transform 1 0 19600 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_176
timestamp 1486834041
transform 1 0 20384 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_178
timestamp 1486834041
transform 1 0 20608 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_193
timestamp 1486834041
transform 1 0 22288 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_201
timestamp 1486834041
transform 1 0 23184 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 23408 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_220
timestamp 1486834041
transform 1 0 25312 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_248
timestamp 1486834041
transform 1 0 28448 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_250
timestamp 1486834041
transform 1 0 28672 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_265
timestamp 1486834041
transform 1 0 30352 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1486834041
transform 1 0 30800 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_271
timestamp 1486834041
transform 1 0 31024 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_274
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_289
timestamp 1486834041
transform 1 0 33040 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_305
timestamp 1486834041
transform 1 0 34832 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_316
timestamp 1486834041
transform 1 0 36064 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_320
timestamp 1486834041
transform 1 0 36512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_322
timestamp 1486834041
transform 1 0 36736 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_337
timestamp 1486834041
transform 1 0 38416 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_339
timestamp 1486834041
transform 1 0 38640 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_342
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_346
timestamp 1486834041
transform 1 0 39424 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_361
timestamp 1486834041
transform 1 0 41104 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_369
timestamp 1486834041
transform 1 0 42000 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_373
timestamp 1486834041
transform 1 0 42448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_390
timestamp 1486834041
transform 1 0 44352 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_418
timestamp 1486834041
transform 1 0 47488 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_433
timestamp 1486834041
transform 1 0 49168 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 50064 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_458
timestamp 1486834041
transform 1 0 51968 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_478
timestamp 1486834041
transform 1 0 54208 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_482
timestamp 1486834041
transform 1 0 54656 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_484
timestamp 1486834041
transform 1 0 54880 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 53424 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 53984 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 54992 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 53424 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 53984 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 54992 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 53424 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 54992 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 54992 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 53424 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 52416 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 54992 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 53984 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 53424 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 54992 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 53984 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 54992 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 53424 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 52416 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 51856 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 53984 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 50848 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 52416 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 50848 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 52416 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 52416 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 53984 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 54992 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 53424 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 53984 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 6272 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform -1 0 33040 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform -1 0 35728 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform -1 0 38416 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform -1 0 41104 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 44352 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 46368 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 49168 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 51968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 52416 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 8288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 9968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 14224 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 16912 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform -1 0 19600 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform -1 0 22288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform -1 0 25312 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform -1 0 27328 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform -1 0 30352 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 22624 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 21952 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 24976 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 25872 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 24192 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 26544 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 25872 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 25760 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 29008 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 29456 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 30576 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 29456 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 30352 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 32928 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 31920 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 33824 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 35392 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 35056 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 42112 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 40880 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 41664 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 43232 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 41664 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 42448 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 36960 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 35952 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 36736 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 38528 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 37744 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 40544 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 39312 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 39312 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 44352 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 48160 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 47152 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 46480 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 48720 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 49504 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 43232 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 41664 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 44352 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 44800 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 43232 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 45584 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 44800 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 2576 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 53984 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal2 s 23968 0 24080 112 0 FreeSans 448 0 0 0 Ci
port 0 nsew signal input
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 57344 0 57456 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 57344 4480 57456 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 57344 4928 57456 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 57344 5376 57456 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 57344 5824 57456 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 57344 6272 57456 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 57344 6720 57456 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 57344 7168 57456 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 57344 7616 57456 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 57344 8064 57456 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 57344 8512 57456 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 57344 448 57456 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 57344 8960 57456 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 57344 9408 57456 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 57344 9856 57456 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 57344 10304 57456 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 57344 10752 57456 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 57344 11200 57456 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 57344 11648 57456 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 57344 12096 57456 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 57344 12544 57456 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 57344 12992 57456 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 57344 896 57456 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 57344 13440 57456 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 57344 13888 57456 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 57344 1344 57456 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 57344 1792 57456 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 57344 2240 57456 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 57344 2688 57456 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 57344 3136 57456 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 57344 3584 57456 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 57344 4032 57456 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 48160 0 48272 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 52640 0 52752 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 53088 0 53200 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 53536 0 53648 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 53984 0 54096 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 54432 0 54544 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 54880 0 54992 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 55328 0 55440 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 55776 0 55888 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 56224 0 56336 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 56672 0 56784 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 48608 0 48720 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 49056 0 49168 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 49504 0 49616 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 49952 0 50064 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 50400 0 50512 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 50848 0 50960 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 51296 0 51408 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 51744 0 51856 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 52192 0 52304 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 4480 14112 4592 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 31360 14112 31472 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 34048 14112 34160 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 36736 14112 36848 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 39424 14112 39536 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 42112 14112 42224 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 44800 14112 44912 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 47488 14112 47600 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 50176 14112 50288 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 52864 14112 52976 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 55552 14112 55664 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 7168 14112 7280 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 9856 14112 9968 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 12544 14112 12656 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 15232 14112 15344 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 17920 14112 18032 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 20608 14112 20720 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 23296 14112 23408 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 25984 14112 26096 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 28672 14112 28784 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 N1END[0]
port 105 nsew signal input
flabel metal2 s 1120 0 1232 112 0 FreeSans 448 0 0 0 N1END[1]
port 106 nsew signal input
flabel metal2 s 1568 0 1680 112 0 FreeSans 448 0 0 0 N1END[2]
port 107 nsew signal input
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 N1END[3]
port 108 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 N2END[0]
port 109 nsew signal input
flabel metal2 s 6496 0 6608 112 0 FreeSans 448 0 0 0 N2END[1]
port 110 nsew signal input
flabel metal2 s 6944 0 7056 112 0 FreeSans 448 0 0 0 N2END[2]
port 111 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 N2END[3]
port 112 nsew signal input
flabel metal2 s 7840 0 7952 112 0 FreeSans 448 0 0 0 N2END[4]
port 113 nsew signal input
flabel metal2 s 8288 0 8400 112 0 FreeSans 448 0 0 0 N2END[5]
port 114 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 N2END[6]
port 115 nsew signal input
flabel metal2 s 9184 0 9296 112 0 FreeSans 448 0 0 0 N2END[7]
port 116 nsew signal input
flabel metal2 s 2464 0 2576 112 0 FreeSans 448 0 0 0 N2MID[0]
port 117 nsew signal input
flabel metal2 s 2912 0 3024 112 0 FreeSans 448 0 0 0 N2MID[1]
port 118 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 N2MID[2]
port 119 nsew signal input
flabel metal2 s 3808 0 3920 112 0 FreeSans 448 0 0 0 N2MID[3]
port 120 nsew signal input
flabel metal2 s 4256 0 4368 112 0 FreeSans 448 0 0 0 N2MID[4]
port 121 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 N2MID[5]
port 122 nsew signal input
flabel metal2 s 5152 0 5264 112 0 FreeSans 448 0 0 0 N2MID[6]
port 123 nsew signal input
flabel metal2 s 5600 0 5712 112 0 FreeSans 448 0 0 0 N2MID[7]
port 124 nsew signal input
flabel metal2 s 9632 0 9744 112 0 FreeSans 448 0 0 0 N4END[0]
port 125 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 N4END[10]
port 126 nsew signal input
flabel metal2 s 14560 0 14672 112 0 FreeSans 448 0 0 0 N4END[11]
port 127 nsew signal input
flabel metal2 s 15008 0 15120 112 0 FreeSans 448 0 0 0 N4END[12]
port 128 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 N4END[13]
port 129 nsew signal input
flabel metal2 s 15904 0 16016 112 0 FreeSans 448 0 0 0 N4END[14]
port 130 nsew signal input
flabel metal2 s 16352 0 16464 112 0 FreeSans 448 0 0 0 N4END[15]
port 131 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 N4END[1]
port 132 nsew signal input
flabel metal2 s 10528 0 10640 112 0 FreeSans 448 0 0 0 N4END[2]
port 133 nsew signal input
flabel metal2 s 10976 0 11088 112 0 FreeSans 448 0 0 0 N4END[3]
port 134 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 N4END[4]
port 135 nsew signal input
flabel metal2 s 11872 0 11984 112 0 FreeSans 448 0 0 0 N4END[5]
port 136 nsew signal input
flabel metal2 s 12320 0 12432 112 0 FreeSans 448 0 0 0 N4END[6]
port 137 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 N4END[7]
port 138 nsew signal input
flabel metal2 s 13216 0 13328 112 0 FreeSans 448 0 0 0 N4END[8]
port 139 nsew signal input
flabel metal2 s 13664 0 13776 112 0 FreeSans 448 0 0 0 N4END[9]
port 140 nsew signal input
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 NN4END[0]
port 141 nsew signal input
flabel metal2 s 21280 0 21392 112 0 FreeSans 448 0 0 0 NN4END[10]
port 142 nsew signal input
flabel metal2 s 21728 0 21840 112 0 FreeSans 448 0 0 0 NN4END[11]
port 143 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 NN4END[12]
port 144 nsew signal input
flabel metal2 s 22624 0 22736 112 0 FreeSans 448 0 0 0 NN4END[13]
port 145 nsew signal input
flabel metal2 s 23072 0 23184 112 0 FreeSans 448 0 0 0 NN4END[14]
port 146 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 NN4END[15]
port 147 nsew signal input
flabel metal2 s 17248 0 17360 112 0 FreeSans 448 0 0 0 NN4END[1]
port 148 nsew signal input
flabel metal2 s 17696 0 17808 112 0 FreeSans 448 0 0 0 NN4END[2]
port 149 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 NN4END[3]
port 150 nsew signal input
flabel metal2 s 18592 0 18704 112 0 FreeSans 448 0 0 0 NN4END[4]
port 151 nsew signal input
flabel metal2 s 19040 0 19152 112 0 FreeSans 448 0 0 0 NN4END[5]
port 152 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 NN4END[6]
port 153 nsew signal input
flabel metal2 s 19936 0 20048 112 0 FreeSans 448 0 0 0 NN4END[7]
port 154 nsew signal input
flabel metal2 s 20384 0 20496 112 0 FreeSans 448 0 0 0 NN4END[8]
port 155 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 NN4END[9]
port 156 nsew signal input
flabel metal2 s 24416 0 24528 112 0 FreeSans 448 0 0 0 S1BEG[0]
port 157 nsew signal output
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 S1BEG[1]
port 158 nsew signal output
flabel metal2 s 25312 0 25424 112 0 FreeSans 448 0 0 0 S1BEG[2]
port 159 nsew signal output
flabel metal2 s 25760 0 25872 112 0 FreeSans 448 0 0 0 S1BEG[3]
port 160 nsew signal output
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 S2BEG[0]
port 161 nsew signal output
flabel metal2 s 26656 0 26768 112 0 FreeSans 448 0 0 0 S2BEG[1]
port 162 nsew signal output
flabel metal2 s 27104 0 27216 112 0 FreeSans 448 0 0 0 S2BEG[2]
port 163 nsew signal output
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 S2BEG[3]
port 164 nsew signal output
flabel metal2 s 28000 0 28112 112 0 FreeSans 448 0 0 0 S2BEG[4]
port 165 nsew signal output
flabel metal2 s 28448 0 28560 112 0 FreeSans 448 0 0 0 S2BEG[5]
port 166 nsew signal output
flabel metal2 s 28896 0 29008 112 0 FreeSans 448 0 0 0 S2BEG[6]
port 167 nsew signal output
flabel metal2 s 29344 0 29456 112 0 FreeSans 448 0 0 0 S2BEG[7]
port 168 nsew signal output
flabel metal2 s 29792 0 29904 112 0 FreeSans 448 0 0 0 S2BEGb[0]
port 169 nsew signal output
flabel metal2 s 30240 0 30352 112 0 FreeSans 448 0 0 0 S2BEGb[1]
port 170 nsew signal output
flabel metal2 s 30688 0 30800 112 0 FreeSans 448 0 0 0 S2BEGb[2]
port 171 nsew signal output
flabel metal2 s 31136 0 31248 112 0 FreeSans 448 0 0 0 S2BEGb[3]
port 172 nsew signal output
flabel metal2 s 31584 0 31696 112 0 FreeSans 448 0 0 0 S2BEGb[4]
port 173 nsew signal output
flabel metal2 s 32032 0 32144 112 0 FreeSans 448 0 0 0 S2BEGb[5]
port 174 nsew signal output
flabel metal2 s 32480 0 32592 112 0 FreeSans 448 0 0 0 S2BEGb[6]
port 175 nsew signal output
flabel metal2 s 32928 0 33040 112 0 FreeSans 448 0 0 0 S2BEGb[7]
port 176 nsew signal output
flabel metal2 s 33376 0 33488 112 0 FreeSans 448 0 0 0 S4BEG[0]
port 177 nsew signal output
flabel metal2 s 37856 0 37968 112 0 FreeSans 448 0 0 0 S4BEG[10]
port 178 nsew signal output
flabel metal2 s 38304 0 38416 112 0 FreeSans 448 0 0 0 S4BEG[11]
port 179 nsew signal output
flabel metal2 s 38752 0 38864 112 0 FreeSans 448 0 0 0 S4BEG[12]
port 180 nsew signal output
flabel metal2 s 39200 0 39312 112 0 FreeSans 448 0 0 0 S4BEG[13]
port 181 nsew signal output
flabel metal2 s 39648 0 39760 112 0 FreeSans 448 0 0 0 S4BEG[14]
port 182 nsew signal output
flabel metal2 s 40096 0 40208 112 0 FreeSans 448 0 0 0 S4BEG[15]
port 183 nsew signal output
flabel metal2 s 33824 0 33936 112 0 FreeSans 448 0 0 0 S4BEG[1]
port 184 nsew signal output
flabel metal2 s 34272 0 34384 112 0 FreeSans 448 0 0 0 S4BEG[2]
port 185 nsew signal output
flabel metal2 s 34720 0 34832 112 0 FreeSans 448 0 0 0 S4BEG[3]
port 186 nsew signal output
flabel metal2 s 35168 0 35280 112 0 FreeSans 448 0 0 0 S4BEG[4]
port 187 nsew signal output
flabel metal2 s 35616 0 35728 112 0 FreeSans 448 0 0 0 S4BEG[5]
port 188 nsew signal output
flabel metal2 s 36064 0 36176 112 0 FreeSans 448 0 0 0 S4BEG[6]
port 189 nsew signal output
flabel metal2 s 36512 0 36624 112 0 FreeSans 448 0 0 0 S4BEG[7]
port 190 nsew signal output
flabel metal2 s 36960 0 37072 112 0 FreeSans 448 0 0 0 S4BEG[8]
port 191 nsew signal output
flabel metal2 s 37408 0 37520 112 0 FreeSans 448 0 0 0 S4BEG[9]
port 192 nsew signal output
flabel metal2 s 40544 0 40656 112 0 FreeSans 448 0 0 0 SS4BEG[0]
port 193 nsew signal output
flabel metal2 s 45024 0 45136 112 0 FreeSans 448 0 0 0 SS4BEG[10]
port 194 nsew signal output
flabel metal2 s 45472 0 45584 112 0 FreeSans 448 0 0 0 SS4BEG[11]
port 195 nsew signal output
flabel metal2 s 45920 0 46032 112 0 FreeSans 448 0 0 0 SS4BEG[12]
port 196 nsew signal output
flabel metal2 s 46368 0 46480 112 0 FreeSans 448 0 0 0 SS4BEG[13]
port 197 nsew signal output
flabel metal2 s 46816 0 46928 112 0 FreeSans 448 0 0 0 SS4BEG[14]
port 198 nsew signal output
flabel metal2 s 47264 0 47376 112 0 FreeSans 448 0 0 0 SS4BEG[15]
port 199 nsew signal output
flabel metal2 s 40992 0 41104 112 0 FreeSans 448 0 0 0 SS4BEG[1]
port 200 nsew signal output
flabel metal2 s 41440 0 41552 112 0 FreeSans 448 0 0 0 SS4BEG[2]
port 201 nsew signal output
flabel metal2 s 41888 0 42000 112 0 FreeSans 448 0 0 0 SS4BEG[3]
port 202 nsew signal output
flabel metal2 s 42336 0 42448 112 0 FreeSans 448 0 0 0 SS4BEG[4]
port 203 nsew signal output
flabel metal2 s 42784 0 42896 112 0 FreeSans 448 0 0 0 SS4BEG[5]
port 204 nsew signal output
flabel metal2 s 43232 0 43344 112 0 FreeSans 448 0 0 0 SS4BEG[6]
port 205 nsew signal output
flabel metal2 s 43680 0 43792 112 0 FreeSans 448 0 0 0 SS4BEG[7]
port 206 nsew signal output
flabel metal2 s 44128 0 44240 112 0 FreeSans 448 0 0 0 SS4BEG[8]
port 207 nsew signal output
flabel metal2 s 44576 0 44688 112 0 FreeSans 448 0 0 0 SS4BEG[9]
port 208 nsew signal output
flabel metal2 s 47712 0 47824 112 0 FreeSans 448 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 1792 14112 1904 14224 0 FreeSans 448 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
rlabel metal1 28728 12544 28728 12544 0 VDD
rlabel metal1 28728 13328 28728 13328 0 VSS
rlabel metal2 13944 1344 13944 1344 0 FrameData[0]
rlabel metal2 10024 4872 10024 4872 0 FrameData[10]
rlabel metal3 4242 4984 4242 4984 0 FrameData[11]
rlabel metal3 2142 5432 2142 5432 0 FrameData[12]
rlabel metal3 3598 5880 3598 5880 0 FrameData[13]
rlabel metal3 1862 6328 1862 6328 0 FrameData[14]
rlabel metal3 2534 6776 2534 6776 0 FrameData[15]
rlabel metal3 854 7224 854 7224 0 FrameData[16]
rlabel metal3 3430 7672 3430 7672 0 FrameData[17]
rlabel metal3 3374 8120 3374 8120 0 FrameData[18]
rlabel metal3 22120 2744 22120 2744 0 FrameData[19]
rlabel metal2 29624 2352 29624 2352 0 FrameData[1]
rlabel metal3 3542 9016 3542 9016 0 FrameData[20]
rlabel metal3 4200 8344 4200 8344 0 FrameData[21]
rlabel metal3 1694 9912 1694 9912 0 FrameData[22]
rlabel metal3 1638 10360 1638 10360 0 FrameData[23]
rlabel metal2 17304 11200 17304 11200 0 FrameData[24]
rlabel metal3 3374 11256 3374 11256 0 FrameData[25]
rlabel metal3 966 11704 966 11704 0 FrameData[26]
rlabel metal3 238 12152 238 12152 0 FrameData[27]
rlabel metal3 854 12600 854 12600 0 FrameData[28]
rlabel metal3 2142 13048 2142 13048 0 FrameData[29]
rlabel metal3 2478 952 2478 952 0 FrameData[2]
rlabel metal2 23576 12824 23576 12824 0 FrameData[30]
rlabel metal3 3710 13944 3710 13944 0 FrameData[31]
rlabel metal2 15288 952 15288 952 0 FrameData[3]
rlabel metal3 1246 1848 1246 1848 0 FrameData[4]
rlabel metal3 854 2296 854 2296 0 FrameData[5]
rlabel metal3 4242 2744 4242 2744 0 FrameData[6]
rlabel metal3 1862 3192 1862 3192 0 FrameData[7]
rlabel metal3 2590 3640 2590 3640 0 FrameData[8]
rlabel metal3 1526 4088 1526 4088 0 FrameData[9]
rlabel metal3 57162 56 57162 56 0 FrameData_O[0]
rlabel metal3 55986 4536 55986 4536 0 FrameData_O[10]
rlabel metal3 55188 5096 55188 5096 0 FrameData_O[11]
rlabel metal2 56168 4984 56168 4984 0 FrameData_O[12]
rlabel metal2 54600 5936 54600 5936 0 FrameData_O[13]
rlabel metal2 55160 6384 55160 6384 0 FrameData_O[14]
rlabel metal2 56168 6440 56168 6440 0 FrameData_O[15]
rlabel metal2 54600 7392 54600 7392 0 FrameData_O[16]
rlabel metal3 56770 7672 56770 7672 0 FrameData_O[17]
rlabel metal3 56658 8120 56658 8120 0 FrameData_O[18]
rlabel metal2 54376 8736 54376 8736 0 FrameData_O[19]
rlabel metal2 53592 3472 53592 3472 0 FrameData_O[1]
rlabel metal3 56770 9016 56770 9016 0 FrameData_O[20]
rlabel metal2 55160 9520 55160 9520 0 FrameData_O[21]
rlabel metal2 54600 10416 54600 10416 0 FrameData_O[22]
rlabel metal3 56658 10360 56658 10360 0 FrameData_O[23]
rlabel metal2 55160 10976 55160 10976 0 FrameData_O[24]
rlabel metal3 56770 11256 56770 11256 0 FrameData_O[25]
rlabel metal3 54908 12040 54908 12040 0 FrameData_O[26]
rlabel metal3 56882 12152 56882 12152 0 FrameData_O[27]
rlabel metal2 53032 10920 53032 10920 0 FrameData_O[28]
rlabel metal3 56000 8344 56000 8344 0 FrameData_O[29]
rlabel metal2 52024 1120 52024 1120 0 FrameData_O[2]
rlabel metal3 56938 13496 56938 13496 0 FrameData_O[30]
rlabel metal3 56602 13944 56602 13944 0 FrameData_O[31]
rlabel metal3 55482 1400 55482 1400 0 FrameData_O[3]
rlabel metal3 55482 1848 55482 1848 0 FrameData_O[4]
rlabel metal2 54936 2184 54936 2184 0 FrameData_O[5]
rlabel metal2 56168 2072 56168 2072 0 FrameData_O[6]
rlabel metal2 54600 3080 54600 3080 0 FrameData_O[7]
rlabel metal3 56154 3640 56154 3640 0 FrameData_O[8]
rlabel metal2 56168 3528 56168 3528 0 FrameData_O[9]
rlabel metal3 47880 7224 47880 7224 0 FrameStrobe[0]
rlabel metal2 52696 1806 52696 1806 0 FrameStrobe[10]
rlabel metal2 53144 574 53144 574 0 FrameStrobe[11]
rlabel metal2 53592 350 53592 350 0 FrameStrobe[12]
rlabel metal2 54040 1022 54040 1022 0 FrameStrobe[13]
rlabel metal2 54488 1750 54488 1750 0 FrameStrobe[14]
rlabel metal2 54936 798 54936 798 0 FrameStrobe[15]
rlabel metal2 55384 1974 55384 1974 0 FrameStrobe[16]
rlabel metal2 55832 2086 55832 2086 0 FrameStrobe[17]
rlabel metal2 56280 2702 56280 2702 0 FrameStrobe[18]
rlabel metal2 51352 3864 51352 3864 0 FrameStrobe[19]
rlabel metal2 48664 406 48664 406 0 FrameStrobe[1]
rlabel metal2 49112 126 49112 126 0 FrameStrobe[2]
rlabel metal2 14840 10472 14840 10472 0 FrameStrobe[3]
rlabel metal2 18760 11088 18760 11088 0 FrameStrobe[4]
rlabel metal2 50456 126 50456 126 0 FrameStrobe[5]
rlabel metal2 50904 1190 50904 1190 0 FrameStrobe[6]
rlabel metal2 51352 854 51352 854 0 FrameStrobe[7]
rlabel metal2 51800 910 51800 910 0 FrameStrobe[8]
rlabel metal2 52248 630 52248 630 0 FrameStrobe[9]
rlabel metal2 4536 14098 4536 14098 0 FrameStrobe_O[0]
rlabel metal2 31416 13482 31416 13482 0 FrameStrobe_O[10]
rlabel metal2 34552 12712 34552 12712 0 FrameStrobe_O[11]
rlabel metal2 36792 13482 36792 13482 0 FrameStrobe_O[12]
rlabel metal2 39480 13482 39480 13482 0 FrameStrobe_O[13]
rlabel metal2 42168 13594 42168 13594 0 FrameStrobe_O[14]
rlabel metal2 44856 14042 44856 14042 0 FrameStrobe_O[15]
rlabel metal2 47544 13482 47544 13482 0 FrameStrobe_O[16]
rlabel metal2 50792 13440 50792 13440 0 FrameStrobe_O[17]
rlabel metal2 52920 13650 52920 13650 0 FrameStrobe_O[18]
rlabel metal2 55608 13258 55608 13258 0 FrameStrobe_O[19]
rlabel metal2 7224 13482 7224 13482 0 FrameStrobe_O[1]
rlabel metal2 9912 13874 9912 13874 0 FrameStrobe_O[2]
rlabel metal2 12600 13482 12600 13482 0 FrameStrobe_O[3]
rlabel metal2 15512 12376 15512 12376 0 FrameStrobe_O[4]
rlabel metal2 17976 13762 17976 13762 0 FrameStrobe_O[5]
rlabel metal2 20664 13482 20664 13482 0 FrameStrobe_O[6]
rlabel metal2 23352 13762 23352 13762 0 FrameStrobe_O[7]
rlabel metal2 26040 13482 26040 13482 0 FrameStrobe_O[8]
rlabel metal2 28728 13482 28728 13482 0 FrameStrobe_O[9]
rlabel metal2 728 1470 728 1470 0 N1END[0]
rlabel metal2 1176 2926 1176 2926 0 N1END[1]
rlabel metal2 1624 686 1624 686 0 N1END[2]
rlabel metal2 2072 2590 2072 2590 0 N1END[3]
rlabel metal2 6104 1414 6104 1414 0 N2END[0]
rlabel metal2 6552 630 6552 630 0 N2END[1]
rlabel metal2 7000 966 7000 966 0 N2END[2]
rlabel metal2 7448 1582 7448 1582 0 N2END[3]
rlabel metal2 7896 854 7896 854 0 N2END[4]
rlabel metal2 8344 1470 8344 1470 0 N2END[5]
rlabel metal2 8792 686 8792 686 0 N2END[6]
rlabel metal2 9240 1918 9240 1918 0 N2END[7]
rlabel metal2 2520 2646 2520 2646 0 N2MID[0]
rlabel metal2 2968 1470 2968 1470 0 N2MID[1]
rlabel metal2 3416 3822 3416 3822 0 N2MID[2]
rlabel metal2 3864 686 3864 686 0 N2MID[3]
rlabel metal2 4312 3990 4312 3990 0 N2MID[4]
rlabel metal2 4760 350 4760 350 0 N2MID[5]
rlabel metal2 5208 518 5208 518 0 N2MID[6]
rlabel metal2 5656 1974 5656 1974 0 N2MID[7]
rlabel metal2 9688 2086 9688 2086 0 N4END[0]
rlabel metal3 28168 3192 28168 3192 0 N4END[10]
rlabel metal2 14616 3430 14616 3430 0 N4END[11]
rlabel metal2 15064 3598 15064 3598 0 N4END[12]
rlabel metal2 36344 3976 36344 3976 0 N4END[13]
rlabel metal2 21672 1624 21672 1624 0 N4END[14]
rlabel metal2 2296 1512 2296 1512 0 N4END[15]
rlabel metal2 10136 1582 10136 1582 0 N4END[1]
rlabel metal2 10584 462 10584 462 0 N4END[2]
rlabel metal2 11032 2534 11032 2534 0 N4END[3]
rlabel metal2 11480 854 11480 854 0 N4END[4]
rlabel metal2 11928 630 11928 630 0 N4END[5]
rlabel metal2 12376 1862 12376 1862 0 N4END[6]
rlabel metal2 12824 126 12824 126 0 N4END[7]
rlabel metal2 13272 406 13272 406 0 N4END[8]
rlabel metal2 13720 630 13720 630 0 N4END[9]
rlabel metal2 6104 3528 6104 3528 0 NN4END[0]
rlabel metal2 21336 1022 21336 1022 0 NN4END[10]
rlabel metal3 22680 3528 22680 3528 0 NN4END[11]
rlabel metal3 23408 3640 23408 3640 0 NN4END[12]
rlabel metal3 23744 5768 23744 5768 0 NN4END[13]
rlabel metal3 24808 5096 24808 5096 0 NN4END[14]
rlabel metal2 23576 1022 23576 1022 0 NN4END[15]
rlabel metal2 5992 6608 5992 6608 0 NN4END[1]
rlabel metal3 13720 7224 13720 7224 0 NN4END[2]
rlabel metal2 18200 350 18200 350 0 NN4END[3]
rlabel metal2 18648 238 18648 238 0 NN4END[4]
rlabel metal2 19096 1078 19096 1078 0 NN4END[5]
rlabel metal2 19544 686 19544 686 0 NN4END[6]
rlabel metal2 19992 854 19992 854 0 NN4END[7]
rlabel metal2 20440 854 20440 854 0 NN4END[8]
rlabel metal2 20888 1022 20888 1022 0 NN4END[9]
rlabel metal2 24472 350 24472 350 0 S1BEG[0]
rlabel metal2 24920 574 24920 574 0 S1BEG[1]
rlabel metal2 25368 1302 25368 1302 0 S1BEG[2]
rlabel metal2 25816 854 25816 854 0 S1BEG[3]
rlabel metal2 26264 574 26264 574 0 S2BEG[0]
rlabel metal2 26712 574 26712 574 0 S2BEG[1]
rlabel metal2 27160 910 27160 910 0 S2BEG[2]
rlabel metal2 27608 686 27608 686 0 S2BEG[3]
rlabel metal2 28056 966 28056 966 0 S2BEG[4]
rlabel metal2 28504 574 28504 574 0 S2BEG[5]
rlabel metal2 28952 462 28952 462 0 S2BEG[6]
rlabel metal2 29400 518 29400 518 0 S2BEG[7]
rlabel metal2 29848 462 29848 462 0 S2BEGb[0]
rlabel metal2 30296 686 30296 686 0 S2BEGb[1]
rlabel metal2 30744 294 30744 294 0 S2BEGb[2]
rlabel metal2 31192 966 31192 966 0 S2BEGb[3]
rlabel metal2 31640 1302 31640 1302 0 S2BEGb[4]
rlabel metal2 32088 350 32088 350 0 S2BEGb[5]
rlabel metal2 32536 910 32536 910 0 S2BEGb[6]
rlabel metal2 32984 854 32984 854 0 S2BEGb[7]
rlabel metal2 33432 518 33432 518 0 S4BEG[0]
rlabel metal2 37912 294 37912 294 0 S4BEG[10]
rlabel metal2 38360 1358 38360 1358 0 S4BEG[11]
rlabel metal2 38808 462 38808 462 0 S4BEG[12]
rlabel metal2 39256 406 39256 406 0 S4BEG[13]
rlabel metal2 39704 854 39704 854 0 S4BEG[14]
rlabel metal2 40152 518 40152 518 0 S4BEG[15]
rlabel metal2 33880 966 33880 966 0 S4BEG[1]
rlabel metal2 34328 854 34328 854 0 S4BEG[2]
rlabel metal2 34776 462 34776 462 0 S4BEG[3]
rlabel metal2 35224 686 35224 686 0 S4BEG[4]
rlabel metal2 35672 910 35672 910 0 S4BEG[5]
rlabel metal2 36120 910 36120 910 0 S4BEG[6]
rlabel metal2 36568 574 36568 574 0 S4BEG[7]
rlabel metal2 37016 1470 37016 1470 0 S4BEG[8]
rlabel metal2 37464 406 37464 406 0 S4BEG[9]
rlabel metal2 40600 574 40600 574 0 SS4BEG[0]
rlabel metal2 45080 238 45080 238 0 SS4BEG[10]
rlabel metal2 45528 462 45528 462 0 SS4BEG[11]
rlabel metal2 45976 910 45976 910 0 SS4BEG[12]
rlabel metal2 46424 686 46424 686 0 SS4BEG[13]
rlabel metal2 46872 686 46872 686 0 SS4BEG[14]
rlabel metal2 47320 182 47320 182 0 SS4BEG[15]
rlabel metal3 43820 1736 43820 1736 0 SS4BEG[1]
rlabel metal2 41496 854 41496 854 0 SS4BEG[2]
rlabel metal2 41944 518 41944 518 0 SS4BEG[3]
rlabel metal2 45752 1008 45752 1008 0 SS4BEG[4]
rlabel metal3 43400 3528 43400 3528 0 SS4BEG[5]
rlabel metal2 44856 2072 44856 2072 0 SS4BEG[6]
rlabel metal2 43736 294 43736 294 0 SS4BEG[7]
rlabel metal2 44184 182 44184 182 0 SS4BEG[8]
rlabel metal2 44632 350 44632 350 0 SS4BEG[9]
rlabel metal3 46368 11928 46368 11928 0 UserCLK
rlabel metal2 2072 13384 2072 13384 0 UserCLKo
rlabel metal3 26040 1232 26040 1232 0 net1
rlabel metal2 55272 8176 55272 8176 0 net10
rlabel metal3 23352 4536 23352 4536 0 net100
rlabel metal2 44296 1568 44296 1568 0 net101
rlabel metal2 46760 1288 46760 1288 0 net102
rlabel metal3 45416 3080 45416 3080 0 net103
rlabel metal2 14280 5096 14280 5096 0 net104
rlabel metal3 4816 10696 4816 10696 0 net105
rlabel metal2 53592 8288 53592 8288 0 net11
rlabel metal2 52584 3696 52584 3696 0 net12
rlabel metal2 55160 10416 55160 10416 0 net13
rlabel metal2 54264 8400 54264 8400 0 net14
rlabel metal2 29848 9408 29848 9408 0 net15
rlabel metal2 55160 11928 55160 11928 0 net16
rlabel metal2 54152 11088 54152 11088 0 net17
rlabel metal2 55048 11032 55048 11032 0 net18
rlabel metal3 41328 12152 41328 12152 0 net19
rlabel metal2 53704 5544 53704 5544 0 net2
rlabel metal2 35224 10640 35224 10640 0 net20
rlabel metal3 43624 10584 43624 10584 0 net21
rlabel metal2 31416 9408 31416 9408 0 net22
rlabel metal2 51016 3304 51016 3304 0 net23
rlabel metal2 24248 10920 24248 10920 0 net24
rlabel metal2 51016 11760 51016 11760 0 net25
rlabel metal2 52808 3472 52808 3472 0 net26
rlabel metal2 52528 2072 52528 2072 0 net27
rlabel metal3 52808 2072 52808 2072 0 net28
rlabel metal3 49448 1904 49448 1904 0 net29
rlabel metal2 54264 5880 54264 5880 0 net3
rlabel metal2 50456 3640 50456 3640 0 net30
rlabel metal2 54152 4144 54152 4144 0 net31
rlabel metal2 55104 2744 55104 2744 0 net32
rlabel metal2 6104 12880 6104 12880 0 net33
rlabel metal3 44184 3584 44184 3584 0 net34
rlabel metal3 36344 12040 36344 12040 0 net35
rlabel metal2 38248 12600 38248 12600 0 net36
rlabel metal3 49000 3304 49000 3304 0 net37
rlabel metal2 51688 4200 51688 4200 0 net38
rlabel metal3 46088 3192 46088 3192 0 net39
rlabel metal3 53704 6888 53704 6888 0 net4
rlabel metal2 49224 8288 49224 8288 0 net40
rlabel metal3 52248 12936 52248 12936 0 net41
rlabel metal2 52472 12936 52472 12936 0 net42
rlabel metal3 51968 3640 51968 3640 0 net43
rlabel metal2 8120 13552 8120 13552 0 net44
rlabel metal2 10416 12264 10416 12264 0 net45
rlabel metal2 14280 12208 14280 12208 0 net46
rlabel metal2 18200 11760 18200 11760 0 net47
rlabel metal3 20048 12264 20048 12264 0 net48
rlabel metal2 22344 12600 22344 12600 0 net49
rlabel metal2 26264 9968 26264 9968 0 net5
rlabel metal3 25816 12264 25816 12264 0 net50
rlabel metal3 27944 10696 27944 10696 0 net51
rlabel metal3 31360 9912 31360 9912 0 net52
rlabel metal3 21476 2072 21476 2072 0 net53
rlabel metal2 17864 1904 17864 1904 0 net54
rlabel metal2 25256 2688 25256 2688 0 net55
rlabel metal3 23744 4088 23744 4088 0 net56
rlabel metal2 24360 2800 24360 2800 0 net57
rlabel metal4 22792 1779 22792 1779 0 net58
rlabel metal2 25984 2072 25984 2072 0 net59
rlabel metal2 54152 6552 54152 6552 0 net6
rlabel metal2 26264 7560 26264 7560 0 net60
rlabel metal2 28896 9128 28896 9128 0 net61
rlabel metal2 29176 2072 29176 2072 0 net62
rlabel metal2 30408 3528 30408 3528 0 net63
rlabel metal2 29568 1176 29568 1176 0 net64
rlabel metal3 29848 1176 29848 1176 0 net65
rlabel metal4 24248 2520 24248 2520 0 net66
rlabel metal2 25704 1624 25704 1624 0 net67
rlabel metal3 30968 2576 30968 2576 0 net68
rlabel metal2 31864 2352 31864 2352 0 net69
rlabel metal2 55384 7896 55384 7896 0 net7
rlabel metal2 33432 3864 33432 3864 0 net70
rlabel metal2 35784 2352 35784 2352 0 net71
rlabel metal3 35280 2744 35280 2744 0 net72
rlabel metal2 1736 3248 1736 3248 0 net73
rlabel metal3 42560 5096 42560 5096 0 net74
rlabel metal3 42224 6552 42224 6552 0 net75
rlabel metal2 41496 2464 41496 2464 0 net76
rlabel metal3 45024 1960 45024 1960 0 net77
rlabel metal2 45304 5824 45304 5824 0 net78
rlabel metal3 43904 4088 43904 4088 0 net79
rlabel metal3 26040 7504 26040 7504 0 net8
rlabel metal3 38024 1960 38024 1960 0 net80
rlabel metal2 36792 4256 36792 4256 0 net81
rlabel metal2 37184 1176 37184 1176 0 net82
rlabel metal2 36288 2744 36288 2744 0 net83
rlabel metal2 38080 1960 38080 1960 0 net84
rlabel metal2 37576 4368 37576 4368 0 net85
rlabel metal2 40096 1176 40096 1176 0 net86
rlabel metal3 39816 2744 39816 2744 0 net87
rlabel metal2 42056 4144 42056 4144 0 net88
rlabel metal2 44184 1344 44184 1344 0 net89
rlabel metal2 55160 8176 55160 8176 0 net9
rlabel metal3 12656 4424 12656 4424 0 net90
rlabel metal3 23128 2856 23128 2856 0 net91
rlabel metal2 10248 4200 10248 4200 0 net92
rlabel metal3 11368 10024 11368 10024 0 net93
rlabel metal3 23688 3248 23688 3248 0 net94
rlabel metal2 49672 2296 49672 2296 0 net95
rlabel metal3 31640 2016 31640 2016 0 net96
rlabel metal2 41832 4704 41832 4704 0 net97
rlabel metal3 37800 784 37800 784 0 net98
rlabel metal2 44968 2352 44968 2352 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 14224
<< end >>
