magic
tech gf180mcuD
magscale 1 10
timestamp 1764972375
<< metal1 >>
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 2158 13186 2210 13198
rect 2158 13122 2210 13134
rect 3726 13186 3778 13198
rect 3726 13122 3778 13134
rect 5966 13186 6018 13198
rect 5966 13122 6018 13134
rect 7534 13186 7586 13198
rect 7534 13122 7586 13134
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 17390 13186 17442 13198
rect 17390 13122 17442 13134
rect 18958 13186 19010 13198
rect 18958 13122 19010 13134
rect 22654 13186 22706 13198
rect 22654 13122 22706 13134
rect 25454 13186 25506 13198
rect 25454 13122 25506 13134
rect 41918 13186 41970 13198
rect 41918 13122 41970 13134
rect 42142 13186 42194 13198
rect 42142 13122 42194 13134
rect 48974 13186 49026 13198
rect 48974 13122 49026 13134
rect 51102 13186 51154 13198
rect 51102 13122 51154 13134
rect 54910 13186 54962 13198
rect 54910 13122 54962 13134
rect 11890 13022 11902 13074
rect 11954 13022 11966 13074
rect 13346 13022 13358 13074
rect 13410 13022 13422 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 23874 13022 23886 13074
rect 23938 13022 23950 13074
rect 48402 13022 48414 13074
rect 48466 13022 48478 13074
rect 52882 13022 52894 13074
rect 52946 13022 52958 13074
rect 31726 12962 31778 12974
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 6290 12910 6302 12962
rect 6354 12910 6366 12962
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 10210 12910 10222 12962
rect 10274 12910 10286 12962
rect 14130 12910 14142 12962
rect 14194 12910 14206 12962
rect 15698 12910 15710 12962
rect 15762 12910 15774 12962
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 19506 12910 19518 12962
rect 19570 12910 19582 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 44930 12910 44942 12962
rect 44994 12910 45006 12962
rect 46834 12910 46846 12962
rect 46898 12910 46910 12962
rect 50754 12910 50766 12962
rect 50818 12910 50830 12962
rect 52322 12910 52334 12962
rect 52386 12910 52398 12962
rect 54562 12910 54574 12962
rect 54626 12910 54638 12962
rect 31726 12898 31778 12910
rect 21534 12850 21586 12862
rect 21534 12786 21586 12798
rect 26014 12850 26066 12862
rect 26014 12786 26066 12798
rect 31390 12850 31442 12862
rect 31390 12786 31442 12798
rect 32286 12850 32338 12862
rect 32286 12786 32338 12798
rect 47854 12850 47906 12862
rect 47854 12786 47906 12798
rect 50094 12850 50146 12862
rect 50094 12786 50146 12798
rect 24446 12738 24498 12750
rect 24446 12674 24498 12686
rect 45950 12738 46002 12750
rect 45950 12674 46002 12686
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 2270 12402 2322 12414
rect 2270 12338 2322 12350
rect 6974 12402 7026 12414
rect 6974 12338 7026 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 12014 12402 12066 12414
rect 12014 12338 12066 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 16382 12402 16434 12414
rect 16382 12338 16434 12350
rect 17950 12402 18002 12414
rect 17950 12338 18002 12350
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 49086 12402 49138 12414
rect 49086 12338 49138 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 54126 12402 54178 12414
rect 54126 12338 54178 12350
rect 55694 12402 55746 12414
rect 55694 12338 55746 12350
rect 13806 12290 13858 12302
rect 20862 12290 20914 12302
rect 31054 12290 31106 12302
rect 3602 12238 3614 12290
rect 3666 12238 3678 12290
rect 5058 12238 5070 12290
rect 5122 12238 5134 12290
rect 8194 12238 8206 12290
rect 8258 12238 8270 12290
rect 19394 12238 19406 12290
rect 19458 12238 19470 12290
rect 22194 12238 22206 12290
rect 22258 12238 22270 12290
rect 13806 12226 13858 12238
rect 20862 12226 20914 12238
rect 31054 12226 31106 12238
rect 36878 12290 36930 12302
rect 41358 12290 41410 12302
rect 37874 12238 37886 12290
rect 37938 12238 37950 12290
rect 36878 12226 36930 12238
rect 41358 12226 41410 12238
rect 42254 12290 42306 12302
rect 46834 12238 46846 12290
rect 46898 12238 46910 12290
rect 42254 12226 42306 12238
rect 20638 12178 20690 12190
rect 2818 12126 2830 12178
rect 2882 12126 2894 12178
rect 4162 12126 4174 12178
rect 4226 12126 4238 12178
rect 8866 12126 8878 12178
rect 8930 12126 8942 12178
rect 10994 12126 11006 12178
rect 11058 12126 11070 12178
rect 15362 12126 15374 12178
rect 15426 12126 15438 12178
rect 16930 12126 16942 12178
rect 16994 12126 17006 12178
rect 18274 12126 18286 12178
rect 18338 12126 18350 12178
rect 20638 12114 20690 12126
rect 21422 12178 21474 12190
rect 32286 12178 32338 12190
rect 22978 12126 22990 12178
rect 23042 12126 23054 12178
rect 26226 12126 26238 12178
rect 26290 12126 26302 12178
rect 31826 12126 31838 12178
rect 31890 12126 31902 12178
rect 21422 12114 21474 12126
rect 32286 12114 32338 12126
rect 36318 12178 36370 12190
rect 41794 12126 41806 12178
rect 41858 12126 41870 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 49970 12126 49982 12178
rect 50034 12126 50046 12178
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 55346 12126 55358 12178
rect 55410 12126 55422 12178
rect 36318 12114 36370 12126
rect 25902 12066 25954 12078
rect 31390 12066 31442 12078
rect 7522 12014 7534 12066
rect 7586 12014 7598 12066
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 20066 12014 20078 12066
rect 20130 12014 20142 12066
rect 24546 12014 24558 12066
rect 24610 12014 24622 12066
rect 27010 12014 27022 12066
rect 27074 12014 27086 12066
rect 25902 12002 25954 12014
rect 31390 12002 31442 12014
rect 32846 12066 32898 12078
rect 44270 12066 44322 12078
rect 38210 12014 38222 12066
rect 38274 12014 38286 12066
rect 32846 12002 32898 12014
rect 44270 12002 44322 12014
rect 44494 12066 44546 12078
rect 44494 12002 44546 12014
rect 45054 12066 45106 12078
rect 45054 12002 45106 12014
rect 45950 12066 46002 12078
rect 50990 12066 51042 12078
rect 48514 12014 48526 12066
rect 48578 12014 48590 12066
rect 53554 12014 53566 12066
rect 53618 12014 53630 12066
rect 45950 12002 46002 12014
rect 50990 12002 51042 12014
rect 5518 11954 5570 11966
rect 5518 11890 5570 11902
rect 5742 11954 5794 11966
rect 5742 11890 5794 11902
rect 13022 11954 13074 11966
rect 13022 11890 13074 11902
rect 13246 11954 13298 11966
rect 13246 11890 13298 11902
rect 25118 11954 25170 11966
rect 25118 11890 25170 11902
rect 25342 11954 25394 11966
rect 25342 11890 25394 11902
rect 37326 11954 37378 11966
rect 37326 11890 37378 11902
rect 39454 11954 39506 11966
rect 39454 11890 39506 11902
rect 45390 11954 45442 11966
rect 45390 11890 45442 11902
rect 46398 11954 46450 11966
rect 46398 11890 46450 11902
rect 50430 11954 50482 11966
rect 50430 11890 50482 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 4622 11618 4674 11630
rect 4622 11554 4674 11566
rect 6190 11618 6242 11630
rect 6190 11554 6242 11566
rect 7758 11618 7810 11630
rect 7758 11554 7810 11566
rect 8878 11618 8930 11630
rect 8878 11554 8930 11566
rect 9214 11618 9266 11630
rect 9214 11554 9266 11566
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 14030 11618 14082 11630
rect 14030 11554 14082 11566
rect 17502 11618 17554 11630
rect 17502 11554 17554 11566
rect 19070 11618 19122 11630
rect 19070 11554 19122 11566
rect 38222 11618 38274 11630
rect 38222 11554 38274 11566
rect 38446 11618 38498 11630
rect 38446 11554 38498 11566
rect 42366 11618 42418 11630
rect 42366 11554 42418 11566
rect 42590 11618 42642 11630
rect 42590 11554 42642 11566
rect 50318 11618 50370 11630
rect 50318 11554 50370 11566
rect 51886 11618 51938 11630
rect 51886 11554 51938 11566
rect 53454 11618 53506 11630
rect 53454 11554 53506 11566
rect 25678 11506 25730 11518
rect 46062 11506 46114 11518
rect 13010 11454 13022 11506
rect 13074 11454 13086 11506
rect 20402 11454 20414 11506
rect 20466 11454 20478 11506
rect 21186 11454 21198 11506
rect 21250 11454 21262 11506
rect 21970 11454 21982 11506
rect 22034 11454 22046 11506
rect 26002 11454 26014 11506
rect 26066 11454 26078 11506
rect 34738 11454 34750 11506
rect 34802 11454 34814 11506
rect 42018 11454 42030 11506
rect 42082 11454 42094 11506
rect 48962 11454 48974 11506
rect 49026 11454 49038 11506
rect 25678 11442 25730 11454
rect 46062 11442 46114 11454
rect 1486 11394 1538 11406
rect 23438 11394 23490 11406
rect 3602 11342 3614 11394
rect 3666 11342 3678 11394
rect 5170 11342 5182 11394
rect 5234 11342 5246 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 8082 11342 8094 11394
rect 8146 11342 8158 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 14578 11342 14590 11394
rect 14642 11342 14654 11394
rect 16146 11342 16158 11394
rect 16210 11342 16222 11394
rect 18050 11342 18062 11394
rect 18114 11342 18126 11394
rect 19618 11342 19630 11394
rect 19682 11342 19694 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 1486 11330 1538 11342
rect 23438 11330 23490 11342
rect 24558 11394 24610 11406
rect 27582 11394 27634 11406
rect 26114 11342 26126 11394
rect 26178 11342 26190 11394
rect 24558 11330 24610 11342
rect 27582 11330 27634 11342
rect 41246 11394 41298 11406
rect 46958 11394 47010 11406
rect 54462 11394 54514 11406
rect 55246 11394 55298 11406
rect 41682 11342 41694 11394
rect 41746 11342 41758 11394
rect 46498 11342 46510 11394
rect 46562 11342 46574 11394
rect 48178 11342 48190 11394
rect 48242 11342 48254 11394
rect 49746 11342 49758 11394
rect 49810 11342 49822 11394
rect 51314 11342 51326 11394
rect 51378 11342 51390 11394
rect 52882 11342 52894 11394
rect 52946 11342 52958 11394
rect 54898 11342 54910 11394
rect 54962 11342 54974 11394
rect 41246 11330 41298 11342
rect 46958 11330 47010 11342
rect 54462 11330 54514 11342
rect 55246 11330 55298 11342
rect 1262 11282 1314 11294
rect 2606 11282 2658 11294
rect 1922 11230 1934 11282
rect 1986 11230 1998 11282
rect 1262 11218 1314 11230
rect 2606 11218 2658 11230
rect 8878 11282 8930 11294
rect 8878 11218 8930 11230
rect 9774 11282 9826 11294
rect 23102 11282 23154 11294
rect 12338 11230 12350 11282
rect 12402 11230 12414 11282
rect 15474 11230 15486 11282
rect 15538 11230 15550 11282
rect 9774 11218 9826 11230
rect 23102 11218 23154 11230
rect 23998 11282 24050 11294
rect 23998 11218 24050 11230
rect 25118 11282 25170 11294
rect 25118 11218 25170 11230
rect 28142 11282 28194 11294
rect 28142 11218 28194 11230
rect 28366 11282 28418 11294
rect 28366 11218 28418 11230
rect 32286 11282 32338 11294
rect 32286 11218 32338 11230
rect 33854 11282 33906 11294
rect 39006 11282 39058 11294
rect 34402 11230 34414 11282
rect 34466 11230 34478 11282
rect 33854 11218 33906 11230
rect 39006 11218 39058 11230
rect 45054 11282 45106 11294
rect 45054 11218 45106 11230
rect 45726 11282 45778 11294
rect 45726 11218 45778 11230
rect 47518 11282 47570 11294
rect 47518 11218 47570 11230
rect 26574 11170 26626 11182
rect 26574 11106 26626 11118
rect 35982 11170 36034 11182
rect 35982 11106 36034 11118
rect 40910 11170 40962 11182
rect 40910 11106 40962 11118
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 3390 10834 3442 10846
rect 3390 10770 3442 10782
rect 6414 10834 6466 10846
rect 6414 10770 6466 10782
rect 7982 10834 8034 10846
rect 7982 10770 8034 10782
rect 14814 10834 14866 10846
rect 14814 10770 14866 10782
rect 41582 10834 41634 10846
rect 41582 10770 41634 10782
rect 49646 10834 49698 10846
rect 49646 10770 49698 10782
rect 50878 10834 50930 10846
rect 50878 10770 50930 10782
rect 52558 10834 52610 10846
rect 52558 10770 52610 10782
rect 18286 10722 18338 10734
rect 2146 10670 2158 10722
rect 2210 10670 2222 10722
rect 13794 10670 13806 10722
rect 13858 10670 13870 10722
rect 16482 10670 16494 10722
rect 16546 10670 16558 10722
rect 18286 10658 18338 10670
rect 19182 10722 19234 10734
rect 19182 10658 19234 10670
rect 19518 10722 19570 10734
rect 19518 10658 19570 10670
rect 20526 10722 20578 10734
rect 25678 10722 25730 10734
rect 21858 10670 21870 10722
rect 21922 10670 21934 10722
rect 20526 10658 20578 10670
rect 25678 10658 25730 10670
rect 42702 10722 42754 10734
rect 42702 10658 42754 10670
rect 46510 10722 46562 10734
rect 46510 10658 46562 10670
rect 54574 10722 54626 10734
rect 54574 10658 54626 10670
rect 56142 10722 56194 10734
rect 56142 10658 56194 10670
rect 34974 10610 35026 10622
rect 47742 10610 47794 10622
rect 8978 10558 8990 10610
rect 9042 10558 9054 10610
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 11666 10558 11678 10610
rect 11730 10558 11742 10610
rect 17490 10558 17502 10610
rect 17554 10558 17566 10610
rect 26226 10558 26238 10610
rect 26290 10558 26302 10610
rect 29922 10558 29934 10610
rect 29986 10558 29998 10610
rect 34514 10558 34526 10610
rect 34578 10558 34590 10610
rect 42354 10558 42366 10610
rect 42418 10558 42430 10610
rect 48738 10558 48750 10610
rect 48802 10558 48814 10610
rect 52098 10558 52110 10610
rect 52162 10558 52174 10610
rect 34974 10546 35026 10558
rect 47742 10546 47794 10558
rect 12126 10498 12178 10510
rect 40798 10498 40850 10510
rect 2818 10446 2830 10498
rect 2882 10446 2894 10498
rect 4386 10446 4398 10498
rect 4450 10446 4462 10498
rect 7410 10446 7422 10498
rect 7474 10446 7486 10498
rect 9874 10446 9886 10498
rect 9938 10446 9950 10498
rect 14242 10446 14254 10498
rect 14306 10446 14318 10498
rect 15810 10446 15822 10498
rect 15874 10446 15886 10498
rect 17714 10446 17726 10498
rect 17778 10446 17790 10498
rect 21074 10446 21086 10498
rect 21138 10446 21150 10498
rect 26562 10446 26574 10498
rect 26626 10446 26638 10498
rect 30370 10446 30382 10498
rect 30434 10446 30446 10498
rect 12126 10434 12178 10446
rect 40798 10434 40850 10446
rect 41246 10498 41298 10510
rect 43038 10498 43090 10510
rect 48302 10498 48354 10510
rect 42130 10446 42142 10498
rect 42194 10446 42206 10498
rect 47394 10446 47406 10498
rect 47458 10446 47470 10498
rect 51426 10446 51438 10498
rect 51490 10446 51502 10498
rect 53554 10446 53566 10498
rect 53618 10446 53630 10498
rect 55122 10446 55134 10498
rect 55186 10446 55198 10498
rect 41246 10434 41298 10446
rect 43038 10434 43090 10446
rect 48302 10434 48354 10446
rect 11118 10386 11170 10398
rect 11118 10322 11170 10334
rect 12686 10386 12738 10398
rect 12686 10322 12738 10334
rect 13134 10386 13186 10398
rect 13134 10322 13186 10334
rect 13358 10386 13410 10398
rect 13358 10322 13410 10334
rect 18622 10386 18674 10398
rect 18622 10322 18674 10334
rect 18958 10386 19010 10398
rect 18958 10322 19010 10334
rect 20078 10386 20130 10398
rect 20078 10322 20130 10334
rect 24222 10386 24274 10398
rect 24222 10322 24274 10334
rect 27806 10386 27858 10398
rect 27806 10322 27858 10334
rect 29598 10386 29650 10398
rect 29598 10322 29650 10334
rect 31614 10386 31666 10398
rect 31614 10322 31666 10334
rect 34078 10386 34130 10398
rect 34078 10322 34130 10334
rect 34414 10386 34466 10398
rect 34414 10322 34466 10334
rect 40462 10386 40514 10398
rect 40462 10322 40514 10334
rect 40686 10386 40738 10398
rect 40686 10322 40738 10334
rect 46622 10386 46674 10398
rect 46622 10322 46674 10334
rect 47070 10386 47122 10398
rect 47070 10322 47122 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 17950 10050 18002 10062
rect 17950 9986 18002 9998
rect 19406 10050 19458 10062
rect 19406 9986 19458 9998
rect 26014 10050 26066 10062
rect 26014 9986 26066 9998
rect 29710 10050 29762 10062
rect 29710 9986 29762 9998
rect 30046 10050 30098 10062
rect 30046 9986 30098 9998
rect 42142 10050 42194 10062
rect 42142 9986 42194 9998
rect 47518 10050 47570 10062
rect 47518 9986 47570 9998
rect 18846 9938 18898 9950
rect 5282 9886 5294 9938
rect 5346 9886 5358 9938
rect 9650 9886 9662 9938
rect 9714 9886 9726 9938
rect 18846 9874 18898 9886
rect 21534 9938 21586 9950
rect 21534 9874 21586 9886
rect 22094 9938 22146 9950
rect 22094 9874 22146 9886
rect 23998 9938 24050 9950
rect 23998 9874 24050 9886
rect 24446 9938 24498 9950
rect 42590 9938 42642 9950
rect 27570 9886 27582 9938
rect 27634 9886 27646 9938
rect 24446 9874 24498 9886
rect 42590 9874 42642 9886
rect 46958 9938 47010 9950
rect 46958 9874 47010 9886
rect 48190 9938 48242 9950
rect 48190 9874 48242 9886
rect 48526 9938 48578 9950
rect 48526 9874 48578 9886
rect 49086 9938 49138 9950
rect 50194 9886 50206 9938
rect 50258 9886 50270 9938
rect 49086 9874 49138 9886
rect 17390 9826 17442 9838
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 7522 9774 7534 9826
rect 7586 9774 7598 9826
rect 10434 9774 10446 9826
rect 10498 9774 10510 9826
rect 12002 9774 12014 9826
rect 12066 9774 12078 9826
rect 13010 9774 13022 9826
rect 13074 9774 13086 9826
rect 15026 9774 15038 9826
rect 15090 9774 15102 9826
rect 17390 9762 17442 9774
rect 18286 9826 18338 9838
rect 18286 9762 18338 9774
rect 20302 9826 20354 9838
rect 20302 9762 20354 9774
rect 21086 9826 21138 9838
rect 46398 9826 46450 9838
rect 27794 9774 27806 9826
rect 27858 9774 27870 9826
rect 49410 9774 49422 9826
rect 49474 9774 49486 9826
rect 50978 9774 50990 9826
rect 51042 9774 51054 9826
rect 52546 9774 52558 9826
rect 52610 9774 52622 9826
rect 54114 9774 54126 9826
rect 54178 9774 54190 9826
rect 21086 9762 21138 9774
rect 46398 9762 46450 9774
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 4286 9714 4338 9726
rect 4286 9650 4338 9662
rect 6526 9714 6578 9726
rect 6526 9650 6578 9662
rect 8878 9714 8930 9726
rect 8878 9650 8930 9662
rect 11006 9714 11058 9726
rect 11006 9650 11058 9662
rect 12574 9714 12626 9726
rect 14142 9714 14194 9726
rect 13346 9662 13358 9714
rect 13410 9662 13422 9714
rect 12574 9650 12626 9662
rect 14142 9650 14194 9662
rect 19182 9714 19234 9726
rect 19182 9650 19234 9662
rect 20526 9714 20578 9726
rect 20526 9650 20578 9662
rect 22318 9714 22370 9726
rect 26350 9714 26402 9726
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 22318 9650 22370 9662
rect 26350 9650 26402 9662
rect 30606 9714 30658 9726
rect 30606 9650 30658 9662
rect 46062 9714 46114 9726
rect 53442 9662 53454 9714
rect 53506 9662 53518 9714
rect 46062 9650 46114 9662
rect 26686 9602 26738 9614
rect 26686 9538 26738 9550
rect 27022 9602 27074 9614
rect 27022 9538 27074 9550
rect 42478 9602 42530 9614
rect 42478 9538 42530 9550
rect 51998 9602 52050 9614
rect 51998 9538 52050 9550
rect 55134 9602 55186 9614
rect 55134 9538 55186 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 2046 9266 2098 9278
rect 2046 9202 2098 9214
rect 11342 9266 11394 9278
rect 11342 9202 11394 9214
rect 31726 9266 31778 9278
rect 31726 9202 31778 9214
rect 51214 9266 51266 9278
rect 51214 9202 51266 9214
rect 53006 9266 53058 9278
rect 53006 9202 53058 9214
rect 12910 9154 12962 9166
rect 12910 9090 12962 9102
rect 18062 9154 18114 9166
rect 18062 9090 18114 9102
rect 18846 9154 18898 9166
rect 18846 9090 18898 9102
rect 20974 9154 21026 9166
rect 20974 9090 21026 9102
rect 24558 9154 24610 9166
rect 24558 9090 24610 9102
rect 24782 9154 24834 9166
rect 24782 9090 24834 9102
rect 25230 9154 25282 9166
rect 25230 9090 25282 9102
rect 28814 9154 28866 9166
rect 28814 9090 28866 9102
rect 30718 9154 30770 9166
rect 30718 9090 30770 9102
rect 30942 9154 30994 9166
rect 35758 9154 35810 9166
rect 33394 9102 33406 9154
rect 33458 9102 33470 9154
rect 30942 9090 30994 9102
rect 35758 9090 35810 9102
rect 38110 9154 38162 9166
rect 38110 9090 38162 9102
rect 48078 9154 48130 9166
rect 48078 9090 48130 9102
rect 48974 9154 49026 9166
rect 48974 9090 49026 9102
rect 18622 9042 18674 9054
rect 22654 9042 22706 9054
rect 25006 9042 25058 9054
rect 11890 8990 11902 9042
rect 11954 8990 11966 9042
rect 21298 8990 21310 9042
rect 21362 8990 21374 9042
rect 21746 8990 21758 9042
rect 21810 8990 21822 9042
rect 23202 8990 23214 9042
rect 23266 8990 23278 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 18622 8978 18674 8990
rect 22654 8978 22706 8990
rect 25006 8978 25058 8990
rect 26686 9042 26738 9054
rect 26686 8978 26738 8990
rect 36318 9042 36370 9054
rect 39454 9042 39506 9054
rect 38546 8990 38558 9042
rect 38610 8990 38622 9042
rect 36318 8978 36370 8990
rect 39454 8978 39506 8990
rect 39902 9042 39954 9054
rect 39902 8978 39954 8990
rect 40014 9042 40066 9054
rect 46062 9042 46114 9054
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 42242 8990 42254 9042
rect 42306 8990 42318 9042
rect 43138 8990 43150 9042
rect 43202 8990 43214 9042
rect 40014 8978 40066 8990
rect 46062 8978 46114 8990
rect 48414 9042 48466 9054
rect 52098 8990 52110 9042
rect 52162 8990 52174 9042
rect 53666 8990 53678 9042
rect 53730 8990 53742 9042
rect 48414 8978 48466 8990
rect 5518 8930 5570 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 5518 8866 5570 8878
rect 10446 8930 10498 8942
rect 27246 8930 27298 8942
rect 39678 8930 39730 8942
rect 12114 8878 12126 8930
rect 12178 8878 12190 8930
rect 31938 8878 31950 8930
rect 32002 8878 32014 8930
rect 32274 8878 32286 8930
rect 32338 8878 32350 8930
rect 33730 8878 33742 8930
rect 33794 8878 33806 8930
rect 10446 8866 10498 8878
rect 27246 8866 27298 8878
rect 39678 8866 39730 8878
rect 40686 8930 40738 8942
rect 49870 8930 49922 8942
rect 41458 8878 41470 8930
rect 41522 8878 41534 8930
rect 42466 8878 42478 8930
rect 42530 8878 42542 8930
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 55122 8878 55134 8930
rect 55186 8878 55198 8930
rect 55906 8878 55918 8930
rect 55970 8878 55982 8930
rect 40686 8866 40738 8878
rect 49870 8866 49922 8878
rect 4510 8818 4562 8830
rect 4510 8754 4562 8766
rect 4958 8818 5010 8830
rect 4958 8754 5010 8766
rect 9662 8818 9714 8830
rect 9662 8754 9714 8766
rect 9886 8818 9938 8830
rect 9886 8754 9938 8766
rect 11006 8818 11058 8830
rect 11006 8754 11058 8766
rect 13470 8818 13522 8830
rect 13470 8754 13522 8766
rect 13806 8818 13858 8830
rect 13806 8754 13858 8766
rect 13918 8818 13970 8830
rect 31390 8818 31442 8830
rect 21970 8766 21982 8818
rect 22034 8766 22046 8818
rect 13918 8754 13970 8766
rect 31390 8754 31442 8766
rect 32846 8818 32898 8830
rect 32846 8754 32898 8766
rect 34974 8818 35026 8830
rect 34974 8754 35026 8766
rect 36878 8818 36930 8830
rect 36878 8754 36930 8766
rect 37774 8818 37826 8830
rect 37774 8754 37826 8766
rect 40798 8818 40850 8830
rect 45278 8818 45330 8830
rect 42018 8766 42030 8818
rect 42082 8766 42094 8818
rect 40798 8754 40850 8766
rect 45278 8754 45330 8766
rect 45502 8818 45554 8830
rect 45502 8754 45554 8766
rect 49310 8818 49362 8830
rect 49310 8754 49362 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 12462 8482 12514 8494
rect 12462 8418 12514 8430
rect 28590 8482 28642 8494
rect 28590 8418 28642 8430
rect 33294 8482 33346 8494
rect 33294 8418 33346 8430
rect 33518 8482 33570 8494
rect 33518 8418 33570 8430
rect 39006 8482 39058 8494
rect 39006 8418 39058 8430
rect 41918 8482 41970 8494
rect 41918 8418 41970 8430
rect 49086 8482 49138 8494
rect 49086 8418 49138 8430
rect 14926 8370 14978 8382
rect 13458 8318 13470 8370
rect 13522 8318 13534 8370
rect 13906 8318 13918 8370
rect 13970 8318 13982 8370
rect 14926 8306 14978 8318
rect 18398 8370 18450 8382
rect 18398 8306 18450 8318
rect 18510 8370 18562 8382
rect 18510 8306 18562 8318
rect 28030 8370 28082 8382
rect 28030 8306 28082 8318
rect 28926 8370 28978 8382
rect 28926 8306 28978 8318
rect 29710 8370 29762 8382
rect 29710 8306 29762 8318
rect 35086 8370 35138 8382
rect 36654 8370 36706 8382
rect 41134 8370 41186 8382
rect 35746 8318 35758 8370
rect 35810 8318 35822 8370
rect 36082 8318 36094 8370
rect 36146 8318 36158 8370
rect 37986 8318 37998 8370
rect 38050 8318 38062 8370
rect 38434 8318 38446 8370
rect 38498 8318 38510 8370
rect 35086 8306 35138 8318
rect 36654 8306 36706 8318
rect 41134 8306 41186 8318
rect 41582 8370 41634 8382
rect 41582 8306 41634 8318
rect 42142 8370 42194 8382
rect 42142 8306 42194 8318
rect 42254 8370 42306 8382
rect 42254 8306 42306 8318
rect 50318 8370 50370 8382
rect 51762 8318 51774 8370
rect 51826 8318 51838 8370
rect 53330 8318 53342 8370
rect 53394 8318 53406 8370
rect 50318 8306 50370 8318
rect 7758 8258 7810 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 7758 8194 7810 8206
rect 14366 8258 14418 8270
rect 14366 8194 14418 8206
rect 18734 8258 18786 8270
rect 18734 8194 18786 8206
rect 19070 8258 19122 8270
rect 37438 8258 37490 8270
rect 29362 8206 29374 8258
rect 29426 8206 29438 8258
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 19070 8194 19122 8206
rect 37438 8194 37490 8206
rect 38670 8258 38722 8270
rect 38670 8194 38722 8206
rect 40798 8258 40850 8270
rect 40798 8194 40850 8206
rect 41022 8258 41074 8270
rect 41022 8194 41074 8206
rect 41358 8258 41410 8270
rect 41358 8194 41410 8206
rect 49758 8258 49810 8270
rect 50978 8206 50990 8258
rect 51042 8206 51054 8258
rect 52546 8206 52558 8258
rect 52610 8206 52622 8258
rect 54114 8206 54126 8258
rect 54178 8206 54190 8258
rect 49758 8194 49810 8206
rect 1262 8146 1314 8158
rect 1262 8082 1314 8094
rect 7422 8146 7474 8158
rect 15150 8146 15202 8158
rect 8194 8094 8206 8146
rect 8258 8094 8270 8146
rect 7422 8082 7474 8094
rect 15150 8082 15202 8094
rect 31166 8146 31218 8158
rect 31166 8082 31218 8094
rect 34078 8146 34130 8158
rect 37214 8146 37266 8158
rect 34626 8094 34638 8146
rect 34690 8094 34702 8146
rect 34078 8082 34130 8094
rect 37214 8082 37266 8094
rect 49422 8146 49474 8158
rect 49422 8082 49474 8094
rect 50542 8146 50594 8158
rect 50542 8082 50594 8094
rect 55134 8146 55186 8158
rect 55134 8082 55186 8094
rect 12798 8034 12850 8046
rect 12798 7970 12850 7982
rect 13134 8034 13186 8046
rect 13134 7970 13186 7982
rect 18958 8034 19010 8046
rect 18958 7970 19010 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 41694 8034 41746 8046
rect 41694 7970 41746 7982
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 19966 7698 20018 7710
rect 19966 7634 20018 7646
rect 28926 7698 28978 7710
rect 28926 7634 28978 7646
rect 53006 7698 53058 7710
rect 53006 7634 53058 7646
rect 56142 7698 56194 7710
rect 56142 7634 56194 7646
rect 7758 7586 7810 7598
rect 14030 7586 14082 7598
rect 8306 7534 8318 7586
rect 8370 7534 8382 7586
rect 7758 7522 7810 7534
rect 14030 7522 14082 7534
rect 14702 7586 14754 7598
rect 30046 7586 30098 7598
rect 16146 7534 16158 7586
rect 16210 7534 16222 7586
rect 19730 7534 19742 7586
rect 19794 7534 19806 7586
rect 14702 7522 14754 7534
rect 30046 7522 30098 7534
rect 30382 7586 30434 7598
rect 30382 7522 30434 7534
rect 34302 7586 34354 7598
rect 34302 7522 34354 7534
rect 34974 7586 35026 7598
rect 34974 7522 35026 7534
rect 35198 7586 35250 7598
rect 35198 7522 35250 7534
rect 35422 7586 35474 7598
rect 35422 7522 35474 7534
rect 35646 7586 35698 7598
rect 35646 7522 35698 7534
rect 35870 7586 35922 7598
rect 35870 7522 35922 7534
rect 49646 7586 49698 7598
rect 49646 7522 49698 7534
rect 54574 7586 54626 7598
rect 54574 7522 54626 7534
rect 12238 7474 12290 7486
rect 14478 7474 14530 7486
rect 13570 7422 13582 7474
rect 13634 7422 13646 7474
rect 12238 7410 12290 7422
rect 14478 7410 14530 7422
rect 18622 7474 18674 7486
rect 18622 7410 18674 7422
rect 18958 7474 19010 7486
rect 49982 7474 50034 7486
rect 19618 7422 19630 7474
rect 19682 7422 19694 7474
rect 36642 7422 36654 7474
rect 36706 7422 36718 7474
rect 37090 7422 37102 7474
rect 37154 7422 37166 7474
rect 38546 7422 38558 7474
rect 38610 7422 38622 7474
rect 39330 7422 39342 7474
rect 39394 7422 39406 7474
rect 18958 7410 19010 7422
rect 49982 7410 50034 7422
rect 50542 7474 50594 7486
rect 50542 7410 50594 7422
rect 50878 7474 50930 7486
rect 55122 7422 55134 7474
rect 55186 7422 55198 7474
rect 50878 7410 50930 7422
rect 17726 7362 17778 7374
rect 8642 7310 8654 7362
rect 8706 7310 8718 7362
rect 16482 7310 16494 7362
rect 16546 7310 16558 7362
rect 17726 7298 17778 7310
rect 18286 7362 18338 7374
rect 18286 7298 18338 7310
rect 19294 7362 19346 7374
rect 36318 7362 36370 7374
rect 29138 7310 29150 7362
rect 29202 7310 29214 7362
rect 29698 7310 29710 7362
rect 29762 7310 29774 7362
rect 19294 7298 19346 7310
rect 36318 7298 36370 7310
rect 37774 7362 37826 7374
rect 37774 7298 37826 7310
rect 42590 7362 42642 7374
rect 42590 7298 42642 7310
rect 51438 7362 51490 7374
rect 51986 7310 51998 7362
rect 52050 7310 52062 7362
rect 53554 7310 53566 7362
rect 53618 7310 53630 7362
rect 51438 7298 51490 7310
rect 9886 7250 9938 7262
rect 9886 7186 9938 7198
rect 11902 7250 11954 7262
rect 11902 7186 11954 7198
rect 12126 7250 12178 7262
rect 12126 7186 12178 7198
rect 14366 7250 14418 7262
rect 14366 7186 14418 7198
rect 15598 7250 15650 7262
rect 15598 7186 15650 7198
rect 18398 7250 18450 7262
rect 18398 7186 18450 7198
rect 18846 7250 18898 7262
rect 18846 7186 18898 7198
rect 28590 7250 28642 7262
rect 42030 7250 42082 7262
rect 37314 7198 37326 7250
rect 37378 7198 37390 7250
rect 28590 7186 28642 7198
rect 42030 7186 42082 7198
rect 42254 7250 42306 7262
rect 42254 7186 42306 7198
rect 43150 7250 43202 7262
rect 43150 7186 43202 7198
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 18622 6914 18674 6926
rect 18622 6850 18674 6862
rect 20750 6914 20802 6926
rect 20750 6850 20802 6862
rect 22878 6914 22930 6926
rect 22878 6850 22930 6862
rect 23998 6914 24050 6926
rect 23998 6850 24050 6862
rect 16718 6802 16770 6814
rect 16718 6738 16770 6750
rect 18734 6802 18786 6814
rect 21634 6750 21646 6802
rect 21698 6750 21710 6802
rect 25218 6750 25230 6802
rect 25282 6750 25294 6802
rect 41794 6750 41806 6802
rect 41858 6750 41870 6802
rect 42018 6750 42030 6802
rect 42082 6750 42094 6802
rect 42242 6750 42254 6802
rect 42306 6750 42318 6802
rect 43362 6750 43374 6802
rect 43426 6750 43438 6802
rect 43698 6750 43710 6802
rect 43762 6750 43774 6802
rect 18734 6738 18786 6750
rect 10558 6690 10610 6702
rect 10558 6626 10610 6638
rect 11006 6690 11058 6702
rect 11006 6626 11058 6638
rect 11118 6690 11170 6702
rect 11118 6626 11170 6638
rect 11230 6690 11282 6702
rect 11230 6626 11282 6638
rect 11566 6690 11618 6702
rect 11566 6626 11618 6638
rect 11790 6690 11842 6702
rect 11790 6626 11842 6638
rect 12126 6690 12178 6702
rect 12126 6626 12178 6638
rect 12350 6690 12402 6702
rect 12350 6626 12402 6638
rect 18286 6690 18338 6702
rect 18286 6626 18338 6638
rect 18846 6690 18898 6702
rect 31838 6690 31890 6702
rect 24770 6638 24782 6690
rect 24834 6638 24846 6690
rect 18846 6626 18898 6638
rect 31838 6626 31890 6638
rect 36094 6690 36146 6702
rect 36094 6626 36146 6638
rect 40686 6690 40738 6702
rect 40686 6626 40738 6638
rect 42814 6690 42866 6702
rect 42814 6626 42866 6638
rect 45614 6690 45666 6702
rect 45614 6626 45666 6638
rect 45838 6690 45890 6702
rect 45838 6626 45890 6638
rect 50206 6690 50258 6702
rect 50206 6626 50258 6638
rect 50542 6690 50594 6702
rect 50542 6626 50594 6638
rect 51102 6690 51154 6702
rect 51102 6626 51154 6638
rect 51438 6690 51490 6702
rect 52658 6638 52670 6690
rect 52722 6638 52734 6690
rect 54226 6638 54238 6690
rect 54290 6638 54302 6690
rect 51438 6626 51490 6638
rect 12014 6578 12066 6590
rect 12014 6514 12066 6526
rect 16270 6578 16322 6590
rect 16270 6514 16322 6526
rect 17278 6578 17330 6590
rect 31278 6578 31330 6590
rect 21298 6526 21310 6578
rect 21362 6526 21374 6578
rect 17278 6514 17330 6526
rect 31278 6514 31330 6526
rect 40462 6578 40514 6590
rect 46274 6526 46286 6578
rect 46338 6526 46350 6578
rect 51874 6526 51886 6578
rect 51938 6526 51950 6578
rect 53218 6526 53230 6578
rect 53282 6526 53294 6578
rect 40462 6514 40514 6526
rect 10670 6466 10722 6478
rect 10670 6402 10722 6414
rect 26350 6466 26402 6478
rect 26350 6402 26402 6414
rect 41134 6466 41186 6478
rect 41134 6402 41186 6414
rect 41470 6466 41522 6478
rect 41470 6402 41522 6414
rect 43150 6466 43202 6478
rect 43150 6402 43202 6414
rect 55134 6466 55186 6478
rect 55134 6402 55186 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 9438 6130 9490 6142
rect 9438 6066 9490 6078
rect 11566 6130 11618 6142
rect 11566 6066 11618 6078
rect 27022 6130 27074 6142
rect 27022 6066 27074 6078
rect 32622 6130 32674 6142
rect 32622 6066 32674 6078
rect 32958 6130 33010 6142
rect 32958 6066 33010 6078
rect 37326 6130 37378 6142
rect 37326 6066 37378 6078
rect 53006 6130 53058 6142
rect 53006 6066 53058 6078
rect 56142 6130 56194 6142
rect 56142 6066 56194 6078
rect 6414 6018 6466 6030
rect 21310 6018 21362 6030
rect 7858 5966 7870 6018
rect 7922 5966 7934 6018
rect 6414 5954 6466 5966
rect 21310 5954 21362 5966
rect 22206 6018 22258 6030
rect 22206 5954 22258 5966
rect 24334 6018 24386 6030
rect 29262 6018 29314 6030
rect 25106 5966 25118 6018
rect 25170 5966 25182 6018
rect 28578 5966 28590 6018
rect 28642 5966 28654 6018
rect 24334 5954 24386 5966
rect 29262 5954 29314 5966
rect 38558 6018 38610 6030
rect 38558 5954 38610 5966
rect 41470 6018 41522 6030
rect 41470 5954 41522 5966
rect 41806 6018 41858 6030
rect 41806 5954 41858 5966
rect 42702 6018 42754 6030
rect 42702 5954 42754 5966
rect 48638 6018 48690 6030
rect 48638 5954 48690 5966
rect 54574 6018 54626 6030
rect 54574 5954 54626 5966
rect 6750 5906 6802 5918
rect 6750 5842 6802 5854
rect 21646 5906 21698 5918
rect 21646 5842 21698 5854
rect 24670 5906 24722 5918
rect 24670 5842 24722 5854
rect 26238 5906 26290 5918
rect 38446 5906 38498 5918
rect 30370 5854 30382 5906
rect 30434 5854 30446 5906
rect 26238 5842 26290 5854
rect 38446 5842 38498 5854
rect 38782 5906 38834 5918
rect 38782 5842 38834 5854
rect 39230 5906 39282 5918
rect 39230 5842 39282 5854
rect 39566 5906 39618 5918
rect 48974 5906 49026 5918
rect 42242 5854 42254 5906
rect 42306 5854 42318 5906
rect 52098 5854 52110 5906
rect 52162 5854 52174 5906
rect 53554 5854 53566 5906
rect 53618 5854 53630 5906
rect 39566 5842 39618 5854
rect 48974 5842 49026 5854
rect 7310 5794 7362 5806
rect 11678 5794 11730 5806
rect 8306 5742 8318 5794
rect 8370 5742 8382 5794
rect 7310 5730 7362 5742
rect 11678 5730 11730 5742
rect 25678 5794 25730 5806
rect 29038 5794 29090 5806
rect 32062 5794 32114 5806
rect 37214 5794 37266 5806
rect 27234 5742 27246 5794
rect 27298 5742 27310 5794
rect 27682 5742 27694 5794
rect 27746 5742 27758 5794
rect 30818 5742 30830 5794
rect 30882 5742 30894 5794
rect 33170 5742 33182 5794
rect 33234 5742 33246 5794
rect 33618 5742 33630 5794
rect 33682 5742 33694 5794
rect 25678 5730 25730 5742
rect 29038 5730 29090 5742
rect 32062 5730 32114 5742
rect 37214 5730 37266 5742
rect 38110 5794 38162 5806
rect 38110 5730 38162 5742
rect 39454 5794 39506 5806
rect 39454 5730 39506 5742
rect 49534 5794 49586 5806
rect 55122 5742 55134 5794
rect 55186 5742 55198 5794
rect 49534 5730 49586 5742
rect 26686 5682 26738 5694
rect 26686 5618 26738 5630
rect 29934 5682 29986 5694
rect 29934 5618 29986 5630
rect 37102 5682 37154 5694
rect 37102 5618 37154 5630
rect 51102 5682 51154 5694
rect 51102 5618 51154 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 7422 5346 7474 5358
rect 7422 5282 7474 5294
rect 12014 5346 12066 5358
rect 12014 5282 12066 5294
rect 15934 5346 15986 5358
rect 15934 5282 15986 5294
rect 16606 5346 16658 5358
rect 16606 5282 16658 5294
rect 23774 5346 23826 5358
rect 23774 5282 23826 5294
rect 26574 5346 26626 5358
rect 26574 5282 26626 5294
rect 28254 5346 28306 5358
rect 28254 5282 28306 5294
rect 28478 5346 28530 5358
rect 28478 5282 28530 5294
rect 30718 5346 30770 5358
rect 30718 5282 30770 5294
rect 30942 5346 30994 5358
rect 30942 5282 30994 5294
rect 31838 5346 31890 5358
rect 31838 5282 31890 5294
rect 32286 5346 32338 5358
rect 32286 5282 32338 5294
rect 35758 5346 35810 5358
rect 35758 5282 35810 5294
rect 39454 5346 39506 5358
rect 39454 5282 39506 5294
rect 53006 5346 53058 5358
rect 53006 5282 53058 5294
rect 53230 5346 53282 5358
rect 53230 5282 53282 5294
rect 12462 5234 12514 5246
rect 13918 5234 13970 5246
rect 31502 5234 31554 5246
rect 13458 5182 13470 5234
rect 13522 5182 13534 5234
rect 22978 5182 22990 5234
rect 23042 5182 23054 5234
rect 23202 5182 23214 5234
rect 23266 5182 23278 5234
rect 23426 5182 23438 5234
rect 23490 5182 23502 5234
rect 12462 5170 12514 5182
rect 13918 5170 13970 5182
rect 31502 5170 31554 5182
rect 33630 5234 33682 5246
rect 38670 5234 38722 5246
rect 34514 5182 34526 5234
rect 34578 5182 34590 5234
rect 33630 5170 33682 5182
rect 38670 5170 38722 5182
rect 39678 5234 39730 5246
rect 54114 5182 54126 5234
rect 54178 5182 54190 5234
rect 39678 5170 39730 5182
rect 20974 5122 21026 5134
rect 11778 5070 11790 5122
rect 11842 5070 11854 5122
rect 12898 5070 12910 5122
rect 12962 5070 12974 5122
rect 13346 5070 13358 5122
rect 13410 5070 13422 5122
rect 14690 5070 14702 5122
rect 14754 5070 14766 5122
rect 15474 5070 15486 5122
rect 15538 5070 15550 5122
rect 20974 5058 21026 5070
rect 21310 5122 21362 5134
rect 21310 5058 21362 5070
rect 21870 5122 21922 5134
rect 21870 5058 21922 5070
rect 22318 5122 22370 5134
rect 22318 5058 22370 5070
rect 38782 5122 38834 5134
rect 38782 5058 38834 5070
rect 39118 5122 39170 5134
rect 39118 5058 39170 5070
rect 39454 5122 39506 5134
rect 39454 5058 39506 5070
rect 51662 5122 51714 5134
rect 51662 5058 51714 5070
rect 51998 5122 52050 5134
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 51998 5058 52050 5070
rect 12126 5010 12178 5022
rect 12126 4946 12178 4958
rect 16158 5010 16210 5022
rect 16158 4946 16210 4958
rect 22654 5010 22706 5022
rect 34178 4958 34190 5010
rect 34242 4958 34254 5010
rect 52434 4958 52446 5010
rect 52498 4958 52510 5010
rect 53666 4958 53678 5010
rect 53730 4958 53742 5010
rect 22654 4946 22706 4958
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 10894 4562 10946 4574
rect 10894 4498 10946 4510
rect 17950 4562 18002 4574
rect 17950 4498 18002 4510
rect 18286 4562 18338 4574
rect 18286 4498 18338 4510
rect 22990 4562 23042 4574
rect 22990 4498 23042 4510
rect 39454 4562 39506 4574
rect 39454 4498 39506 4510
rect 54574 4562 54626 4574
rect 54574 4498 54626 4510
rect 56142 4562 56194 4574
rect 56142 4498 56194 4510
rect 8766 4450 8818 4462
rect 12686 4450 12738 4462
rect 9314 4398 9326 4450
rect 9378 4398 9390 4450
rect 11778 4398 11790 4450
rect 11842 4398 11854 4450
rect 8766 4386 8818 4398
rect 12686 4386 12738 4398
rect 13470 4450 13522 4462
rect 13470 4386 13522 4398
rect 14254 4450 14306 4462
rect 14254 4386 14306 4398
rect 16046 4450 16098 4462
rect 16046 4386 16098 4398
rect 16158 4450 16210 4462
rect 16158 4386 16210 4398
rect 19406 4450 19458 4462
rect 19406 4386 19458 4398
rect 19630 4450 19682 4462
rect 19630 4386 19682 4398
rect 20862 4450 20914 4462
rect 34078 4450 34130 4462
rect 21410 4398 21422 4450
rect 21474 4398 21486 4450
rect 20862 4386 20914 4398
rect 34078 4386 34130 4398
rect 44158 4450 44210 4462
rect 49534 4450 49586 4462
rect 52334 4450 52386 4462
rect 44930 4398 44942 4450
rect 44994 4398 45006 4450
rect 50306 4398 50318 4450
rect 50370 4398 50382 4450
rect 44158 4386 44210 4398
rect 49534 4386 49586 4398
rect 52334 4386 52386 4398
rect 12238 4338 12290 4350
rect 12238 4274 12290 4286
rect 14030 4338 14082 4350
rect 27582 4338 27634 4350
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 14030 4274 14082 4286
rect 27582 4274 27634 4286
rect 28478 4338 28530 4350
rect 39566 4338 39618 4350
rect 34514 4286 34526 4338
rect 34578 4286 34590 4338
rect 28478 4274 28530 4286
rect 39566 4274 39618 4286
rect 44494 4338 44546 4350
rect 44494 4274 44546 4286
rect 49870 4338 49922 4350
rect 49870 4274 49922 4286
rect 52670 4338 52722 4350
rect 55122 4286 55134 4338
rect 55186 4286 55198 4338
rect 52670 4274 52722 4286
rect 15150 4226 15202 4238
rect 9762 4174 9774 4226
rect 9826 4174 9838 4226
rect 15150 4162 15202 4174
rect 15710 4226 15762 4238
rect 27022 4226 27074 4238
rect 18834 4174 18846 4226
rect 18898 4174 18910 4226
rect 21746 4174 21758 4226
rect 21810 4174 21822 4226
rect 15710 4162 15762 4174
rect 27022 4162 27074 4174
rect 27246 4226 27298 4238
rect 27246 4162 27298 4174
rect 34974 4226 35026 4238
rect 34974 4162 35026 4174
rect 53230 4226 53282 4238
rect 53554 4174 53566 4226
rect 53618 4174 53630 4226
rect 53230 4162 53282 4174
rect 27470 4114 27522 4126
rect 27470 4050 27522 4062
rect 28590 4114 28642 4126
rect 28590 4050 28642 4062
rect 28814 4114 28866 4126
rect 28814 4050 28866 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 9102 3778 9154 3790
rect 9102 3714 9154 3726
rect 9326 3778 9378 3790
rect 9326 3714 9378 3726
rect 18510 3778 18562 3790
rect 18510 3714 18562 3726
rect 18846 3778 18898 3790
rect 18846 3714 18898 3726
rect 19966 3778 20018 3790
rect 19966 3714 20018 3726
rect 26910 3778 26962 3790
rect 26910 3714 26962 3726
rect 27246 3778 27298 3790
rect 27246 3714 27298 3726
rect 32398 3778 32450 3790
rect 32398 3714 32450 3726
rect 35198 3778 35250 3790
rect 35198 3714 35250 3726
rect 51438 3778 51490 3790
rect 51438 3714 51490 3726
rect 51662 3778 51714 3790
rect 51662 3714 51714 3726
rect 17950 3666 18002 3678
rect 17950 3602 18002 3614
rect 19070 3666 19122 3678
rect 19070 3602 19122 3614
rect 27358 3666 27410 3678
rect 27358 3602 27410 3614
rect 28702 3666 28754 3678
rect 28702 3602 28754 3614
rect 29710 3666 29762 3678
rect 52222 3666 52274 3678
rect 36082 3614 36094 3666
rect 36146 3614 36158 3666
rect 52546 3614 52558 3666
rect 52610 3614 52622 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 29710 3602 29762 3614
rect 52222 3602 52274 3614
rect 26798 3554 26850 3566
rect 19506 3502 19518 3554
rect 19570 3502 19582 3554
rect 26798 3490 26850 3502
rect 28926 3554 28978 3566
rect 28926 3490 28978 3502
rect 29262 3554 29314 3566
rect 35634 3502 35646 3554
rect 35698 3502 35710 3554
rect 54114 3502 54126 3554
rect 54178 3502 54190 3554
rect 29262 3490 29314 3502
rect 9886 3442 9938 3454
rect 9886 3378 9938 3390
rect 28814 3442 28866 3454
rect 53566 3442 53618 3454
rect 29586 3390 29598 3442
rect 29650 3390 29662 3442
rect 28814 3378 28866 3390
rect 53566 3378 53618 3390
rect 29934 3330 29986 3342
rect 29934 3266 29986 3278
rect 37326 3330 37378 3342
rect 37326 3266 37378 3278
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 26910 2994 26962 3006
rect 26910 2930 26962 2942
rect 38222 2994 38274 3006
rect 38222 2930 38274 2942
rect 54574 2994 54626 3006
rect 54574 2930 54626 2942
rect 56142 2994 56194 3006
rect 56142 2930 56194 2942
rect 21198 2882 21250 2894
rect 21198 2818 21250 2830
rect 24782 2882 24834 2894
rect 24782 2818 24834 2830
rect 28366 2882 28418 2894
rect 28366 2818 28418 2830
rect 28702 2882 28754 2894
rect 28702 2818 28754 2830
rect 28926 2882 28978 2894
rect 28926 2818 28978 2830
rect 33294 2882 33346 2894
rect 33294 2818 33346 2830
rect 34862 2882 34914 2894
rect 40574 2882 40626 2894
rect 35634 2830 35646 2882
rect 35698 2830 35710 2882
rect 34862 2818 34914 2830
rect 40574 2818 40626 2830
rect 41582 2882 41634 2894
rect 41582 2818 41634 2830
rect 48414 2882 48466 2894
rect 48414 2818 48466 2830
rect 50542 2882 50594 2894
rect 50542 2818 50594 2830
rect 21534 2770 21586 2782
rect 30382 2770 30434 2782
rect 32510 2770 32562 2782
rect 25218 2718 25230 2770
rect 25282 2718 25294 2770
rect 29250 2718 29262 2770
rect 29314 2718 29326 2770
rect 29698 2718 29710 2770
rect 29762 2718 29774 2770
rect 30930 2718 30942 2770
rect 30994 2718 31006 2770
rect 32050 2718 32062 2770
rect 32114 2718 32126 2770
rect 21534 2706 21586 2718
rect 30382 2706 30434 2718
rect 32510 2706 32562 2718
rect 35198 2770 35250 2782
rect 50878 2770 50930 2782
rect 36530 2718 36542 2770
rect 36594 2718 36606 2770
rect 52098 2718 52110 2770
rect 52162 2718 52174 2770
rect 53554 2718 53566 2770
rect 53618 2718 53630 2770
rect 55122 2718 55134 2770
rect 55186 2718 55198 2770
rect 35198 2706 35250 2718
rect 50878 2706 50930 2718
rect 22094 2658 22146 2670
rect 33070 2658 33122 2670
rect 51438 2658 51490 2670
rect 25666 2606 25678 2658
rect 25730 2606 25742 2658
rect 29922 2606 29934 2658
rect 29986 2606 29998 2658
rect 36978 2606 36990 2658
rect 37042 2606 37054 2658
rect 52770 2606 52782 2658
rect 52834 2606 52846 2658
rect 22094 2594 22146 2606
rect 33070 2594 33122 2606
rect 51438 2594 51490 2606
rect 39790 2546 39842 2558
rect 39790 2482 39842 2494
rect 40014 2546 40066 2558
rect 40014 2482 40066 2494
rect 42142 2546 42194 2558
rect 42142 2482 42194 2494
rect 42478 2546 42530 2558
rect 42478 2482 42530 2494
rect 47630 2546 47682 2558
rect 47630 2482 47682 2494
rect 47854 2546 47906 2558
rect 47854 2482 47906 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 23102 2210 23154 2222
rect 23102 2146 23154 2158
rect 23438 2210 23490 2222
rect 23438 2146 23490 2158
rect 26350 2210 26402 2222
rect 26350 2146 26402 2158
rect 28702 2210 28754 2222
rect 28702 2146 28754 2158
rect 29038 2210 29090 2222
rect 29038 2146 29090 2158
rect 30158 2210 30210 2222
rect 30158 2146 30210 2158
rect 30494 2210 30546 2222
rect 30494 2146 30546 2158
rect 32398 2210 32450 2222
rect 32398 2146 32450 2158
rect 36206 2210 36258 2222
rect 36206 2146 36258 2158
rect 36430 2210 36482 2222
rect 36430 2146 36482 2158
rect 36654 2210 36706 2222
rect 36654 2146 36706 2158
rect 40910 2210 40962 2222
rect 40910 2146 40962 2158
rect 41134 2210 41186 2222
rect 49074 2158 49086 2210
rect 49138 2158 49150 2210
rect 41134 2146 41186 2158
rect 41694 2098 41746 2110
rect 12898 2046 12910 2098
rect 12962 2046 12974 2098
rect 25106 2046 25118 2098
rect 25170 2046 25182 2098
rect 41694 2034 41746 2046
rect 47518 2098 47570 2110
rect 47518 2034 47570 2046
rect 50430 2098 50482 2110
rect 50430 2034 50482 2046
rect 51326 2098 51378 2110
rect 51326 2034 51378 2046
rect 52222 2098 52274 2110
rect 52546 2046 52558 2098
rect 52610 2046 52622 2098
rect 54114 2046 54126 2098
rect 54178 2046 54190 2098
rect 54898 2046 54910 2098
rect 54962 2046 54974 2098
rect 52222 2034 52274 2046
rect 28142 1986 28194 1998
rect 24770 1934 24782 1986
rect 24834 1934 24846 1986
rect 28142 1922 28194 1934
rect 38446 1986 38498 1998
rect 38446 1922 38498 1934
rect 46958 1986 47010 1998
rect 49870 1986 49922 1998
rect 49298 1934 49310 1986
rect 49362 1934 49374 1986
rect 46958 1922 47010 1934
rect 49870 1922 49922 1934
rect 50766 1986 50818 1998
rect 50766 1922 50818 1934
rect 51662 1986 51714 1998
rect 51662 1922 51714 1934
rect 23998 1874 24050 1886
rect 23998 1810 24050 1822
rect 29598 1874 29650 1886
rect 29598 1810 29650 1822
rect 37214 1874 37266 1886
rect 38670 1874 38722 1886
rect 37986 1822 37998 1874
rect 38050 1822 38062 1874
rect 37214 1810 37266 1822
rect 38670 1810 38722 1822
rect 46734 1874 46786 1886
rect 46734 1810 46786 1822
rect 48750 1874 48802 1886
rect 48750 1810 48802 1822
rect 53566 1874 53618 1886
rect 53566 1810 53618 1822
rect 11902 1762 11954 1774
rect 11902 1698 11954 1710
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 53566 1426 53618 1438
rect 53566 1362 53618 1374
rect 56142 1426 56194 1438
rect 56142 1362 56194 1374
rect 5518 1314 5570 1326
rect 9886 1314 9938 1326
rect 7410 1262 7422 1314
rect 7474 1262 7486 1314
rect 5518 1250 5570 1262
rect 9886 1250 9938 1262
rect 13918 1314 13970 1326
rect 13918 1250 13970 1262
rect 24334 1314 24386 1326
rect 24334 1250 24386 1262
rect 25230 1314 25282 1326
rect 25230 1250 25282 1262
rect 26126 1314 26178 1326
rect 26126 1250 26178 1262
rect 50430 1314 50482 1326
rect 50430 1250 50482 1262
rect 50654 1314 50706 1326
rect 50654 1250 50706 1262
rect 51998 1314 52050 1326
rect 51998 1250 52050 1262
rect 6514 1150 6526 1202
rect 6578 1150 6590 1202
rect 8082 1150 8094 1202
rect 8146 1150 8158 1202
rect 10882 1150 10894 1202
rect 10946 1150 10958 1202
rect 14802 1150 14814 1202
rect 14866 1150 14878 1202
rect 25666 1150 25678 1202
rect 25730 1150 25742 1202
rect 50978 1150 50990 1202
rect 51042 1150 51054 1202
rect 52546 1150 52558 1202
rect 52610 1150 52622 1202
rect 55122 1038 55134 1090
rect 55186 1038 55198 1090
rect 49534 978 49586 990
rect 49534 914 49586 926
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 2158 13134 2210 13186
rect 3726 13134 3778 13186
rect 5966 13134 6018 13186
rect 7534 13134 7586 13186
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 17390 13134 17442 13186
rect 18958 13134 19010 13186
rect 22654 13134 22706 13186
rect 25454 13134 25506 13186
rect 41918 13134 41970 13186
rect 42142 13134 42194 13186
rect 48974 13134 49026 13186
rect 51102 13134 51154 13186
rect 54910 13134 54962 13186
rect 11902 13022 11954 13074
rect 13358 13022 13410 13074
rect 14926 13022 14978 13074
rect 23886 13022 23938 13074
rect 48414 13022 48466 13074
rect 52894 13022 52946 13074
rect 2718 12910 2770 12962
rect 4286 12910 4338 12962
rect 6302 12910 6354 12962
rect 8094 12910 8146 12962
rect 10222 12910 10274 12962
rect 14142 12910 14194 12962
rect 15710 12910 15762 12962
rect 17838 12910 17890 12962
rect 19518 12910 19570 12962
rect 20526 12910 20578 12962
rect 22094 12910 22146 12962
rect 31726 12910 31778 12962
rect 44942 12910 44994 12962
rect 46846 12910 46898 12962
rect 50766 12910 50818 12962
rect 52334 12910 52386 12962
rect 54574 12910 54626 12962
rect 21534 12798 21586 12850
rect 26014 12798 26066 12850
rect 31390 12798 31442 12850
rect 32286 12798 32338 12850
rect 47854 12798 47906 12850
rect 50094 12798 50146 12850
rect 24446 12686 24498 12738
rect 45950 12686 46002 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 2270 12350 2322 12402
rect 6974 12350 7026 12402
rect 10110 12350 10162 12402
rect 12014 12350 12066 12402
rect 14814 12350 14866 12402
rect 16382 12350 16434 12402
rect 17950 12350 18002 12402
rect 23550 12350 23602 12402
rect 47966 12350 48018 12402
rect 49086 12350 49138 12402
rect 52558 12350 52610 12402
rect 54126 12350 54178 12402
rect 55694 12350 55746 12402
rect 3614 12238 3666 12290
rect 5070 12238 5122 12290
rect 8206 12238 8258 12290
rect 13806 12238 13858 12290
rect 19406 12238 19458 12290
rect 20862 12238 20914 12290
rect 22206 12238 22258 12290
rect 31054 12238 31106 12290
rect 36878 12238 36930 12290
rect 37886 12238 37938 12290
rect 41358 12238 41410 12290
rect 42254 12238 42306 12290
rect 46846 12238 46898 12290
rect 2830 12126 2882 12178
rect 4174 12126 4226 12178
rect 8878 12126 8930 12178
rect 11006 12126 11058 12178
rect 15374 12126 15426 12178
rect 16942 12126 16994 12178
rect 18286 12126 18338 12178
rect 20638 12126 20690 12178
rect 21422 12126 21474 12178
rect 22990 12126 23042 12178
rect 26238 12126 26290 12178
rect 31838 12126 31890 12178
rect 32286 12126 32338 12178
rect 36318 12126 36370 12178
rect 41806 12126 41858 12178
rect 42702 12126 42754 12178
rect 49982 12126 50034 12178
rect 52222 12126 52274 12178
rect 55358 12126 55410 12178
rect 7534 12014 7586 12066
rect 10670 12014 10722 12066
rect 20078 12014 20130 12066
rect 24558 12014 24610 12066
rect 25902 12014 25954 12066
rect 27022 12014 27074 12066
rect 31390 12014 31442 12066
rect 32846 12014 32898 12066
rect 38222 12014 38274 12066
rect 44270 12014 44322 12066
rect 44494 12014 44546 12066
rect 45054 12014 45106 12066
rect 45950 12014 46002 12066
rect 48526 12014 48578 12066
rect 50990 12014 51042 12066
rect 53566 12014 53618 12066
rect 5518 11902 5570 11954
rect 5742 11902 5794 11954
rect 13022 11902 13074 11954
rect 13246 11902 13298 11954
rect 25118 11902 25170 11954
rect 25342 11902 25394 11954
rect 37326 11902 37378 11954
rect 39454 11902 39506 11954
rect 45390 11902 45442 11954
rect 46398 11902 46450 11954
rect 50430 11902 50482 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 4622 11566 4674 11618
rect 6190 11566 6242 11618
rect 7758 11566 7810 11618
rect 8878 11566 8930 11618
rect 9214 11566 9266 11618
rect 10894 11566 10946 11618
rect 14030 11566 14082 11618
rect 17502 11566 17554 11618
rect 19070 11566 19122 11618
rect 38222 11566 38274 11618
rect 38446 11566 38498 11618
rect 42366 11566 42418 11618
rect 42590 11566 42642 11618
rect 50318 11566 50370 11618
rect 51886 11566 51938 11618
rect 53454 11566 53506 11618
rect 13022 11454 13074 11506
rect 20414 11454 20466 11506
rect 21198 11454 21250 11506
rect 21982 11454 22034 11506
rect 25678 11454 25730 11506
rect 26014 11454 26066 11506
rect 34750 11454 34802 11506
rect 42030 11454 42082 11506
rect 46062 11454 46114 11506
rect 48974 11454 49026 11506
rect 1486 11342 1538 11394
rect 3614 11342 3666 11394
rect 5182 11342 5234 11394
rect 6638 11342 6690 11394
rect 8094 11342 8146 11394
rect 11454 11342 11506 11394
rect 14590 11342 14642 11394
rect 16158 11342 16210 11394
rect 18062 11342 18114 11394
rect 19630 11342 19682 11394
rect 22766 11342 22818 11394
rect 23438 11342 23490 11394
rect 24558 11342 24610 11394
rect 26126 11342 26178 11394
rect 27582 11342 27634 11394
rect 41246 11342 41298 11394
rect 41694 11342 41746 11394
rect 46510 11342 46562 11394
rect 46958 11342 47010 11394
rect 48190 11342 48242 11394
rect 49758 11342 49810 11394
rect 51326 11342 51378 11394
rect 52894 11342 52946 11394
rect 54462 11342 54514 11394
rect 54910 11342 54962 11394
rect 55246 11342 55298 11394
rect 1262 11230 1314 11282
rect 1934 11230 1986 11282
rect 2606 11230 2658 11282
rect 8878 11230 8930 11282
rect 9774 11230 9826 11282
rect 12350 11230 12402 11282
rect 15486 11230 15538 11282
rect 23102 11230 23154 11282
rect 23998 11230 24050 11282
rect 25118 11230 25170 11282
rect 28142 11230 28194 11282
rect 28366 11230 28418 11282
rect 32286 11230 32338 11282
rect 33854 11230 33906 11282
rect 34414 11230 34466 11282
rect 39006 11230 39058 11282
rect 45054 11230 45106 11282
rect 45726 11230 45778 11282
rect 47518 11230 47570 11282
rect 26574 11118 26626 11170
rect 35982 11118 36034 11170
rect 40910 11118 40962 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 3390 10782 3442 10834
rect 6414 10782 6466 10834
rect 7982 10782 8034 10834
rect 14814 10782 14866 10834
rect 41582 10782 41634 10834
rect 49646 10782 49698 10834
rect 50878 10782 50930 10834
rect 52558 10782 52610 10834
rect 2158 10670 2210 10722
rect 13806 10670 13858 10722
rect 16494 10670 16546 10722
rect 18286 10670 18338 10722
rect 19182 10670 19234 10722
rect 19518 10670 19570 10722
rect 20526 10670 20578 10722
rect 21870 10670 21922 10722
rect 25678 10670 25730 10722
rect 42702 10670 42754 10722
rect 46510 10670 46562 10722
rect 54574 10670 54626 10722
rect 56142 10670 56194 10722
rect 8990 10558 9042 10610
rect 9550 10558 9602 10610
rect 11678 10558 11730 10610
rect 17502 10558 17554 10610
rect 26238 10558 26290 10610
rect 29934 10558 29986 10610
rect 34526 10558 34578 10610
rect 34974 10558 35026 10610
rect 42366 10558 42418 10610
rect 47742 10558 47794 10610
rect 48750 10558 48802 10610
rect 52110 10558 52162 10610
rect 2830 10446 2882 10498
rect 4398 10446 4450 10498
rect 7422 10446 7474 10498
rect 9886 10446 9938 10498
rect 12126 10446 12178 10498
rect 14254 10446 14306 10498
rect 15822 10446 15874 10498
rect 17726 10446 17778 10498
rect 21086 10446 21138 10498
rect 26574 10446 26626 10498
rect 30382 10446 30434 10498
rect 40798 10446 40850 10498
rect 41246 10446 41298 10498
rect 42142 10446 42194 10498
rect 43038 10446 43090 10498
rect 47406 10446 47458 10498
rect 48302 10446 48354 10498
rect 51438 10446 51490 10498
rect 53566 10446 53618 10498
rect 55134 10446 55186 10498
rect 11118 10334 11170 10386
rect 12686 10334 12738 10386
rect 13134 10334 13186 10386
rect 13358 10334 13410 10386
rect 18622 10334 18674 10386
rect 18958 10334 19010 10386
rect 20078 10334 20130 10386
rect 24222 10334 24274 10386
rect 27806 10334 27858 10386
rect 29598 10334 29650 10386
rect 31614 10334 31666 10386
rect 34078 10334 34130 10386
rect 34414 10334 34466 10386
rect 40462 10334 40514 10386
rect 40686 10334 40738 10386
rect 46622 10334 46674 10386
rect 47070 10334 47122 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 17950 9998 18002 10050
rect 19406 9998 19458 10050
rect 26014 9998 26066 10050
rect 29710 9998 29762 10050
rect 30046 9998 30098 10050
rect 42142 9998 42194 10050
rect 47518 9998 47570 10050
rect 5294 9886 5346 9938
rect 9662 9886 9714 9938
rect 18846 9886 18898 9938
rect 21534 9886 21586 9938
rect 22094 9886 22146 9938
rect 23998 9886 24050 9938
rect 24446 9886 24498 9938
rect 27582 9886 27634 9938
rect 42590 9886 42642 9938
rect 46958 9886 47010 9938
rect 48190 9886 48242 9938
rect 48526 9886 48578 9938
rect 49086 9886 49138 9938
rect 50206 9886 50258 9938
rect 3054 9774 3106 9826
rect 7534 9774 7586 9826
rect 10446 9774 10498 9826
rect 12014 9774 12066 9826
rect 13022 9774 13074 9826
rect 15038 9774 15090 9826
rect 17390 9774 17442 9826
rect 18286 9774 18338 9826
rect 20302 9774 20354 9826
rect 21086 9774 21138 9826
rect 27806 9774 27858 9826
rect 46398 9774 46450 9826
rect 49422 9774 49474 9826
rect 50990 9774 51042 9826
rect 52558 9774 52610 9826
rect 54126 9774 54178 9826
rect 2046 9662 2098 9714
rect 4286 9662 4338 9714
rect 6526 9662 6578 9714
rect 8878 9662 8930 9714
rect 11006 9662 11058 9714
rect 12574 9662 12626 9714
rect 13358 9662 13410 9714
rect 14142 9662 14194 9714
rect 19182 9662 19234 9714
rect 20526 9662 20578 9714
rect 22318 9662 22370 9714
rect 23550 9662 23602 9714
rect 26350 9662 26402 9714
rect 30606 9662 30658 9714
rect 46062 9662 46114 9714
rect 53454 9662 53506 9714
rect 26686 9550 26738 9602
rect 27022 9550 27074 9602
rect 42478 9550 42530 9602
rect 51998 9550 52050 9602
rect 55134 9550 55186 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 2046 9214 2098 9266
rect 11342 9214 11394 9266
rect 31726 9214 31778 9266
rect 51214 9214 51266 9266
rect 53006 9214 53058 9266
rect 12910 9102 12962 9154
rect 18062 9102 18114 9154
rect 18846 9102 18898 9154
rect 20974 9102 21026 9154
rect 24558 9102 24610 9154
rect 24782 9102 24834 9154
rect 25230 9102 25282 9154
rect 28814 9102 28866 9154
rect 30718 9102 30770 9154
rect 30942 9102 30994 9154
rect 33406 9102 33458 9154
rect 35758 9102 35810 9154
rect 38110 9102 38162 9154
rect 48078 9102 48130 9154
rect 48974 9102 49026 9154
rect 11902 8990 11954 9042
rect 18622 8990 18674 9042
rect 21310 8990 21362 9042
rect 21758 8990 21810 9042
rect 22654 8990 22706 9042
rect 23214 8990 23266 9042
rect 24110 8990 24162 9042
rect 25006 8990 25058 9042
rect 26686 8990 26738 9042
rect 36318 8990 36370 9042
rect 38558 8990 38610 9042
rect 39454 8990 39506 9042
rect 39902 8990 39954 9042
rect 40014 8990 40066 9042
rect 41806 8990 41858 9042
rect 42254 8990 42306 9042
rect 43150 8990 43202 9042
rect 46062 8990 46114 9042
rect 48414 8990 48466 9042
rect 52110 8990 52162 9042
rect 53678 8990 53730 9042
rect 2606 8878 2658 8930
rect 5518 8878 5570 8930
rect 10446 8878 10498 8930
rect 12126 8878 12178 8930
rect 27246 8878 27298 8930
rect 31950 8878 32002 8930
rect 32286 8878 32338 8930
rect 33742 8878 33794 8930
rect 39678 8878 39730 8930
rect 40686 8878 40738 8930
rect 41470 8878 41522 8930
rect 42478 8878 42530 8930
rect 49870 8878 49922 8930
rect 50206 8878 50258 8930
rect 54350 8878 54402 8930
rect 55134 8878 55186 8930
rect 55918 8878 55970 8930
rect 4510 8766 4562 8818
rect 4958 8766 5010 8818
rect 9662 8766 9714 8818
rect 9886 8766 9938 8818
rect 11006 8766 11058 8818
rect 13470 8766 13522 8818
rect 13806 8766 13858 8818
rect 13918 8766 13970 8818
rect 21982 8766 22034 8818
rect 31390 8766 31442 8818
rect 32846 8766 32898 8818
rect 34974 8766 35026 8818
rect 36878 8766 36930 8818
rect 37774 8766 37826 8818
rect 40798 8766 40850 8818
rect 42030 8766 42082 8818
rect 45278 8766 45330 8818
rect 45502 8766 45554 8818
rect 49310 8766 49362 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 12462 8430 12514 8482
rect 28590 8430 28642 8482
rect 33294 8430 33346 8482
rect 33518 8430 33570 8482
rect 39006 8430 39058 8482
rect 41918 8430 41970 8482
rect 49086 8430 49138 8482
rect 13470 8318 13522 8370
rect 13918 8318 13970 8370
rect 14926 8318 14978 8370
rect 18398 8318 18450 8370
rect 18510 8318 18562 8370
rect 28030 8318 28082 8370
rect 28926 8318 28978 8370
rect 29710 8318 29762 8370
rect 35086 8318 35138 8370
rect 35758 8318 35810 8370
rect 36094 8318 36146 8370
rect 36654 8318 36706 8370
rect 37998 8318 38050 8370
rect 38446 8318 38498 8370
rect 41134 8318 41186 8370
rect 41582 8318 41634 8370
rect 42142 8318 42194 8370
rect 42254 8318 42306 8370
rect 50318 8318 50370 8370
rect 51774 8318 51826 8370
rect 53342 8318 53394 8370
rect 2270 8206 2322 8258
rect 7758 8206 7810 8258
rect 14366 8206 14418 8258
rect 18734 8206 18786 8258
rect 19070 8206 19122 8258
rect 29374 8206 29426 8258
rect 31614 8206 31666 8258
rect 37438 8206 37490 8258
rect 38670 8206 38722 8258
rect 40798 8206 40850 8258
rect 41022 8206 41074 8258
rect 41358 8206 41410 8258
rect 49758 8206 49810 8258
rect 50990 8206 51042 8258
rect 52558 8206 52610 8258
rect 54126 8206 54178 8258
rect 1262 8094 1314 8146
rect 7422 8094 7474 8146
rect 8206 8094 8258 8146
rect 15150 8094 15202 8146
rect 31166 8094 31218 8146
rect 34078 8094 34130 8146
rect 34638 8094 34690 8146
rect 37214 8094 37266 8146
rect 49422 8094 49474 8146
rect 50542 8094 50594 8146
rect 55134 8094 55186 8146
rect 12798 7982 12850 8034
rect 13134 7982 13186 8034
rect 18958 7982 19010 8034
rect 36318 7982 36370 8034
rect 41694 7982 41746 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 19966 7646 20018 7698
rect 28926 7646 28978 7698
rect 53006 7646 53058 7698
rect 56142 7646 56194 7698
rect 7758 7534 7810 7586
rect 8318 7534 8370 7586
rect 14030 7534 14082 7586
rect 14702 7534 14754 7586
rect 16158 7534 16210 7586
rect 19742 7534 19794 7586
rect 30046 7534 30098 7586
rect 30382 7534 30434 7586
rect 34302 7534 34354 7586
rect 34974 7534 35026 7586
rect 35198 7534 35250 7586
rect 35422 7534 35474 7586
rect 35646 7534 35698 7586
rect 35870 7534 35922 7586
rect 49646 7534 49698 7586
rect 54574 7534 54626 7586
rect 12238 7422 12290 7474
rect 13582 7422 13634 7474
rect 14478 7422 14530 7474
rect 18622 7422 18674 7474
rect 18958 7422 19010 7474
rect 19630 7422 19682 7474
rect 36654 7422 36706 7474
rect 37102 7422 37154 7474
rect 38558 7422 38610 7474
rect 39342 7422 39394 7474
rect 49982 7422 50034 7474
rect 50542 7422 50594 7474
rect 50878 7422 50930 7474
rect 55134 7422 55186 7474
rect 8654 7310 8706 7362
rect 16494 7310 16546 7362
rect 17726 7310 17778 7362
rect 18286 7310 18338 7362
rect 19294 7310 19346 7362
rect 29150 7310 29202 7362
rect 29710 7310 29762 7362
rect 36318 7310 36370 7362
rect 37774 7310 37826 7362
rect 42590 7310 42642 7362
rect 51438 7310 51490 7362
rect 51998 7310 52050 7362
rect 53566 7310 53618 7362
rect 9886 7198 9938 7250
rect 11902 7198 11954 7250
rect 12126 7198 12178 7250
rect 14366 7198 14418 7250
rect 15598 7198 15650 7250
rect 18398 7198 18450 7250
rect 18846 7198 18898 7250
rect 28590 7198 28642 7250
rect 37326 7198 37378 7250
rect 42030 7198 42082 7250
rect 42254 7198 42306 7250
rect 43150 7198 43202 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 18622 6862 18674 6914
rect 20750 6862 20802 6914
rect 22878 6862 22930 6914
rect 23998 6862 24050 6914
rect 16718 6750 16770 6802
rect 18734 6750 18786 6802
rect 21646 6750 21698 6802
rect 25230 6750 25282 6802
rect 41806 6750 41858 6802
rect 42030 6750 42082 6802
rect 42254 6750 42306 6802
rect 43374 6750 43426 6802
rect 43710 6750 43762 6802
rect 10558 6638 10610 6690
rect 11006 6638 11058 6690
rect 11118 6638 11170 6690
rect 11230 6638 11282 6690
rect 11566 6638 11618 6690
rect 11790 6638 11842 6690
rect 12126 6638 12178 6690
rect 12350 6638 12402 6690
rect 18286 6638 18338 6690
rect 18846 6638 18898 6690
rect 24782 6638 24834 6690
rect 31838 6638 31890 6690
rect 36094 6638 36146 6690
rect 40686 6638 40738 6690
rect 42814 6638 42866 6690
rect 45614 6638 45666 6690
rect 45838 6638 45890 6690
rect 50206 6638 50258 6690
rect 50542 6638 50594 6690
rect 51102 6638 51154 6690
rect 51438 6638 51490 6690
rect 52670 6638 52722 6690
rect 54238 6638 54290 6690
rect 12014 6526 12066 6578
rect 16270 6526 16322 6578
rect 17278 6526 17330 6578
rect 21310 6526 21362 6578
rect 31278 6526 31330 6578
rect 40462 6526 40514 6578
rect 46286 6526 46338 6578
rect 51886 6526 51938 6578
rect 53230 6526 53282 6578
rect 10670 6414 10722 6466
rect 26350 6414 26402 6466
rect 41134 6414 41186 6466
rect 41470 6414 41522 6466
rect 43150 6414 43202 6466
rect 55134 6414 55186 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 9438 6078 9490 6130
rect 11566 6078 11618 6130
rect 27022 6078 27074 6130
rect 32622 6078 32674 6130
rect 32958 6078 33010 6130
rect 37326 6078 37378 6130
rect 53006 6078 53058 6130
rect 56142 6078 56194 6130
rect 6414 5966 6466 6018
rect 7870 5966 7922 6018
rect 21310 5966 21362 6018
rect 22206 5966 22258 6018
rect 24334 5966 24386 6018
rect 25118 5966 25170 6018
rect 28590 5966 28642 6018
rect 29262 5966 29314 6018
rect 38558 5966 38610 6018
rect 41470 5966 41522 6018
rect 41806 5966 41858 6018
rect 42702 5966 42754 6018
rect 48638 5966 48690 6018
rect 54574 5966 54626 6018
rect 6750 5854 6802 5906
rect 21646 5854 21698 5906
rect 24670 5854 24722 5906
rect 26238 5854 26290 5906
rect 30382 5854 30434 5906
rect 38446 5854 38498 5906
rect 38782 5854 38834 5906
rect 39230 5854 39282 5906
rect 39566 5854 39618 5906
rect 42254 5854 42306 5906
rect 48974 5854 49026 5906
rect 52110 5854 52162 5906
rect 53566 5854 53618 5906
rect 7310 5742 7362 5794
rect 8318 5742 8370 5794
rect 11678 5742 11730 5794
rect 25678 5742 25730 5794
rect 27246 5742 27298 5794
rect 27694 5742 27746 5794
rect 29038 5742 29090 5794
rect 30830 5742 30882 5794
rect 32062 5742 32114 5794
rect 33182 5742 33234 5794
rect 33630 5742 33682 5794
rect 37214 5742 37266 5794
rect 38110 5742 38162 5794
rect 39454 5742 39506 5794
rect 49534 5742 49586 5794
rect 55134 5742 55186 5794
rect 26686 5630 26738 5682
rect 29934 5630 29986 5682
rect 37102 5630 37154 5682
rect 51102 5630 51154 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 7422 5294 7474 5346
rect 12014 5294 12066 5346
rect 15934 5294 15986 5346
rect 16606 5294 16658 5346
rect 23774 5294 23826 5346
rect 26574 5294 26626 5346
rect 28254 5294 28306 5346
rect 28478 5294 28530 5346
rect 30718 5294 30770 5346
rect 30942 5294 30994 5346
rect 31838 5294 31890 5346
rect 32286 5294 32338 5346
rect 35758 5294 35810 5346
rect 39454 5294 39506 5346
rect 53006 5294 53058 5346
rect 53230 5294 53282 5346
rect 12462 5182 12514 5234
rect 13470 5182 13522 5234
rect 13918 5182 13970 5234
rect 22990 5182 23042 5234
rect 23214 5182 23266 5234
rect 23438 5182 23490 5234
rect 31502 5182 31554 5234
rect 33630 5182 33682 5234
rect 34526 5182 34578 5234
rect 38670 5182 38722 5234
rect 39678 5182 39730 5234
rect 54126 5182 54178 5234
rect 11790 5070 11842 5122
rect 12910 5070 12962 5122
rect 13358 5070 13410 5122
rect 14702 5070 14754 5122
rect 15486 5070 15538 5122
rect 20974 5070 21026 5122
rect 21310 5070 21362 5122
rect 21870 5070 21922 5122
rect 22318 5070 22370 5122
rect 38782 5070 38834 5122
rect 39118 5070 39170 5122
rect 39454 5070 39506 5122
rect 51662 5070 51714 5122
rect 51998 5070 52050 5122
rect 54910 5070 54962 5122
rect 12126 4958 12178 5010
rect 16158 4958 16210 5010
rect 22654 4958 22706 5010
rect 34190 4958 34242 5010
rect 52446 4958 52498 5010
rect 53678 4958 53730 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 10894 4510 10946 4562
rect 17950 4510 18002 4562
rect 18286 4510 18338 4562
rect 22990 4510 23042 4562
rect 39454 4510 39506 4562
rect 54574 4510 54626 4562
rect 56142 4510 56194 4562
rect 8766 4398 8818 4450
rect 9326 4398 9378 4450
rect 11790 4398 11842 4450
rect 12686 4398 12738 4450
rect 13470 4398 13522 4450
rect 14254 4398 14306 4450
rect 16046 4398 16098 4450
rect 16158 4398 16210 4450
rect 19406 4398 19458 4450
rect 19630 4398 19682 4450
rect 20862 4398 20914 4450
rect 21422 4398 21474 4450
rect 34078 4398 34130 4450
rect 44158 4398 44210 4450
rect 44942 4398 44994 4450
rect 49534 4398 49586 4450
rect 50318 4398 50370 4450
rect 52334 4398 52386 4450
rect 12238 4286 12290 4338
rect 14030 4286 14082 4338
rect 19070 4286 19122 4338
rect 21310 4286 21362 4338
rect 27582 4286 27634 4338
rect 28478 4286 28530 4338
rect 34526 4286 34578 4338
rect 39566 4286 39618 4338
rect 44494 4286 44546 4338
rect 49870 4286 49922 4338
rect 52670 4286 52722 4338
rect 55134 4286 55186 4338
rect 9774 4174 9826 4226
rect 15150 4174 15202 4226
rect 15710 4174 15762 4226
rect 18846 4174 18898 4226
rect 21758 4174 21810 4226
rect 27022 4174 27074 4226
rect 27246 4174 27298 4226
rect 34974 4174 35026 4226
rect 53230 4174 53282 4226
rect 53566 4174 53618 4226
rect 27470 4062 27522 4114
rect 28590 4062 28642 4114
rect 28814 4062 28866 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 9102 3726 9154 3778
rect 9326 3726 9378 3778
rect 18510 3726 18562 3778
rect 18846 3726 18898 3778
rect 19966 3726 20018 3778
rect 26910 3726 26962 3778
rect 27246 3726 27298 3778
rect 32398 3726 32450 3778
rect 35198 3726 35250 3778
rect 51438 3726 51490 3778
rect 51662 3726 51714 3778
rect 17950 3614 18002 3666
rect 19070 3614 19122 3666
rect 27358 3614 27410 3666
rect 28702 3614 28754 3666
rect 29710 3614 29762 3666
rect 36094 3614 36146 3666
rect 52222 3614 52274 3666
rect 52558 3614 52610 3666
rect 54910 3614 54962 3666
rect 19518 3502 19570 3554
rect 26798 3502 26850 3554
rect 28926 3502 28978 3554
rect 29262 3502 29314 3554
rect 35646 3502 35698 3554
rect 54126 3502 54178 3554
rect 9886 3390 9938 3442
rect 28814 3390 28866 3442
rect 29598 3390 29650 3442
rect 53566 3390 53618 3442
rect 29934 3278 29986 3330
rect 37326 3278 37378 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 26910 2942 26962 2994
rect 38222 2942 38274 2994
rect 54574 2942 54626 2994
rect 56142 2942 56194 2994
rect 21198 2830 21250 2882
rect 24782 2830 24834 2882
rect 28366 2830 28418 2882
rect 28702 2830 28754 2882
rect 28926 2830 28978 2882
rect 33294 2830 33346 2882
rect 34862 2830 34914 2882
rect 35646 2830 35698 2882
rect 40574 2830 40626 2882
rect 41582 2830 41634 2882
rect 48414 2830 48466 2882
rect 50542 2830 50594 2882
rect 21534 2718 21586 2770
rect 25230 2718 25282 2770
rect 29262 2718 29314 2770
rect 29710 2718 29762 2770
rect 30382 2718 30434 2770
rect 30942 2718 30994 2770
rect 32062 2718 32114 2770
rect 32510 2718 32562 2770
rect 35198 2718 35250 2770
rect 36542 2718 36594 2770
rect 50878 2718 50930 2770
rect 52110 2718 52162 2770
rect 53566 2718 53618 2770
rect 55134 2718 55186 2770
rect 22094 2606 22146 2658
rect 25678 2606 25730 2658
rect 29934 2606 29986 2658
rect 33070 2606 33122 2658
rect 36990 2606 37042 2658
rect 51438 2606 51490 2658
rect 52782 2606 52834 2658
rect 39790 2494 39842 2546
rect 40014 2494 40066 2546
rect 42142 2494 42194 2546
rect 42478 2494 42530 2546
rect 47630 2494 47682 2546
rect 47854 2494 47906 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 23102 2158 23154 2210
rect 23438 2158 23490 2210
rect 26350 2158 26402 2210
rect 28702 2158 28754 2210
rect 29038 2158 29090 2210
rect 30158 2158 30210 2210
rect 30494 2158 30546 2210
rect 32398 2158 32450 2210
rect 36206 2158 36258 2210
rect 36430 2158 36482 2210
rect 36654 2158 36706 2210
rect 40910 2158 40962 2210
rect 41134 2158 41186 2210
rect 49086 2158 49138 2210
rect 12910 2046 12962 2098
rect 25118 2046 25170 2098
rect 41694 2046 41746 2098
rect 47518 2046 47570 2098
rect 50430 2046 50482 2098
rect 51326 2046 51378 2098
rect 52222 2046 52274 2098
rect 52558 2046 52610 2098
rect 54126 2046 54178 2098
rect 54910 2046 54962 2098
rect 24782 1934 24834 1986
rect 28142 1934 28194 1986
rect 38446 1934 38498 1986
rect 46958 1934 47010 1986
rect 49310 1934 49362 1986
rect 49870 1934 49922 1986
rect 50766 1934 50818 1986
rect 51662 1934 51714 1986
rect 23998 1822 24050 1874
rect 29598 1822 29650 1874
rect 37214 1822 37266 1874
rect 37998 1822 38050 1874
rect 38670 1822 38722 1874
rect 46734 1822 46786 1874
rect 48750 1822 48802 1874
rect 53566 1822 53618 1874
rect 11902 1710 11954 1762
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 53566 1374 53618 1426
rect 56142 1374 56194 1426
rect 5518 1262 5570 1314
rect 7422 1262 7474 1314
rect 9886 1262 9938 1314
rect 13918 1262 13970 1314
rect 24334 1262 24386 1314
rect 25230 1262 25282 1314
rect 26126 1262 26178 1314
rect 50430 1262 50482 1314
rect 50654 1262 50706 1314
rect 51998 1262 52050 1314
rect 6526 1150 6578 1202
rect 8094 1150 8146 1202
rect 10894 1150 10946 1202
rect 14814 1150 14866 1202
rect 25678 1150 25730 1202
rect 50990 1150 51042 1202
rect 52558 1150 52610 1202
rect 55134 1038 55186 1090
rect 49534 926 49586 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 672 14112 784 14224
rect 1120 14112 1232 14224
rect 1568 14112 1680 14224
rect 2016 14112 2128 14224
rect 2464 14112 2576 14224
rect 2912 14112 3024 14224
rect 3360 14112 3472 14224
rect 3808 14112 3920 14224
rect 4256 14112 4368 14224
rect 4704 14112 4816 14224
rect 5152 14112 5264 14224
rect 5600 14112 5712 14224
rect 6048 14112 6160 14224
rect 6496 14112 6608 14224
rect 6944 14112 7056 14224
rect 7392 14112 7504 14224
rect 7840 14112 7952 14224
rect 8288 14112 8400 14224
rect 8736 14112 8848 14224
rect 9184 14112 9296 14224
rect 9632 14112 9744 14224
rect 10080 14112 10192 14224
rect 10528 14112 10640 14224
rect 10976 14112 11088 14224
rect 11424 14112 11536 14224
rect 11872 14112 11984 14224
rect 12320 14112 12432 14224
rect 12768 14112 12880 14224
rect 13216 14112 13328 14224
rect 13664 14112 13776 14224
rect 14112 14112 14224 14224
rect 14560 14112 14672 14224
rect 15008 14112 15120 14224
rect 15456 14112 15568 14224
rect 15904 14112 16016 14224
rect 16352 14112 16464 14224
rect 16800 14112 16912 14224
rect 17052 14196 17108 14206
rect 476 13972 532 13982
rect 140 13524 196 13534
rect 140 9268 196 13468
rect 364 12628 420 12638
rect 140 9202 196 9212
rect 252 11284 308 11294
rect 252 6468 308 11228
rect 252 6402 308 6412
rect 364 4900 420 12572
rect 476 11172 532 13916
rect 588 12180 644 12190
rect 588 11396 644 12124
rect 588 11330 644 11340
rect 700 11284 756 14112
rect 1148 11844 1204 14112
rect 1148 11778 1204 11788
rect 1484 13076 1540 13086
rect 1484 11620 1540 13020
rect 1596 11956 1652 14112
rect 1932 12068 1988 12078
rect 1596 11900 1764 11956
rect 1484 11554 1540 11564
rect 1484 11394 1540 11406
rect 1484 11342 1486 11394
rect 1538 11342 1540 11394
rect 1260 11284 1316 11294
rect 1484 11284 1540 11342
rect 700 11228 1204 11284
rect 476 11106 532 11116
rect 1036 9940 1092 9950
rect 1036 7700 1092 9884
rect 1148 8428 1204 11228
rect 1260 11282 1540 11284
rect 1260 11230 1262 11282
rect 1314 11230 1540 11282
rect 1260 11228 1540 11230
rect 1260 11218 1316 11228
rect 1372 10388 1428 10398
rect 1148 8372 1316 8428
rect 1260 8146 1316 8372
rect 1260 8094 1262 8146
rect 1314 8094 1316 8146
rect 1260 8082 1316 8094
rect 1036 7644 1204 7700
rect 1036 7476 1092 7486
rect 1036 6356 1092 7420
rect 1148 6580 1204 7644
rect 1148 6514 1204 6524
rect 1036 6290 1092 6300
rect 1372 6020 1428 10332
rect 1484 7588 1540 11228
rect 1708 9716 1764 11900
rect 1932 11282 1988 12012
rect 2044 11620 2100 14112
rect 2268 13636 2324 13646
rect 2156 13300 2212 13310
rect 2156 13186 2212 13244
rect 2156 13134 2158 13186
rect 2210 13134 2212 13186
rect 2156 13122 2212 13134
rect 2268 12402 2324 13580
rect 2268 12350 2270 12402
rect 2322 12350 2324 12402
rect 2268 12338 2324 12350
rect 2268 11844 2324 11854
rect 2044 11564 2212 11620
rect 1932 11230 1934 11282
rect 1986 11230 1988 11282
rect 1932 11218 1988 11230
rect 2156 10722 2212 11564
rect 2156 10670 2158 10722
rect 2210 10670 2212 10722
rect 2156 10658 2212 10670
rect 2044 9716 2100 9726
rect 1708 9714 2100 9716
rect 1708 9662 2046 9714
rect 2098 9662 2100 9714
rect 1708 9660 2100 9662
rect 2044 9650 2100 9660
rect 1932 9492 1988 9502
rect 2268 9492 2324 11788
rect 2492 11284 2548 14112
rect 2716 12962 2772 12974
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2604 11284 2660 11294
rect 2492 11282 2660 11284
rect 2492 11230 2606 11282
rect 2658 11230 2660 11282
rect 2492 11228 2660 11230
rect 2604 11218 2660 11228
rect 2716 9716 2772 12910
rect 2828 12404 2884 12414
rect 2828 12178 2884 12348
rect 2940 12292 2996 14112
rect 3388 13636 3444 14112
rect 3388 13570 3444 13580
rect 3612 13524 3668 13534
rect 2940 12236 3444 12292
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 2828 12114 2884 12126
rect 2940 11620 2996 11630
rect 2716 9650 2772 9660
rect 2828 10498 2884 10510
rect 2828 10446 2830 10498
rect 2882 10446 2884 10498
rect 1484 7522 1540 7532
rect 1596 9268 1652 9278
rect 1596 7252 1652 9212
rect 1596 7186 1652 7196
rect 1708 8820 1764 8830
rect 1372 5954 1428 5964
rect 1148 5908 1204 5918
rect 364 4834 420 4844
rect 924 5012 980 5022
rect 924 644 980 4956
rect 1148 2884 1204 5852
rect 1708 5124 1764 8764
rect 1932 6916 1988 9436
rect 2044 9436 2324 9492
rect 2044 9266 2100 9436
rect 2044 9214 2046 9266
rect 2098 9214 2100 9266
rect 2044 9202 2100 9214
rect 2604 8930 2660 8942
rect 2604 8878 2606 8930
rect 2658 8878 2660 8930
rect 2604 8484 2660 8878
rect 2604 8418 2660 8428
rect 1932 6850 1988 6860
rect 2268 8258 2324 8270
rect 2268 8206 2270 8258
rect 2322 8206 2324 8258
rect 2268 5236 2324 8206
rect 2828 5796 2884 10446
rect 2940 7252 2996 11564
rect 3388 10834 3444 12236
rect 3612 12290 3668 13468
rect 3724 13188 3780 13198
rect 3724 13094 3780 13132
rect 3836 12740 3892 14112
rect 4284 13300 4340 14112
rect 4732 13524 4788 14112
rect 4732 13458 4788 13468
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4284 13234 4340 13244
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 3836 12684 4340 12740
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 3612 12238 3614 12290
rect 3666 12238 3668 12290
rect 3612 12226 3668 12238
rect 4172 12178 4228 12190
rect 4172 12126 4174 12178
rect 4226 12126 4228 12178
rect 3388 10782 3390 10834
rect 3442 10782 3444 10834
rect 3388 10770 3444 10782
rect 3612 11394 3668 11406
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3276 10500 3332 10510
rect 2940 7186 2996 7196
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 2828 5730 2884 5740
rect 2268 5170 2324 5180
rect 1148 2818 1204 2828
rect 1484 5068 1764 5124
rect 924 578 980 588
rect 1372 1428 1428 1438
rect 1372 112 1428 1372
rect 1484 980 1540 5068
rect 1596 4452 1652 4462
rect 1596 2772 1652 4396
rect 1596 2706 1652 2716
rect 1484 914 1540 924
rect 3052 980 3108 9774
rect 3276 9044 3332 10444
rect 3276 8978 3332 8988
rect 3276 8596 3332 8606
rect 3276 4900 3332 8540
rect 3276 4834 3332 4844
rect 3276 4116 3332 4126
rect 3276 2324 3332 4060
rect 3612 3668 3668 11342
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4172 8932 4228 12126
rect 4284 9714 4340 12684
rect 5068 12290 5124 12302
rect 5068 12238 5070 12290
rect 5122 12238 5124 12290
rect 5068 12180 5124 12238
rect 5068 12114 5124 12124
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4620 11620 4676 11630
rect 4620 11526 4676 11564
rect 5180 11620 5236 14112
rect 5628 13188 5684 14112
rect 5628 13122 5684 13132
rect 5964 13188 6020 13198
rect 5964 13094 6020 13132
rect 6076 13076 6132 14112
rect 6524 13188 6580 14112
rect 6076 13010 6132 13020
rect 6412 13132 6580 13188
rect 5852 12964 5908 12974
rect 5516 11956 5572 11966
rect 5740 11956 5796 11966
rect 5516 11954 5796 11956
rect 5516 11902 5518 11954
rect 5570 11902 5742 11954
rect 5794 11902 5796 11954
rect 5516 11900 5796 11902
rect 5516 11890 5572 11900
rect 5740 11844 5796 11900
rect 5740 11778 5796 11788
rect 5180 11554 5236 11564
rect 5180 11394 5236 11406
rect 5180 11342 5182 11394
rect 5234 11342 5236 11394
rect 4956 10836 5012 10846
rect 4396 10498 4452 10510
rect 4396 10446 4398 10498
rect 4450 10446 4452 10498
rect 4396 10388 4452 10446
rect 4396 10322 4452 10332
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4956 10052 5012 10780
rect 4956 9986 5012 9996
rect 4284 9662 4286 9714
rect 4338 9662 4340 9714
rect 4284 9650 4340 9662
rect 4172 8866 4228 8876
rect 4508 8820 4564 8858
rect 4508 8754 4564 8764
rect 4956 8820 5012 8830
rect 4956 8726 5012 8764
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 5180 7364 5236 11342
rect 5292 10836 5348 10846
rect 5292 9938 5348 10780
rect 5292 9886 5294 9938
rect 5346 9886 5348 9938
rect 5292 9874 5348 9886
rect 5516 8930 5572 8942
rect 5516 8878 5518 8930
rect 5570 8878 5572 8930
rect 5180 7308 5348 7364
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4956 5236 5012 5246
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 3612 3602 3668 3612
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 3276 2258 3332 2268
rect 4956 2212 5012 5180
rect 5180 4340 5236 4350
rect 4956 2146 5012 2156
rect 5068 4228 5124 4238
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 3052 914 3108 924
rect 3388 1316 3444 1326
rect 3388 112 3444 1260
rect 5068 868 5124 4172
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 5068 802 5124 812
rect 4464 746 4728 756
rect 5180 532 5236 4284
rect 5292 2660 5348 7308
rect 5292 2594 5348 2604
rect 5516 1540 5572 8878
rect 5852 4788 5908 12908
rect 6300 12962 6356 12974
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6188 11620 6244 11630
rect 6188 11526 6244 11564
rect 6300 8260 6356 12910
rect 6412 10834 6468 13132
rect 6412 10782 6414 10834
rect 6466 10782 6468 10834
rect 6412 10770 6468 10782
rect 6524 12964 6580 12974
rect 6524 9714 6580 12908
rect 6972 12740 7028 14112
rect 7420 13188 7476 14112
rect 7420 13122 7476 13132
rect 7532 13300 7588 13310
rect 7532 13186 7588 13244
rect 7532 13134 7534 13186
rect 7586 13134 7588 13186
rect 7532 13122 7588 13134
rect 6860 12684 7028 12740
rect 6860 11620 6916 12684
rect 6972 12404 7028 12414
rect 6972 12310 7028 12348
rect 7532 12068 7588 12078
rect 7532 12066 7700 12068
rect 7532 12014 7534 12066
rect 7586 12014 7700 12066
rect 7532 12012 7700 12014
rect 7532 12002 7588 12012
rect 6860 11554 6916 11564
rect 6524 9662 6526 9714
rect 6578 9662 6580 9714
rect 6524 9650 6580 9662
rect 6636 11394 6692 11406
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6300 8194 6356 8204
rect 5852 4722 5908 4732
rect 6076 7140 6132 7150
rect 6076 3388 6132 7084
rect 6524 6132 6580 6142
rect 6412 6020 6468 6030
rect 6412 5926 6468 5964
rect 5964 3332 6132 3388
rect 5516 1474 5572 1484
rect 5628 2884 5684 2894
rect 5516 1316 5572 1326
rect 5180 466 5236 476
rect 5404 1314 5572 1316
rect 5404 1262 5518 1314
rect 5570 1262 5572 1314
rect 5404 1260 5572 1262
rect 5404 112 5460 1260
rect 5516 1250 5572 1260
rect 5628 756 5684 2828
rect 5964 1316 6020 3332
rect 5964 1250 6020 1260
rect 6524 1202 6580 6076
rect 6636 2100 6692 11342
rect 7420 10498 7476 10510
rect 7420 10446 7422 10498
rect 7474 10446 7476 10498
rect 7420 10276 7476 10446
rect 7420 10210 7476 10220
rect 7532 9826 7588 9838
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 7308 9604 7364 9614
rect 6860 7476 6916 7486
rect 6860 6804 6916 7420
rect 7308 7364 7364 9548
rect 7420 8148 7476 8158
rect 7420 8054 7476 8092
rect 7308 7298 7364 7308
rect 6860 6738 6916 6748
rect 6748 6020 6804 6030
rect 6748 5906 6804 5964
rect 7420 6020 7476 6030
rect 6748 5854 6750 5906
rect 6802 5854 6804 5906
rect 6748 5842 6804 5854
rect 6972 5908 7028 5918
rect 6860 5236 6916 5246
rect 6748 3892 6804 3902
rect 6748 3332 6804 3836
rect 6748 3266 6804 3276
rect 6636 2034 6692 2044
rect 6860 1428 6916 5180
rect 6972 1764 7028 5852
rect 7308 5794 7364 5806
rect 7308 5742 7310 5794
rect 7362 5742 7364 5794
rect 7308 2772 7364 5742
rect 7420 5346 7476 5964
rect 7420 5294 7422 5346
rect 7474 5294 7476 5346
rect 7420 5282 7476 5294
rect 7308 2706 7364 2716
rect 7532 2436 7588 9774
rect 7644 8932 7700 12012
rect 7756 11620 7812 11630
rect 7756 11526 7812 11564
rect 7868 10836 7924 14112
rect 8204 13076 8260 13086
rect 8092 12962 8148 12974
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 8092 11620 8148 12910
rect 8204 12290 8260 13020
rect 8316 12404 8372 14112
rect 8764 12740 8820 14112
rect 9212 12964 9268 14112
rect 9660 13300 9716 14112
rect 9660 13234 9716 13244
rect 9772 13972 9828 13982
rect 9772 13186 9828 13916
rect 9772 13134 9774 13186
rect 9826 13134 9828 13186
rect 9772 13122 9828 13134
rect 10108 13076 10164 14112
rect 10108 13010 10164 13020
rect 9212 12908 9716 12964
rect 9324 12740 9380 12750
rect 8764 12684 9044 12740
rect 8316 12338 8372 12348
rect 8204 12238 8206 12290
rect 8258 12238 8260 12290
rect 8204 12226 8260 12238
rect 8876 12180 8932 12190
rect 8540 12178 8932 12180
rect 8540 12126 8878 12178
rect 8930 12126 8932 12178
rect 8540 12124 8932 12126
rect 8428 11956 8484 11966
rect 8092 11564 8260 11620
rect 8092 11394 8148 11406
rect 8092 11342 8094 11394
rect 8146 11342 8148 11394
rect 7980 10836 8036 10846
rect 7868 10834 8036 10836
rect 7868 10782 7982 10834
rect 8034 10782 8036 10834
rect 7868 10780 8036 10782
rect 7980 10770 8036 10780
rect 7644 8866 7700 8876
rect 7756 8258 7812 8270
rect 7756 8206 7758 8258
rect 7810 8206 7812 8258
rect 7756 8148 7812 8206
rect 7756 7586 7812 8092
rect 7756 7534 7758 7586
rect 7810 7534 7812 7586
rect 7756 7364 7812 7534
rect 7756 7298 7812 7308
rect 7980 7588 8036 7598
rect 7980 6580 8036 7532
rect 7980 6514 8036 6524
rect 7868 6244 7924 6254
rect 7868 6018 7924 6188
rect 7868 5966 7870 6018
rect 7922 5966 7924 6018
rect 7868 5954 7924 5966
rect 7532 2370 7588 2380
rect 8092 1988 8148 11342
rect 8204 8372 8260 11564
rect 8316 10052 8372 10062
rect 8428 10052 8484 11900
rect 8372 9996 8484 10052
rect 8316 9986 8372 9996
rect 8204 8316 8372 8372
rect 8204 8146 8260 8158
rect 8204 8094 8206 8146
rect 8258 8094 8260 8146
rect 8204 2884 8260 8094
rect 8316 7924 8372 8316
rect 8316 7858 8372 7868
rect 8428 8036 8484 8046
rect 8316 7588 8372 7598
rect 8428 7588 8484 7980
rect 8316 7586 8484 7588
rect 8316 7534 8318 7586
rect 8370 7534 8484 7586
rect 8316 7532 8484 7534
rect 8316 6244 8372 7532
rect 8316 6178 8372 6188
rect 8316 6020 8372 6030
rect 8316 5794 8372 5964
rect 8316 5742 8318 5794
rect 8370 5742 8372 5794
rect 8316 5730 8372 5742
rect 8204 2818 8260 2828
rect 8428 3556 8484 3566
rect 8092 1922 8148 1932
rect 6972 1698 7028 1708
rect 6860 1362 6916 1372
rect 6524 1150 6526 1202
rect 6578 1150 6580 1202
rect 6524 1138 6580 1150
rect 7420 1314 7476 1326
rect 7420 1262 7422 1314
rect 7474 1262 7476 1314
rect 5628 690 5684 700
rect 7420 112 7476 1262
rect 8092 1204 8148 1214
rect 8428 1204 8484 3500
rect 8092 1202 8484 1204
rect 8092 1150 8094 1202
rect 8146 1150 8484 1202
rect 8092 1148 8484 1150
rect 8092 1138 8148 1148
rect 8540 420 8596 12124
rect 8876 12114 8932 12124
rect 8988 11844 9044 12684
rect 8764 11788 9044 11844
rect 8764 11620 8820 11788
rect 8764 11554 8820 11564
rect 8876 11620 8932 11630
rect 9212 11620 9268 11630
rect 8876 11618 9268 11620
rect 8876 11566 8878 11618
rect 8930 11566 9214 11618
rect 9266 11566 9268 11618
rect 8876 11564 9268 11566
rect 8876 11554 8932 11564
rect 9212 11554 9268 11564
rect 8876 11282 8932 11294
rect 8876 11230 8878 11282
rect 8930 11230 8932 11282
rect 8876 10500 8932 11230
rect 9324 11284 9380 12684
rect 9324 11218 9380 11228
rect 9436 12068 9492 12078
rect 9436 10948 9492 12012
rect 9436 10882 9492 10892
rect 8988 10724 9044 10734
rect 8988 10610 9044 10668
rect 9548 10612 9604 10622
rect 8988 10558 8990 10610
rect 9042 10558 9044 10610
rect 8988 10546 9044 10558
rect 9324 10610 9604 10612
rect 9324 10558 9550 10610
rect 9602 10558 9604 10610
rect 9324 10556 9604 10558
rect 8876 9714 8932 10444
rect 8876 9662 8878 9714
rect 8930 9662 8932 9714
rect 8876 7700 8932 9662
rect 9324 8036 9380 10556
rect 9548 10546 9604 10556
rect 9324 7970 9380 7980
rect 9548 9940 9604 9950
rect 8876 7634 8932 7644
rect 8652 7364 8708 7374
rect 8652 7270 8708 7308
rect 9324 6244 9380 6254
rect 8764 4900 8820 4910
rect 8764 4452 8820 4844
rect 8764 4450 9156 4452
rect 8764 4398 8766 4450
rect 8818 4398 9156 4450
rect 8764 4396 9156 4398
rect 8764 4386 8820 4396
rect 9100 4228 9156 4396
rect 9324 4450 9380 6188
rect 9436 6132 9492 6142
rect 9548 6132 9604 9884
rect 9660 9938 9716 12908
rect 10220 12962 10276 12974
rect 10220 12910 10222 12962
rect 10274 12910 10276 12962
rect 10108 12404 10164 12414
rect 10108 12310 10164 12348
rect 10108 11844 10164 11854
rect 9772 11284 9828 11294
rect 9772 11282 10052 11284
rect 9772 11230 9774 11282
rect 9826 11230 10052 11282
rect 9772 11228 10052 11230
rect 9772 11218 9828 11228
rect 9884 10500 9940 10510
rect 9884 10406 9940 10444
rect 9660 9886 9662 9938
rect 9714 9886 9716 9938
rect 9660 9874 9716 9886
rect 9436 6130 9604 6132
rect 9436 6078 9438 6130
rect 9490 6078 9604 6130
rect 9436 6076 9604 6078
rect 9660 8820 9716 8830
rect 9884 8820 9940 8830
rect 9660 8818 9940 8820
rect 9660 8766 9662 8818
rect 9714 8766 9886 8818
rect 9938 8766 9940 8818
rect 9660 8764 9940 8766
rect 9436 6066 9492 6076
rect 9324 4398 9326 4450
rect 9378 4398 9380 4450
rect 9324 4386 9380 4398
rect 9100 3780 9156 4172
rect 9324 3780 9380 3790
rect 9100 3778 9380 3780
rect 9100 3726 9102 3778
rect 9154 3726 9326 3778
rect 9378 3726 9380 3778
rect 9100 3724 9380 3726
rect 9100 3714 9156 3724
rect 9324 3714 9380 3724
rect 9660 3388 9716 8764
rect 9884 8754 9940 8764
rect 9996 8484 10052 11228
rect 10108 11172 10164 11788
rect 10108 11106 10164 11116
rect 10220 9716 10276 12910
rect 10220 9650 10276 9660
rect 10332 10052 10388 10062
rect 10220 9156 10276 9166
rect 10220 8820 10276 9100
rect 10220 8754 10276 8764
rect 9996 8428 10276 8484
rect 9772 8148 9828 8158
rect 9772 5348 9828 8092
rect 9884 7252 9940 7262
rect 9884 7158 9940 7196
rect 9772 5282 9828 5292
rect 10108 6916 10164 6926
rect 10108 4788 10164 6860
rect 10108 4722 10164 4732
rect 9772 4228 9828 4238
rect 9772 4134 9828 4172
rect 10220 3780 10276 8428
rect 10220 3714 10276 3724
rect 9884 3442 9940 3454
rect 9884 3390 9886 3442
rect 9938 3390 9940 3442
rect 9660 3332 9828 3388
rect 9772 1876 9828 3332
rect 9772 1810 9828 1820
rect 9884 1652 9940 3390
rect 10332 2996 10388 9996
rect 10444 9826 10500 9838
rect 10444 9774 10446 9826
rect 10498 9774 10500 9826
rect 10444 9156 10500 9774
rect 10556 9716 10612 14112
rect 11004 12404 11060 14112
rect 11340 13188 11396 13198
rect 11340 13094 11396 13132
rect 11004 12338 11060 12348
rect 11452 12292 11508 14112
rect 11900 13972 11956 14112
rect 11900 13906 11956 13916
rect 11900 13748 11956 13758
rect 11900 13074 11956 13692
rect 11900 13022 11902 13074
rect 11954 13022 11956 13074
rect 11900 13010 11956 13022
rect 12012 12404 12068 12414
rect 12012 12310 12068 12348
rect 11116 12236 11508 12292
rect 11004 12180 11060 12190
rect 11004 12086 11060 12124
rect 10668 12068 10724 12078
rect 10668 11974 10724 12012
rect 11116 11956 11172 12236
rect 10892 11900 11172 11956
rect 11564 12180 11620 12190
rect 10892 11618 10948 11900
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 11452 11394 11508 11406
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11340 10612 11396 10622
rect 11116 10386 11172 10398
rect 11116 10334 11118 10386
rect 11170 10334 11172 10386
rect 11116 10164 11172 10334
rect 11116 10098 11172 10108
rect 11004 9716 11060 9726
rect 10556 9714 11060 9716
rect 10556 9662 11006 9714
rect 11058 9662 11060 9714
rect 10556 9660 11060 9662
rect 11004 9650 11060 9660
rect 11340 9266 11396 10556
rect 11340 9214 11342 9266
rect 11394 9214 11396 9266
rect 11340 9202 11396 9214
rect 10444 9090 10500 9100
rect 10444 8930 10500 8942
rect 10444 8878 10446 8930
rect 10498 8878 10500 8930
rect 10444 3220 10500 8878
rect 11004 8818 11060 8830
rect 11004 8766 11006 8818
rect 11058 8766 11060 8818
rect 10556 7252 10612 7262
rect 10556 6690 10612 7196
rect 10556 6638 10558 6690
rect 10610 6638 10612 6690
rect 10556 6626 10612 6638
rect 11004 6690 11060 8766
rect 11340 7700 11396 7710
rect 11004 6638 11006 6690
rect 11058 6638 11060 6690
rect 11004 6626 11060 6638
rect 11116 6692 11172 6702
rect 11116 6598 11172 6636
rect 11228 6690 11284 6702
rect 11228 6638 11230 6690
rect 11282 6638 11284 6690
rect 10668 6468 10724 6478
rect 11228 6468 11284 6638
rect 10668 6466 11284 6468
rect 10668 6414 10670 6466
rect 10722 6414 11284 6466
rect 10668 6412 11284 6414
rect 10668 6402 10724 6412
rect 10892 5124 10948 5134
rect 10892 4562 10948 5068
rect 10892 4510 10894 4562
rect 10946 4510 10948 4562
rect 10892 4498 10948 4510
rect 11340 3388 11396 7644
rect 10444 3154 10500 3164
rect 10892 3332 11396 3388
rect 11452 3388 11508 11342
rect 11564 9604 11620 12124
rect 12348 11282 12404 14112
rect 12796 12404 12852 14112
rect 12796 12338 12852 12348
rect 12908 13972 12964 13982
rect 12908 12068 12964 13916
rect 13244 13188 13300 14112
rect 13244 13122 13300 13132
rect 13356 13300 13412 13310
rect 13356 13074 13412 13244
rect 13356 13022 13358 13074
rect 13410 13022 13412 13074
rect 13356 13010 13412 13022
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 11218 12404 11230
rect 12796 12012 12964 12068
rect 13468 12516 13524 12526
rect 11676 10612 11732 10622
rect 11676 10518 11732 10556
rect 12572 10612 12628 10622
rect 11900 10500 11956 10510
rect 12124 10500 12180 10510
rect 11956 10444 12068 10500
rect 11900 10434 11956 10444
rect 12012 10276 12068 10444
rect 12124 10406 12180 10444
rect 12572 10388 12628 10556
rect 12684 10388 12740 10398
rect 12572 10386 12740 10388
rect 12572 10334 12686 10386
rect 12738 10334 12740 10386
rect 12572 10332 12740 10334
rect 12012 10220 12292 10276
rect 11900 10164 11956 10174
rect 11564 9538 11620 9548
rect 11676 9716 11732 9726
rect 11564 6690 11620 6702
rect 11564 6638 11566 6690
rect 11618 6638 11620 6690
rect 11564 6130 11620 6638
rect 11676 6468 11732 9660
rect 11788 9156 11844 9166
rect 11788 6916 11844 9100
rect 11900 9042 11956 10108
rect 11900 8990 11902 9042
rect 11954 8990 11956 9042
rect 11900 8372 11956 8990
rect 12012 9826 12068 9838
rect 12012 9774 12014 9826
rect 12066 9774 12068 9826
rect 12012 9044 12068 9774
rect 12012 8978 12068 8988
rect 12124 8930 12180 8942
rect 12124 8878 12126 8930
rect 12178 8878 12180 8930
rect 12124 8484 12180 8878
rect 12124 8418 12180 8428
rect 11900 8306 11956 8316
rect 12236 8260 12292 10220
rect 12124 8204 12292 8260
rect 12348 10164 12404 10174
rect 12124 7588 12180 8204
rect 12348 8148 12404 10108
rect 12572 9714 12628 10332
rect 12684 10322 12740 10332
rect 12572 9662 12574 9714
rect 12626 9662 12628 9714
rect 12460 8484 12516 8494
rect 12460 8390 12516 8428
rect 12572 8260 12628 9662
rect 12796 8260 12852 12012
rect 13020 11956 13076 11966
rect 13244 11956 13300 11966
rect 12908 11954 13300 11956
rect 12908 11902 13022 11954
rect 13074 11902 13246 11954
rect 13298 11902 13300 11954
rect 12908 11900 13300 11902
rect 12908 10052 12964 11900
rect 13020 11890 13076 11900
rect 13244 11890 13300 11900
rect 13020 11508 13076 11518
rect 13468 11508 13524 12460
rect 13020 11506 13524 11508
rect 13020 11454 13022 11506
rect 13074 11454 13524 11506
rect 13020 11452 13524 11454
rect 13580 12068 13636 12078
rect 13020 11442 13076 11452
rect 13580 11060 13636 12012
rect 13692 11956 13748 14112
rect 13804 13412 13860 13422
rect 13804 12290 13860 13356
rect 14140 13188 14196 14112
rect 13804 12238 13806 12290
rect 13858 12238 13860 12290
rect 13804 12226 13860 12238
rect 14028 13132 14196 13188
rect 14364 13636 14420 13646
rect 13692 11900 13972 11956
rect 13580 10994 13636 11004
rect 13804 10724 13860 10734
rect 13580 10722 13860 10724
rect 13580 10670 13806 10722
rect 13858 10670 13860 10722
rect 13580 10668 13860 10670
rect 13132 10388 13188 10398
rect 13356 10388 13412 10398
rect 13132 10386 13412 10388
rect 13132 10334 13134 10386
rect 13186 10334 13358 10386
rect 13410 10334 13412 10386
rect 13132 10332 13412 10334
rect 13132 10164 13188 10332
rect 13356 10322 13412 10332
rect 13132 10098 13188 10108
rect 13356 10164 13412 10174
rect 12908 9986 12964 9996
rect 13020 9826 13076 9838
rect 13020 9774 13022 9826
rect 13074 9774 13076 9826
rect 12908 9156 12964 9166
rect 12908 9062 12964 9100
rect 13020 8484 13076 9774
rect 13020 8418 13076 8428
rect 13244 9716 13300 9726
rect 12348 8082 12404 8092
rect 12460 8204 12628 8260
rect 12684 8204 12852 8260
rect 12908 8372 12964 8382
rect 12124 7522 12180 7532
rect 12236 7812 12292 7822
rect 12236 7474 12292 7756
rect 12236 7422 12238 7474
rect 12290 7422 12292 7474
rect 12236 7410 12292 7422
rect 11900 7252 11956 7262
rect 12124 7252 12180 7262
rect 11900 7250 12068 7252
rect 11900 7198 11902 7250
rect 11954 7198 12068 7250
rect 11900 7196 12068 7198
rect 11900 7186 11956 7196
rect 11788 6860 11956 6916
rect 11788 6692 11844 6702
rect 11788 6598 11844 6636
rect 11676 6412 11844 6468
rect 11788 6244 11844 6412
rect 11788 6178 11844 6188
rect 11564 6078 11566 6130
rect 11618 6078 11620 6130
rect 11564 6066 11620 6078
rect 11676 5796 11732 5806
rect 11676 5794 11844 5796
rect 11676 5742 11678 5794
rect 11730 5742 11844 5794
rect 11676 5740 11844 5742
rect 11676 5730 11732 5740
rect 11788 5124 11844 5740
rect 11788 5058 11844 5068
rect 11676 5012 11732 5022
rect 11452 3332 11620 3388
rect 10332 2930 10388 2940
rect 9884 1586 9940 1596
rect 10780 2324 10836 2334
rect 8540 354 8596 364
rect 9884 1314 9940 1326
rect 9884 1262 9886 1314
rect 9938 1262 9940 1314
rect 9436 196 9492 206
rect 9436 112 9492 140
rect 9884 196 9940 1262
rect 9884 130 9940 140
rect 1344 0 1456 112
rect 3360 0 3472 112
rect 5376 0 5488 112
rect 7392 0 7504 112
rect 9408 0 9520 112
rect 10780 84 10836 2268
rect 10892 1202 10948 3332
rect 10892 1150 10894 1202
rect 10946 1150 10948 1202
rect 10892 1138 10948 1150
rect 11564 1204 11620 3332
rect 11676 1428 11732 4956
rect 11788 4452 11844 4462
rect 11900 4452 11956 6860
rect 12012 6804 12068 7196
rect 12124 7158 12180 7196
rect 12012 6748 12180 6804
rect 12124 6690 12180 6748
rect 12348 6692 12404 6702
rect 12124 6638 12126 6690
rect 12178 6638 12180 6690
rect 12124 6626 12180 6638
rect 12236 6690 12404 6692
rect 12236 6638 12350 6690
rect 12402 6638 12404 6690
rect 12236 6636 12404 6638
rect 12012 6578 12068 6590
rect 12012 6526 12014 6578
rect 12066 6526 12068 6578
rect 12012 6132 12068 6526
rect 12012 6066 12068 6076
rect 12236 5796 12292 6636
rect 12348 6626 12404 6636
rect 12460 6468 12516 8204
rect 12684 7140 12740 8204
rect 12796 8034 12852 8046
rect 12796 7982 12798 8034
rect 12850 7982 12852 8034
rect 12796 7812 12852 7982
rect 12796 7746 12852 7756
rect 12684 7074 12740 7084
rect 12796 7476 12852 7486
rect 12012 5740 12292 5796
rect 12348 6412 12516 6468
rect 12012 5346 12068 5740
rect 12012 5294 12014 5346
rect 12066 5294 12068 5346
rect 12012 5282 12068 5294
rect 12236 5124 12292 5134
rect 12124 5012 12180 5022
rect 12124 4918 12180 4956
rect 11788 4450 11956 4452
rect 11788 4398 11790 4450
rect 11842 4398 11956 4450
rect 11788 4396 11956 4398
rect 11788 4386 11844 4396
rect 12236 4338 12292 5068
rect 12236 4286 12238 4338
rect 12290 4286 12292 4338
rect 12236 4274 12292 4286
rect 12348 2548 12404 6412
rect 12460 6132 12516 6142
rect 12460 5236 12516 6076
rect 12460 5234 12740 5236
rect 12460 5182 12462 5234
rect 12514 5182 12740 5234
rect 12460 5180 12740 5182
rect 12460 5124 12516 5180
rect 12460 5058 12516 5068
rect 12684 4450 12740 5180
rect 12684 4398 12686 4450
rect 12738 4398 12740 4450
rect 12684 4386 12740 4398
rect 12796 3444 12852 7420
rect 12908 5122 12964 8316
rect 13132 8034 13188 8046
rect 13132 7982 13134 8034
rect 13186 7982 13188 8034
rect 13132 7476 13188 7982
rect 13132 7410 13188 7420
rect 13132 7140 13188 7150
rect 12908 5070 12910 5122
rect 12962 5070 12964 5122
rect 12908 5058 12964 5070
rect 13020 6804 13076 6814
rect 13020 3892 13076 6748
rect 13020 3826 13076 3836
rect 13132 3388 13188 7084
rect 12796 3378 12852 3388
rect 12348 2482 12404 2492
rect 12908 3332 13188 3388
rect 12908 2098 12964 3332
rect 12908 2046 12910 2098
rect 12962 2046 12964 2098
rect 12908 2034 12964 2046
rect 11676 1362 11732 1372
rect 11900 1762 11956 1774
rect 11900 1710 11902 1762
rect 11954 1710 11956 1762
rect 11564 1138 11620 1148
rect 11452 196 11508 206
rect 11452 112 11508 140
rect 11900 196 11956 1710
rect 13244 644 13300 9660
rect 13356 9714 13412 10108
rect 13356 9662 13358 9714
rect 13410 9662 13412 9714
rect 13356 9650 13412 9662
rect 13580 9044 13636 10668
rect 13804 10658 13860 10668
rect 13916 9828 13972 11900
rect 14028 11618 14084 13132
rect 14028 11566 14030 11618
rect 14082 11566 14084 11618
rect 14028 11554 14084 11566
rect 14140 12962 14196 12974
rect 14140 12910 14142 12962
rect 14194 12910 14196 12962
rect 14140 9940 14196 12910
rect 14252 12180 14308 12190
rect 14252 11956 14308 12124
rect 14252 11890 14308 11900
rect 14252 10500 14308 10510
rect 14252 10406 14308 10444
rect 14140 9884 14308 9940
rect 13916 9772 14196 9828
rect 14140 9714 14196 9772
rect 14140 9662 14142 9714
rect 14194 9662 14196 9714
rect 14140 9650 14196 9662
rect 13580 8988 14196 9044
rect 13468 8820 13524 8830
rect 13804 8820 13860 8830
rect 13468 8818 13860 8820
rect 13468 8766 13470 8818
rect 13522 8766 13806 8818
rect 13858 8766 13860 8818
rect 13468 8764 13860 8766
rect 13468 8754 13524 8764
rect 13468 8372 13524 8382
rect 13468 8278 13524 8316
rect 13356 8036 13412 8046
rect 13356 6804 13412 7980
rect 13580 7476 13636 7486
rect 13580 7382 13636 7420
rect 13356 6738 13412 6748
rect 13468 5234 13524 5246
rect 13468 5182 13470 5234
rect 13522 5182 13524 5234
rect 13356 5124 13412 5134
rect 13356 5030 13412 5068
rect 13468 5012 13524 5182
rect 13468 4946 13524 4956
rect 13468 4676 13524 4686
rect 13468 4450 13524 4620
rect 13468 4398 13470 4450
rect 13522 4398 13524 4450
rect 13468 4386 13524 4398
rect 13804 4228 13860 8764
rect 13916 8820 13972 8830
rect 13916 8818 14084 8820
rect 13916 8766 13918 8818
rect 13970 8766 14084 8818
rect 13916 8764 14084 8766
rect 13916 8754 13972 8764
rect 14028 8484 14084 8764
rect 14028 8418 14084 8428
rect 13916 8372 13972 8382
rect 13916 8278 13972 8316
rect 14028 7812 14084 7822
rect 14028 7586 14084 7756
rect 14028 7534 14030 7586
rect 14082 7534 14084 7586
rect 14028 7522 14084 7534
rect 13916 7252 13972 7262
rect 13916 5234 13972 7196
rect 14140 6356 14196 8988
rect 14252 7028 14308 9884
rect 14364 9156 14420 13580
rect 14364 9090 14420 9100
rect 14476 12852 14532 12862
rect 14364 8372 14420 8382
rect 14364 8258 14420 8316
rect 14364 8206 14366 8258
rect 14418 8206 14420 8258
rect 14364 7252 14420 8206
rect 14476 7812 14532 12796
rect 14588 12292 14644 14112
rect 14812 13860 14868 13870
rect 14812 12852 14868 13804
rect 15036 13300 15092 14112
rect 15036 13234 15092 13244
rect 14924 13076 14980 13086
rect 14924 12982 14980 13020
rect 14812 12796 14980 12852
rect 14812 12404 14868 12414
rect 14812 12310 14868 12348
rect 14588 12236 14756 12292
rect 14476 7746 14532 7756
rect 14588 11394 14644 11406
rect 14588 11342 14590 11394
rect 14642 11342 14644 11394
rect 14476 7476 14532 7486
rect 14476 7382 14532 7420
rect 14364 7158 14420 7196
rect 14252 6972 14420 7028
rect 14140 6290 14196 6300
rect 13916 5182 13918 5234
rect 13970 5182 13972 5234
rect 13916 5170 13972 5182
rect 14252 5908 14308 5918
rect 14252 5124 14308 5852
rect 14252 4452 14308 5068
rect 14028 4450 14308 4452
rect 14028 4398 14254 4450
rect 14306 4398 14308 4450
rect 14028 4396 14308 4398
rect 14028 4338 14084 4396
rect 14252 4386 14308 4396
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 13804 4162 13860 4172
rect 13356 3668 13412 3678
rect 13356 3332 13412 3612
rect 13356 3266 13412 3276
rect 13244 578 13300 588
rect 13916 1314 13972 1326
rect 13916 1262 13918 1314
rect 13970 1262 13972 1314
rect 11900 130 11956 140
rect 13468 196 13524 206
rect 13468 112 13524 140
rect 13916 196 13972 1262
rect 14364 532 14420 6972
rect 14588 5796 14644 11342
rect 14700 10836 14756 12236
rect 14812 10836 14868 10846
rect 14700 10834 14868 10836
rect 14700 10782 14814 10834
rect 14866 10782 14868 10834
rect 14700 10780 14868 10782
rect 14812 10770 14868 10780
rect 14812 9380 14868 9390
rect 14700 8596 14756 8606
rect 14700 7586 14756 8540
rect 14700 7534 14702 7586
rect 14754 7534 14756 7586
rect 14700 7476 14756 7534
rect 14700 7410 14756 7420
rect 14588 5730 14644 5740
rect 14700 5236 14756 5246
rect 14700 5122 14756 5180
rect 14700 5070 14702 5122
rect 14754 5070 14756 5122
rect 14700 5058 14756 5070
rect 14812 1202 14868 9324
rect 14924 8370 14980 12796
rect 15260 12628 15316 12638
rect 15148 12180 15204 12190
rect 15148 11508 15204 12124
rect 15148 11442 15204 11452
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14924 8306 14980 8318
rect 15036 9826 15092 9838
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 14924 4564 14980 4574
rect 14924 2884 14980 4508
rect 15036 4340 15092 9774
rect 15260 9492 15316 12572
rect 15372 12180 15428 12190
rect 15372 12086 15428 12124
rect 15484 11282 15540 14112
rect 15820 13300 15876 13310
rect 15708 12962 15764 12974
rect 15708 12910 15710 12962
rect 15762 12910 15764 12962
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15484 11218 15540 11230
rect 15596 12740 15652 12750
rect 15260 9436 15428 9492
rect 15260 9268 15316 9278
rect 15148 8146 15204 8158
rect 15148 8094 15150 8146
rect 15202 8094 15204 8146
rect 15148 7140 15204 8094
rect 15148 7074 15204 7084
rect 15260 7028 15316 9212
rect 15372 7364 15428 9436
rect 15596 9268 15652 12684
rect 15708 11620 15764 12910
rect 15708 11554 15764 11564
rect 15820 10724 15876 13244
rect 15932 12404 15988 14112
rect 16380 13748 16436 14112
rect 16380 13692 16548 13748
rect 15932 12338 15988 12348
rect 16380 12404 16436 12414
rect 16380 12310 16436 12348
rect 15596 9202 15652 9212
rect 15708 10668 15876 10724
rect 16156 11394 16212 11406
rect 16156 11342 16158 11394
rect 16210 11342 16212 11394
rect 15372 7298 15428 7308
rect 15484 9044 15540 9054
rect 15260 6962 15316 6972
rect 15484 6244 15540 8988
rect 15596 7250 15652 7262
rect 15596 7198 15598 7250
rect 15650 7198 15652 7250
rect 15596 6468 15652 7198
rect 15596 6402 15652 6412
rect 15484 6188 15652 6244
rect 15484 5348 15540 5358
rect 15484 5122 15540 5292
rect 15484 5070 15486 5122
rect 15538 5070 15540 5122
rect 15484 5058 15540 5070
rect 15484 4676 15540 4686
rect 15036 4274 15092 4284
rect 15260 4564 15316 4574
rect 15148 4226 15204 4238
rect 15148 4174 15150 4226
rect 15202 4174 15204 4226
rect 15148 3892 15204 4174
rect 15148 3826 15204 3836
rect 15036 3780 15092 3790
rect 15036 2996 15092 3724
rect 15036 2930 15092 2940
rect 14924 2818 14980 2828
rect 15260 2436 15316 4508
rect 15260 2370 15316 2380
rect 15372 4452 15428 4462
rect 15372 2212 15428 4396
rect 15484 3332 15540 4620
rect 15484 3266 15540 3276
rect 15372 2146 15428 2156
rect 14812 1150 14814 1202
rect 14866 1150 14868 1202
rect 14812 1138 14868 1150
rect 15484 1764 15540 1774
rect 14364 466 14420 476
rect 13916 130 13972 140
rect 15484 112 15540 1708
rect 15596 1540 15652 6188
rect 15708 5908 15764 10668
rect 15820 10498 15876 10510
rect 15820 10446 15822 10498
rect 15874 10446 15876 10498
rect 15820 10164 15876 10446
rect 15820 10098 15876 10108
rect 16044 9940 16100 9950
rect 16044 9604 16100 9884
rect 16044 9538 16100 9548
rect 16156 8484 16212 11342
rect 16492 10722 16548 13692
rect 16828 13076 16884 14112
rect 16828 13010 16884 13020
rect 16492 10670 16494 10722
rect 16546 10670 16548 10722
rect 16492 10658 16548 10670
rect 16828 12516 16884 12526
rect 16156 8418 16212 8428
rect 16604 10612 16660 10622
rect 16604 8036 16660 10556
rect 16828 10164 16884 12460
rect 16940 12180 16996 12190
rect 17052 12180 17108 14140
rect 17248 14112 17360 14224
rect 17696 14112 17808 14224
rect 18144 14112 18256 14224
rect 18592 14112 18704 14224
rect 19040 14112 19152 14224
rect 19488 14112 19600 14224
rect 19936 14112 20048 14224
rect 20384 14112 20496 14224
rect 20832 14112 20944 14224
rect 21280 14112 21392 14224
rect 21728 14112 21840 14224
rect 22176 14112 22288 14224
rect 22624 14112 22736 14224
rect 23072 14112 23184 14224
rect 23520 14112 23632 14224
rect 23968 14112 24080 14224
rect 24416 14112 24528 14224
rect 24864 14112 24976 14224
rect 25312 14112 25424 14224
rect 25760 14112 25872 14224
rect 26208 14112 26320 14224
rect 26656 14112 26768 14224
rect 27104 14112 27216 14224
rect 27552 14112 27664 14224
rect 28000 14112 28112 14224
rect 28448 14112 28560 14224
rect 28896 14112 29008 14224
rect 29344 14112 29456 14224
rect 29792 14112 29904 14224
rect 30044 14196 30100 14206
rect 16940 12178 17108 12180
rect 16940 12126 16942 12178
rect 16994 12126 17108 12178
rect 16940 12124 17108 12126
rect 17164 13076 17220 13086
rect 16940 12114 16996 12124
rect 16716 10108 16884 10164
rect 16940 11732 16996 11742
rect 16716 9828 16772 10108
rect 16716 9762 16772 9772
rect 16716 8820 16772 8830
rect 16716 8260 16772 8764
rect 16716 8194 16772 8204
rect 16604 7970 16660 7980
rect 16380 7924 16436 7934
rect 15708 5842 15764 5852
rect 15820 7812 15876 7822
rect 15820 7588 15876 7756
rect 15820 5124 15876 7532
rect 16044 7812 16100 7822
rect 15932 6132 15988 6142
rect 15932 5346 15988 6076
rect 16044 6020 16100 7756
rect 16156 7588 16212 7598
rect 16156 7494 16212 7532
rect 16380 6804 16436 7868
rect 16380 6738 16436 6748
rect 16492 7362 16548 7374
rect 16492 7310 16494 7362
rect 16546 7310 16548 7362
rect 16492 6804 16548 7310
rect 16716 6804 16772 6814
rect 16492 6802 16772 6804
rect 16492 6750 16718 6802
rect 16770 6750 16772 6802
rect 16492 6748 16772 6750
rect 16268 6580 16324 6590
rect 16492 6580 16548 6748
rect 16716 6738 16772 6748
rect 16268 6578 16548 6580
rect 16268 6526 16270 6578
rect 16322 6526 16548 6578
rect 16268 6524 16548 6526
rect 16268 6468 16324 6524
rect 16268 6402 16324 6412
rect 16716 6468 16772 6478
rect 16716 6244 16772 6412
rect 16716 6178 16772 6188
rect 16044 5954 16100 5964
rect 16268 5908 16324 5918
rect 15932 5294 15934 5346
rect 15986 5294 15988 5346
rect 15932 5282 15988 5294
rect 16044 5572 16100 5582
rect 16044 5348 16100 5516
rect 15820 5058 15876 5068
rect 16044 4450 16100 5292
rect 16268 5124 16324 5852
rect 16940 5684 16996 11676
rect 17164 10500 17220 13020
rect 17276 12404 17332 14112
rect 17388 13188 17444 13198
rect 17388 13094 17444 13132
rect 17724 12628 17780 14112
rect 17276 12338 17332 12348
rect 17500 12572 17780 12628
rect 17836 12962 17892 12974
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17500 11618 17556 12572
rect 17500 11566 17502 11618
rect 17554 11566 17556 11618
rect 17500 11554 17556 11566
rect 17164 10434 17220 10444
rect 17500 10610 17556 10622
rect 17500 10558 17502 10610
rect 17554 10558 17556 10610
rect 17388 9828 17444 9838
rect 17388 9734 17444 9772
rect 17500 9604 17556 10558
rect 17500 9538 17556 9548
rect 17724 10498 17780 10510
rect 17724 10446 17726 10498
rect 17778 10446 17780 10498
rect 17724 9492 17780 10446
rect 17836 10164 17892 12910
rect 17948 12404 18004 12414
rect 18172 12404 18228 14112
rect 18620 13188 18676 14112
rect 18620 13122 18676 13132
rect 18956 13188 19012 13198
rect 18956 13094 19012 13132
rect 17948 12402 18228 12404
rect 17948 12350 17950 12402
rect 18002 12350 18228 12402
rect 17948 12348 18228 12350
rect 17948 12338 18004 12348
rect 18284 12178 18340 12190
rect 18284 12126 18286 12178
rect 18338 12126 18340 12178
rect 18172 11956 18228 11966
rect 18060 11396 18116 11406
rect 18060 11302 18116 11340
rect 18172 11172 18228 11900
rect 18284 11732 18340 12126
rect 18284 11666 18340 11676
rect 18396 12180 18452 12190
rect 18396 11284 18452 12124
rect 19068 11618 19124 14112
rect 19516 13188 19572 14112
rect 19404 13132 19572 13188
rect 19964 13188 20020 14112
rect 19068 11566 19070 11618
rect 19122 11566 19124 11618
rect 19068 11554 19124 11566
rect 19292 12740 19348 12750
rect 18396 11218 18452 11228
rect 18172 11106 18228 11116
rect 18284 10724 18340 10734
rect 18060 10668 18284 10724
rect 18060 10276 18116 10668
rect 18284 10630 18340 10668
rect 19180 10724 19236 10734
rect 19180 10630 19236 10668
rect 19292 10612 19348 12684
rect 19404 12290 19460 13132
rect 19964 13122 20020 13132
rect 19404 12238 19406 12290
rect 19458 12238 19460 12290
rect 19404 12226 19460 12238
rect 19516 12962 19572 12974
rect 19516 12910 19518 12962
rect 19570 12910 19572 12962
rect 19516 11844 19572 12910
rect 19516 11778 19572 11788
rect 19964 12068 20020 12078
rect 19516 11508 19572 11518
rect 19516 11060 19572 11452
rect 19964 11508 20020 12012
rect 20076 12068 20132 12078
rect 20076 12066 20244 12068
rect 20076 12014 20078 12066
rect 20130 12014 20244 12066
rect 20076 12012 20244 12014
rect 20076 12002 20132 12012
rect 19964 11442 20020 11452
rect 19628 11396 19684 11406
rect 19628 11394 19908 11396
rect 19628 11342 19630 11394
rect 19682 11342 19908 11394
rect 19628 11340 19908 11342
rect 19628 11330 19684 11340
rect 19516 11004 19684 11060
rect 19516 10836 19572 10846
rect 19292 10546 19348 10556
rect 19404 10724 19460 10734
rect 18732 10500 18788 10510
rect 18620 10388 18676 10398
rect 17836 10098 17892 10108
rect 17948 10220 18116 10276
rect 18396 10386 18676 10388
rect 18396 10334 18622 10386
rect 18674 10334 18676 10386
rect 18396 10332 18676 10334
rect 17948 10050 18004 10220
rect 17948 9998 17950 10050
rect 18002 9998 18004 10050
rect 17948 9986 18004 9998
rect 18060 10052 18116 10062
rect 17724 9426 17780 9436
rect 18060 9154 18116 9996
rect 18284 9826 18340 9838
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 18284 9492 18340 9774
rect 18284 9426 18340 9436
rect 18060 9102 18062 9154
rect 18114 9102 18116 9154
rect 18060 9090 18116 9102
rect 18284 9268 18340 9278
rect 17836 8484 17892 8494
rect 17724 7364 17780 7374
rect 17724 7270 17780 7308
rect 17724 6804 17780 6814
rect 16940 5618 16996 5628
rect 17052 6692 17108 6702
rect 16604 5348 16660 5358
rect 16156 5068 16324 5124
rect 16380 5292 16604 5348
rect 16380 5236 16436 5292
rect 16604 5254 16660 5292
rect 16156 5010 16212 5068
rect 16156 4958 16158 5010
rect 16210 4958 16212 5010
rect 16156 4946 16212 4958
rect 16044 4398 16046 4450
rect 16098 4398 16100 4450
rect 16044 4386 16100 4398
rect 16156 4452 16212 4462
rect 16380 4452 16436 5180
rect 17052 5236 17108 6636
rect 17052 5170 17108 5180
rect 17276 6578 17332 6590
rect 17276 6526 17278 6578
rect 17330 6526 17332 6578
rect 16156 4450 16436 4452
rect 16156 4398 16158 4450
rect 16210 4398 16436 4450
rect 16156 4396 16436 4398
rect 15708 4228 15764 4238
rect 16156 4228 16212 4396
rect 15708 4226 16212 4228
rect 15708 4174 15710 4226
rect 15762 4174 16212 4226
rect 15708 4172 16212 4174
rect 15708 4162 15764 4172
rect 15596 1474 15652 1484
rect 17276 644 17332 6526
rect 17612 6020 17668 6030
rect 17612 2884 17668 5964
rect 17724 5012 17780 6748
rect 17724 4946 17780 4956
rect 17836 3668 17892 8428
rect 18284 8484 18340 9212
rect 18284 8418 18340 8428
rect 18396 8370 18452 10332
rect 18620 10322 18676 10332
rect 18732 9828 18788 10444
rect 18956 10386 19012 10398
rect 18956 10334 18958 10386
rect 19010 10334 19012 10386
rect 18844 10052 18900 10062
rect 18844 9938 18900 9996
rect 18844 9886 18846 9938
rect 18898 9886 18900 9938
rect 18844 9874 18900 9886
rect 18732 9762 18788 9772
rect 18956 9492 19012 10334
rect 19404 10050 19460 10668
rect 19516 10722 19572 10780
rect 19516 10670 19518 10722
rect 19570 10670 19572 10722
rect 19516 10658 19572 10670
rect 19404 9998 19406 10050
rect 19458 9998 19460 10050
rect 19404 9986 19460 9998
rect 18956 9426 19012 9436
rect 19180 9714 19236 9726
rect 19180 9662 19182 9714
rect 19234 9662 19236 9714
rect 19180 9492 19236 9662
rect 19180 9426 19236 9436
rect 19292 9604 19348 9614
rect 18844 9268 18900 9278
rect 18844 9156 18900 9212
rect 18620 9154 18900 9156
rect 18620 9102 18846 9154
rect 18898 9102 18900 9154
rect 18620 9100 18900 9102
rect 18620 9042 18676 9100
rect 18844 9090 18900 9100
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18620 8978 18676 8990
rect 18620 8596 18676 8606
rect 18396 8318 18398 8370
rect 18450 8318 18452 8370
rect 18396 8306 18452 8318
rect 18508 8370 18564 8382
rect 18508 8318 18510 8370
rect 18562 8318 18564 8370
rect 18508 8036 18564 8318
rect 18508 7970 18564 7980
rect 18620 7812 18676 8540
rect 18732 8260 18788 8270
rect 19068 8260 19124 8270
rect 18732 8258 18900 8260
rect 18732 8206 18734 8258
rect 18786 8206 18900 8258
rect 18732 8204 18900 8206
rect 18732 8194 18788 8204
rect 18508 7756 18676 7812
rect 18284 7588 18340 7598
rect 18284 7364 18340 7532
rect 18284 7270 18340 7308
rect 18396 7250 18452 7262
rect 18396 7198 18398 7250
rect 18450 7198 18452 7250
rect 18284 6692 18340 6702
rect 17948 6690 18340 6692
rect 17948 6638 18286 6690
rect 18338 6638 18340 6690
rect 17948 6636 18340 6638
rect 17948 4562 18004 6636
rect 18284 6626 18340 6636
rect 18396 6692 18452 7198
rect 18396 6626 18452 6636
rect 18508 6580 18564 7756
rect 18732 7700 18788 7710
rect 18620 7474 18676 7486
rect 18620 7422 18622 7474
rect 18674 7422 18676 7474
rect 18620 6914 18676 7422
rect 18732 7252 18788 7644
rect 18844 7476 18900 8204
rect 19068 8258 19236 8260
rect 19068 8206 19070 8258
rect 19122 8206 19236 8258
rect 19068 8204 19236 8206
rect 19068 8194 19124 8204
rect 18956 8036 19012 8046
rect 19180 8036 19236 8204
rect 18956 8034 19124 8036
rect 18956 7982 18958 8034
rect 19010 7982 19124 8034
rect 18956 7980 19124 7982
rect 18956 7970 19012 7980
rect 18956 7476 19012 7486
rect 18844 7474 19012 7476
rect 18844 7422 18958 7474
rect 19010 7422 19012 7474
rect 18844 7420 19012 7422
rect 18956 7410 19012 7420
rect 18844 7252 18900 7262
rect 18732 7250 18900 7252
rect 18732 7198 18846 7250
rect 18898 7198 18900 7250
rect 18732 7196 18900 7198
rect 18844 7186 18900 7196
rect 19068 7028 19124 7980
rect 19180 7970 19236 7980
rect 19292 7700 19348 9548
rect 19628 7812 19684 11004
rect 19628 7746 19684 7756
rect 18620 6862 18622 6914
rect 18674 6862 18676 6914
rect 18620 6850 18676 6862
rect 18732 6972 19124 7028
rect 19180 7644 19348 7700
rect 19404 7700 19460 7710
rect 18732 6802 18788 6972
rect 18732 6750 18734 6802
rect 18786 6750 18788 6802
rect 18732 6738 18788 6750
rect 18844 6692 18900 6702
rect 18844 6598 18900 6636
rect 18508 6524 18788 6580
rect 18508 6132 18564 6142
rect 18396 5124 18452 5134
rect 17948 4510 17950 4562
rect 18002 4510 18004 4562
rect 17948 4498 18004 4510
rect 18284 5012 18340 5022
rect 18284 4562 18340 4956
rect 18284 4510 18286 4562
rect 18338 4510 18340 4562
rect 17836 3602 17892 3612
rect 17948 4340 18004 4350
rect 17948 3666 18004 4284
rect 18284 4116 18340 4510
rect 18396 4340 18452 5068
rect 18508 4676 18564 6076
rect 18508 4610 18564 4620
rect 18396 4274 18452 4284
rect 18284 4060 18564 4116
rect 18508 3780 18564 4060
rect 18732 4004 18788 6524
rect 18844 5124 18900 5134
rect 18844 4226 18900 5068
rect 19068 4340 19124 4350
rect 19180 4340 19236 7644
rect 19292 7364 19348 7402
rect 19292 7298 19348 7308
rect 19404 6244 19460 7644
rect 19516 7588 19572 7598
rect 19572 7532 19684 7588
rect 19516 7522 19572 7532
rect 19628 7474 19684 7532
rect 19628 7422 19630 7474
rect 19682 7422 19684 7474
rect 19628 7410 19684 7422
rect 19740 7586 19796 7598
rect 19740 7534 19742 7586
rect 19794 7534 19796 7586
rect 19740 7364 19796 7534
rect 19852 7476 19908 11340
rect 20188 10612 20244 12012
rect 20412 11506 20468 14112
rect 20636 13972 20692 13982
rect 20524 12962 20580 12974
rect 20524 12910 20526 12962
rect 20578 12910 20580 12962
rect 20524 12852 20580 12910
rect 20524 12786 20580 12796
rect 20636 12404 20692 13916
rect 20860 12516 20916 14112
rect 21308 12740 21364 14112
rect 21308 12674 21364 12684
rect 21420 12964 21476 12974
rect 21420 12628 21476 12908
rect 21756 12898 21812 14112
rect 21532 12850 21812 12898
rect 21532 12798 21534 12850
rect 21586 12842 21812 12850
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 21586 12798 21588 12842
rect 21532 12786 21588 12798
rect 21980 12740 22036 12750
rect 21420 12572 21700 12628
rect 20860 12450 20916 12460
rect 20412 11454 20414 11506
rect 20466 11454 20468 11506
rect 20412 11442 20468 11454
rect 20524 12348 20692 12404
rect 20188 10546 20244 10556
rect 20412 10948 20468 10958
rect 20076 10388 20132 10398
rect 20076 10294 20132 10332
rect 19964 10164 20020 10174
rect 20020 10108 20244 10164
rect 19964 10098 20020 10108
rect 20188 9380 20244 10108
rect 20300 9828 20356 9838
rect 20300 9734 20356 9772
rect 20188 9324 20356 9380
rect 20188 9156 20244 9166
rect 19964 8820 20020 8830
rect 19964 7698 20020 8764
rect 20188 8484 20244 9100
rect 20300 9044 20356 9324
rect 20300 8978 20356 8988
rect 20188 8418 20244 8428
rect 19964 7646 19966 7698
rect 20018 7646 20020 7698
rect 19964 7634 20020 7646
rect 20076 7700 20132 7710
rect 19852 7420 20020 7476
rect 19740 7298 19796 7308
rect 19964 7364 20020 7420
rect 19964 7298 20020 7308
rect 20076 6916 20132 7644
rect 20076 6850 20132 6860
rect 19404 6178 19460 6188
rect 19404 5908 19460 5918
rect 19404 5124 19460 5852
rect 19404 4452 19460 5068
rect 19628 5012 19684 5022
rect 19628 4676 19684 4956
rect 19404 4450 19572 4452
rect 19404 4398 19406 4450
rect 19458 4398 19572 4450
rect 19404 4396 19572 4398
rect 19404 4386 19460 4396
rect 19068 4338 19236 4340
rect 19068 4286 19070 4338
rect 19122 4286 19236 4338
rect 19068 4284 19236 4286
rect 19068 4274 19124 4284
rect 18844 4174 18846 4226
rect 18898 4174 18900 4226
rect 18844 4162 18900 4174
rect 18732 3938 18788 3948
rect 18956 4116 19012 4126
rect 18844 3780 18900 3790
rect 18508 3778 18900 3780
rect 18508 3726 18510 3778
rect 18562 3726 18846 3778
rect 18898 3726 18900 3778
rect 18508 3724 18900 3726
rect 18508 3714 18564 3724
rect 18844 3714 18900 3724
rect 17948 3614 17950 3666
rect 18002 3614 18004 3666
rect 17948 3602 18004 3614
rect 18396 3556 18452 3566
rect 18396 3388 18452 3500
rect 18620 3444 18676 3454
rect 18396 3332 18564 3388
rect 17276 578 17332 588
rect 17500 2828 17668 2884
rect 17500 112 17556 2828
rect 18508 2548 18564 3332
rect 18620 2772 18676 3388
rect 18620 2706 18676 2716
rect 18732 3108 18788 3118
rect 18508 2482 18564 2492
rect 18396 2212 18452 2222
rect 18396 756 18452 2156
rect 18508 2100 18564 2110
rect 18508 1652 18564 2044
rect 18508 1586 18564 1596
rect 18732 868 18788 3052
rect 18732 802 18788 812
rect 18396 690 18452 700
rect 18956 196 19012 4060
rect 19180 4116 19236 4126
rect 19068 3668 19124 3678
rect 19068 3574 19124 3612
rect 19180 3220 19236 4060
rect 19516 3780 19572 4396
rect 19628 4450 19684 4620
rect 19628 4398 19630 4450
rect 19682 4398 19684 4450
rect 19628 4386 19684 4398
rect 20076 4900 20132 4910
rect 19964 3780 20020 3790
rect 19516 3778 20020 3780
rect 19516 3726 19966 3778
rect 20018 3726 20020 3778
rect 19516 3724 20020 3726
rect 19516 3554 19572 3724
rect 19964 3714 20020 3724
rect 19516 3502 19518 3554
rect 19570 3502 19572 3554
rect 19516 3490 19572 3502
rect 19180 3154 19236 3164
rect 19964 2324 20020 2334
rect 20076 2324 20132 4844
rect 20188 4788 20244 4798
rect 20188 3220 20244 4732
rect 20412 4676 20468 10892
rect 20524 10722 20580 12348
rect 20860 12292 20916 12302
rect 20860 12198 20916 12236
rect 20636 12180 20692 12190
rect 20636 12086 20692 12124
rect 21420 12180 21476 12190
rect 21420 12086 21476 12124
rect 20524 10670 20526 10722
rect 20578 10670 20580 10722
rect 20524 10388 20580 10670
rect 20524 10322 20580 10332
rect 20636 11844 20692 11854
rect 20524 9714 20580 9726
rect 20524 9662 20526 9714
rect 20578 9662 20580 9714
rect 20524 8932 20580 9662
rect 20524 8866 20580 8876
rect 20412 4610 20468 4620
rect 20524 6692 20580 6702
rect 20188 3154 20244 3164
rect 20020 2268 20132 2324
rect 19964 2258 20020 2268
rect 20524 2212 20580 6636
rect 20636 3444 20692 11788
rect 21196 11844 21252 11854
rect 21084 11732 21140 11742
rect 21084 11172 21140 11676
rect 21196 11506 21252 11788
rect 21196 11454 21198 11506
rect 21250 11454 21252 11506
rect 21196 11442 21252 11454
rect 21308 11732 21364 11742
rect 21084 11116 21252 11172
rect 21084 10500 21140 10510
rect 21084 10406 21140 10444
rect 21084 9828 21140 9838
rect 20860 9380 20916 9390
rect 20748 7812 20804 7822
rect 20748 6914 20804 7756
rect 20860 7588 20916 9324
rect 20972 9156 21028 9166
rect 21084 9156 21140 9772
rect 20972 9154 21140 9156
rect 20972 9102 20974 9154
rect 21026 9102 21140 9154
rect 20972 9100 21140 9102
rect 20972 9090 21028 9100
rect 20860 7522 20916 7532
rect 20748 6862 20750 6914
rect 20802 6862 20804 6914
rect 20748 6244 20804 6862
rect 20748 6178 20804 6188
rect 20860 6916 20916 6926
rect 20748 5460 20804 5470
rect 20748 5012 20804 5404
rect 20748 4946 20804 4956
rect 20860 4452 20916 6860
rect 21196 6916 21252 11116
rect 21308 10948 21364 11676
rect 21308 10882 21364 10892
rect 21420 10500 21476 10510
rect 21308 9604 21364 9614
rect 21308 9042 21364 9548
rect 21420 9268 21476 10444
rect 21532 9940 21588 9950
rect 21532 9846 21588 9884
rect 21420 9202 21476 9212
rect 21644 9268 21700 12572
rect 21868 12516 21924 12526
rect 21756 11396 21812 11406
rect 21756 9604 21812 11340
rect 21868 10722 21924 12460
rect 21980 11506 22036 12684
rect 21980 11454 21982 11506
rect 22034 11454 22036 11506
rect 21980 11442 22036 11454
rect 21868 10670 21870 10722
rect 21922 10670 21924 10722
rect 21868 10658 21924 10670
rect 21756 9538 21812 9548
rect 21868 10388 21924 10398
rect 21644 9202 21700 9212
rect 21308 8990 21310 9042
rect 21362 8990 21364 9042
rect 21308 8978 21364 8990
rect 21532 9044 21588 9054
rect 21196 6850 21252 6860
rect 21308 6580 21364 6590
rect 21308 6578 21476 6580
rect 21308 6526 21310 6578
rect 21362 6526 21476 6578
rect 21308 6524 21476 6526
rect 21308 6514 21364 6524
rect 21308 6244 21364 6254
rect 21308 6018 21364 6188
rect 21308 5966 21310 6018
rect 21362 5966 21364 6018
rect 21308 5954 21364 5966
rect 20972 5348 21028 5358
rect 20972 5124 21028 5292
rect 20972 5030 21028 5068
rect 21308 5124 21364 5134
rect 21308 5030 21364 5068
rect 21420 4788 21476 6524
rect 20860 4450 21252 4452
rect 20860 4398 20862 4450
rect 20914 4398 21252 4450
rect 20860 4396 21252 4398
rect 20860 4386 20916 4396
rect 20636 3378 20692 3388
rect 21196 4116 21252 4396
rect 21420 4450 21476 4732
rect 21532 4676 21588 8988
rect 21756 9044 21812 9054
rect 21756 8950 21812 8988
rect 21868 8484 21924 10332
rect 22092 10164 22148 12910
rect 22204 12290 22260 14112
rect 22204 12238 22206 12290
rect 22258 12238 22260 12290
rect 22204 12226 22260 12238
rect 22540 13188 22596 13198
rect 22428 11284 22484 11294
rect 22092 10098 22148 10108
rect 22204 10276 22260 10286
rect 22092 9940 22148 9950
rect 22092 9846 22148 9884
rect 21980 8820 22036 8830
rect 21980 8726 22036 8764
rect 22204 8820 22260 10220
rect 22316 9940 22372 9950
rect 22316 9714 22372 9884
rect 22316 9662 22318 9714
rect 22370 9662 22372 9714
rect 22316 9044 22372 9662
rect 22316 8978 22372 8988
rect 22428 8932 22484 11228
rect 22428 8866 22484 8876
rect 22204 8754 22260 8764
rect 21644 8428 21924 8484
rect 21644 8260 21700 8428
rect 21644 8194 21700 8204
rect 22092 8148 22148 8158
rect 21756 8092 22092 8148
rect 21644 7252 21700 7262
rect 21644 7028 21700 7196
rect 21644 6962 21700 6972
rect 21644 6802 21700 6814
rect 21644 6750 21646 6802
rect 21698 6750 21700 6802
rect 21644 6244 21700 6750
rect 21644 5906 21700 6188
rect 21756 6020 21812 8092
rect 22092 8082 22148 8092
rect 22204 7812 22260 7822
rect 21868 7252 21924 7262
rect 21868 6580 21924 7196
rect 22204 7140 22260 7756
rect 22204 7074 22260 7084
rect 21868 6514 21924 6524
rect 21756 5954 21812 5964
rect 22204 6020 22260 6030
rect 22204 5926 22260 5964
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5842 21700 5854
rect 22540 5684 22596 13132
rect 22652 13186 22708 14112
rect 22652 13134 22654 13186
rect 22706 13134 22708 13186
rect 22652 13122 22708 13134
rect 22988 12740 23044 12750
rect 22988 12178 23044 12684
rect 23100 12404 23156 14112
rect 23548 13524 23604 14112
rect 23884 13860 23940 13870
rect 23548 13468 23716 13524
rect 23100 12338 23156 12348
rect 23548 12404 23604 12414
rect 23548 12310 23604 12348
rect 23660 12292 23716 13468
rect 23884 13074 23940 13804
rect 23996 13524 24052 14112
rect 24444 13524 24500 14112
rect 23996 13458 24052 13468
rect 24332 13468 24500 13524
rect 23884 13022 23886 13074
rect 23938 13022 23940 13074
rect 23884 13010 23940 13022
rect 24108 13188 24164 13198
rect 24108 13076 24164 13132
rect 24108 13020 24276 13076
rect 24220 12628 24276 13020
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24220 12562 24276 12572
rect 23804 12506 24068 12516
rect 23996 12292 24052 12302
rect 23660 12236 23996 12292
rect 23996 12226 24052 12236
rect 22988 12126 22990 12178
rect 23042 12126 23044 12178
rect 22988 12114 23044 12126
rect 23548 11956 23604 11966
rect 23324 11844 23380 11854
rect 23324 11620 23380 11788
rect 23436 11620 23492 11630
rect 23324 11564 23436 11620
rect 23436 11554 23492 11564
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22652 9042 22708 9054
rect 22652 8990 22654 9042
rect 22706 8990 22708 9042
rect 22652 8036 22708 8990
rect 22764 8372 22820 11342
rect 23436 11394 23492 11406
rect 23436 11342 23438 11394
rect 23490 11342 23492 11394
rect 23100 11284 23156 11294
rect 23436 11284 23492 11342
rect 23548 11396 23604 11900
rect 23548 11330 23604 11340
rect 23100 11282 23492 11284
rect 23100 11230 23102 11282
rect 23154 11230 23492 11282
rect 23100 11228 23492 11230
rect 23996 11284 24052 11294
rect 23100 9716 23156 11228
rect 23996 11190 24052 11228
rect 24220 11060 24276 11070
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 24220 10386 24276 11004
rect 24220 10334 24222 10386
rect 24274 10334 24276 10386
rect 23324 10276 23380 10286
rect 23100 9650 23156 9660
rect 23212 9940 23268 9950
rect 22764 8306 22820 8316
rect 22876 9492 22932 9502
rect 22652 6916 22708 7980
rect 22876 8036 22932 9436
rect 23212 9042 23268 9884
rect 23212 8990 23214 9042
rect 23266 8990 23268 9042
rect 23212 8978 23268 8990
rect 22876 7970 22932 7980
rect 23212 8260 23268 8270
rect 22876 6916 22932 6926
rect 22652 6914 22932 6916
rect 22652 6862 22878 6914
rect 22930 6862 22932 6914
rect 22652 6860 22932 6862
rect 22876 6850 22932 6860
rect 22540 5618 22596 5628
rect 22652 6580 22708 6590
rect 22652 5348 22708 6524
rect 23212 6244 23268 8204
rect 23212 6178 23268 6188
rect 22428 5236 22484 5246
rect 21868 5124 21924 5134
rect 21868 5030 21924 5068
rect 22316 5124 22372 5134
rect 22316 5030 22372 5068
rect 21532 4610 21588 4620
rect 21420 4398 21422 4450
rect 21474 4398 21476 4450
rect 21420 4386 21476 4398
rect 21308 4340 21364 4350
rect 21308 4246 21364 4284
rect 21868 4340 21924 4350
rect 21756 4226 21812 4238
rect 21756 4174 21758 4226
rect 21810 4174 21812 4226
rect 21756 4116 21812 4174
rect 21196 4060 21812 4116
rect 21196 2884 21252 4060
rect 21644 3780 21700 3790
rect 21196 2882 21588 2884
rect 21196 2830 21198 2882
rect 21250 2830 21588 2882
rect 21196 2828 21588 2830
rect 21196 2818 21252 2828
rect 21532 2770 21588 2828
rect 21532 2718 21534 2770
rect 21586 2718 21588 2770
rect 21532 2706 21588 2718
rect 20524 2146 20580 2156
rect 21644 1428 21700 3724
rect 21756 3556 21812 3566
rect 21868 3556 21924 4284
rect 21812 3500 21924 3556
rect 21756 3490 21812 3500
rect 21756 3220 21812 3230
rect 21756 2884 21812 3164
rect 21756 2818 21812 2828
rect 22092 2658 22148 2670
rect 22092 2606 22094 2658
rect 22146 2606 22148 2658
rect 22092 2436 22148 2606
rect 22092 2370 22148 2380
rect 22428 2212 22484 5180
rect 22540 5124 22596 5134
rect 22540 4340 22596 5068
rect 22652 5010 22708 5292
rect 22652 4958 22654 5010
rect 22706 4958 22708 5010
rect 22652 4946 22708 4958
rect 22988 5234 23044 5246
rect 22988 5182 22990 5234
rect 23042 5182 23044 5234
rect 22988 4562 23044 5182
rect 23212 5234 23268 5246
rect 23212 5182 23214 5234
rect 23266 5182 23268 5234
rect 23212 5012 23268 5182
rect 23212 4946 23268 4956
rect 22988 4510 22990 4562
rect 23042 4510 23044 4562
rect 22988 4498 23044 4510
rect 22540 4274 22596 4284
rect 23324 3892 23380 10220
rect 24220 10276 24276 10334
rect 24220 10210 24276 10220
rect 24220 10052 24276 10062
rect 23996 9940 24052 9950
rect 23996 9846 24052 9884
rect 23548 9714 23604 9726
rect 23548 9662 23550 9714
rect 23602 9662 23604 9714
rect 23548 8708 23604 9662
rect 24220 9492 24276 9996
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24220 9426 24276 9436
rect 23804 9370 24068 9380
rect 24332 9268 24388 13468
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24444 12738 24500 12750
rect 24444 12686 24446 12738
rect 24498 12686 24500 12738
rect 24444 12292 24500 12686
rect 24444 12226 24500 12236
rect 24556 12066 24612 12078
rect 24556 12014 24558 12066
rect 24610 12014 24612 12066
rect 24556 11956 24612 12014
rect 24556 11890 24612 11900
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24556 11394 24612 11406
rect 24556 11342 24558 11394
rect 24610 11342 24612 11394
rect 24556 11060 24612 11342
rect 24556 10994 24612 11004
rect 24892 10948 24948 14112
rect 25340 14084 25396 14112
rect 25340 14018 25396 14028
rect 25452 13524 25508 13534
rect 25228 13412 25284 13422
rect 25116 11956 25172 11966
rect 24892 10882 24948 10892
rect 25004 11954 25172 11956
rect 25004 11902 25118 11954
rect 25170 11902 25172 11954
rect 25004 11900 25172 11902
rect 25004 11844 25060 11900
rect 25116 11890 25172 11900
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 25004 10018 25060 11788
rect 24668 9962 25060 10018
rect 25116 11282 25172 11294
rect 25116 11230 25118 11282
rect 25170 11230 25172 11282
rect 24444 9940 24500 9950
rect 24444 9846 24500 9884
rect 23548 8642 23604 8652
rect 23660 9212 24388 9268
rect 24556 9716 24612 9726
rect 23548 8260 23604 8270
rect 23548 7924 23604 8204
rect 23548 7858 23604 7868
rect 23660 6468 23716 9212
rect 24556 9156 24612 9660
rect 24108 9154 24612 9156
rect 24108 9102 24558 9154
rect 24610 9102 24612 9154
rect 24108 9100 24612 9102
rect 24108 9042 24164 9100
rect 24556 9090 24612 9100
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 24108 8978 24164 8990
rect 24668 8820 24724 9962
rect 24780 9828 24836 9838
rect 24780 9604 24836 9772
rect 25116 9828 25172 11230
rect 25228 10948 25284 13356
rect 25452 13186 25508 13468
rect 25452 13134 25454 13186
rect 25506 13134 25508 13186
rect 25452 13122 25508 13134
rect 25788 12516 25844 14112
rect 25900 13636 25956 13646
rect 25900 13300 25956 13580
rect 25900 13234 25956 13244
rect 25788 12450 25844 12460
rect 26012 12850 26068 12862
rect 26012 12798 26014 12850
rect 26066 12798 26068 12850
rect 25452 12292 25508 12302
rect 25340 11954 25396 11966
rect 25340 11902 25342 11954
rect 25394 11902 25396 11954
rect 25340 11844 25396 11902
rect 25340 11778 25396 11788
rect 25228 10892 25396 10948
rect 25116 9762 25172 9772
rect 25228 10724 25284 10734
rect 25228 9604 25284 10668
rect 25340 10500 25396 10892
rect 25340 10434 25396 10444
rect 24780 9548 25284 9604
rect 25340 10052 25396 10062
rect 24780 9154 24836 9548
rect 24780 9102 24782 9154
rect 24834 9102 24836 9154
rect 24780 9090 24836 9102
rect 24892 9380 24948 9390
rect 24332 8764 24724 8820
rect 24892 8820 24948 9324
rect 25004 9268 25060 9278
rect 25228 9268 25284 9278
rect 25060 9212 25172 9268
rect 25004 9202 25060 9212
rect 25004 9044 25060 9054
rect 25004 8950 25060 8988
rect 25116 8932 25172 9212
rect 25228 9154 25284 9212
rect 25228 9102 25230 9154
rect 25282 9102 25284 9154
rect 25228 9090 25284 9102
rect 25228 8932 25284 8942
rect 25116 8876 25228 8932
rect 25228 8866 25284 8876
rect 24892 8764 25060 8820
rect 24220 8260 24276 8270
rect 24220 7924 24276 8204
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24220 7858 24276 7868
rect 23804 7802 24068 7812
rect 24332 7700 24388 8764
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24892 8596 24948 8606
rect 23884 7644 24388 7700
rect 24444 8036 24500 8046
rect 24444 7700 24500 7980
rect 23884 6804 23940 7644
rect 24444 7634 24500 7644
rect 24668 8036 24724 8046
rect 23996 7476 24052 7486
rect 23996 6916 24052 7420
rect 24668 7252 24724 7980
rect 24332 7196 24724 7252
rect 24332 7140 24388 7196
rect 24332 7074 24388 7084
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 23996 6914 24388 6916
rect 23996 6862 23998 6914
rect 24050 6862 24388 6914
rect 23996 6860 24388 6862
rect 23996 6850 24052 6860
rect 23884 6738 23940 6748
rect 24332 6804 24388 6860
rect 23436 6412 23716 6468
rect 23436 5348 23492 6412
rect 23804 6300 24068 6310
rect 23548 6244 23604 6254
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24220 6244 24276 6254
rect 23548 6020 23604 6188
rect 23548 5964 23940 6020
rect 23772 5348 23828 5358
rect 23436 5346 23828 5348
rect 23436 5294 23774 5346
rect 23826 5294 23828 5346
rect 23436 5292 23828 5294
rect 23884 5348 23940 5964
rect 24220 5460 24276 6188
rect 24332 6020 24388 6748
rect 24780 6692 24836 6702
rect 24892 6692 24948 8540
rect 25004 7140 25060 8764
rect 25004 7074 25060 7084
rect 24780 6690 24948 6692
rect 24780 6638 24782 6690
rect 24834 6638 24948 6690
rect 24780 6636 24948 6638
rect 24780 6626 24836 6636
rect 24332 6018 24724 6020
rect 24332 5966 24334 6018
rect 24386 5966 24724 6018
rect 24332 5964 24724 5966
rect 24332 5954 24388 5964
rect 24668 5906 24724 5964
rect 24668 5854 24670 5906
rect 24722 5854 24724 5906
rect 24668 5842 24724 5854
rect 24220 5394 24276 5404
rect 24332 5572 24388 5582
rect 23996 5348 24052 5358
rect 23884 5292 23996 5348
rect 23436 5234 23492 5292
rect 23772 5282 23828 5292
rect 23996 5282 24052 5292
rect 23436 5182 23438 5234
rect 23490 5182 23492 5234
rect 23436 5170 23492 5182
rect 23548 5012 23604 5022
rect 23324 3826 23380 3836
rect 23436 4340 23492 4350
rect 23436 3332 23492 4284
rect 23436 3266 23492 3276
rect 22428 2146 22484 2156
rect 22988 3220 23044 3230
rect 21644 1362 21700 1372
rect 22988 1204 23044 3164
rect 23324 2324 23380 2334
rect 23100 2212 23156 2222
rect 23100 2118 23156 2156
rect 22988 1138 23044 1148
rect 23324 1204 23380 2268
rect 23436 2212 23492 2222
rect 23436 2118 23492 2156
rect 23436 1764 23492 1774
rect 23548 1764 23604 4956
rect 24332 4788 24388 5516
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23804 4732 24068 4742
rect 23660 4676 23716 4686
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24332 4722 24388 4732
rect 24668 4900 24724 4910
rect 23804 4666 24068 4676
rect 23660 4564 23716 4620
rect 24444 4564 24500 4574
rect 23660 4508 24444 4564
rect 24444 4498 24500 4508
rect 24668 4340 24724 4844
rect 24332 4284 24724 4340
rect 24220 4228 24276 4238
rect 23660 3668 23716 3678
rect 23660 3108 23716 3612
rect 24220 3220 24276 4172
rect 24332 4004 24388 4284
rect 24332 3938 24388 3948
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24220 3154 24276 3164
rect 24892 3388 24948 6636
rect 25116 6916 25172 6926
rect 25116 6018 25172 6860
rect 25228 6804 25284 6814
rect 25228 6710 25284 6748
rect 25116 5966 25118 6018
rect 25170 5966 25172 6018
rect 25116 5954 25172 5966
rect 25340 5012 25396 9996
rect 25452 9940 25508 12236
rect 26012 12180 26068 12798
rect 26236 12628 26292 14112
rect 26236 12562 26292 12572
rect 26460 14084 26516 14094
rect 26236 12180 26292 12190
rect 26012 12178 26292 12180
rect 26012 12126 26238 12178
rect 26290 12126 26292 12178
rect 26012 12124 26292 12126
rect 25900 12068 25956 12078
rect 25900 11974 25956 12012
rect 25564 11508 25620 11518
rect 25564 10724 25620 11452
rect 25676 11508 25732 11518
rect 26012 11508 26068 12124
rect 26236 12114 26292 12124
rect 25676 11506 26068 11508
rect 25676 11454 25678 11506
rect 25730 11454 26014 11506
rect 26066 11454 26068 11506
rect 25676 11452 26068 11454
rect 25676 11442 25732 11452
rect 26012 11442 26068 11452
rect 26348 11956 26404 11966
rect 26124 11394 26180 11406
rect 26124 11342 26126 11394
rect 26178 11342 26180 11394
rect 25676 10948 25732 10958
rect 26012 10948 26068 10958
rect 25732 10892 25844 10948
rect 25676 10882 25732 10892
rect 25676 10724 25732 10734
rect 25564 10722 25732 10724
rect 25564 10670 25678 10722
rect 25730 10670 25732 10722
rect 25564 10668 25732 10670
rect 25676 10500 25732 10668
rect 25676 10434 25732 10444
rect 25452 9268 25508 9884
rect 25452 9202 25508 9212
rect 25340 4946 25396 4956
rect 25452 8932 25508 8942
rect 25452 3388 25508 8876
rect 25788 7476 25844 10892
rect 26012 10050 26068 10892
rect 26012 9998 26014 10050
rect 26066 9998 26068 10050
rect 26012 9716 26068 9998
rect 26012 9650 26068 9660
rect 26124 9492 26180 11342
rect 26236 10610 26292 10622
rect 26236 10558 26238 10610
rect 26290 10558 26292 10610
rect 26236 10276 26292 10558
rect 26236 10210 26292 10220
rect 26348 9940 26404 11900
rect 26460 11620 26516 14028
rect 26572 13972 26628 13982
rect 26572 11732 26628 13916
rect 26684 13748 26740 14112
rect 26684 13682 26740 13692
rect 26796 13972 26852 13982
rect 26796 13300 26852 13916
rect 26796 13234 26852 13244
rect 27132 12292 27188 14112
rect 27356 13748 27412 13758
rect 27132 12226 27188 12236
rect 27244 12516 27300 12526
rect 27020 12068 27076 12078
rect 27020 12066 27188 12068
rect 27020 12014 27022 12066
rect 27074 12014 27188 12066
rect 27020 12012 27188 12014
rect 27020 12002 27076 12012
rect 26572 11676 26964 11732
rect 26460 11564 26852 11620
rect 26796 11284 26852 11564
rect 26684 11228 26852 11284
rect 26572 11172 26628 11182
rect 26460 11170 26628 11172
rect 26460 11118 26574 11170
rect 26626 11118 26628 11170
rect 26460 11116 26628 11118
rect 26460 10276 26516 11116
rect 26572 11106 26628 11116
rect 26572 10500 26628 10510
rect 26572 10406 26628 10444
rect 26460 10210 26516 10220
rect 26684 9940 26740 11228
rect 26348 9884 26516 9940
rect 26348 9716 26404 9726
rect 26236 9714 26404 9716
rect 26236 9662 26350 9714
rect 26402 9662 26404 9714
rect 26236 9660 26404 9662
rect 26236 9604 26292 9660
rect 26348 9650 26404 9660
rect 26236 9538 26292 9548
rect 26012 9436 26180 9492
rect 26012 8148 26068 9436
rect 26012 8082 26068 8092
rect 26124 8932 26180 8942
rect 25788 7410 25844 7420
rect 25676 5796 25732 5806
rect 25676 5702 25732 5740
rect 25676 5572 25732 5582
rect 25676 5236 25732 5516
rect 25676 5170 25732 5180
rect 26012 3892 26068 3902
rect 24892 3332 25060 3388
rect 25452 3332 25620 3388
rect 24892 3276 25284 3332
rect 23804 3098 24068 3108
rect 23660 3042 23716 3052
rect 24780 2884 24836 2894
rect 24780 2790 24836 2828
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24332 2212 24388 2222
rect 23996 1876 24052 1886
rect 23996 1874 24276 1876
rect 23996 1822 23998 1874
rect 24050 1822 24276 1874
rect 23996 1820 24276 1822
rect 23996 1810 24052 1820
rect 23492 1708 23604 1764
rect 23436 1698 23492 1708
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 23324 1138 23380 1148
rect 23548 1428 23604 1438
rect 18956 130 19012 140
rect 19516 1092 19572 1102
rect 19516 112 19572 1036
rect 21532 1092 21588 1102
rect 21532 112 21588 1036
rect 23548 112 23604 1372
rect 23996 980 24052 990
rect 23996 308 24052 924
rect 24220 980 24276 1820
rect 24332 1314 24388 2156
rect 24780 1988 24836 1998
rect 24892 1988 24948 3276
rect 25116 2772 25172 2782
rect 25116 2548 25172 2716
rect 25228 2770 25284 3276
rect 25228 2718 25230 2770
rect 25282 2718 25284 2770
rect 25228 2706 25284 2718
rect 25116 2492 25284 2548
rect 25116 2212 25172 2222
rect 25116 2098 25172 2156
rect 25116 2046 25118 2098
rect 25170 2046 25172 2098
rect 25116 2034 25172 2046
rect 24780 1986 24948 1988
rect 24780 1934 24782 1986
rect 24834 1934 24948 1986
rect 24780 1932 24948 1934
rect 24780 1922 24836 1932
rect 25228 1652 25284 2492
rect 25564 2324 25620 3332
rect 26012 3332 26068 3836
rect 26012 3266 26068 3276
rect 25564 2258 25620 2268
rect 25676 2884 25732 2894
rect 25676 2658 25732 2828
rect 25676 2606 25678 2658
rect 25730 2606 25732 2658
rect 25228 1586 25284 1596
rect 24332 1262 24334 1314
rect 24386 1262 24388 1314
rect 24332 1250 24388 1262
rect 25228 1316 25284 1326
rect 25676 1316 25732 2606
rect 26012 2884 26068 2894
rect 25788 1764 25844 1774
rect 25788 1428 25844 1708
rect 26012 1540 26068 2828
rect 26012 1474 26068 1484
rect 25788 1362 25844 1372
rect 25228 1314 25732 1316
rect 25228 1262 25230 1314
rect 25282 1262 25732 1314
rect 25228 1260 25732 1262
rect 25228 1250 25284 1260
rect 25676 1202 25732 1260
rect 26124 1314 26180 8876
rect 26460 8036 26516 9884
rect 26572 9884 26740 9940
rect 26572 9044 26628 9884
rect 26572 8978 26628 8988
rect 26684 9602 26740 9614
rect 26684 9550 26686 9602
rect 26738 9550 26740 9602
rect 26684 9042 26740 9550
rect 26684 8990 26686 9042
rect 26738 8990 26740 9042
rect 26684 8978 26740 8990
rect 26796 9044 26852 9054
rect 26460 7970 26516 7980
rect 26460 6580 26516 6590
rect 26348 6466 26404 6478
rect 26348 6414 26350 6466
rect 26402 6414 26404 6466
rect 26236 5908 26292 5918
rect 26236 5814 26292 5852
rect 26348 5796 26404 6414
rect 26460 6020 26516 6524
rect 26796 6132 26852 8988
rect 26908 6692 26964 11676
rect 27020 11172 27076 11182
rect 27020 10948 27076 11116
rect 27020 10882 27076 10892
rect 27020 9604 27076 9614
rect 27020 9510 27076 9548
rect 27132 9268 27188 12012
rect 27244 9492 27300 12460
rect 27244 9426 27300 9436
rect 27356 9380 27412 13692
rect 27468 12628 27524 12638
rect 27468 11620 27524 12572
rect 27580 11844 27636 14112
rect 28028 13860 28084 14112
rect 28028 13794 28084 13804
rect 27580 11778 27636 11788
rect 27692 13524 27748 13534
rect 27468 11554 27524 11564
rect 27580 11394 27636 11406
rect 27580 11342 27582 11394
rect 27634 11342 27636 11394
rect 27580 10500 27636 11342
rect 27580 10434 27636 10444
rect 27580 9938 27636 9950
rect 27580 9886 27582 9938
rect 27634 9886 27636 9938
rect 27580 9716 27636 9886
rect 27580 9650 27636 9660
rect 27356 9314 27412 9324
rect 27020 9212 27188 9268
rect 27020 8596 27076 9212
rect 27020 8530 27076 8540
rect 27244 8930 27300 8942
rect 27244 8878 27246 8930
rect 27298 8878 27300 8930
rect 27244 8484 27300 8878
rect 27244 8418 27300 8428
rect 27692 7924 27748 13468
rect 28252 13188 28308 13198
rect 28140 11282 28196 11294
rect 28140 11230 28142 11282
rect 28194 11230 28196 11282
rect 28140 11172 28196 11230
rect 28140 11106 28196 11116
rect 27804 10386 27860 10398
rect 27804 10334 27806 10386
rect 27858 10334 27860 10386
rect 27804 9826 27860 10334
rect 28252 10018 28308 13132
rect 28476 12180 28532 14112
rect 28924 13412 28980 14112
rect 28924 13346 28980 13356
rect 28476 12114 28532 12124
rect 28700 12516 28756 12526
rect 28364 11282 28420 11294
rect 28364 11230 28366 11282
rect 28418 11230 28420 11282
rect 28364 10500 28420 11230
rect 28700 10724 28756 12460
rect 29372 12292 29428 14112
rect 29372 12226 29428 12236
rect 29484 12180 29540 12190
rect 29260 11844 29316 11854
rect 28700 10658 28756 10668
rect 28924 11732 28980 11742
rect 28364 10434 28420 10444
rect 28588 10276 28644 10286
rect 28588 10052 28644 10220
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 28140 9962 28308 10018
rect 28364 9996 28644 10052
rect 28028 8372 28084 8382
rect 28028 8278 28084 8316
rect 27692 7858 27748 7868
rect 27020 6692 27076 6702
rect 26908 6636 27020 6692
rect 27020 6626 27076 6636
rect 26796 6066 26852 6076
rect 27020 6132 27076 6142
rect 28140 6132 28196 9962
rect 28252 9828 28308 9838
rect 28252 6916 28308 9772
rect 28252 6850 28308 6860
rect 28364 6804 28420 9996
rect 28812 9380 28868 9390
rect 28812 9156 28868 9324
rect 28588 9154 28868 9156
rect 28588 9102 28814 9154
rect 28866 9102 28868 9154
rect 28588 9100 28868 9102
rect 28588 8482 28644 9100
rect 28588 8430 28590 8482
rect 28642 8430 28644 8482
rect 28588 8418 28644 8430
rect 28700 8708 28756 8718
rect 28476 8372 28532 8382
rect 28476 7028 28532 8316
rect 28476 6962 28532 6972
rect 28588 7250 28644 7262
rect 28588 7198 28590 7250
rect 28642 7198 28644 7250
rect 28364 6738 28420 6748
rect 28588 6804 28644 7198
rect 28588 6738 28644 6748
rect 28476 6692 28532 6702
rect 28476 6468 28532 6636
rect 28476 6402 28532 6412
rect 27020 6130 27188 6132
rect 27020 6078 27022 6130
rect 27074 6078 27188 6130
rect 27020 6076 27188 6078
rect 27020 6066 27076 6076
rect 27132 6020 27188 6076
rect 27580 6076 28532 6132
rect 27132 5964 27412 6020
rect 26460 5954 26516 5964
rect 26348 5730 26404 5740
rect 26572 5908 26628 5918
rect 26236 5348 26292 5358
rect 26236 3108 26292 5292
rect 26572 5346 26628 5852
rect 27356 5908 27412 5964
rect 27356 5842 27412 5852
rect 27580 5908 27636 6076
rect 27580 5842 27636 5852
rect 27132 5796 27188 5806
rect 26572 5294 26574 5346
rect 26626 5294 26628 5346
rect 26572 5282 26628 5294
rect 26684 5682 26740 5694
rect 26684 5630 26686 5682
rect 26738 5630 26740 5682
rect 26684 5124 26740 5630
rect 27132 5684 27188 5740
rect 27244 5794 27300 5806
rect 27244 5742 27246 5794
rect 27298 5742 27300 5794
rect 27244 5684 27300 5742
rect 27132 5628 27300 5684
rect 27692 5794 27748 5806
rect 27692 5742 27694 5794
rect 27746 5742 27748 5794
rect 27692 5684 27748 5742
rect 27692 5618 27748 5628
rect 28252 5796 28308 5806
rect 28252 5346 28308 5740
rect 28252 5294 28254 5346
rect 28306 5294 28308 5346
rect 28252 5282 28308 5294
rect 28364 5684 28420 5694
rect 26684 5058 26740 5068
rect 27580 5124 27636 5134
rect 27804 5124 27860 5134
rect 27468 5012 27524 5022
rect 26908 4900 26964 4910
rect 26908 4788 26964 4844
rect 27468 4788 27524 4956
rect 26908 4732 27524 4788
rect 27580 4338 27636 5068
rect 27580 4286 27582 4338
rect 27634 4286 27636 4338
rect 27580 4274 27636 4286
rect 27692 5068 27804 5124
rect 26572 4228 26628 4238
rect 26236 3042 26292 3052
rect 26348 3556 26404 3566
rect 26348 2210 26404 3500
rect 26348 2158 26350 2210
rect 26402 2158 26404 2210
rect 26348 2146 26404 2158
rect 26124 1262 26126 1314
rect 26178 1262 26180 1314
rect 26124 1250 26180 1262
rect 25676 1150 25678 1202
rect 25730 1150 25732 1202
rect 25676 1138 25732 1150
rect 24220 914 24276 924
rect 25564 868 25620 878
rect 24464 812 24728 822
rect 24332 756 24388 766
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24892 756 24948 766
rect 24332 644 24388 700
rect 24892 644 24948 700
rect 24332 588 24948 644
rect 23996 242 24052 252
rect 25564 112 25620 812
rect 26572 308 26628 4172
rect 27020 4226 27076 4238
rect 27020 4174 27022 4226
rect 27074 4174 27076 4226
rect 26908 3780 26964 3790
rect 27020 3780 27076 4174
rect 26908 3778 27076 3780
rect 26908 3726 26910 3778
rect 26962 3726 27076 3778
rect 26908 3724 27076 3726
rect 27244 4226 27300 4238
rect 27244 4174 27246 4226
rect 27298 4174 27300 4226
rect 27244 3778 27300 4174
rect 27244 3726 27246 3778
rect 27298 3726 27300 3778
rect 26908 3714 26964 3724
rect 27244 3714 27300 3726
rect 27356 4116 27412 4126
rect 27356 3666 27412 4060
rect 27356 3614 27358 3666
rect 27410 3614 27412 3666
rect 26796 3556 26852 3566
rect 26796 3462 26852 3500
rect 26684 3444 26740 3454
rect 27356 3388 27412 3614
rect 27468 4114 27524 4126
rect 27692 4116 27748 5068
rect 27804 5058 27860 5068
rect 27468 4062 27470 4114
rect 27522 4062 27524 4114
rect 27468 3668 27524 4062
rect 27468 3602 27524 3612
rect 27580 4060 27748 4116
rect 27804 4228 27860 4238
rect 26684 2772 26740 3388
rect 26908 3332 27412 3388
rect 26908 2994 26964 3332
rect 26908 2942 26910 2994
rect 26962 2942 26964 2994
rect 26908 2930 26964 2942
rect 27020 3220 27076 3230
rect 27020 2772 27076 3164
rect 26684 2716 27076 2772
rect 26796 2100 26852 2110
rect 26796 1092 26852 2044
rect 26796 1026 26852 1036
rect 26572 242 26628 252
rect 27580 112 27636 4060
rect 27804 4004 27860 4172
rect 27692 3948 27860 4004
rect 27692 2996 27748 3948
rect 27692 2930 27748 2940
rect 27804 3780 27860 3790
rect 27804 196 27860 3724
rect 28364 3108 28420 5628
rect 28476 5346 28532 6076
rect 28588 6020 28644 6030
rect 28700 6020 28756 8652
rect 28812 7700 28868 9100
rect 28924 8370 28980 11676
rect 29260 9828 29316 11788
rect 29260 9762 29316 9772
rect 29372 10500 29428 10510
rect 28924 8318 28926 8370
rect 28978 8318 28980 8370
rect 28924 8306 28980 8318
rect 29372 8372 29428 10444
rect 29484 9268 29540 12124
rect 29820 11956 29876 14112
rect 30044 13860 30100 14140
rect 30240 14112 30352 14224
rect 30688 14112 30800 14224
rect 31136 14112 31248 14224
rect 31584 14112 31696 14224
rect 32032 14112 32144 14224
rect 32480 14112 32592 14224
rect 32928 14112 33040 14224
rect 33376 14112 33488 14224
rect 33824 14112 33936 14224
rect 34272 14112 34384 14224
rect 34720 14112 34832 14224
rect 35168 14112 35280 14224
rect 35616 14112 35728 14224
rect 36064 14112 36176 14224
rect 36512 14112 36624 14224
rect 36960 14112 37072 14224
rect 37408 14112 37520 14224
rect 37856 14112 37968 14224
rect 38304 14112 38416 14224
rect 38752 14112 38864 14224
rect 39200 14112 39312 14224
rect 39648 14112 39760 14224
rect 40096 14112 40208 14224
rect 40544 14112 40656 14224
rect 40992 14112 41104 14224
rect 41440 14112 41552 14224
rect 41888 14112 42000 14224
rect 42336 14112 42448 14224
rect 42784 14112 42896 14224
rect 43232 14112 43344 14224
rect 43680 14112 43792 14224
rect 44128 14112 44240 14224
rect 44576 14112 44688 14224
rect 45024 14112 45136 14224
rect 45472 14112 45584 14224
rect 45920 14112 46032 14224
rect 46368 14112 46480 14224
rect 46816 14112 46928 14224
rect 47264 14112 47376 14224
rect 47712 14112 47824 14224
rect 48160 14112 48272 14224
rect 48608 14112 48720 14224
rect 49056 14112 49168 14224
rect 49504 14112 49616 14224
rect 49952 14112 50064 14224
rect 50400 14112 50512 14224
rect 50848 14112 50960 14224
rect 51296 14112 51408 14224
rect 51744 14112 51856 14224
rect 52192 14112 52304 14224
rect 52640 14112 52752 14224
rect 53088 14112 53200 14224
rect 53536 14112 53648 14224
rect 53984 14112 54096 14224
rect 54432 14112 54544 14224
rect 54880 14112 54992 14224
rect 55328 14112 55440 14224
rect 55776 14112 55888 14224
rect 56224 14112 56336 14224
rect 56672 14112 56784 14224
rect 30044 13794 30100 13804
rect 29820 11890 29876 11900
rect 30156 12404 30212 12414
rect 29820 10948 29876 10958
rect 29596 10388 29652 10398
rect 29596 10386 29764 10388
rect 29596 10334 29598 10386
rect 29650 10334 29764 10386
rect 29596 10332 29764 10334
rect 29596 10322 29652 10332
rect 29708 10276 29764 10332
rect 29708 10050 29764 10220
rect 29708 9998 29710 10050
rect 29762 9998 29764 10050
rect 29708 9986 29764 9998
rect 29484 9202 29540 9212
rect 29820 9044 29876 10892
rect 30156 10724 30212 12348
rect 30156 10658 30212 10668
rect 29932 10610 29988 10622
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29932 9940 29988 10558
rect 30044 10276 30100 10286
rect 30044 10050 30100 10220
rect 30044 9998 30046 10050
rect 30098 9998 30100 10050
rect 30044 9986 30100 9998
rect 29932 9874 29988 9884
rect 30156 9940 30212 9950
rect 29820 8978 29876 8988
rect 29708 8372 29764 8382
rect 29372 8370 29764 8372
rect 29372 8318 29710 8370
rect 29762 8318 29764 8370
rect 29372 8316 29764 8318
rect 29372 8258 29428 8316
rect 29372 8206 29374 8258
rect 29426 8206 29428 8258
rect 29372 8194 29428 8206
rect 29596 7812 29652 7822
rect 28924 7700 28980 7710
rect 28812 7698 28980 7700
rect 28812 7646 28926 7698
rect 28978 7646 28980 7698
rect 28812 7644 28980 7646
rect 28924 7634 28980 7644
rect 28588 6018 28756 6020
rect 28588 5966 28590 6018
rect 28642 5966 28756 6018
rect 28588 5964 28756 5966
rect 28812 7476 28868 7486
rect 28588 5954 28644 5964
rect 28812 5908 28868 7420
rect 29148 7362 29204 7374
rect 29148 7310 29150 7362
rect 29202 7310 29204 7362
rect 28476 5294 28478 5346
rect 28530 5294 28532 5346
rect 28476 5282 28532 5294
rect 28700 5852 28868 5908
rect 28924 6804 28980 6814
rect 28700 5124 28756 5852
rect 28476 5012 28532 5022
rect 28476 4338 28532 4956
rect 28476 4286 28478 4338
rect 28530 4286 28532 4338
rect 28476 4274 28532 4286
rect 28588 4116 28644 4126
rect 28588 4022 28644 4060
rect 28700 3892 28756 5068
rect 28812 5684 28868 5694
rect 28812 4340 28868 5628
rect 28924 5012 28980 6748
rect 29148 5908 29204 7310
rect 29036 5796 29092 5806
rect 29036 5702 29092 5740
rect 28924 4946 28980 4956
rect 28812 4274 28868 4284
rect 28812 4116 28868 4126
rect 28812 4114 28980 4116
rect 28812 4062 28814 4114
rect 28866 4062 28980 4114
rect 28812 4060 28980 4062
rect 28812 4050 28868 4060
rect 28364 2882 28420 3052
rect 28364 2830 28366 2882
rect 28418 2830 28420 2882
rect 28364 2818 28420 2830
rect 28588 3836 28756 3892
rect 28588 2884 28644 3836
rect 28700 3668 28756 3678
rect 28700 3574 28756 3612
rect 28924 3554 28980 4060
rect 28924 3502 28926 3554
rect 28978 3502 28980 3554
rect 28924 3490 28980 3502
rect 28812 3442 28868 3454
rect 28812 3390 28814 3442
rect 28866 3390 28868 3442
rect 28700 2884 28756 2894
rect 28588 2882 28756 2884
rect 28588 2830 28702 2882
rect 28754 2830 28756 2882
rect 28588 2828 28756 2830
rect 28700 2818 28756 2828
rect 28812 2436 28868 3390
rect 28812 2370 28868 2380
rect 28924 2884 28980 2894
rect 28700 2212 28756 2222
rect 28924 2212 28980 2828
rect 29148 2772 29204 5852
rect 29260 7364 29316 7374
rect 29260 6018 29316 7308
rect 29260 5966 29262 6018
rect 29314 5966 29316 6018
rect 29260 5796 29316 5966
rect 29260 5730 29316 5740
rect 29596 4340 29652 7756
rect 29708 7588 29764 8316
rect 30044 7588 30100 7598
rect 29708 7586 30100 7588
rect 29708 7534 30046 7586
rect 30098 7534 30100 7586
rect 29708 7532 30100 7534
rect 29708 7362 29764 7532
rect 30044 7522 30100 7532
rect 29708 7310 29710 7362
rect 29762 7310 29764 7362
rect 29708 7298 29764 7310
rect 30044 6916 30100 6926
rect 29820 5908 29876 5918
rect 29708 5796 29764 5806
rect 29708 5124 29764 5740
rect 29708 5058 29764 5068
rect 29596 4274 29652 4284
rect 29708 3666 29764 3678
rect 29708 3614 29710 3666
rect 29762 3614 29764 3666
rect 29260 3554 29316 3566
rect 29260 3502 29262 3554
rect 29314 3502 29316 3554
rect 29260 3444 29316 3502
rect 29708 3556 29764 3614
rect 29708 3490 29764 3500
rect 29596 3444 29652 3454
rect 29260 3442 29652 3444
rect 29260 3390 29598 3442
rect 29650 3390 29652 3442
rect 29260 3388 29652 3390
rect 29596 3378 29652 3388
rect 29484 2996 29540 3006
rect 29260 2772 29316 2782
rect 29148 2770 29316 2772
rect 29148 2718 29262 2770
rect 29314 2718 29316 2770
rect 29148 2716 29316 2718
rect 29260 2706 29316 2716
rect 29036 2212 29092 2222
rect 28700 2210 29092 2212
rect 28700 2158 28702 2210
rect 28754 2158 29038 2210
rect 29090 2158 29092 2210
rect 28700 2156 29092 2158
rect 28700 2146 28756 2156
rect 29036 2146 29092 2156
rect 28140 1988 28196 1998
rect 28140 1894 28196 1932
rect 28476 1988 28532 1998
rect 28476 1204 28532 1932
rect 29484 1428 29540 2940
rect 29820 2884 29876 5852
rect 29932 5684 29988 5694
rect 29932 5590 29988 5628
rect 29820 2818 29876 2828
rect 29932 3330 29988 3342
rect 29932 3278 29934 3330
rect 29986 3278 29988 3330
rect 29708 2770 29764 2782
rect 29708 2718 29710 2770
rect 29762 2718 29764 2770
rect 29708 2212 29764 2718
rect 29932 2658 29988 3278
rect 30044 2884 30100 6860
rect 30156 5348 30212 9884
rect 30268 5908 30324 14112
rect 30716 12516 30772 14112
rect 30940 13860 30996 13870
rect 30716 12450 30772 12460
rect 30828 13412 30884 13422
rect 30492 11620 30548 11630
rect 30380 10498 30436 10510
rect 30380 10446 30382 10498
rect 30434 10446 30436 10498
rect 30380 10276 30436 10446
rect 30380 10210 30436 10220
rect 30380 9380 30436 9390
rect 30380 7586 30436 9324
rect 30380 7534 30382 7586
rect 30434 7534 30436 7586
rect 30380 7522 30436 7534
rect 30492 7364 30548 11564
rect 30604 9716 30660 9726
rect 30604 9622 30660 9660
rect 30716 9492 30772 9502
rect 30716 9154 30772 9436
rect 30828 9380 30884 13356
rect 30940 10500 30996 13804
rect 31052 12292 31108 12302
rect 31052 12198 31108 12236
rect 30940 10434 30996 10444
rect 31164 10276 31220 14112
rect 31612 13636 31668 14112
rect 31612 13570 31668 13580
rect 31724 12962 31780 12974
rect 31724 12910 31726 12962
rect 31778 12910 31780 12962
rect 31388 12852 31444 12862
rect 31388 12758 31444 12796
rect 31724 12852 31780 12910
rect 31724 12786 31780 12796
rect 31836 12178 31892 12190
rect 31836 12126 31838 12178
rect 31890 12126 31892 12178
rect 31388 12066 31444 12078
rect 31388 12014 31390 12066
rect 31442 12014 31444 12066
rect 31388 11844 31444 12014
rect 31388 11778 31444 11788
rect 31836 11284 31892 12126
rect 32060 11508 32116 14112
rect 32508 14084 32564 14112
rect 32508 14018 32564 14028
rect 32284 12852 32340 12862
rect 32284 12758 32340 12796
rect 32508 12516 32564 12526
rect 32284 12292 32340 12302
rect 32284 12178 32340 12236
rect 32284 12126 32286 12178
rect 32338 12126 32340 12178
rect 32284 12114 32340 12126
rect 32060 11452 32452 11508
rect 32284 11284 32340 11294
rect 31836 11282 32340 11284
rect 31836 11230 32286 11282
rect 32338 11230 32340 11282
rect 31836 11228 32340 11230
rect 32172 11060 32228 11070
rect 31612 10388 31668 10398
rect 31612 10386 31892 10388
rect 31612 10334 31614 10386
rect 31666 10334 31892 10386
rect 31612 10332 31892 10334
rect 31612 10322 31668 10332
rect 31164 10210 31220 10220
rect 31276 10052 31332 10062
rect 30828 9314 30884 9324
rect 30940 9604 30996 9614
rect 30716 9102 30718 9154
rect 30770 9102 30772 9154
rect 30716 9044 30772 9102
rect 30940 9154 30996 9548
rect 30940 9102 30942 9154
rect 30994 9102 30996 9154
rect 30940 9090 30996 9102
rect 30716 8978 30772 8988
rect 31276 8932 31332 9996
rect 31276 8866 31332 8876
rect 31724 9604 31780 9614
rect 31724 9266 31780 9548
rect 31724 9214 31726 9266
rect 31778 9214 31780 9266
rect 31388 8820 31444 8830
rect 31388 8818 31668 8820
rect 31388 8766 31390 8818
rect 31442 8766 31668 8818
rect 31388 8764 31668 8766
rect 31388 8754 31444 8764
rect 31500 8596 31556 8606
rect 31164 8148 31220 8158
rect 31164 8054 31220 8092
rect 30492 7298 30548 7308
rect 31388 7028 31444 7038
rect 31276 6578 31332 6590
rect 31276 6526 31278 6578
rect 31330 6526 31332 6578
rect 30268 5842 30324 5852
rect 30380 5906 30436 5918
rect 30380 5854 30382 5906
rect 30434 5854 30436 5906
rect 30380 5572 30436 5854
rect 30828 5794 30884 5806
rect 30828 5742 30830 5794
rect 30882 5742 30884 5794
rect 30380 5506 30436 5516
rect 30716 5684 30772 5694
rect 30828 5684 30884 5742
rect 30772 5628 30884 5684
rect 30156 5292 30324 5348
rect 30156 5124 30212 5134
rect 30156 4564 30212 5068
rect 30156 4498 30212 4508
rect 30268 4340 30324 5292
rect 30716 5346 30772 5628
rect 30716 5294 30718 5346
rect 30770 5294 30772 5346
rect 30716 5282 30772 5294
rect 30828 5348 30884 5628
rect 30940 5348 30996 5358
rect 30828 5346 30996 5348
rect 30828 5294 30942 5346
rect 30994 5294 30996 5346
rect 30828 5292 30996 5294
rect 30940 5282 30996 5292
rect 31276 5348 31332 6526
rect 31388 5460 31444 6972
rect 31500 6468 31556 8540
rect 31612 8258 31668 8764
rect 31612 8206 31614 8258
rect 31666 8206 31668 8258
rect 31612 8194 31668 8206
rect 31724 6692 31780 9214
rect 31836 8932 31892 10332
rect 31948 8932 32004 8942
rect 31836 8930 32004 8932
rect 31836 8878 31950 8930
rect 32002 8878 32004 8930
rect 31836 8876 32004 8878
rect 31948 8866 32004 8876
rect 32172 7476 32228 11004
rect 32284 9492 32340 11228
rect 32284 9426 32340 9436
rect 32284 9044 32340 9054
rect 32284 8930 32340 8988
rect 32284 8878 32286 8930
rect 32338 8878 32340 8930
rect 32284 8866 32340 8878
rect 32396 7476 32452 11452
rect 32508 10836 32564 12460
rect 32844 12066 32900 12078
rect 32844 12014 32846 12066
rect 32898 12014 32900 12066
rect 32508 10770 32564 10780
rect 32620 11732 32676 11742
rect 32508 9604 32564 9614
rect 32508 8820 32564 9548
rect 32508 8754 32564 8764
rect 32620 7700 32676 11676
rect 32844 10948 32900 12014
rect 32956 11788 33012 14112
rect 32956 11732 33348 11788
rect 32844 10882 32900 10892
rect 33292 10948 33348 11732
rect 33292 10882 33348 10892
rect 33404 10612 33460 14112
rect 33852 11620 33908 14112
rect 33852 11554 33908 11564
rect 33852 11284 33908 11294
rect 34300 11284 34356 14112
rect 34748 11732 34804 14112
rect 34748 11666 34804 11676
rect 34860 12068 34916 12078
rect 34748 11506 34804 11518
rect 34748 11454 34750 11506
rect 34802 11454 34804 11506
rect 33852 11282 34020 11284
rect 33852 11230 33854 11282
rect 33906 11230 34020 11282
rect 33852 11228 34020 11230
rect 33852 11218 33908 11228
rect 32844 10556 33460 10612
rect 33628 11060 33684 11070
rect 32844 9156 32900 10556
rect 33628 10052 33684 11004
rect 33964 10388 34020 11228
rect 34300 11218 34356 11228
rect 34412 11282 34468 11294
rect 34412 11230 34414 11282
rect 34466 11230 34468 11282
rect 34412 11060 34468 11230
rect 34412 10994 34468 11004
rect 34524 10612 34580 10622
rect 34748 10612 34804 11454
rect 34524 10610 34804 10612
rect 34524 10558 34526 10610
rect 34578 10558 34804 10610
rect 34524 10556 34804 10558
rect 34524 10546 34580 10556
rect 34076 10388 34132 10398
rect 34412 10388 34468 10398
rect 33964 10386 34468 10388
rect 33964 10334 34078 10386
rect 34130 10334 34414 10386
rect 34466 10334 34468 10386
rect 33964 10332 34468 10334
rect 33404 9996 33908 10052
rect 33068 9268 33124 9278
rect 33068 9156 33124 9212
rect 33404 9156 33460 9996
rect 33068 9154 33460 9156
rect 33068 9102 33406 9154
rect 33458 9102 33460 9154
rect 33068 9100 33460 9102
rect 32844 9090 32900 9100
rect 33404 9090 33460 9100
rect 33628 9380 33684 9390
rect 33628 9156 33684 9324
rect 33628 9090 33684 9100
rect 33516 9044 33572 9054
rect 32844 8820 32900 8830
rect 32844 8818 33012 8820
rect 32844 8766 32846 8818
rect 32898 8766 33012 8818
rect 32844 8764 33012 8766
rect 32844 8754 32900 8764
rect 32956 8484 33012 8764
rect 33516 8708 33572 8988
rect 33404 8652 33572 8708
rect 33740 8930 33796 8942
rect 33740 8878 33742 8930
rect 33794 8878 33796 8930
rect 32956 8418 33012 8428
rect 33292 8484 33348 8494
rect 33292 8390 33348 8428
rect 33404 8260 33460 8652
rect 33516 8484 33572 8494
rect 33740 8484 33796 8878
rect 33572 8428 33796 8484
rect 33516 8390 33572 8428
rect 33404 8194 33460 8204
rect 32620 7634 32676 7644
rect 32396 7420 32900 7476
rect 32172 7410 32228 7420
rect 32732 7140 32788 7150
rect 31724 6626 31780 6636
rect 31836 6690 31892 6702
rect 31836 6638 31838 6690
rect 31890 6638 31892 6690
rect 31500 6412 31668 6468
rect 31388 5394 31444 5404
rect 31276 5282 31332 5292
rect 31500 5348 31556 5358
rect 31500 5234 31556 5292
rect 31500 5182 31502 5234
rect 31554 5182 31556 5234
rect 31500 5170 31556 5182
rect 30044 2818 30100 2828
rect 30156 4284 30324 4340
rect 29932 2606 29934 2658
rect 29986 2606 29988 2658
rect 29932 2594 29988 2606
rect 30156 2436 30212 4284
rect 30380 4116 30436 4126
rect 30380 2770 30436 4060
rect 31500 4116 31556 4126
rect 31500 3668 31556 4060
rect 31500 3602 31556 3612
rect 30380 2718 30382 2770
rect 30434 2718 30436 2770
rect 30380 2706 30436 2718
rect 30940 3108 30996 3118
rect 30940 2770 30996 3052
rect 30940 2718 30942 2770
rect 30994 2718 30996 2770
rect 30940 2706 30996 2718
rect 29708 2146 29764 2156
rect 29932 2380 30212 2436
rect 29596 1876 29652 1886
rect 29596 1782 29652 1820
rect 29484 1362 29540 1372
rect 29596 1540 29652 1550
rect 28476 1138 28532 1148
rect 27804 130 27860 140
rect 29596 112 29652 1484
rect 29932 868 29988 2380
rect 30156 2212 30212 2222
rect 30156 2118 30212 2156
rect 30492 2212 30548 2222
rect 30492 2118 30548 2156
rect 30156 1876 30212 1886
rect 29932 802 29988 812
rect 30044 1764 30100 1774
rect 30044 420 30100 1708
rect 30156 756 30212 1820
rect 30156 690 30212 700
rect 30044 354 30100 364
rect 31612 112 31668 6412
rect 31836 6132 31892 6638
rect 31836 6066 31892 6076
rect 32284 6692 32340 6702
rect 32060 5796 32116 5806
rect 32060 5702 32116 5740
rect 31836 5572 31892 5582
rect 31836 5346 31892 5516
rect 32060 5572 32116 5582
rect 31836 5294 31838 5346
rect 31890 5294 31892 5346
rect 31836 5282 31892 5294
rect 31948 5460 32004 5470
rect 31836 4228 31892 4238
rect 31948 4228 32004 5404
rect 31892 4172 32004 4228
rect 31836 4162 31892 4172
rect 31836 3668 31892 3678
rect 31836 2324 31892 3612
rect 32060 2770 32116 5516
rect 32284 5346 32340 6636
rect 32620 6132 32676 6142
rect 32620 6038 32676 6076
rect 32284 5294 32286 5346
rect 32338 5294 32340 5346
rect 32284 5282 32340 5294
rect 32396 5908 32452 5918
rect 32396 3778 32452 5852
rect 32396 3726 32398 3778
rect 32450 3726 32452 3778
rect 32396 3714 32452 3726
rect 32620 5908 32676 5918
rect 32060 2718 32062 2770
rect 32114 2718 32116 2770
rect 32060 2706 32116 2718
rect 32508 3108 32564 3118
rect 32508 2770 32564 3052
rect 32508 2718 32510 2770
rect 32562 2718 32564 2770
rect 31836 2258 31892 2268
rect 32396 2212 32452 2222
rect 32508 2212 32564 2718
rect 32396 2210 32564 2212
rect 32396 2158 32398 2210
rect 32450 2158 32564 2210
rect 32396 2156 32564 2158
rect 32396 2146 32452 2156
rect 32620 1988 32676 5852
rect 32732 5684 32788 7084
rect 32732 5618 32788 5628
rect 32732 4900 32788 4910
rect 32732 2548 32788 4844
rect 32844 3388 32900 7420
rect 33068 6916 33124 6926
rect 32956 6692 33012 6702
rect 32956 6130 33012 6636
rect 32956 6078 32958 6130
rect 33010 6078 33012 6130
rect 32956 6066 33012 6078
rect 33068 4900 33124 6860
rect 33628 6580 33684 6590
rect 33628 6132 33684 6524
rect 33852 6132 33908 9996
rect 33964 6356 34020 10332
rect 34076 10322 34132 10332
rect 34412 10322 34468 10332
rect 34860 10276 34916 12012
rect 34972 10612 35028 10622
rect 34972 10518 35028 10556
rect 34748 10220 34916 10276
rect 34524 9828 34580 9838
rect 34412 9380 34468 9390
rect 34076 8148 34132 8158
rect 34076 8054 34132 8092
rect 34300 7588 34356 7598
rect 34300 7494 34356 7532
rect 33964 6290 34020 6300
rect 33852 6076 34244 6132
rect 33628 6066 33684 6076
rect 33180 5796 33236 5806
rect 33180 5702 33236 5740
rect 33628 5794 33684 5806
rect 33628 5742 33630 5794
rect 33682 5742 33684 5794
rect 33628 5572 33684 5742
rect 33628 5506 33684 5516
rect 34188 5572 34244 6076
rect 33628 5236 33684 5246
rect 33628 5142 33684 5180
rect 34076 5236 34132 5246
rect 33068 4834 33124 4844
rect 33516 5012 33572 5022
rect 32844 3332 33348 3388
rect 33292 2882 33348 3332
rect 33516 3220 33572 4956
rect 34076 4450 34132 5180
rect 34188 5010 34244 5516
rect 34188 4958 34190 5010
rect 34242 4958 34244 5010
rect 34188 4946 34244 4958
rect 34076 4398 34078 4450
rect 34130 4398 34132 4450
rect 34076 4386 34132 4398
rect 33516 3154 33572 3164
rect 33628 3892 33684 3902
rect 33292 2830 33294 2882
rect 33346 2830 33348 2882
rect 33068 2660 33124 2670
rect 33068 2566 33124 2604
rect 32732 2482 32788 2492
rect 33292 2212 33348 2830
rect 33292 2146 33348 2156
rect 32620 1922 32676 1932
rect 32844 1988 32900 1998
rect 32844 644 32900 1932
rect 33628 756 33684 3836
rect 33628 690 33684 700
rect 33740 2436 33796 2446
rect 32844 578 32900 588
rect 33740 420 33796 2380
rect 33964 2100 34020 2110
rect 33852 1764 33908 1774
rect 33852 1540 33908 1708
rect 33852 1474 33908 1484
rect 33964 532 34020 2044
rect 33964 466 34020 476
rect 33740 354 33796 364
rect 33628 196 33684 206
rect 33628 112 33684 140
rect 34412 196 34468 9324
rect 34524 8036 34580 9772
rect 34524 7970 34580 7980
rect 34636 8146 34692 8158
rect 34636 8094 34638 8146
rect 34690 8094 34692 8146
rect 34524 5236 34580 5246
rect 34524 4338 34580 5180
rect 34636 4676 34692 8094
rect 34748 5348 34804 10220
rect 34972 8820 35028 8830
rect 34972 8726 35028 8764
rect 35196 8596 35252 14112
rect 35308 13748 35364 13758
rect 35308 13076 35364 13692
rect 35644 13188 35700 14112
rect 36092 13972 36148 14112
rect 36092 13906 36148 13916
rect 35644 13122 35700 13132
rect 35308 13010 35364 13020
rect 36204 12852 36260 12862
rect 35308 12292 35364 12302
rect 35308 11060 35364 12236
rect 35868 11844 35924 11854
rect 35308 10994 35364 11004
rect 35532 11060 35588 11070
rect 34860 8540 35252 8596
rect 34860 5908 34916 8540
rect 35084 8372 35140 8382
rect 34972 7588 35028 7598
rect 35084 7588 35140 8316
rect 35420 8036 35476 8046
rect 35308 7812 35364 7822
rect 35028 7532 35140 7588
rect 35196 7700 35252 7710
rect 35196 7586 35252 7644
rect 35196 7534 35198 7586
rect 35250 7534 35252 7586
rect 34972 7494 35028 7532
rect 35196 7522 35252 7534
rect 34860 5842 34916 5852
rect 35308 5348 35364 7756
rect 35420 7586 35476 7980
rect 35420 7534 35422 7586
rect 35474 7534 35476 7586
rect 35420 7522 35476 7534
rect 35308 5292 35476 5348
rect 34748 5282 34804 5292
rect 34636 4610 34692 4620
rect 34860 5236 34916 5246
rect 34524 4286 34526 4338
rect 34578 4286 34580 4338
rect 34524 4274 34580 4286
rect 34860 4228 34916 5180
rect 35308 5124 35364 5134
rect 35196 4340 35252 4350
rect 34860 4162 34916 4172
rect 34972 4226 35028 4238
rect 34972 4174 34974 4226
rect 35026 4174 35028 4226
rect 34972 4116 35028 4174
rect 34972 4050 35028 4060
rect 35196 3778 35252 4284
rect 35308 4228 35364 5068
rect 35308 4162 35364 4172
rect 35196 3726 35198 3778
rect 35250 3726 35252 3778
rect 35196 3332 35252 3726
rect 35420 3780 35476 5292
rect 35420 3714 35476 3724
rect 34860 2884 34916 2894
rect 35196 2884 35252 3276
rect 34860 2882 35252 2884
rect 34860 2830 34862 2882
rect 34914 2830 35252 2882
rect 34860 2828 35252 2830
rect 35532 2884 35588 11004
rect 35756 10276 35812 10286
rect 35756 9154 35812 10220
rect 35756 9102 35758 9154
rect 35810 9102 35812 9154
rect 35756 8372 35812 9102
rect 35756 7700 35812 8316
rect 35868 7812 35924 11788
rect 35980 11170 36036 11182
rect 35980 11118 35982 11170
rect 36034 11118 36036 11170
rect 35980 10948 36036 11118
rect 35980 10882 36036 10892
rect 35980 10276 36036 10286
rect 35980 8708 36036 10220
rect 35980 8642 36036 8652
rect 36092 8370 36148 8382
rect 36092 8318 36094 8370
rect 36146 8318 36148 8370
rect 36092 7924 36148 8318
rect 36092 7858 36148 7868
rect 35868 7756 36036 7812
rect 35644 7588 35700 7598
rect 35756 7588 35812 7644
rect 35868 7588 35924 7598
rect 35756 7586 35924 7588
rect 35756 7534 35870 7586
rect 35922 7534 35924 7586
rect 35756 7532 35924 7534
rect 35644 7494 35700 7532
rect 35868 7364 35924 7532
rect 35868 7298 35924 7308
rect 35756 6356 35812 6366
rect 35644 5572 35700 5582
rect 35644 3554 35700 5516
rect 35756 5346 35812 6300
rect 35980 5572 36036 7756
rect 36092 7252 36148 7262
rect 36092 6690 36148 7196
rect 36092 6638 36094 6690
rect 36146 6638 36148 6690
rect 36092 6626 36148 6638
rect 35980 5506 36036 5516
rect 35756 5294 35758 5346
rect 35810 5294 35812 5346
rect 35756 5282 35812 5294
rect 35756 5124 35812 5134
rect 35756 4788 35812 5068
rect 35756 4722 35812 4732
rect 36204 4004 36260 12796
rect 36316 12292 36372 12302
rect 36316 12178 36372 12236
rect 36316 12126 36318 12178
rect 36370 12126 36372 12178
rect 36316 12114 36372 12126
rect 36540 11396 36596 14112
rect 36988 13300 37044 14112
rect 36988 13234 37044 13244
rect 36876 13076 36932 13086
rect 36876 12290 36932 13020
rect 36876 12238 36878 12290
rect 36930 12238 36932 12290
rect 36876 12226 36932 12238
rect 36988 12404 37044 12414
rect 36540 11330 36596 11340
rect 36764 11732 36820 11742
rect 36540 10948 36596 10958
rect 36316 9044 36372 9054
rect 36316 8950 36372 8988
rect 36428 8260 36484 8270
rect 36316 8034 36372 8046
rect 36316 7982 36318 8034
rect 36370 7982 36372 8034
rect 36316 7588 36372 7982
rect 36316 7522 36372 7532
rect 36316 7364 36372 7374
rect 36316 7270 36372 7308
rect 36428 7252 36484 8204
rect 36540 7476 36596 10892
rect 36652 9044 36708 9054
rect 36652 8370 36708 8988
rect 36652 8318 36654 8370
rect 36706 8318 36708 8370
rect 36652 8306 36708 8318
rect 36652 7476 36708 7486
rect 36540 7474 36708 7476
rect 36540 7422 36654 7474
rect 36706 7422 36708 7474
rect 36540 7420 36708 7422
rect 36652 7364 36708 7420
rect 36652 7298 36708 7308
rect 36428 7186 36484 7196
rect 36764 6692 36820 11676
rect 36876 8818 36932 8830
rect 36876 8766 36878 8818
rect 36930 8766 36932 8818
rect 36876 8372 36932 8766
rect 36876 8306 36932 8316
rect 36988 8148 37044 12348
rect 37324 11954 37380 11966
rect 37324 11902 37326 11954
rect 37378 11902 37380 11954
rect 37324 11844 37380 11902
rect 37324 10388 37380 11788
rect 37436 10724 37492 14112
rect 37884 12740 37940 14112
rect 38332 13636 38388 14112
rect 38332 13570 38388 13580
rect 38780 12964 38836 14112
rect 38780 12898 38836 12908
rect 37884 12684 38052 12740
rect 37884 12292 37940 12302
rect 37884 12198 37940 12236
rect 37884 11396 37940 11406
rect 37436 10668 37604 10724
rect 37324 10322 37380 10332
rect 37436 8260 37492 8270
rect 37436 8166 37492 8204
rect 36764 6626 36820 6636
rect 36876 8092 37044 8148
rect 37212 8146 37268 8158
rect 37212 8094 37214 8146
rect 37266 8094 37268 8146
rect 36876 5236 36932 8092
rect 37212 8036 37268 8094
rect 37212 7970 37268 7980
rect 37100 7588 37156 7598
rect 37100 7474 37156 7532
rect 37100 7422 37102 7474
rect 37154 7422 37156 7474
rect 37100 7410 37156 7422
rect 37324 7250 37380 7262
rect 37324 7198 37326 7250
rect 37378 7198 37380 7250
rect 37324 6130 37380 7198
rect 37548 7252 37604 10668
rect 37772 8818 37828 8830
rect 37772 8766 37774 8818
rect 37826 8766 37828 8818
rect 37772 8260 37828 8766
rect 37772 8036 37828 8204
rect 37772 7970 37828 7980
rect 37548 7186 37604 7196
rect 37772 7362 37828 7374
rect 37772 7310 37774 7362
rect 37826 7310 37828 7362
rect 37772 6692 37828 7310
rect 37772 6356 37828 6636
rect 37884 6356 37940 11340
rect 37996 11284 38052 12684
rect 38220 12066 38276 12078
rect 38220 12014 38222 12066
rect 38274 12014 38276 12066
rect 38220 11844 38276 12014
rect 38220 11620 38276 11788
rect 38444 11620 38500 11630
rect 38220 11618 38500 11620
rect 38220 11566 38222 11618
rect 38274 11566 38446 11618
rect 38498 11566 38500 11618
rect 38220 11564 38500 11566
rect 38220 11554 38276 11564
rect 38444 11554 38500 11564
rect 37996 11218 38052 11228
rect 38332 11396 38388 11406
rect 38108 9268 38164 9278
rect 38108 9154 38164 9212
rect 38108 9102 38110 9154
rect 38162 9102 38164 9154
rect 38108 9090 38164 9102
rect 38220 9156 38276 9166
rect 37996 8372 38052 8382
rect 37996 8036 38052 8316
rect 37996 7970 38052 7980
rect 37996 6356 38052 6366
rect 37884 6300 37996 6356
rect 37772 6290 37828 6300
rect 37996 6290 38052 6300
rect 37324 6078 37326 6130
rect 37378 6078 37380 6130
rect 37324 6066 37380 6078
rect 37212 5796 37268 5806
rect 38108 5796 38164 5806
rect 37212 5794 38164 5796
rect 37212 5742 37214 5794
rect 37266 5742 38110 5794
rect 38162 5742 38164 5794
rect 37212 5740 38164 5742
rect 37212 5730 37268 5740
rect 38108 5730 38164 5740
rect 36876 5170 36932 5180
rect 37100 5682 37156 5694
rect 37100 5630 37102 5682
rect 37154 5630 37156 5682
rect 37100 5236 37156 5630
rect 37100 5170 37156 5180
rect 37436 5572 37492 5582
rect 38220 5572 38276 9100
rect 38332 7812 38388 11340
rect 39004 11282 39060 11294
rect 39004 11230 39006 11282
rect 39058 11230 39060 11282
rect 39004 9828 39060 11230
rect 39004 9762 39060 9772
rect 38556 9042 38612 9054
rect 38556 8990 38558 9042
rect 38610 8990 38612 9042
rect 38332 7746 38388 7756
rect 38444 8370 38500 8382
rect 38444 8318 38446 8370
rect 38498 8318 38500 8370
rect 38444 7924 38500 8318
rect 38444 7252 38500 7868
rect 38556 8260 38612 8990
rect 39004 8484 39060 8494
rect 39004 8390 39060 8428
rect 38668 8260 38724 8270
rect 38612 8258 38724 8260
rect 38612 8206 38670 8258
rect 38722 8206 38724 8258
rect 38612 8204 38724 8206
rect 38556 7474 38612 8204
rect 38668 8194 38724 8204
rect 38780 8260 38836 8270
rect 38780 7924 38836 8204
rect 38780 7858 38836 7868
rect 39228 7924 39284 14112
rect 39452 11954 39508 11966
rect 39452 11902 39454 11954
rect 39506 11902 39508 11954
rect 39452 10052 39508 11902
rect 39676 11060 39732 14112
rect 40124 13748 40180 14112
rect 40012 13692 40180 13748
rect 39900 12292 39956 12302
rect 39900 11732 39956 12236
rect 39900 11666 39956 11676
rect 39676 10994 39732 11004
rect 40012 10724 40068 13692
rect 40012 10658 40068 10668
rect 40124 13524 40180 13534
rect 39452 9986 39508 9996
rect 39900 10052 39956 10062
rect 39452 9044 39508 9054
rect 39452 8950 39508 8988
rect 39900 9042 39956 9996
rect 39900 8990 39902 9042
rect 39954 8990 39956 9042
rect 39900 8978 39956 8990
rect 40012 9042 40068 9054
rect 40012 8990 40014 9042
rect 40066 8990 40068 9042
rect 39676 8932 39732 8942
rect 39676 8838 39732 8876
rect 40012 8820 40068 8990
rect 40012 8754 40068 8764
rect 39564 8596 39620 8606
rect 39228 7858 39284 7868
rect 39340 8036 39396 8046
rect 38556 7422 38558 7474
rect 38610 7422 38612 7474
rect 38556 7410 38612 7422
rect 39340 7474 39396 7980
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39340 7410 39396 7422
rect 37436 4676 37492 5516
rect 37436 4610 37492 4620
rect 37996 5516 38276 5572
rect 38332 7196 38500 7252
rect 36204 3938 36260 3948
rect 37660 3780 37716 3790
rect 35644 3502 35646 3554
rect 35698 3502 35700 3554
rect 35644 3388 35700 3502
rect 36092 3666 36148 3678
rect 36092 3614 36094 3666
rect 36146 3614 36148 3666
rect 35644 3332 36036 3388
rect 35980 3108 36036 3332
rect 36092 3332 36148 3614
rect 36092 3266 36148 3276
rect 37324 3332 37380 3342
rect 37324 3238 37380 3276
rect 36764 3108 36820 3118
rect 35980 3052 36596 3108
rect 35644 2884 35700 2894
rect 35532 2882 35700 2884
rect 35532 2830 35646 2882
rect 35698 2830 35700 2882
rect 35532 2828 35700 2830
rect 34860 2818 34916 2828
rect 35196 2770 35252 2828
rect 35644 2818 35700 2828
rect 35196 2718 35198 2770
rect 35250 2718 35252 2770
rect 35196 2706 35252 2718
rect 36540 2770 36596 3052
rect 36540 2718 36542 2770
rect 36594 2718 36596 2770
rect 36540 2706 36596 2718
rect 36764 2772 36820 3052
rect 36764 2706 36820 2716
rect 36988 2658 37044 2670
rect 36988 2606 36990 2658
rect 37042 2606 37044 2658
rect 36204 2324 36260 2334
rect 36204 2212 36260 2268
rect 36428 2212 36484 2222
rect 36652 2212 36708 2222
rect 36988 2212 37044 2606
rect 36204 2210 37044 2212
rect 36204 2158 36206 2210
rect 36258 2158 36430 2210
rect 36482 2158 36654 2210
rect 36706 2158 37044 2210
rect 36204 2156 37044 2158
rect 36204 2146 36260 2156
rect 36428 2146 36484 2156
rect 36652 2146 36708 2156
rect 37100 2100 37156 2110
rect 37100 1652 37156 2044
rect 37100 1586 37156 1596
rect 37212 1874 37268 1886
rect 37212 1822 37214 1874
rect 37266 1822 37268 1874
rect 34412 130 34468 140
rect 35644 1540 35700 1550
rect 35644 112 35700 1484
rect 37212 868 37268 1822
rect 37660 1316 37716 3724
rect 37996 1874 38052 5516
rect 38220 5236 38276 5246
rect 38220 2994 38276 5180
rect 38332 3332 38388 7196
rect 38668 6916 38724 6926
rect 38556 6244 38612 6254
rect 38556 6018 38612 6188
rect 38556 5966 38558 6018
rect 38610 5966 38612 6018
rect 38556 5954 38612 5966
rect 38444 5908 38500 5918
rect 38444 5814 38500 5852
rect 38668 5796 38724 6860
rect 39452 6692 39508 6702
rect 38780 5908 38836 5918
rect 39228 5908 39284 5918
rect 38780 5906 39172 5908
rect 38780 5854 38782 5906
rect 38834 5854 39172 5906
rect 38780 5852 39172 5854
rect 38780 5842 38836 5852
rect 38668 5730 38724 5740
rect 39116 5460 39172 5852
rect 39228 5814 39284 5852
rect 39452 5794 39508 6636
rect 39564 5906 39620 8540
rect 40124 8372 40180 13468
rect 40572 11396 40628 14112
rect 41020 13860 41076 14112
rect 41020 13794 41076 13804
rect 41356 12628 41412 12638
rect 41356 12290 41412 12572
rect 41356 12238 41358 12290
rect 41410 12238 41412 12290
rect 41356 12226 41412 12238
rect 40572 11330 40628 11340
rect 41244 12180 41300 12190
rect 41244 11396 41300 12124
rect 41468 11620 41524 14112
rect 41804 13188 41860 13198
rect 41804 12180 41860 13132
rect 41916 13188 41972 14112
rect 42140 13188 42196 13198
rect 41916 13186 42084 13188
rect 41916 13134 41918 13186
rect 41970 13134 42084 13186
rect 41916 13132 42084 13134
rect 41916 13122 41972 13132
rect 41804 12086 41860 12124
rect 42028 12180 42084 13132
rect 42140 13094 42196 13132
rect 42252 12740 42308 12750
rect 42252 12290 42308 12684
rect 42364 12404 42420 14112
rect 42812 13412 42868 14112
rect 42812 13346 42868 13356
rect 42588 13188 42644 13198
rect 42364 12338 42420 12348
rect 42476 12964 42532 12974
rect 42252 12238 42254 12290
rect 42306 12238 42308 12290
rect 42252 12226 42308 12238
rect 41468 11554 41524 11564
rect 42028 11620 42084 12124
rect 42364 11620 42420 11630
rect 42028 11618 42420 11620
rect 42028 11566 42366 11618
rect 42418 11566 42420 11618
rect 42028 11564 42420 11566
rect 41916 11508 41972 11518
rect 41244 11394 41636 11396
rect 41244 11342 41246 11394
rect 41298 11342 41636 11394
rect 41244 11340 41636 11342
rect 41244 11330 41300 11340
rect 40908 11172 40964 11182
rect 40572 11170 40964 11172
rect 40572 11118 40910 11170
rect 40962 11118 40964 11170
rect 40572 11116 40964 11118
rect 40460 10388 40516 10398
rect 40460 10294 40516 10332
rect 40124 8306 40180 8316
rect 40236 9492 40292 9502
rect 40124 7700 40180 7710
rect 39564 5854 39566 5906
rect 39618 5854 39620 5906
rect 39564 5842 39620 5854
rect 39788 6244 39844 6254
rect 39452 5742 39454 5794
rect 39506 5742 39508 5794
rect 39452 5572 39508 5742
rect 39452 5516 39620 5572
rect 39116 5404 39508 5460
rect 39452 5346 39508 5404
rect 39452 5294 39454 5346
rect 39506 5294 39508 5346
rect 39452 5282 39508 5294
rect 38668 5236 38724 5246
rect 38668 5142 38724 5180
rect 38780 5124 38836 5134
rect 39116 5124 39172 5134
rect 38780 5122 39172 5124
rect 38780 5070 38782 5122
rect 38834 5070 39118 5122
rect 39170 5070 39172 5122
rect 38780 5068 39172 5070
rect 38780 5058 38836 5068
rect 39116 5058 39172 5068
rect 39452 5122 39508 5134
rect 39452 5070 39454 5122
rect 39506 5070 39508 5122
rect 39452 4562 39508 5070
rect 39452 4510 39454 4562
rect 39506 4510 39508 4562
rect 39452 4498 39508 4510
rect 38332 3266 38388 3276
rect 38444 4340 38500 4350
rect 38220 2942 38222 2994
rect 38274 2942 38276 2994
rect 38220 2930 38276 2942
rect 38444 2212 38500 4284
rect 39564 4338 39620 5516
rect 39676 5236 39732 5246
rect 39676 5142 39732 5180
rect 39564 4286 39566 4338
rect 39618 4286 39620 4338
rect 39564 4274 39620 4286
rect 39788 3388 39844 6188
rect 40124 6020 40180 7644
rect 40236 6692 40292 9436
rect 40572 8596 40628 11116
rect 40908 11106 40964 11116
rect 41580 10834 41636 11340
rect 41580 10782 41582 10834
rect 41634 10782 41636 10834
rect 41580 10770 41636 10782
rect 41692 11394 41748 11406
rect 41692 11342 41694 11394
rect 41746 11342 41748 11394
rect 40796 10500 40852 10510
rect 41244 10500 41300 10510
rect 40796 10498 41300 10500
rect 40796 10446 40798 10498
rect 40850 10446 41246 10498
rect 41298 10446 41300 10498
rect 40796 10444 41300 10446
rect 40796 10434 40852 10444
rect 41244 10434 41300 10444
rect 40684 10386 40740 10398
rect 40684 10334 40686 10386
rect 40738 10334 40740 10386
rect 40684 10052 40740 10334
rect 40684 9986 40740 9996
rect 40908 10276 40964 10286
rect 40684 8930 40740 8942
rect 40684 8878 40686 8930
rect 40738 8878 40740 8930
rect 40684 8820 40740 8878
rect 40684 8754 40740 8764
rect 40796 8818 40852 8830
rect 40796 8766 40798 8818
rect 40850 8766 40852 8818
rect 40572 8530 40628 8540
rect 40684 8372 40740 8382
rect 40684 7140 40740 8316
rect 40796 8258 40852 8766
rect 40796 8206 40798 8258
rect 40850 8206 40852 8258
rect 40796 8194 40852 8206
rect 40908 8036 40964 10220
rect 41580 10052 41636 10062
rect 41132 9044 41188 9054
rect 41132 8370 41188 8988
rect 41468 8932 41524 8942
rect 41468 8838 41524 8876
rect 41132 8318 41134 8370
rect 41186 8318 41188 8370
rect 41132 8306 41188 8318
rect 41244 8372 41300 8382
rect 40908 7970 40964 7980
rect 41020 8258 41076 8270
rect 41020 8206 41022 8258
rect 41074 8206 41076 8258
rect 40684 7074 40740 7084
rect 40796 7924 40852 7934
rect 40236 6626 40292 6636
rect 40684 6804 40740 6814
rect 40684 6690 40740 6748
rect 40684 6638 40686 6690
rect 40738 6638 40740 6690
rect 40684 6626 40740 6638
rect 40460 6578 40516 6590
rect 40460 6526 40462 6578
rect 40514 6526 40516 6578
rect 40460 6356 40516 6526
rect 40460 6290 40516 6300
rect 40124 5954 40180 5964
rect 40572 5908 40628 5918
rect 39676 3332 39844 3388
rect 40348 3892 40404 3902
rect 39004 3220 39060 3230
rect 37996 1822 37998 1874
rect 38050 1822 38052 1874
rect 37996 1810 38052 1822
rect 38332 2156 38500 2212
rect 38892 2212 38948 2222
rect 38332 1764 38388 2156
rect 38444 1986 38500 1998
rect 38444 1934 38446 1986
rect 38498 1934 38500 1986
rect 38444 1876 38500 1934
rect 38780 1988 38836 1998
rect 38668 1876 38724 1886
rect 38444 1874 38724 1876
rect 38444 1822 38670 1874
rect 38722 1822 38724 1874
rect 38444 1820 38724 1822
rect 38332 1698 38388 1708
rect 38668 1764 38724 1820
rect 38668 1698 38724 1708
rect 37884 1316 37940 1326
rect 37660 1250 37716 1260
rect 37772 1260 37884 1316
rect 37212 802 37268 812
rect 37772 644 37828 1260
rect 37884 1250 37940 1260
rect 38780 980 38836 1932
rect 38780 914 38836 924
rect 37660 588 37828 644
rect 38892 644 38948 2156
rect 37660 112 37716 588
rect 38892 578 38948 588
rect 39004 420 39060 3164
rect 39004 354 39060 364
rect 39676 112 39732 3332
rect 40348 2772 40404 3836
rect 40572 2882 40628 5852
rect 40684 5796 40740 5806
rect 40684 4900 40740 5740
rect 40684 4834 40740 4844
rect 40572 2830 40574 2882
rect 40626 2830 40628 2882
rect 40572 2818 40628 2830
rect 40684 4676 40740 4686
rect 40684 2884 40740 4620
rect 40684 2818 40740 2828
rect 40348 2706 40404 2716
rect 39788 2548 39844 2558
rect 40012 2548 40068 2558
rect 39788 2546 40068 2548
rect 39788 2494 39790 2546
rect 39842 2494 40014 2546
rect 40066 2494 40068 2546
rect 39788 2492 40068 2494
rect 39788 1540 39844 2492
rect 40012 2482 40068 2492
rect 40348 1876 40404 1886
rect 39788 1474 39844 1484
rect 40236 1764 40292 1774
rect 40236 756 40292 1708
rect 40348 980 40404 1820
rect 40796 1540 40852 7868
rect 41020 7924 41076 8206
rect 41020 7858 41076 7868
rect 41132 6466 41188 6478
rect 41132 6414 41134 6466
rect 41186 6414 41188 6466
rect 41132 5236 41188 6414
rect 41244 5348 41300 8316
rect 41580 8370 41636 9996
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 41692 8372 41748 11342
rect 41916 10052 41972 11452
rect 42028 11506 42084 11564
rect 42028 11454 42030 11506
rect 42082 11454 42084 11506
rect 42028 11442 42084 11454
rect 42140 10498 42196 11564
rect 42364 11554 42420 11564
rect 42140 10446 42142 10498
rect 42194 10446 42196 10498
rect 42140 10434 42196 10446
rect 42364 10610 42420 10622
rect 42364 10558 42366 10610
rect 42418 10558 42420 10610
rect 42252 10388 42308 10398
rect 42140 10052 42196 10062
rect 41916 9996 42140 10052
rect 42140 9958 42196 9996
rect 41804 9042 41860 9054
rect 41804 8990 41806 9042
rect 41858 8990 41860 9042
rect 41804 8484 41860 8990
rect 42252 9042 42308 10332
rect 42364 10276 42420 10558
rect 42364 10210 42420 10220
rect 42476 10164 42532 12908
rect 42588 11618 42644 13132
rect 43260 12516 43316 14112
rect 43708 13188 43764 14112
rect 43708 13122 43764 13132
rect 43260 12450 43316 12460
rect 43484 12964 43540 12974
rect 43260 12292 43316 12302
rect 42588 11566 42590 11618
rect 42642 11566 42644 11618
rect 42588 10500 42644 11566
rect 42700 12180 42756 12190
rect 42700 10722 42756 12124
rect 42700 10670 42702 10722
rect 42754 10670 42756 10722
rect 42700 10658 42756 10670
rect 43148 11060 43204 11070
rect 43036 10500 43092 10510
rect 42588 10498 43092 10500
rect 42588 10446 43038 10498
rect 43090 10446 43092 10498
rect 42588 10444 43092 10446
rect 43036 10434 43092 10444
rect 42476 10098 42532 10108
rect 42588 10052 42644 10062
rect 42588 9938 42644 9996
rect 42588 9886 42590 9938
rect 42642 9886 42644 9938
rect 42588 9874 42644 9886
rect 42476 9602 42532 9614
rect 42476 9550 42478 9602
rect 42530 9550 42532 9602
rect 42252 8990 42254 9042
rect 42306 8990 42308 9042
rect 42252 8978 42308 8990
rect 42364 9268 42420 9278
rect 42028 8820 42084 8830
rect 42028 8726 42084 8764
rect 41916 8484 41972 8494
rect 41804 8482 41972 8484
rect 41804 8430 41918 8482
rect 41970 8430 41972 8482
rect 41804 8428 41972 8430
rect 41916 8418 41972 8428
rect 42252 8484 42308 8494
rect 41692 8316 41860 8372
rect 41356 8258 41412 8270
rect 41356 8206 41358 8258
rect 41410 8206 41412 8258
rect 41356 6916 41412 8206
rect 41692 8034 41748 8046
rect 41692 7982 41694 8034
rect 41746 7982 41748 8034
rect 41692 7924 41748 7982
rect 41692 7858 41748 7868
rect 41356 6850 41412 6860
rect 41804 7364 41860 8316
rect 42140 8370 42196 8382
rect 42140 8318 42142 8370
rect 42194 8318 42196 8370
rect 42140 7924 42196 8318
rect 42252 8370 42308 8428
rect 42252 8318 42254 8370
rect 42306 8318 42308 8370
rect 42252 8306 42308 8318
rect 42140 7858 42196 7868
rect 41804 6802 41860 7308
rect 42028 7252 42084 7262
rect 42252 7252 42308 7262
rect 42028 7250 42196 7252
rect 42028 7198 42030 7250
rect 42082 7198 42196 7250
rect 42028 7196 42196 7198
rect 42028 7186 42084 7196
rect 41804 6750 41806 6802
rect 41858 6750 41860 6802
rect 41804 6738 41860 6750
rect 42028 6804 42084 6814
rect 42028 6710 42084 6748
rect 41468 6692 41524 6702
rect 41524 6636 41636 6692
rect 41468 6626 41524 6636
rect 41468 6466 41524 6478
rect 41468 6414 41470 6466
rect 41522 6414 41524 6466
rect 41468 6356 41524 6414
rect 41468 6018 41524 6300
rect 41468 5966 41470 6018
rect 41522 5966 41524 6018
rect 41468 5954 41524 5966
rect 41580 5460 41636 6636
rect 42140 6356 42196 7196
rect 42252 6802 42308 7196
rect 42252 6750 42254 6802
rect 42306 6750 42308 6802
rect 42252 6738 42308 6750
rect 42364 6804 42420 9212
rect 42476 8930 42532 9550
rect 43148 9268 43204 11004
rect 43148 9202 43204 9212
rect 43148 9044 43204 9054
rect 43148 8950 43204 8988
rect 42476 8878 42478 8930
rect 42530 8878 42532 8930
rect 42476 8866 42532 8878
rect 43260 8932 43316 12236
rect 43260 8866 43316 8876
rect 43372 10276 43428 10286
rect 43372 8260 43428 10220
rect 42364 6738 42420 6748
rect 42588 7362 42644 7374
rect 42588 7310 42590 7362
rect 42642 7310 42644 7362
rect 42252 6356 42308 6366
rect 42140 6300 42252 6356
rect 41804 6020 41860 6030
rect 41804 5926 41860 5964
rect 42252 5906 42308 6300
rect 42252 5854 42254 5906
rect 42306 5854 42308 5906
rect 42252 5842 42308 5854
rect 42140 5460 42196 5470
rect 41580 5404 42140 5460
rect 42140 5394 42196 5404
rect 41244 5282 41300 5292
rect 41132 5170 41188 5180
rect 42028 5124 42084 5134
rect 41916 5012 41972 5022
rect 41692 3892 41748 3902
rect 41580 2884 41636 2894
rect 41580 2790 41636 2828
rect 40908 2212 40964 2222
rect 40908 2118 40964 2156
rect 41132 2212 41188 2222
rect 41132 2118 41188 2156
rect 41692 2098 41748 3836
rect 41692 2046 41694 2098
rect 41746 2046 41748 2098
rect 41692 2034 41748 2046
rect 41916 1876 41972 4956
rect 42028 4340 42084 5068
rect 42588 4676 42644 7310
rect 42700 7252 42756 7262
rect 42700 6018 42756 7196
rect 43148 7252 43204 7262
rect 43148 7158 43204 7196
rect 42812 6916 42868 6926
rect 42812 6690 42868 6860
rect 43372 6802 43428 8204
rect 43372 6750 43374 6802
rect 43426 6750 43428 6802
rect 43372 6738 43428 6750
rect 42812 6638 42814 6690
rect 42866 6638 42868 6690
rect 42812 6626 42868 6638
rect 43148 6466 43204 6478
rect 43148 6414 43150 6466
rect 43202 6414 43204 6466
rect 43148 6356 43204 6414
rect 43148 6290 43204 6300
rect 42700 5966 42702 6018
rect 42754 5966 42756 6018
rect 42700 5954 42756 5966
rect 42588 4610 42644 4620
rect 42700 5012 42756 5022
rect 42028 4274 42084 4284
rect 42476 4004 42532 4014
rect 42476 3556 42532 3948
rect 42476 3490 42532 3500
rect 42700 3388 42756 4956
rect 42588 3332 42756 3388
rect 42140 2548 42196 2558
rect 42476 2548 42532 2558
rect 42140 2546 42532 2548
rect 42140 2494 42142 2546
rect 42194 2494 42478 2546
rect 42530 2494 42532 2546
rect 42140 2492 42532 2494
rect 42140 2482 42196 2492
rect 41916 1810 41972 1820
rect 40796 1474 40852 1484
rect 40348 914 40404 924
rect 41916 1428 41972 1438
rect 40236 690 40292 700
rect 41692 196 41748 206
rect 41692 112 41748 140
rect 41916 196 41972 1372
rect 42476 420 42532 2492
rect 42588 868 42644 3332
rect 43372 2884 43428 2894
rect 43484 2884 43540 12908
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 44156 12180 44212 14112
rect 44604 13524 44660 14112
rect 44604 13468 44884 13524
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 44156 12114 44212 12124
rect 44268 12068 44324 12078
rect 44492 12068 44548 12078
rect 44324 12066 44548 12068
rect 44324 12014 44494 12066
rect 44546 12014 44548 12066
rect 44324 12012 44548 12014
rect 44268 11974 44324 12012
rect 44492 12002 44548 12012
rect 44828 11844 44884 13468
rect 44940 12962 44996 12974
rect 44940 12910 44942 12962
rect 44994 12910 44996 12962
rect 44940 12852 44996 12910
rect 44940 12786 44996 12796
rect 45052 12292 45108 14112
rect 45052 12226 45108 12236
rect 45052 12068 45108 12078
rect 45052 11974 45108 12012
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44828 11778 44884 11788
rect 45388 11954 45444 11966
rect 45388 11902 45390 11954
rect 45442 11902 45444 11954
rect 45388 11732 45444 11902
rect 44464 11722 44728 11732
rect 45276 11676 45444 11732
rect 45052 11284 45108 11294
rect 45276 11284 45332 11676
rect 45052 11282 45332 11284
rect 45052 11230 45054 11282
rect 45106 11230 45332 11282
rect 45052 11228 45332 11230
rect 45388 11284 45444 11294
rect 45052 11218 45108 11228
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44828 10724 44884 10734
rect 43596 10388 43652 10398
rect 43596 6356 43652 10332
rect 44464 10220 44728 10230
rect 44156 10164 44212 10174
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44828 10164 44884 10668
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 43708 7252 43764 7262
rect 43708 6802 43764 7196
rect 43820 7140 43876 7150
rect 43820 6916 43876 7084
rect 43820 6850 43876 6860
rect 43708 6750 43710 6802
rect 43762 6750 43764 6802
rect 43708 6738 43764 6750
rect 43596 6290 43652 6300
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 43596 6132 43652 6142
rect 43596 4564 43652 6076
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 43596 4498 43652 4508
rect 44156 4452 44212 10108
rect 44828 10098 44884 10108
rect 44268 8932 44324 8942
rect 44268 8148 44324 8876
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44268 8082 44324 8092
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44268 5908 44324 5918
rect 44268 4900 44324 5852
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 44268 4834 44324 4844
rect 44940 4564 44996 4574
rect 44156 4450 44548 4452
rect 44156 4398 44158 4450
rect 44210 4398 44548 4450
rect 44156 4396 44548 4398
rect 44156 4386 44212 4396
rect 44492 4338 44548 4396
rect 44940 4450 44996 4508
rect 44940 4398 44942 4450
rect 44994 4398 44996 4450
rect 44940 4386 44996 4398
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44492 4274 44548 4286
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 45164 3388 45220 11228
rect 45388 10724 45444 11228
rect 45388 10658 45444 10668
rect 45500 9716 45556 14112
rect 45836 13636 45892 13646
rect 45500 9650 45556 9660
rect 45612 11508 45668 11518
rect 45276 8820 45332 8830
rect 45500 8820 45556 8830
rect 45276 8818 45556 8820
rect 45276 8766 45278 8818
rect 45330 8766 45502 8818
rect 45554 8766 45556 8818
rect 45276 8764 45556 8766
rect 45276 8484 45332 8764
rect 45500 8754 45556 8764
rect 45276 8418 45332 8428
rect 45612 8372 45668 11452
rect 45724 11284 45780 11294
rect 45724 9604 45780 11228
rect 45724 9538 45780 9548
rect 45612 8306 45668 8316
rect 45388 7812 45444 7822
rect 45388 6804 45444 7756
rect 45388 6738 45444 6748
rect 45612 6692 45668 6702
rect 45836 6692 45892 13580
rect 45948 13300 46004 14112
rect 45948 13234 46004 13244
rect 45948 12738 46004 12750
rect 45948 12686 45950 12738
rect 46002 12686 46004 12738
rect 45948 12516 46004 12686
rect 45948 12450 46004 12460
rect 46396 12180 46452 14112
rect 46844 13188 46900 14112
rect 46732 13132 46900 13188
rect 46396 12124 46564 12180
rect 45948 12066 46004 12078
rect 45948 12014 45950 12066
rect 46002 12014 46004 12066
rect 45948 8484 46004 12014
rect 46060 11956 46116 11966
rect 46060 11506 46116 11900
rect 46060 11454 46062 11506
rect 46114 11454 46116 11506
rect 46060 11442 46116 11454
rect 46396 11954 46452 11966
rect 46396 11902 46398 11954
rect 46450 11902 46452 11954
rect 46396 11284 46452 11902
rect 46396 11218 46452 11228
rect 46508 11394 46564 12124
rect 46508 11342 46510 11394
rect 46562 11342 46564 11394
rect 46508 10722 46564 11342
rect 46508 10670 46510 10722
rect 46562 10670 46564 10722
rect 46508 10658 46564 10670
rect 46620 10388 46676 10398
rect 46620 10294 46676 10332
rect 46620 10164 46676 10174
rect 46396 9826 46452 9838
rect 46396 9774 46398 9826
rect 46450 9774 46452 9826
rect 46060 9714 46116 9726
rect 46060 9662 46062 9714
rect 46114 9662 46116 9714
rect 46060 9604 46116 9662
rect 46060 9538 46116 9548
rect 46396 9604 46452 9774
rect 46396 9538 46452 9548
rect 46060 9044 46116 9054
rect 46060 8950 46116 8988
rect 45948 8418 46004 8428
rect 45612 6690 45892 6692
rect 45612 6638 45614 6690
rect 45666 6638 45838 6690
rect 45890 6638 45892 6690
rect 45612 6636 45892 6638
rect 45612 6626 45668 6636
rect 45836 6626 45892 6636
rect 46396 8260 46452 8270
rect 46284 6578 46340 6590
rect 46284 6526 46286 6578
rect 46338 6526 46340 6578
rect 45724 5348 45780 5358
rect 45052 3332 45220 3388
rect 45500 3892 45556 3902
rect 43804 3164 44068 3174
rect 43428 2828 43540 2884
rect 43596 3108 43652 3118
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 43596 2884 43652 3052
rect 43372 2818 43428 2828
rect 43596 2818 43652 2828
rect 43932 2660 43988 2670
rect 43708 2324 43764 2334
rect 43708 1988 43764 2268
rect 43708 1922 43764 1932
rect 43932 1988 43988 2604
rect 44156 2660 44212 2670
rect 44156 2436 44212 2604
rect 45052 2660 45108 3332
rect 45052 2594 45108 2604
rect 44156 2370 44212 2380
rect 44464 2380 44728 2390
rect 44268 2324 44324 2334
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 44828 2324 44884 2334
rect 44268 2212 44324 2268
rect 44828 2212 44884 2268
rect 44268 2156 44884 2212
rect 43932 1922 43988 1932
rect 43596 1652 43652 1662
rect 43596 1428 43652 1596
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 43596 1372 43764 1428
rect 42588 802 42644 812
rect 42476 354 42532 364
rect 41916 130 41972 140
rect 43708 112 43764 1372
rect 45500 980 45556 3836
rect 45724 2996 45780 5292
rect 45724 2930 45780 2940
rect 46284 2772 46340 6526
rect 46396 5012 46452 8204
rect 46620 5796 46676 10108
rect 46732 6020 46788 13132
rect 46844 12964 46900 12974
rect 46844 12870 46900 12908
rect 46844 12290 46900 12302
rect 46844 12238 46846 12290
rect 46898 12238 46900 12290
rect 46844 10836 46900 12238
rect 47180 12068 47236 12078
rect 46844 10770 46900 10780
rect 46956 11394 47012 11406
rect 46956 11342 46958 11394
rect 47010 11342 47012 11394
rect 46844 10388 46900 10398
rect 46956 10388 47012 11342
rect 46900 10332 47012 10388
rect 47068 10388 47124 10398
rect 46844 10322 46900 10332
rect 47068 10294 47124 10332
rect 46956 10164 47012 10174
rect 46956 9938 47012 10108
rect 46956 9886 46958 9938
rect 47010 9886 47012 9938
rect 46956 9874 47012 9886
rect 46956 8596 47012 8606
rect 46956 7700 47012 8540
rect 46956 7634 47012 7644
rect 46732 5954 46788 5964
rect 46620 5740 46788 5796
rect 46396 4946 46452 4956
rect 46620 5236 46676 5246
rect 46620 2884 46676 5180
rect 46732 4564 46788 5740
rect 46732 4498 46788 4508
rect 47180 3388 47236 12012
rect 47292 7924 47348 14112
rect 47740 12292 47796 14112
rect 47852 13412 47908 13422
rect 47852 12850 47908 13356
rect 48188 13188 48244 14112
rect 48188 13122 48244 13132
rect 48412 13076 48468 13086
rect 48412 12982 48468 13020
rect 47852 12798 47854 12850
rect 47906 12798 47908 12850
rect 47852 12786 47908 12798
rect 47964 12964 48020 12974
rect 48636 12964 48692 14112
rect 49084 13636 49140 14112
rect 49084 13570 49140 13580
rect 48972 13188 49028 13198
rect 48972 13094 49028 13132
rect 48636 12908 49140 12964
rect 47964 12402 48020 12908
rect 47964 12350 47966 12402
rect 48018 12350 48020 12402
rect 47964 12338 48020 12350
rect 49084 12402 49140 12908
rect 49084 12350 49086 12402
rect 49138 12350 49140 12402
rect 49084 12338 49140 12350
rect 47404 12236 47796 12292
rect 48076 12292 48132 12302
rect 47404 10498 47460 12236
rect 47740 11844 47796 11854
rect 47516 11284 47572 11294
rect 47516 11190 47572 11228
rect 47740 10612 47796 11788
rect 47404 10446 47406 10498
rect 47458 10446 47460 10498
rect 47404 10434 47460 10446
rect 47516 10610 47796 10612
rect 47516 10558 47742 10610
rect 47794 10558 47796 10610
rect 47516 10556 47796 10558
rect 47516 10050 47572 10556
rect 47740 10546 47796 10556
rect 47516 9998 47518 10050
rect 47570 9998 47572 10050
rect 47516 9986 47572 9998
rect 48076 9156 48132 12236
rect 49420 12180 49476 12190
rect 48524 12066 48580 12078
rect 48524 12014 48526 12066
rect 48578 12014 48580 12066
rect 48188 11394 48244 11406
rect 48188 11342 48190 11394
rect 48242 11342 48244 11394
rect 48188 10612 48244 11342
rect 48524 11396 48580 12014
rect 48972 11508 49028 11518
rect 48972 11414 49028 11452
rect 48524 11330 48580 11340
rect 48188 10546 48244 10556
rect 48748 11172 48804 11182
rect 48748 10610 48804 11116
rect 48748 10558 48750 10610
rect 48802 10558 48804 10610
rect 48748 10546 48804 10558
rect 48972 11060 49028 11070
rect 48300 10500 48356 10510
rect 48300 10406 48356 10444
rect 48860 10388 48916 10398
rect 48188 9940 48244 9950
rect 48188 9846 48244 9884
rect 48524 9940 48580 9950
rect 48524 9846 48580 9884
rect 48076 9154 48468 9156
rect 48076 9102 48078 9154
rect 48130 9102 48468 9154
rect 48076 9100 48468 9102
rect 48076 9090 48132 9100
rect 48412 9042 48468 9100
rect 48412 8990 48414 9042
rect 48466 8990 48468 9042
rect 48412 8978 48468 8990
rect 48524 9044 48580 9054
rect 47292 7858 47348 7868
rect 47964 8484 48020 8494
rect 47068 3332 47236 3388
rect 47404 4788 47460 4798
rect 47068 2996 47124 3332
rect 47068 2930 47124 2940
rect 46620 2818 46676 2828
rect 46284 2706 46340 2716
rect 46956 1986 47012 1998
rect 46956 1934 46958 1986
rect 47010 1934 47012 1986
rect 46732 1876 46788 1886
rect 46956 1876 47012 1934
rect 46732 1874 47012 1876
rect 46732 1822 46734 1874
rect 46786 1822 47012 1874
rect 46732 1820 47012 1822
rect 46732 1428 46788 1820
rect 46732 1362 46788 1372
rect 47068 1540 47124 1550
rect 45500 914 45556 924
rect 45724 980 45780 990
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 45724 112 45780 924
rect 10780 18 10836 28
rect 11424 0 11536 112
rect 13440 0 13552 112
rect 15456 0 15568 112
rect 17472 0 17584 112
rect 19488 0 19600 112
rect 21504 0 21616 112
rect 23520 0 23632 112
rect 25536 0 25648 112
rect 27552 0 27664 112
rect 29568 0 29680 112
rect 31584 0 31696 112
rect 33600 0 33712 112
rect 35616 0 35728 112
rect 37632 0 37744 112
rect 39648 0 39760 112
rect 41664 0 41776 112
rect 43680 0 43792 112
rect 45696 0 45808 112
rect 47068 84 47124 1484
rect 47404 1428 47460 4732
rect 47964 2772 48020 8428
rect 48300 7812 48356 7822
rect 48076 6804 48132 6814
rect 48076 3220 48132 6748
rect 48076 3154 48132 3164
rect 47964 2706 48020 2716
rect 47628 2548 47684 2558
rect 47852 2548 47908 2558
rect 47628 2546 47908 2548
rect 47628 2494 47630 2546
rect 47682 2494 47854 2546
rect 47906 2494 47908 2546
rect 47628 2492 47908 2494
rect 47516 2212 47572 2222
rect 47516 2098 47572 2156
rect 47516 2046 47518 2098
rect 47570 2046 47572 2098
rect 47516 2034 47572 2046
rect 47628 1540 47684 2492
rect 47852 2482 47908 2492
rect 48300 1988 48356 7756
rect 48412 2884 48468 2894
rect 48524 2884 48580 8988
rect 48748 7588 48804 7598
rect 48748 6580 48804 7532
rect 48748 6514 48804 6524
rect 48636 6020 48692 6030
rect 48636 5926 48692 5964
rect 48412 2882 48580 2884
rect 48412 2830 48414 2882
rect 48466 2830 48580 2882
rect 48412 2828 48580 2830
rect 48412 2818 48468 2828
rect 48860 2212 48916 10332
rect 48972 9154 49028 11004
rect 49084 10052 49140 10062
rect 49420 10052 49476 12124
rect 49532 11620 49588 14112
rect 49532 11554 49588 11564
rect 49868 13300 49924 13310
rect 49756 11394 49812 11406
rect 49756 11342 49758 11394
rect 49810 11342 49812 11394
rect 49644 11060 49700 11070
rect 49644 10834 49700 11004
rect 49644 10782 49646 10834
rect 49698 10782 49700 10834
rect 49644 10770 49700 10782
rect 49756 10164 49812 11342
rect 49756 10098 49812 10108
rect 49420 9996 49588 10052
rect 49084 9938 49140 9996
rect 49084 9886 49086 9938
rect 49138 9886 49140 9938
rect 49084 9874 49140 9886
rect 49420 9828 49476 9838
rect 49420 9734 49476 9772
rect 48972 9102 48974 9154
rect 49026 9102 49028 9154
rect 48972 9090 49028 9102
rect 49308 8818 49364 8830
rect 49308 8766 49310 8818
rect 49362 8766 49364 8818
rect 49084 8596 49140 8606
rect 49308 8596 49364 8766
rect 49140 8540 49364 8596
rect 49084 8482 49140 8540
rect 49084 8430 49086 8482
rect 49138 8430 49140 8482
rect 49084 8418 49140 8430
rect 49420 8148 49476 8158
rect 49420 7028 49476 8092
rect 49420 6962 49476 6972
rect 48972 6020 49028 6030
rect 49532 6020 49588 9996
rect 49868 9828 49924 13244
rect 49980 13076 50036 14112
rect 49980 13010 50036 13020
rect 50092 12852 50148 12862
rect 50092 12850 50260 12852
rect 50092 12798 50094 12850
rect 50146 12798 50260 12850
rect 50092 12796 50260 12798
rect 50092 12786 50148 12796
rect 49980 12178 50036 12190
rect 49980 12126 49982 12178
rect 50034 12126 50036 12178
rect 49980 9940 50036 12126
rect 50204 11956 50260 12796
rect 50428 12404 50484 14112
rect 50428 12338 50484 12348
rect 50764 12962 50820 12974
rect 50764 12910 50766 12962
rect 50818 12910 50820 12962
rect 50204 11890 50260 11900
rect 50428 11956 50484 11966
rect 50428 11862 50484 11900
rect 50316 11620 50372 11630
rect 50316 11526 50372 11564
rect 50540 10724 50596 10734
rect 49980 9874 50036 9884
rect 50204 10276 50260 10286
rect 50204 9938 50260 10220
rect 50204 9886 50206 9938
rect 50258 9886 50260 9938
rect 50204 9874 50260 9886
rect 49868 9762 49924 9772
rect 50428 9268 50484 9278
rect 49868 8932 49924 8942
rect 50204 8932 50260 8942
rect 49868 8930 50036 8932
rect 49868 8878 49870 8930
rect 49922 8878 50036 8930
rect 49868 8876 50036 8878
rect 49868 8866 49924 8876
rect 49756 8258 49812 8270
rect 49756 8206 49758 8258
rect 49810 8206 49812 8258
rect 49756 8148 49812 8206
rect 49756 8082 49812 8092
rect 49644 7924 49700 7934
rect 49644 7586 49700 7868
rect 49980 7812 50036 8876
rect 50204 8838 50260 8876
rect 50316 8372 50372 8382
rect 50316 8278 50372 8316
rect 49980 7756 50372 7812
rect 49644 7534 49646 7586
rect 49698 7534 49700 7586
rect 49644 7476 49700 7534
rect 49980 7476 50036 7486
rect 49644 7474 50036 7476
rect 49644 7422 49982 7474
rect 50034 7422 50036 7474
rect 49644 7420 50036 7422
rect 49980 7410 50036 7420
rect 50204 6692 50260 6702
rect 50204 6598 50260 6636
rect 50316 6020 50372 7756
rect 49532 5964 49700 6020
rect 48972 5906 49028 5964
rect 48972 5854 48974 5906
rect 49026 5854 49028 5906
rect 48972 5842 49028 5854
rect 49532 5796 49588 5806
rect 49532 5702 49588 5740
rect 49532 4452 49588 4462
rect 49644 4452 49700 5964
rect 50204 5964 50372 6020
rect 49532 4450 49924 4452
rect 49532 4398 49534 4450
rect 49586 4398 49924 4450
rect 49532 4396 49924 4398
rect 49532 4386 49588 4396
rect 49868 4338 49924 4396
rect 49868 4286 49870 4338
rect 49922 4286 49924 4338
rect 49868 4274 49924 4286
rect 50204 3332 50260 5964
rect 50316 4450 50372 4462
rect 50316 4398 50318 4450
rect 50370 4398 50372 4450
rect 50316 3892 50372 4398
rect 50428 4452 50484 9212
rect 50540 8148 50596 10668
rect 50764 9492 50820 12910
rect 50876 11620 50932 14112
rect 51100 13636 51156 13646
rect 51100 13186 51156 13580
rect 51100 13134 51102 13186
rect 51154 13134 51156 13186
rect 51100 13122 51156 13134
rect 50988 12068 51044 12078
rect 50988 12066 51156 12068
rect 50988 12014 50990 12066
rect 51042 12014 51156 12066
rect 50988 12012 51156 12014
rect 50988 12002 51044 12012
rect 50876 11554 50932 11564
rect 50876 11172 50932 11182
rect 50876 10834 50932 11116
rect 50876 10782 50878 10834
rect 50930 10782 50932 10834
rect 50876 10770 50932 10782
rect 50764 9426 50820 9436
rect 50988 9826 51044 9838
rect 50988 9774 50990 9826
rect 51042 9774 51044 9826
rect 50988 8820 51044 9774
rect 50988 8754 51044 8764
rect 50988 8260 51044 8270
rect 50988 8166 51044 8204
rect 50540 8146 50708 8148
rect 50540 8094 50542 8146
rect 50594 8094 50708 8146
rect 50540 8092 50708 8094
rect 50540 8082 50596 8092
rect 50540 7476 50596 7486
rect 50652 7476 50708 8092
rect 50876 7476 50932 7486
rect 50652 7474 50932 7476
rect 50652 7422 50878 7474
rect 50930 7422 50932 7474
rect 50652 7420 50932 7422
rect 50540 7382 50596 7420
rect 50876 7410 50932 7420
rect 50652 7028 50708 7038
rect 50540 6692 50596 6702
rect 50540 6598 50596 6636
rect 50540 6356 50596 6366
rect 50540 4900 50596 6300
rect 50540 4834 50596 4844
rect 50428 4396 50596 4452
rect 50316 3826 50372 3836
rect 50204 3266 50260 3276
rect 50428 3332 50484 3342
rect 49084 2212 49140 2222
rect 48860 2210 49140 2212
rect 48860 2158 49086 2210
rect 49138 2158 49140 2210
rect 48860 2156 49140 2158
rect 49084 2146 49140 2156
rect 50428 2098 50484 3276
rect 50540 2884 50596 4396
rect 50652 4116 50708 6972
rect 51100 6916 51156 12012
rect 51324 11732 51380 14112
rect 51772 12740 51828 14112
rect 52220 13188 52276 14112
rect 52220 13122 52276 13132
rect 51772 12674 51828 12684
rect 52332 12962 52388 12974
rect 52332 12910 52334 12962
rect 52386 12910 52388 12962
rect 51324 11666 51380 11676
rect 51996 12628 52052 12638
rect 51884 11620 51940 11630
rect 51884 11526 51940 11564
rect 51324 11394 51380 11406
rect 51324 11342 51326 11394
rect 51378 11342 51380 11394
rect 51324 10948 51380 11342
rect 51324 10882 51380 10892
rect 51436 10500 51492 10510
rect 51436 10498 51716 10500
rect 51436 10446 51438 10498
rect 51490 10446 51716 10498
rect 51436 10444 51716 10446
rect 51436 10434 51492 10444
rect 51548 9828 51604 9838
rect 51212 9380 51268 9390
rect 51212 9266 51268 9324
rect 51212 9214 51214 9266
rect 51266 9214 51268 9266
rect 51212 9202 51268 9214
rect 51436 7364 51492 7374
rect 51436 7270 51492 7308
rect 51100 6850 51156 6860
rect 51100 6692 51156 6702
rect 51100 6598 51156 6636
rect 51436 6690 51492 6702
rect 51436 6638 51438 6690
rect 51490 6638 51492 6690
rect 50652 4050 50708 4060
rect 51100 5684 51156 5694
rect 51436 5684 51492 6638
rect 51100 5682 51492 5684
rect 51100 5630 51102 5682
rect 51154 5630 51492 5682
rect 51100 5628 51492 5630
rect 50540 2882 50932 2884
rect 50540 2830 50542 2882
rect 50594 2830 50932 2882
rect 50540 2828 50932 2830
rect 50540 2818 50596 2828
rect 50876 2770 50932 2828
rect 50876 2718 50878 2770
rect 50930 2718 50932 2770
rect 50876 2706 50932 2718
rect 50428 2046 50430 2098
rect 50482 2046 50484 2098
rect 50428 2034 50484 2046
rect 48300 1922 48356 1932
rect 49308 1986 49364 1998
rect 49308 1934 49310 1986
rect 49362 1934 49364 1986
rect 48748 1876 48804 1886
rect 48748 1782 48804 1820
rect 49308 1876 49364 1934
rect 49308 1810 49364 1820
rect 49868 1986 49924 1998
rect 49868 1934 49870 1986
rect 49922 1934 49924 1986
rect 47628 1474 47684 1484
rect 47404 1362 47460 1372
rect 49532 980 49588 990
rect 49868 980 49924 1934
rect 50764 1986 50820 1998
rect 50764 1934 50766 1986
rect 50818 1934 50820 1986
rect 50652 1652 50708 1662
rect 50428 1316 50484 1326
rect 50428 1222 50484 1260
rect 50652 1314 50708 1596
rect 50652 1262 50654 1314
rect 50706 1262 50708 1314
rect 50652 1250 50708 1262
rect 50764 1316 50820 1934
rect 50764 1250 50820 1260
rect 50988 1204 51044 1214
rect 50988 1110 51044 1148
rect 49532 978 49924 980
rect 49532 926 49534 978
rect 49586 926 49924 978
rect 49532 924 49924 926
rect 51100 980 51156 5628
rect 51436 3780 51492 3790
rect 51548 3780 51604 9772
rect 51660 6580 51716 10444
rect 51996 9828 52052 12572
rect 52220 12178 52276 12190
rect 52220 12126 52222 12178
rect 52274 12126 52276 12178
rect 52108 10836 52164 10846
rect 52108 10610 52164 10780
rect 52108 10558 52110 10610
rect 52162 10558 52164 10610
rect 52108 10546 52164 10558
rect 51772 9772 52052 9828
rect 51772 8370 51828 9772
rect 51996 9604 52052 9614
rect 51996 9510 52052 9548
rect 51772 8318 51774 8370
rect 51826 8318 51828 8370
rect 51772 8306 51828 8318
rect 51884 9492 51940 9502
rect 51884 6804 51940 9436
rect 52108 9156 52164 9166
rect 52108 9042 52164 9100
rect 52108 8990 52110 9042
rect 52162 8990 52164 9042
rect 52108 8978 52164 8990
rect 52220 8372 52276 12126
rect 52332 10052 52388 12910
rect 52668 12964 52724 14112
rect 53116 13300 53172 14112
rect 53116 13234 53172 13244
rect 52892 13076 52948 13086
rect 52892 12982 52948 13020
rect 52668 12908 52836 12964
rect 52556 12404 52612 12414
rect 52556 12310 52612 12348
rect 52556 11732 52612 11742
rect 52556 10834 52612 11676
rect 52780 11620 52836 12908
rect 53564 12292 53620 14112
rect 53788 13076 53844 13086
rect 53564 12236 53732 12292
rect 53564 12066 53620 12078
rect 53564 12014 53566 12066
rect 53618 12014 53620 12066
rect 53452 11620 53508 11630
rect 52780 11618 53508 11620
rect 52780 11566 53454 11618
rect 53506 11566 53508 11618
rect 52780 11564 53508 11566
rect 53452 11554 53508 11564
rect 52892 11396 52948 11406
rect 52556 10782 52558 10834
rect 52610 10782 52612 10834
rect 52556 10770 52612 10782
rect 52780 11394 52948 11396
rect 52780 11342 52894 11394
rect 52946 11342 52948 11394
rect 52780 11340 52948 11342
rect 52332 9986 52388 9996
rect 52556 9826 52612 9838
rect 52556 9774 52558 9826
rect 52610 9774 52612 9826
rect 52556 9044 52612 9774
rect 52556 8978 52612 8988
rect 52220 8306 52276 8316
rect 52556 8258 52612 8270
rect 52556 8206 52558 8258
rect 52610 8206 52612 8258
rect 51996 7362 52052 7374
rect 51996 7310 51998 7362
rect 52050 7310 52052 7362
rect 51996 7028 52052 7310
rect 51996 6962 52052 6972
rect 52444 6916 52500 6926
rect 51884 6748 52052 6804
rect 51884 6580 51940 6590
rect 51660 6578 51940 6580
rect 51660 6526 51886 6578
rect 51938 6526 51940 6578
rect 51660 6524 51940 6526
rect 51884 6514 51940 6524
rect 51996 6356 52052 6748
rect 52444 6468 52500 6860
rect 52556 6804 52612 8206
rect 52556 6738 52612 6748
rect 52668 6690 52724 6702
rect 52668 6638 52670 6690
rect 52722 6638 52724 6690
rect 52444 6412 52612 6468
rect 51884 6300 52052 6356
rect 51660 5124 51716 5134
rect 51660 5030 51716 5068
rect 51660 3780 51716 3790
rect 51436 3778 51716 3780
rect 51436 3726 51438 3778
rect 51490 3726 51662 3778
rect 51714 3726 51716 3778
rect 51436 3724 51716 3726
rect 51436 3714 51492 3724
rect 51660 3714 51716 3724
rect 51884 3332 51940 6300
rect 52108 5906 52164 5918
rect 52108 5854 52110 5906
rect 52162 5854 52164 5906
rect 52108 5348 52164 5854
rect 52108 5282 52164 5292
rect 51996 5124 52052 5134
rect 51996 5030 52052 5068
rect 52444 5010 52500 5022
rect 52444 4958 52446 5010
rect 52498 4958 52500 5010
rect 52332 4564 52388 4574
rect 52220 4452 52276 4462
rect 52220 3666 52276 4396
rect 52332 4450 52388 4508
rect 52332 4398 52334 4450
rect 52386 4398 52388 4450
rect 52332 4386 52388 4398
rect 52220 3614 52222 3666
rect 52274 3614 52276 3666
rect 52220 3602 52276 3614
rect 51884 3266 51940 3276
rect 51324 3220 51380 3230
rect 51324 2098 51380 3164
rect 52108 2772 52164 2782
rect 52108 2678 52164 2716
rect 51324 2046 51326 2098
rect 51378 2046 51380 2098
rect 51324 2034 51380 2046
rect 51436 2658 51492 2670
rect 51436 2606 51438 2658
rect 51490 2606 51492 2658
rect 51436 2100 51492 2606
rect 51436 2034 51492 2044
rect 52220 2100 52276 2110
rect 52220 2006 52276 2044
rect 51660 1986 51716 1998
rect 51660 1934 51662 1986
rect 51714 1934 51716 1986
rect 51660 1652 51716 1934
rect 51660 1586 51716 1596
rect 49532 644 49588 924
rect 51100 914 51156 924
rect 51772 1428 51828 1438
rect 49532 578 49588 588
rect 49756 756 49812 766
rect 47740 420 47796 430
rect 47740 112 47796 364
rect 49756 112 49812 700
rect 51772 112 51828 1372
rect 51996 1314 52052 1326
rect 51996 1262 51998 1314
rect 52050 1262 52052 1314
rect 51996 980 52052 1262
rect 52444 1204 52500 4958
rect 52556 3666 52612 6412
rect 52668 5908 52724 6638
rect 52668 5842 52724 5852
rect 52668 4564 52724 4574
rect 52668 4338 52724 4508
rect 52668 4286 52670 4338
rect 52722 4286 52724 4338
rect 52668 4274 52724 4286
rect 52556 3614 52558 3666
rect 52610 3614 52612 3666
rect 52556 3602 52612 3614
rect 52780 3220 52836 11340
rect 52892 11330 52948 11340
rect 53564 10836 53620 12014
rect 52892 10780 53620 10836
rect 52892 6692 52948 10780
rect 53676 10724 53732 12236
rect 53788 11060 53844 13020
rect 53788 10994 53844 11004
rect 53452 10668 53732 10724
rect 53788 10836 53844 10846
rect 53228 10500 53284 10510
rect 53116 9716 53172 9726
rect 53004 9268 53060 9278
rect 53004 9174 53060 9212
rect 53004 7924 53060 7934
rect 53004 7698 53060 7868
rect 53004 7646 53006 7698
rect 53058 7646 53060 7698
rect 53004 7634 53060 7646
rect 52892 6626 52948 6636
rect 53004 6132 53060 6142
rect 53004 6038 53060 6076
rect 53004 5348 53060 5358
rect 53116 5348 53172 9660
rect 53228 6578 53284 10444
rect 53452 9714 53508 10668
rect 53452 9662 53454 9714
rect 53506 9662 53508 9714
rect 53452 9650 53508 9662
rect 53564 10498 53620 10510
rect 53564 10446 53566 10498
rect 53618 10446 53620 10498
rect 53564 8428 53620 10446
rect 53788 9604 53844 10780
rect 53788 9538 53844 9548
rect 54012 9268 54068 14112
rect 54124 12740 54180 12750
rect 54124 12402 54180 12684
rect 54124 12350 54126 12402
rect 54178 12350 54180 12402
rect 54124 12338 54180 12350
rect 54460 12292 54516 14112
rect 54684 13524 54740 13534
rect 54348 12236 54516 12292
rect 54572 12962 54628 12974
rect 54572 12910 54574 12962
rect 54626 12910 54628 12962
rect 54236 11508 54292 11518
rect 54012 9202 54068 9212
rect 54124 9826 54180 9838
rect 54124 9774 54126 9826
rect 54178 9774 54180 9826
rect 53340 8372 53396 8382
rect 53340 8278 53396 8316
rect 53452 8372 53620 8428
rect 53676 9042 53732 9054
rect 53676 8990 53678 9042
rect 53730 8990 53732 9042
rect 53228 6526 53230 6578
rect 53282 6526 53284 6578
rect 53228 6514 53284 6526
rect 53228 5348 53284 5358
rect 53004 5346 53284 5348
rect 53004 5294 53006 5346
rect 53058 5294 53230 5346
rect 53282 5294 53284 5346
rect 53004 5292 53284 5294
rect 53004 5282 53060 5292
rect 53228 5282 53284 5292
rect 53228 4228 53284 4238
rect 53228 4134 53284 4172
rect 52780 3154 52836 3164
rect 52556 2884 52612 2894
rect 52556 2098 52612 2828
rect 52780 2660 52836 2670
rect 52780 2566 52836 2604
rect 53452 2324 53508 8372
rect 53564 7362 53620 7374
rect 53564 7310 53566 7362
rect 53618 7310 53620 7362
rect 53564 7252 53620 7310
rect 53564 7186 53620 7196
rect 53564 6580 53620 6590
rect 53564 5906 53620 6524
rect 53564 5854 53566 5906
rect 53618 5854 53620 5906
rect 53564 5842 53620 5854
rect 53676 5460 53732 8990
rect 54124 8708 54180 9774
rect 54236 9380 54292 11452
rect 54348 11172 54404 12236
rect 54460 11396 54516 11406
rect 54460 11302 54516 11340
rect 54348 11106 54404 11116
rect 54572 10948 54628 12910
rect 54236 9314 54292 9324
rect 54460 10892 54628 10948
rect 54124 8642 54180 8652
rect 54348 8930 54404 8942
rect 54348 8878 54350 8930
rect 54402 8878 54404 8930
rect 54348 8596 54404 8878
rect 54348 8530 54404 8540
rect 54460 8428 54516 10892
rect 54572 10722 54628 10734
rect 54572 10670 54574 10722
rect 54626 10670 54628 10722
rect 54572 10164 54628 10670
rect 54684 10276 54740 13468
rect 54908 13412 54964 14112
rect 54908 13346 54964 13356
rect 54908 13188 54964 13198
rect 54908 13094 54964 13132
rect 55356 12964 55412 14112
rect 55356 12898 55412 12908
rect 55692 13300 55748 13310
rect 55692 12402 55748 13244
rect 55692 12350 55694 12402
rect 55746 12350 55748 12402
rect 55692 12338 55748 12350
rect 55356 12178 55412 12190
rect 55356 12126 55358 12178
rect 55410 12126 55412 12178
rect 54908 11396 54964 11406
rect 55244 11396 55300 11406
rect 54684 10210 54740 10220
rect 54796 11394 55300 11396
rect 54796 11342 54910 11394
rect 54962 11342 55246 11394
rect 55298 11342 55300 11394
rect 54796 11340 55300 11342
rect 54572 10098 54628 10108
rect 53900 8372 54516 8428
rect 53900 6244 53956 8372
rect 54124 8258 54180 8270
rect 54124 8206 54126 8258
rect 54178 8206 54180 8258
rect 54124 7812 54180 8206
rect 54124 7746 54180 7756
rect 54572 7586 54628 7598
rect 54572 7534 54574 7586
rect 54626 7534 54628 7586
rect 54572 7252 54628 7534
rect 54572 7186 54628 7196
rect 53900 6178 53956 6188
rect 54236 6690 54292 6702
rect 54236 6638 54238 6690
rect 54290 6638 54292 6690
rect 53564 5404 53732 5460
rect 54124 5684 54180 5694
rect 53564 5012 53620 5404
rect 54124 5234 54180 5628
rect 54124 5182 54126 5234
rect 54178 5182 54180 5234
rect 54124 5170 54180 5182
rect 54236 5236 54292 6638
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 5908 54628 5966
rect 54572 5842 54628 5852
rect 54236 5170 54292 5180
rect 53564 4946 53620 4956
rect 53676 5010 53732 5022
rect 53676 4958 53678 5010
rect 53730 4958 53732 5010
rect 53564 4226 53620 4238
rect 53564 4174 53566 4226
rect 53618 4174 53620 4226
rect 53564 3780 53620 4174
rect 53564 3714 53620 3724
rect 53676 3668 53732 4958
rect 54572 4564 54628 4574
rect 54572 4470 54628 4508
rect 53676 3602 53732 3612
rect 54124 3556 54180 3566
rect 54124 3462 54180 3500
rect 53564 3444 53620 3454
rect 53564 3350 53620 3388
rect 54572 3220 54628 3230
rect 53564 3108 53620 3118
rect 53564 2770 53620 3052
rect 54572 2994 54628 3164
rect 54572 2942 54574 2994
rect 54626 2942 54628 2994
rect 54572 2930 54628 2942
rect 53564 2718 53566 2770
rect 53618 2718 53620 2770
rect 53564 2706 53620 2718
rect 53452 2258 53508 2268
rect 54124 2548 54180 2558
rect 52556 2046 52558 2098
rect 52610 2046 52612 2098
rect 52556 2034 52612 2046
rect 54124 2098 54180 2492
rect 54124 2046 54126 2098
rect 54178 2046 54180 2098
rect 54124 2034 54180 2046
rect 53564 1876 53620 1886
rect 53564 1782 53620 1820
rect 53564 1428 53620 1438
rect 53564 1334 53620 1372
rect 52556 1204 52612 1214
rect 52444 1202 52612 1204
rect 52444 1150 52558 1202
rect 52610 1150 52612 1202
rect 52444 1148 52612 1150
rect 52556 1138 52612 1148
rect 51996 914 52052 924
rect 53788 868 53844 878
rect 53788 112 53844 812
rect 54796 756 54852 11340
rect 54908 11330 54964 11340
rect 55244 11330 55300 11340
rect 55356 11284 55412 12126
rect 55356 11218 55412 11228
rect 55580 11284 55636 11294
rect 55132 10500 55188 10510
rect 54908 10498 55188 10500
rect 54908 10446 55134 10498
rect 55186 10446 55188 10498
rect 54908 10444 55188 10446
rect 54908 7140 54964 10444
rect 55132 10434 55188 10444
rect 55468 10388 55524 10398
rect 55132 9602 55188 9614
rect 55132 9550 55134 9602
rect 55186 9550 55188 9602
rect 55132 9492 55188 9550
rect 55132 9426 55188 9436
rect 55132 8932 55188 8942
rect 55020 8930 55188 8932
rect 55020 8878 55134 8930
rect 55186 8878 55188 8930
rect 55020 8876 55188 8878
rect 55020 8484 55076 8876
rect 55132 8866 55188 8876
rect 55020 8418 55076 8428
rect 55468 8372 55524 10332
rect 55132 8316 55524 8372
rect 55580 8372 55636 11228
rect 55804 10500 55860 14112
rect 56252 12516 56308 14112
rect 56252 12450 56308 12460
rect 55804 10434 55860 10444
rect 56140 10722 56196 10734
rect 56140 10670 56142 10722
rect 56194 10670 56196 10722
rect 56140 9044 56196 10670
rect 56140 8978 56196 8988
rect 55132 8146 55188 8316
rect 55580 8306 55636 8316
rect 55916 8930 55972 8942
rect 55916 8878 55918 8930
rect 55970 8878 55972 8930
rect 55132 8094 55134 8146
rect 55186 8094 55188 8146
rect 55132 8082 55188 8094
rect 55916 8148 55972 8878
rect 55916 8082 55972 8092
rect 55132 7700 55188 7710
rect 55132 7474 55188 7644
rect 56140 7700 56196 7710
rect 56140 7606 56196 7644
rect 55132 7422 55134 7474
rect 55186 7422 55188 7474
rect 55132 7410 55188 7422
rect 54908 7074 54964 7084
rect 56140 6804 56196 6814
rect 55132 6466 55188 6478
rect 55132 6414 55134 6466
rect 55186 6414 55188 6466
rect 55132 6356 55188 6414
rect 55132 6290 55188 6300
rect 56140 6130 56196 6748
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 56700 6132 56756 14112
rect 57036 13972 57092 13982
rect 57036 11508 57092 13916
rect 57036 11442 57092 11452
rect 57260 12180 57316 12190
rect 57260 7924 57316 12124
rect 57260 7858 57316 7868
rect 56700 6066 56756 6076
rect 55132 5794 55188 5806
rect 55132 5742 55134 5794
rect 55186 5742 55188 5794
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 55132 4900 55188 5742
rect 55132 4834 55188 4844
rect 56140 5460 56196 5470
rect 56140 4562 56196 5404
rect 56140 4510 56142 4562
rect 56194 4510 56196 4562
rect 56140 4498 56196 4510
rect 55132 4340 55188 4350
rect 55132 4246 55188 4284
rect 56140 4116 56196 4126
rect 54908 3668 54964 3678
rect 54908 3574 54964 3612
rect 55132 2996 55188 3006
rect 55132 2770 55188 2940
rect 56140 2994 56196 4060
rect 56140 2942 56142 2994
rect 56194 2942 56196 2994
rect 56140 2930 56196 2942
rect 56700 3444 56756 3454
rect 55132 2718 55134 2770
rect 55186 2718 55188 2770
rect 55132 2706 55188 2718
rect 56140 2772 56196 2782
rect 54908 2324 54964 2334
rect 54908 2098 54964 2268
rect 54908 2046 54910 2098
rect 54962 2046 54964 2098
rect 54908 2034 54964 2046
rect 56140 1426 56196 2716
rect 56140 1374 56142 1426
rect 56194 1374 56196 1426
rect 56140 1362 56196 1374
rect 56476 2660 56532 2670
rect 55132 1092 55188 1102
rect 55132 998 55188 1036
rect 54796 690 54852 700
rect 56476 532 56532 2604
rect 56476 466 56532 476
rect 55804 196 55860 206
rect 55804 112 55860 140
rect 47068 18 47124 28
rect 47712 0 47824 112
rect 49728 0 49840 112
rect 51744 0 51856 112
rect 53760 0 53872 112
rect 55776 0 55888 112
rect 56700 84 56756 3388
rect 56700 18 56756 28
<< via2 >>
rect 17052 14140 17108 14196
rect 476 13916 532 13972
rect 140 13468 196 13524
rect 364 12572 420 12628
rect 140 9212 196 9268
rect 252 11228 308 11284
rect 252 6412 308 6468
rect 588 12124 644 12180
rect 588 11340 644 11396
rect 1148 11788 1204 11844
rect 1484 13020 1540 13076
rect 1932 12012 1988 12068
rect 1484 11564 1540 11620
rect 476 11116 532 11172
rect 1036 9884 1092 9940
rect 1372 10332 1428 10388
rect 1036 7420 1092 7476
rect 1148 6524 1204 6580
rect 1036 6300 1092 6356
rect 2268 13580 2324 13636
rect 2156 13244 2212 13300
rect 2268 11788 2324 11844
rect 2828 12348 2884 12404
rect 3388 13580 3444 13636
rect 3612 13468 3668 13524
rect 2940 11564 2996 11620
rect 2716 9660 2772 9716
rect 1932 9436 1988 9492
rect 1484 7532 1540 7588
rect 1596 9212 1652 9268
rect 1596 7196 1652 7252
rect 1708 8764 1764 8820
rect 1372 5964 1428 6020
rect 1148 5852 1204 5908
rect 364 4844 420 4900
rect 924 4956 980 5012
rect 2604 8428 2660 8484
rect 1932 6860 1988 6916
rect 3724 13186 3780 13188
rect 3724 13134 3726 13186
rect 3726 13134 3778 13186
rect 3778 13134 3780 13186
rect 3724 13132 3780 13134
rect 4732 13468 4788 13524
rect 4284 13244 4340 13300
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 3276 10444 3332 10500
rect 2940 7196 2996 7252
rect 2828 5740 2884 5796
rect 2268 5180 2324 5236
rect 1148 2828 1204 2884
rect 924 588 980 644
rect 1372 1372 1428 1428
rect 1596 4396 1652 4452
rect 1596 2716 1652 2772
rect 1484 924 1540 980
rect 3276 8988 3332 9044
rect 3276 8540 3332 8596
rect 3276 4844 3332 4900
rect 3276 4060 3332 4116
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 5068 12124 5124 12180
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4620 11618 4676 11620
rect 4620 11566 4622 11618
rect 4622 11566 4674 11618
rect 4674 11566 4676 11618
rect 4620 11564 4676 11566
rect 5628 13132 5684 13188
rect 5964 13186 6020 13188
rect 5964 13134 5966 13186
rect 5966 13134 6018 13186
rect 6018 13134 6020 13186
rect 5964 13132 6020 13134
rect 6076 13020 6132 13076
rect 5852 12908 5908 12964
rect 5740 11788 5796 11844
rect 5180 11564 5236 11620
rect 4956 10780 5012 10836
rect 4396 10332 4452 10388
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4956 9996 5012 10052
rect 4172 8876 4228 8932
rect 4508 8818 4564 8820
rect 4508 8766 4510 8818
rect 4510 8766 4562 8818
rect 4562 8766 4564 8818
rect 4508 8764 4564 8766
rect 4956 8818 5012 8820
rect 4956 8766 4958 8818
rect 4958 8766 5010 8818
rect 5010 8766 5012 8818
rect 4956 8764 5012 8766
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 5292 10780 5348 10836
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4956 5180 5012 5236
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 3612 3612 3668 3668
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 3276 2268 3332 2324
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 5180 4284 5236 4340
rect 4956 2156 5012 2212
rect 5068 4172 5124 4228
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 3052 924 3108 980
rect 3388 1260 3444 1316
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 5068 812 5124 868
rect 4672 756 4728 758
rect 5292 2604 5348 2660
rect 6188 11618 6244 11620
rect 6188 11566 6190 11618
rect 6190 11566 6242 11618
rect 6242 11566 6244 11618
rect 6188 11564 6244 11566
rect 6524 12908 6580 12964
rect 7420 13132 7476 13188
rect 7532 13244 7588 13300
rect 6972 12402 7028 12404
rect 6972 12350 6974 12402
rect 6974 12350 7026 12402
rect 7026 12350 7028 12402
rect 6972 12348 7028 12350
rect 6860 11564 6916 11620
rect 6300 8204 6356 8260
rect 5852 4732 5908 4788
rect 6076 7084 6132 7140
rect 6524 6076 6580 6132
rect 6412 6018 6468 6020
rect 6412 5966 6414 6018
rect 6414 5966 6466 6018
rect 6466 5966 6468 6018
rect 6412 5964 6468 5966
rect 5516 1484 5572 1540
rect 5628 2828 5684 2884
rect 5180 476 5236 532
rect 5964 1260 6020 1316
rect 7420 10220 7476 10276
rect 7308 9548 7364 9604
rect 6860 7420 6916 7476
rect 7420 8146 7476 8148
rect 7420 8094 7422 8146
rect 7422 8094 7474 8146
rect 7474 8094 7476 8146
rect 7420 8092 7476 8094
rect 7308 7308 7364 7364
rect 6860 6748 6916 6804
rect 6748 5964 6804 6020
rect 7420 5964 7476 6020
rect 6972 5852 7028 5908
rect 6860 5180 6916 5236
rect 6748 3836 6804 3892
rect 6748 3276 6804 3332
rect 6636 2044 6692 2100
rect 7308 2716 7364 2772
rect 7756 11618 7812 11620
rect 7756 11566 7758 11618
rect 7758 11566 7810 11618
rect 7810 11566 7812 11618
rect 7756 11564 7812 11566
rect 8204 13020 8260 13076
rect 9660 13244 9716 13300
rect 9772 13916 9828 13972
rect 10108 13020 10164 13076
rect 8316 12348 8372 12404
rect 8428 11900 8484 11956
rect 7644 8876 7700 8932
rect 7756 8092 7812 8148
rect 7756 7308 7812 7364
rect 7980 7532 8036 7588
rect 7980 6524 8036 6580
rect 7868 6188 7924 6244
rect 7532 2380 7588 2436
rect 8316 9996 8372 10052
rect 8316 7868 8372 7924
rect 8428 7980 8484 8036
rect 8316 6188 8372 6244
rect 8316 5964 8372 6020
rect 8204 2828 8260 2884
rect 8428 3500 8484 3556
rect 8092 1932 8148 1988
rect 6972 1708 7028 1764
rect 6860 1372 6916 1428
rect 5628 700 5684 756
rect 9324 12684 9380 12740
rect 8764 11564 8820 11620
rect 9324 11228 9380 11284
rect 9436 12012 9492 12068
rect 9436 10892 9492 10948
rect 8988 10668 9044 10724
rect 8876 10444 8932 10500
rect 9324 7980 9380 8036
rect 9548 9884 9604 9940
rect 8876 7644 8932 7700
rect 8652 7362 8708 7364
rect 8652 7310 8654 7362
rect 8654 7310 8706 7362
rect 8706 7310 8708 7362
rect 8652 7308 8708 7310
rect 9324 6188 9380 6244
rect 8764 4844 8820 4900
rect 10108 12402 10164 12404
rect 10108 12350 10110 12402
rect 10110 12350 10162 12402
rect 10162 12350 10164 12402
rect 10108 12348 10164 12350
rect 10108 11788 10164 11844
rect 9884 10498 9940 10500
rect 9884 10446 9886 10498
rect 9886 10446 9938 10498
rect 9938 10446 9940 10498
rect 9884 10444 9940 10446
rect 9100 4172 9156 4228
rect 10108 11116 10164 11172
rect 10220 9660 10276 9716
rect 10332 9996 10388 10052
rect 10220 9100 10276 9156
rect 10220 8764 10276 8820
rect 9772 8092 9828 8148
rect 9884 7250 9940 7252
rect 9884 7198 9886 7250
rect 9886 7198 9938 7250
rect 9938 7198 9940 7250
rect 9884 7196 9940 7198
rect 9772 5292 9828 5348
rect 10108 6860 10164 6916
rect 10108 4732 10164 4788
rect 9772 4226 9828 4228
rect 9772 4174 9774 4226
rect 9774 4174 9826 4226
rect 9826 4174 9828 4226
rect 9772 4172 9828 4174
rect 10220 3724 10276 3780
rect 9772 1820 9828 1876
rect 11340 13186 11396 13188
rect 11340 13134 11342 13186
rect 11342 13134 11394 13186
rect 11394 13134 11396 13186
rect 11340 13132 11396 13134
rect 11004 12348 11060 12404
rect 11900 13916 11956 13972
rect 11900 13692 11956 13748
rect 12012 12402 12068 12404
rect 12012 12350 12014 12402
rect 12014 12350 12066 12402
rect 12066 12350 12068 12402
rect 12012 12348 12068 12350
rect 11004 12178 11060 12180
rect 11004 12126 11006 12178
rect 11006 12126 11058 12178
rect 11058 12126 11060 12178
rect 11004 12124 11060 12126
rect 10668 12066 10724 12068
rect 10668 12014 10670 12066
rect 10670 12014 10722 12066
rect 10722 12014 10724 12066
rect 10668 12012 10724 12014
rect 11564 12124 11620 12180
rect 11340 10556 11396 10612
rect 11116 10108 11172 10164
rect 10444 9100 10500 9156
rect 10556 7196 10612 7252
rect 11340 7644 11396 7700
rect 11116 6690 11172 6692
rect 11116 6638 11118 6690
rect 11118 6638 11170 6690
rect 11170 6638 11172 6690
rect 11116 6636 11172 6638
rect 10892 5068 10948 5124
rect 10444 3164 10500 3220
rect 12796 12348 12852 12404
rect 12908 13916 12964 13972
rect 13244 13132 13300 13188
rect 13356 13244 13412 13300
rect 13468 12460 13524 12516
rect 11676 10610 11732 10612
rect 11676 10558 11678 10610
rect 11678 10558 11730 10610
rect 11730 10558 11732 10610
rect 11676 10556 11732 10558
rect 12572 10556 12628 10612
rect 11900 10444 11956 10500
rect 12124 10498 12180 10500
rect 12124 10446 12126 10498
rect 12126 10446 12178 10498
rect 12178 10446 12180 10498
rect 12124 10444 12180 10446
rect 11900 10108 11956 10164
rect 11564 9548 11620 9604
rect 11676 9660 11732 9716
rect 11788 9100 11844 9156
rect 12012 8988 12068 9044
rect 12124 8428 12180 8484
rect 11900 8316 11956 8372
rect 12348 10108 12404 10164
rect 12460 8482 12516 8484
rect 12460 8430 12462 8482
rect 12462 8430 12514 8482
rect 12514 8430 12516 8482
rect 12460 8428 12516 8430
rect 13580 12012 13636 12068
rect 13804 13356 13860 13412
rect 14364 13580 14420 13636
rect 13580 11004 13636 11060
rect 13132 10108 13188 10164
rect 13356 10108 13412 10164
rect 12908 9996 12964 10052
rect 12908 9154 12964 9156
rect 12908 9102 12910 9154
rect 12910 9102 12962 9154
rect 12962 9102 12964 9154
rect 12908 9100 12964 9102
rect 13020 8428 13076 8484
rect 13244 9660 13300 9716
rect 12348 8092 12404 8148
rect 12908 8316 12964 8372
rect 12124 7532 12180 7588
rect 12236 7756 12292 7812
rect 11788 6690 11844 6692
rect 11788 6638 11790 6690
rect 11790 6638 11842 6690
rect 11842 6638 11844 6690
rect 11788 6636 11844 6638
rect 11788 6188 11844 6244
rect 11788 5122 11844 5124
rect 11788 5070 11790 5122
rect 11790 5070 11842 5122
rect 11842 5070 11844 5122
rect 11788 5068 11844 5070
rect 11676 4956 11732 5012
rect 10332 2940 10388 2996
rect 9884 1596 9940 1652
rect 10780 2268 10836 2324
rect 8540 364 8596 420
rect 9436 140 9492 196
rect 9884 140 9940 196
rect 12124 7250 12180 7252
rect 12124 7198 12126 7250
rect 12126 7198 12178 7250
rect 12178 7198 12180 7250
rect 12124 7196 12180 7198
rect 12012 6076 12068 6132
rect 12796 7756 12852 7812
rect 12684 7084 12740 7140
rect 12796 7420 12852 7476
rect 12236 5068 12292 5124
rect 12124 5010 12180 5012
rect 12124 4958 12126 5010
rect 12126 4958 12178 5010
rect 12178 4958 12180 5010
rect 12124 4956 12180 4958
rect 12460 6076 12516 6132
rect 12460 5068 12516 5124
rect 13132 7420 13188 7476
rect 13132 7084 13188 7140
rect 13020 6748 13076 6804
rect 13020 3836 13076 3892
rect 12796 3388 12852 3444
rect 12348 2492 12404 2548
rect 11676 1372 11732 1428
rect 11564 1148 11620 1204
rect 11452 140 11508 196
rect 14252 12124 14308 12180
rect 14252 11900 14308 11956
rect 14252 10498 14308 10500
rect 14252 10446 14254 10498
rect 14254 10446 14306 10498
rect 14306 10446 14308 10498
rect 14252 10444 14308 10446
rect 13468 8370 13524 8372
rect 13468 8318 13470 8370
rect 13470 8318 13522 8370
rect 13522 8318 13524 8370
rect 13468 8316 13524 8318
rect 13356 7980 13412 8036
rect 13580 7474 13636 7476
rect 13580 7422 13582 7474
rect 13582 7422 13634 7474
rect 13634 7422 13636 7474
rect 13580 7420 13636 7422
rect 13356 6748 13412 6804
rect 13356 5122 13412 5124
rect 13356 5070 13358 5122
rect 13358 5070 13410 5122
rect 13410 5070 13412 5122
rect 13356 5068 13412 5070
rect 13468 4956 13524 5012
rect 13468 4620 13524 4676
rect 14028 8428 14084 8484
rect 13916 8370 13972 8372
rect 13916 8318 13918 8370
rect 13918 8318 13970 8370
rect 13970 8318 13972 8370
rect 13916 8316 13972 8318
rect 14028 7756 14084 7812
rect 13916 7196 13972 7252
rect 14364 9100 14420 9156
rect 14476 12796 14532 12852
rect 14364 8316 14420 8372
rect 14812 13804 14868 13860
rect 15036 13244 15092 13300
rect 14924 13074 14980 13076
rect 14924 13022 14926 13074
rect 14926 13022 14978 13074
rect 14978 13022 14980 13074
rect 14924 13020 14980 13022
rect 14812 12402 14868 12404
rect 14812 12350 14814 12402
rect 14814 12350 14866 12402
rect 14866 12350 14868 12402
rect 14812 12348 14868 12350
rect 14476 7756 14532 7812
rect 14476 7474 14532 7476
rect 14476 7422 14478 7474
rect 14478 7422 14530 7474
rect 14530 7422 14532 7474
rect 14476 7420 14532 7422
rect 14364 7250 14420 7252
rect 14364 7198 14366 7250
rect 14366 7198 14418 7250
rect 14418 7198 14420 7250
rect 14364 7196 14420 7198
rect 14140 6300 14196 6356
rect 14252 5852 14308 5908
rect 14252 5068 14308 5124
rect 13804 4172 13860 4228
rect 13356 3612 13412 3668
rect 13356 3276 13412 3332
rect 13244 588 13300 644
rect 11900 140 11956 196
rect 13468 140 13524 196
rect 14812 9324 14868 9380
rect 14700 8540 14756 8596
rect 14700 7420 14756 7476
rect 14588 5740 14644 5796
rect 14700 5180 14756 5236
rect 15260 12572 15316 12628
rect 15148 12124 15204 12180
rect 15148 11452 15204 11508
rect 14924 4508 14980 4564
rect 15372 12178 15428 12180
rect 15372 12126 15374 12178
rect 15374 12126 15426 12178
rect 15426 12126 15428 12178
rect 15372 12124 15428 12126
rect 15820 13244 15876 13300
rect 15596 12684 15652 12740
rect 15260 9212 15316 9268
rect 15148 7084 15204 7140
rect 15708 11564 15764 11620
rect 15932 12348 15988 12404
rect 16380 12402 16436 12404
rect 16380 12350 16382 12402
rect 16382 12350 16434 12402
rect 16434 12350 16436 12402
rect 16380 12348 16436 12350
rect 15596 9212 15652 9268
rect 15372 7308 15428 7364
rect 15484 8988 15540 9044
rect 15260 6972 15316 7028
rect 15596 6412 15652 6468
rect 15484 5292 15540 5348
rect 15484 4620 15540 4676
rect 15036 4284 15092 4340
rect 15260 4508 15316 4564
rect 15148 3836 15204 3892
rect 15036 3724 15092 3780
rect 15036 2940 15092 2996
rect 14924 2828 14980 2884
rect 15260 2380 15316 2436
rect 15372 4396 15428 4452
rect 15484 3276 15540 3332
rect 15372 2156 15428 2212
rect 15484 1708 15540 1764
rect 14364 476 14420 532
rect 13916 140 13972 196
rect 15820 10108 15876 10164
rect 16044 9884 16100 9940
rect 16044 9548 16100 9604
rect 16828 13020 16884 13076
rect 16828 12460 16884 12516
rect 16156 8428 16212 8484
rect 16604 10556 16660 10612
rect 30044 14140 30100 14196
rect 17164 13020 17220 13076
rect 16940 11676 16996 11732
rect 16716 9772 16772 9828
rect 16716 8764 16772 8820
rect 16716 8204 16772 8260
rect 16604 7980 16660 8036
rect 16380 7868 16436 7924
rect 15708 5852 15764 5908
rect 15820 7756 15876 7812
rect 15820 7532 15876 7588
rect 16044 7756 16100 7812
rect 15932 6076 15988 6132
rect 16156 7586 16212 7588
rect 16156 7534 16158 7586
rect 16158 7534 16210 7586
rect 16210 7534 16212 7586
rect 16156 7532 16212 7534
rect 16380 6748 16436 6804
rect 16268 6412 16324 6468
rect 16716 6412 16772 6468
rect 16716 6188 16772 6244
rect 16044 5964 16100 6020
rect 16268 5852 16324 5908
rect 16044 5516 16100 5572
rect 16044 5292 16100 5348
rect 15820 5068 15876 5124
rect 17388 13186 17444 13188
rect 17388 13134 17390 13186
rect 17390 13134 17442 13186
rect 17442 13134 17444 13186
rect 17388 13132 17444 13134
rect 17276 12348 17332 12404
rect 17164 10444 17220 10500
rect 17388 9826 17444 9828
rect 17388 9774 17390 9826
rect 17390 9774 17442 9826
rect 17442 9774 17444 9826
rect 17388 9772 17444 9774
rect 17500 9548 17556 9604
rect 18620 13132 18676 13188
rect 18956 13186 19012 13188
rect 18956 13134 18958 13186
rect 18958 13134 19010 13186
rect 19010 13134 19012 13186
rect 18956 13132 19012 13134
rect 18172 11900 18228 11956
rect 18060 11394 18116 11396
rect 18060 11342 18062 11394
rect 18062 11342 18114 11394
rect 18114 11342 18116 11394
rect 18060 11340 18116 11342
rect 18284 11676 18340 11732
rect 18396 12124 18452 12180
rect 19964 13132 20020 13188
rect 19292 12684 19348 12740
rect 18396 11228 18452 11284
rect 18172 11116 18228 11172
rect 18284 10722 18340 10724
rect 18284 10670 18286 10722
rect 18286 10670 18338 10722
rect 18338 10670 18340 10722
rect 18284 10668 18340 10670
rect 19180 10722 19236 10724
rect 19180 10670 19182 10722
rect 19182 10670 19234 10722
rect 19234 10670 19236 10722
rect 19180 10668 19236 10670
rect 19516 11788 19572 11844
rect 19964 12012 20020 12068
rect 19516 11452 19572 11508
rect 19964 11452 20020 11508
rect 19516 10780 19572 10836
rect 19292 10556 19348 10612
rect 19404 10668 19460 10724
rect 18732 10444 18788 10500
rect 17836 10108 17892 10164
rect 18060 9996 18116 10052
rect 17724 9436 17780 9492
rect 18284 9436 18340 9492
rect 18284 9212 18340 9268
rect 17836 8428 17892 8484
rect 17724 7362 17780 7364
rect 17724 7310 17726 7362
rect 17726 7310 17778 7362
rect 17778 7310 17780 7362
rect 17724 7308 17780 7310
rect 17724 6748 17780 6804
rect 16940 5628 16996 5684
rect 17052 6636 17108 6692
rect 16604 5346 16660 5348
rect 16604 5294 16606 5346
rect 16606 5294 16658 5346
rect 16658 5294 16660 5346
rect 16604 5292 16660 5294
rect 16380 5180 16436 5236
rect 17052 5180 17108 5236
rect 15596 1484 15652 1540
rect 17612 5964 17668 6020
rect 17724 4956 17780 5012
rect 18284 8428 18340 8484
rect 18844 9996 18900 10052
rect 18732 9772 18788 9828
rect 18956 9436 19012 9492
rect 19180 9436 19236 9492
rect 19292 9548 19348 9604
rect 18844 9212 18900 9268
rect 18620 8540 18676 8596
rect 18508 7980 18564 8036
rect 18284 7532 18340 7588
rect 18284 7362 18340 7364
rect 18284 7310 18286 7362
rect 18286 7310 18338 7362
rect 18338 7310 18340 7362
rect 18284 7308 18340 7310
rect 18396 6636 18452 6692
rect 18732 7644 18788 7700
rect 19180 7980 19236 8036
rect 19628 7756 19684 7812
rect 19404 7644 19460 7700
rect 18844 6690 18900 6692
rect 18844 6638 18846 6690
rect 18846 6638 18898 6690
rect 18898 6638 18900 6690
rect 18844 6636 18900 6638
rect 18508 6076 18564 6132
rect 18396 5068 18452 5124
rect 18284 4956 18340 5012
rect 17836 3612 17892 3668
rect 17948 4284 18004 4340
rect 18508 4620 18564 4676
rect 18396 4284 18452 4340
rect 18844 5068 18900 5124
rect 19292 7362 19348 7364
rect 19292 7310 19294 7362
rect 19294 7310 19346 7362
rect 19346 7310 19348 7362
rect 19292 7308 19348 7310
rect 19516 7532 19572 7588
rect 20636 13916 20692 13972
rect 20524 12796 20580 12852
rect 21308 12684 21364 12740
rect 21420 12908 21476 12964
rect 21980 12684 22036 12740
rect 20860 12460 20916 12516
rect 20188 10556 20244 10612
rect 20412 10892 20468 10948
rect 20076 10386 20132 10388
rect 20076 10334 20078 10386
rect 20078 10334 20130 10386
rect 20130 10334 20132 10386
rect 20076 10332 20132 10334
rect 19964 10108 20020 10164
rect 20300 9826 20356 9828
rect 20300 9774 20302 9826
rect 20302 9774 20354 9826
rect 20354 9774 20356 9826
rect 20300 9772 20356 9774
rect 20188 9100 20244 9156
rect 19964 8764 20020 8820
rect 20300 8988 20356 9044
rect 20188 8428 20244 8484
rect 20076 7644 20132 7700
rect 19740 7308 19796 7364
rect 19964 7308 20020 7364
rect 20076 6860 20132 6916
rect 19404 6188 19460 6244
rect 19404 5852 19460 5908
rect 19404 5068 19460 5124
rect 19628 4956 19684 5012
rect 19628 4620 19684 4676
rect 18732 3948 18788 4004
rect 18956 4060 19012 4116
rect 18396 3500 18452 3556
rect 18620 3388 18676 3444
rect 17276 588 17332 644
rect 18620 2716 18676 2772
rect 18732 3052 18788 3108
rect 18508 2492 18564 2548
rect 18396 2156 18452 2212
rect 18508 2044 18564 2100
rect 18508 1596 18564 1652
rect 18732 812 18788 868
rect 18396 700 18452 756
rect 19180 4060 19236 4116
rect 19068 3666 19124 3668
rect 19068 3614 19070 3666
rect 19070 3614 19122 3666
rect 19122 3614 19124 3666
rect 19068 3612 19124 3614
rect 20076 4844 20132 4900
rect 19180 3164 19236 3220
rect 20188 4732 20244 4788
rect 20860 12290 20916 12292
rect 20860 12238 20862 12290
rect 20862 12238 20914 12290
rect 20914 12238 20916 12290
rect 20860 12236 20916 12238
rect 20636 12178 20692 12180
rect 20636 12126 20638 12178
rect 20638 12126 20690 12178
rect 20690 12126 20692 12178
rect 20636 12124 20692 12126
rect 21420 12178 21476 12180
rect 21420 12126 21422 12178
rect 21422 12126 21474 12178
rect 21474 12126 21476 12178
rect 21420 12124 21476 12126
rect 20524 10332 20580 10388
rect 20636 11788 20692 11844
rect 20524 8876 20580 8932
rect 20412 4620 20468 4676
rect 20524 6636 20580 6692
rect 20188 3164 20244 3220
rect 19964 2268 20020 2324
rect 21196 11788 21252 11844
rect 21084 11676 21140 11732
rect 21308 11676 21364 11732
rect 21084 10498 21140 10500
rect 21084 10446 21086 10498
rect 21086 10446 21138 10498
rect 21138 10446 21140 10498
rect 21084 10444 21140 10446
rect 21084 9826 21140 9828
rect 21084 9774 21086 9826
rect 21086 9774 21138 9826
rect 21138 9774 21140 9826
rect 21084 9772 21140 9774
rect 20860 9324 20916 9380
rect 20748 7756 20804 7812
rect 20860 7532 20916 7588
rect 20748 6188 20804 6244
rect 20860 6860 20916 6916
rect 20748 5404 20804 5460
rect 20748 4956 20804 5012
rect 21308 10892 21364 10948
rect 21420 10444 21476 10500
rect 21308 9548 21364 9604
rect 21532 9938 21588 9940
rect 21532 9886 21534 9938
rect 21534 9886 21586 9938
rect 21586 9886 21588 9938
rect 21532 9884 21588 9886
rect 21420 9212 21476 9268
rect 21868 12460 21924 12516
rect 21756 11340 21812 11396
rect 21756 9548 21812 9604
rect 21868 10332 21924 10388
rect 21644 9212 21700 9268
rect 21532 8988 21588 9044
rect 21196 6860 21252 6916
rect 21308 6188 21364 6244
rect 20972 5292 21028 5348
rect 20972 5122 21028 5124
rect 20972 5070 20974 5122
rect 20974 5070 21026 5122
rect 21026 5070 21028 5122
rect 20972 5068 21028 5070
rect 21308 5122 21364 5124
rect 21308 5070 21310 5122
rect 21310 5070 21362 5122
rect 21362 5070 21364 5122
rect 21308 5068 21364 5070
rect 21420 4732 21476 4788
rect 20636 3388 20692 3444
rect 21756 9042 21812 9044
rect 21756 8990 21758 9042
rect 21758 8990 21810 9042
rect 21810 8990 21812 9042
rect 21756 8988 21812 8990
rect 22540 13132 22596 13188
rect 22428 11228 22484 11284
rect 22092 10108 22148 10164
rect 22204 10220 22260 10276
rect 22092 9938 22148 9940
rect 22092 9886 22094 9938
rect 22094 9886 22146 9938
rect 22146 9886 22148 9938
rect 22092 9884 22148 9886
rect 21980 8818 22036 8820
rect 21980 8766 21982 8818
rect 21982 8766 22034 8818
rect 22034 8766 22036 8818
rect 21980 8764 22036 8766
rect 22316 9884 22372 9940
rect 22316 8988 22372 9044
rect 22428 8876 22484 8932
rect 22204 8764 22260 8820
rect 21644 8204 21700 8260
rect 22092 8092 22148 8148
rect 21644 7196 21700 7252
rect 21644 6972 21700 7028
rect 21644 6188 21700 6244
rect 22204 7756 22260 7812
rect 21868 7196 21924 7252
rect 22204 7084 22260 7140
rect 21868 6524 21924 6580
rect 21756 5964 21812 6020
rect 22204 6018 22260 6020
rect 22204 5966 22206 6018
rect 22206 5966 22258 6018
rect 22258 5966 22260 6018
rect 22204 5964 22260 5966
rect 22988 12684 23044 12740
rect 23884 13804 23940 13860
rect 23100 12348 23156 12404
rect 23548 12402 23604 12404
rect 23548 12350 23550 12402
rect 23550 12350 23602 12402
rect 23602 12350 23604 12402
rect 23548 12348 23604 12350
rect 23996 13468 24052 13524
rect 24108 13132 24164 13188
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24220 12572 24276 12628
rect 24012 12516 24068 12518
rect 23996 12236 24052 12292
rect 23548 11900 23604 11956
rect 23324 11788 23380 11844
rect 23436 11564 23492 11620
rect 23548 11340 23604 11396
rect 23996 11282 24052 11284
rect 23996 11230 23998 11282
rect 23998 11230 24050 11282
rect 24050 11230 24052 11282
rect 23996 11228 24052 11230
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 24220 11004 24276 11060
rect 23324 10220 23380 10276
rect 23100 9660 23156 9716
rect 23212 9884 23268 9940
rect 22764 8316 22820 8372
rect 22876 9436 22932 9492
rect 22652 7980 22708 8036
rect 22876 7980 22932 8036
rect 23212 8204 23268 8260
rect 22540 5628 22596 5684
rect 22652 6524 22708 6580
rect 23212 6188 23268 6244
rect 22652 5292 22708 5348
rect 22428 5180 22484 5236
rect 21868 5122 21924 5124
rect 21868 5070 21870 5122
rect 21870 5070 21922 5122
rect 21922 5070 21924 5122
rect 21868 5068 21924 5070
rect 22316 5122 22372 5124
rect 22316 5070 22318 5122
rect 22318 5070 22370 5122
rect 22370 5070 22372 5122
rect 22316 5068 22372 5070
rect 21532 4620 21588 4676
rect 21308 4338 21364 4340
rect 21308 4286 21310 4338
rect 21310 4286 21362 4338
rect 21362 4286 21364 4338
rect 21308 4284 21364 4286
rect 21868 4284 21924 4340
rect 21644 3724 21700 3780
rect 20524 2156 20580 2212
rect 21756 3500 21812 3556
rect 21756 3164 21812 3220
rect 21756 2828 21812 2884
rect 22092 2380 22148 2436
rect 22540 5068 22596 5124
rect 23212 4956 23268 5012
rect 22540 4284 22596 4340
rect 24220 10220 24276 10276
rect 24220 9996 24276 10052
rect 23996 9938 24052 9940
rect 23996 9886 23998 9938
rect 23998 9886 24050 9938
rect 24050 9886 24052 9938
rect 23996 9884 24052 9886
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24220 9436 24276 9492
rect 24012 9380 24068 9382
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 24444 12236 24500 12292
rect 24556 11900 24612 11956
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 24556 11004 24612 11060
rect 25340 14028 25396 14084
rect 25452 13468 25508 13524
rect 25228 13356 25284 13412
rect 24892 10892 24948 10948
rect 25004 11788 25060 11844
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24444 9938 24500 9940
rect 24444 9886 24446 9938
rect 24446 9886 24498 9938
rect 24498 9886 24500 9938
rect 24444 9884 24500 9886
rect 23548 8652 23604 8708
rect 24556 9660 24612 9716
rect 23548 8204 23604 8260
rect 23548 7868 23604 7924
rect 24780 9772 24836 9828
rect 25900 13580 25956 13636
rect 25900 13244 25956 13300
rect 25788 12460 25844 12516
rect 25452 12236 25508 12292
rect 25340 11788 25396 11844
rect 25116 9772 25172 9828
rect 25228 10668 25284 10724
rect 25340 10444 25396 10500
rect 25340 9996 25396 10052
rect 24892 9324 24948 9380
rect 25004 9212 25060 9268
rect 25004 9042 25060 9044
rect 25004 8990 25006 9042
rect 25006 8990 25058 9042
rect 25058 8990 25060 9042
rect 25004 8988 25060 8990
rect 25228 9212 25284 9268
rect 25228 8876 25284 8932
rect 24220 8204 24276 8260
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24220 7868 24276 7924
rect 24012 7812 24068 7814
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24892 8540 24948 8596
rect 24444 7980 24500 8036
rect 24444 7644 24500 7700
rect 24668 7980 24724 8036
rect 23996 7420 24052 7476
rect 24332 7084 24388 7140
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 23884 6748 23940 6804
rect 24332 6748 24388 6804
rect 23804 6298 23860 6300
rect 23548 6188 23604 6244
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24220 6188 24276 6244
rect 25004 7084 25060 7140
rect 24220 5404 24276 5460
rect 24332 5516 24388 5572
rect 23996 5292 24052 5348
rect 23548 4956 23604 5012
rect 23324 3836 23380 3892
rect 23436 4284 23492 4340
rect 23436 3276 23492 3332
rect 22428 2156 22484 2212
rect 22988 3164 23044 3220
rect 21644 1372 21700 1428
rect 23324 2268 23380 2324
rect 23100 2210 23156 2212
rect 23100 2158 23102 2210
rect 23102 2158 23154 2210
rect 23154 2158 23156 2210
rect 23100 2156 23156 2158
rect 22988 1148 23044 1204
rect 23436 2210 23492 2212
rect 23436 2158 23438 2210
rect 23438 2158 23490 2210
rect 23490 2158 23492 2210
rect 23436 2156 23492 2158
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23660 4620 23716 4676
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24332 4732 24388 4788
rect 24668 4844 24724 4900
rect 24012 4676 24068 4678
rect 24444 4508 24500 4564
rect 24220 4172 24276 4228
rect 23660 3612 23716 3668
rect 24332 3948 24388 4004
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 23660 3052 23716 3108
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24220 3164 24276 3220
rect 25116 6860 25172 6916
rect 25228 6802 25284 6804
rect 25228 6750 25230 6802
rect 25230 6750 25282 6802
rect 25282 6750 25284 6802
rect 25228 6748 25284 6750
rect 26236 12572 26292 12628
rect 26460 14028 26516 14084
rect 25900 12066 25956 12068
rect 25900 12014 25902 12066
rect 25902 12014 25954 12066
rect 25954 12014 25956 12066
rect 25900 12012 25956 12014
rect 25564 11452 25620 11508
rect 26348 11900 26404 11956
rect 25676 10892 25732 10948
rect 25676 10444 25732 10500
rect 25452 9884 25508 9940
rect 25452 9212 25508 9268
rect 25340 4956 25396 5012
rect 25452 8876 25508 8932
rect 26012 10892 26068 10948
rect 26012 9660 26068 9716
rect 26236 10220 26292 10276
rect 26572 13916 26628 13972
rect 26684 13692 26740 13748
rect 26796 13916 26852 13972
rect 26796 13244 26852 13300
rect 27356 13692 27412 13748
rect 27132 12236 27188 12292
rect 27244 12460 27300 12516
rect 26572 10498 26628 10500
rect 26572 10446 26574 10498
rect 26574 10446 26626 10498
rect 26626 10446 26628 10498
rect 26572 10444 26628 10446
rect 26460 10220 26516 10276
rect 26236 9548 26292 9604
rect 26012 8092 26068 8148
rect 26124 8876 26180 8932
rect 25788 7420 25844 7476
rect 25676 5794 25732 5796
rect 25676 5742 25678 5794
rect 25678 5742 25730 5794
rect 25730 5742 25732 5794
rect 25676 5740 25732 5742
rect 25676 5516 25732 5572
rect 25676 5180 25732 5236
rect 26012 3836 26068 3892
rect 24012 3108 24068 3110
rect 24780 2882 24836 2884
rect 24780 2830 24782 2882
rect 24782 2830 24834 2882
rect 24834 2830 24836 2882
rect 24780 2828 24836 2830
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24332 2156 24388 2212
rect 23436 1708 23492 1764
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 23324 1148 23380 1204
rect 23548 1372 23604 1428
rect 18956 140 19012 196
rect 19516 1036 19572 1092
rect 21532 1036 21588 1092
rect 23996 924 24052 980
rect 25116 2716 25172 2772
rect 25116 2156 25172 2212
rect 26012 3276 26068 3332
rect 25564 2268 25620 2324
rect 25676 2828 25732 2884
rect 25228 1596 25284 1652
rect 26012 2828 26068 2884
rect 25788 1708 25844 1764
rect 26012 1484 26068 1540
rect 25788 1372 25844 1428
rect 26572 8988 26628 9044
rect 26796 8988 26852 9044
rect 26460 7980 26516 8036
rect 26460 6524 26516 6580
rect 26236 5906 26292 5908
rect 26236 5854 26238 5906
rect 26238 5854 26290 5906
rect 26290 5854 26292 5906
rect 26236 5852 26292 5854
rect 27020 11116 27076 11172
rect 27020 10892 27076 10948
rect 27020 9602 27076 9604
rect 27020 9550 27022 9602
rect 27022 9550 27074 9602
rect 27074 9550 27076 9602
rect 27020 9548 27076 9550
rect 27244 9436 27300 9492
rect 27468 12572 27524 12628
rect 28028 13804 28084 13860
rect 27580 11788 27636 11844
rect 27692 13468 27748 13524
rect 27468 11564 27524 11620
rect 27580 10444 27636 10500
rect 27580 9660 27636 9716
rect 27356 9324 27412 9380
rect 27020 8540 27076 8596
rect 27244 8428 27300 8484
rect 28252 13132 28308 13188
rect 28140 11116 28196 11172
rect 28924 13356 28980 13412
rect 28476 12124 28532 12180
rect 28700 12460 28756 12516
rect 29372 12236 29428 12292
rect 29484 12124 29540 12180
rect 29260 11788 29316 11844
rect 28700 10668 28756 10724
rect 28924 11676 28980 11732
rect 28364 10444 28420 10500
rect 28588 10220 28644 10276
rect 28028 8370 28084 8372
rect 28028 8318 28030 8370
rect 28030 8318 28082 8370
rect 28082 8318 28084 8370
rect 28028 8316 28084 8318
rect 27692 7868 27748 7924
rect 27020 6636 27076 6692
rect 26796 6076 26852 6132
rect 28252 9772 28308 9828
rect 28252 6860 28308 6916
rect 28812 9324 28868 9380
rect 28700 8652 28756 8708
rect 28476 8316 28532 8372
rect 28476 6972 28532 7028
rect 28364 6748 28420 6804
rect 28588 6748 28644 6804
rect 28476 6636 28532 6692
rect 28476 6412 28532 6468
rect 26460 5964 26516 6020
rect 26348 5740 26404 5796
rect 26572 5852 26628 5908
rect 26236 5292 26292 5348
rect 27356 5852 27412 5908
rect 27580 5852 27636 5908
rect 27132 5740 27188 5796
rect 27692 5628 27748 5684
rect 28252 5740 28308 5796
rect 28364 5628 28420 5684
rect 26684 5068 26740 5124
rect 27580 5068 27636 5124
rect 27468 4956 27524 5012
rect 26908 4844 26964 4900
rect 27804 5068 27860 5124
rect 26572 4172 26628 4228
rect 26236 3052 26292 3108
rect 26348 3500 26404 3556
rect 24220 924 24276 980
rect 24464 810 24520 812
rect 24332 700 24388 756
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 25564 812 25620 868
rect 24672 756 24728 758
rect 24892 700 24948 756
rect 23996 252 24052 308
rect 27356 4060 27412 4116
rect 26796 3554 26852 3556
rect 26796 3502 26798 3554
rect 26798 3502 26850 3554
rect 26850 3502 26852 3554
rect 26796 3500 26852 3502
rect 26684 3388 26740 3444
rect 27468 3612 27524 3668
rect 27804 4172 27860 4228
rect 27020 3164 27076 3220
rect 26796 2044 26852 2100
rect 26796 1036 26852 1092
rect 26572 252 26628 308
rect 27692 2940 27748 2996
rect 27804 3724 27860 3780
rect 29260 9772 29316 9828
rect 29372 10444 29428 10500
rect 30044 13804 30100 13860
rect 29820 11900 29876 11956
rect 30156 12348 30212 12404
rect 29820 10892 29876 10948
rect 29708 10220 29764 10276
rect 29484 9212 29540 9268
rect 30156 10668 30212 10724
rect 30044 10220 30100 10276
rect 29932 9884 29988 9940
rect 30156 9884 30212 9940
rect 29820 8988 29876 9044
rect 29596 7756 29652 7812
rect 28812 7420 28868 7476
rect 28924 6748 28980 6804
rect 28700 5068 28756 5124
rect 28476 4956 28532 5012
rect 28588 4114 28644 4116
rect 28588 4062 28590 4114
rect 28590 4062 28642 4114
rect 28642 4062 28644 4114
rect 28588 4060 28644 4062
rect 28812 5628 28868 5684
rect 29148 5852 29204 5908
rect 29036 5794 29092 5796
rect 29036 5742 29038 5794
rect 29038 5742 29090 5794
rect 29090 5742 29092 5794
rect 29036 5740 29092 5742
rect 28924 4956 28980 5012
rect 28812 4284 28868 4340
rect 28364 3052 28420 3108
rect 28700 3666 28756 3668
rect 28700 3614 28702 3666
rect 28702 3614 28754 3666
rect 28754 3614 28756 3666
rect 28700 3612 28756 3614
rect 28812 2380 28868 2436
rect 28924 2882 28980 2884
rect 28924 2830 28926 2882
rect 28926 2830 28978 2882
rect 28978 2830 28980 2882
rect 28924 2828 28980 2830
rect 29260 7308 29316 7364
rect 29260 5740 29316 5796
rect 30044 6860 30100 6916
rect 29820 5852 29876 5908
rect 29708 5740 29764 5796
rect 29708 5068 29764 5124
rect 29596 4284 29652 4340
rect 29708 3500 29764 3556
rect 29484 2940 29540 2996
rect 28140 1986 28196 1988
rect 28140 1934 28142 1986
rect 28142 1934 28194 1986
rect 28194 1934 28196 1986
rect 28140 1932 28196 1934
rect 28476 1932 28532 1988
rect 29932 5682 29988 5684
rect 29932 5630 29934 5682
rect 29934 5630 29986 5682
rect 29986 5630 29988 5682
rect 29932 5628 29988 5630
rect 29820 2828 29876 2884
rect 30940 13804 30996 13860
rect 30716 12460 30772 12516
rect 30828 13356 30884 13412
rect 30492 11564 30548 11620
rect 30380 10220 30436 10276
rect 30380 9324 30436 9380
rect 30604 9714 30660 9716
rect 30604 9662 30606 9714
rect 30606 9662 30658 9714
rect 30658 9662 30660 9714
rect 30604 9660 30660 9662
rect 30716 9436 30772 9492
rect 31052 12290 31108 12292
rect 31052 12238 31054 12290
rect 31054 12238 31106 12290
rect 31106 12238 31108 12290
rect 31052 12236 31108 12238
rect 30940 10444 30996 10500
rect 31612 13580 31668 13636
rect 31388 12850 31444 12852
rect 31388 12798 31390 12850
rect 31390 12798 31442 12850
rect 31442 12798 31444 12850
rect 31388 12796 31444 12798
rect 31724 12796 31780 12852
rect 31388 11788 31444 11844
rect 32508 14028 32564 14084
rect 32284 12850 32340 12852
rect 32284 12798 32286 12850
rect 32286 12798 32338 12850
rect 32338 12798 32340 12850
rect 32284 12796 32340 12798
rect 32508 12460 32564 12516
rect 32284 12236 32340 12292
rect 32172 11004 32228 11060
rect 31164 10220 31220 10276
rect 31276 9996 31332 10052
rect 30828 9324 30884 9380
rect 30940 9548 30996 9604
rect 30716 8988 30772 9044
rect 31276 8876 31332 8932
rect 31724 9548 31780 9604
rect 31500 8540 31556 8596
rect 31164 8146 31220 8148
rect 31164 8094 31166 8146
rect 31166 8094 31218 8146
rect 31218 8094 31220 8146
rect 31164 8092 31220 8094
rect 30492 7308 30548 7364
rect 31388 6972 31444 7028
rect 30268 5852 30324 5908
rect 30380 5516 30436 5572
rect 30716 5628 30772 5684
rect 30156 5068 30212 5124
rect 30156 4508 30212 4564
rect 32284 9436 32340 9492
rect 32284 8988 32340 9044
rect 32172 7420 32228 7476
rect 32508 10780 32564 10836
rect 32620 11676 32676 11732
rect 32508 9548 32564 9604
rect 32508 8764 32564 8820
rect 32844 10892 32900 10948
rect 33292 10892 33348 10948
rect 33852 11564 33908 11620
rect 34748 11676 34804 11732
rect 34860 12012 34916 12068
rect 33628 11004 33684 11060
rect 34300 11228 34356 11284
rect 34412 11004 34468 11060
rect 32844 9100 32900 9156
rect 33068 9212 33124 9268
rect 33628 9324 33684 9380
rect 33628 9100 33684 9156
rect 33516 8988 33572 9044
rect 32956 8428 33012 8484
rect 33292 8482 33348 8484
rect 33292 8430 33294 8482
rect 33294 8430 33346 8482
rect 33346 8430 33348 8482
rect 33292 8428 33348 8430
rect 33516 8482 33572 8484
rect 33516 8430 33518 8482
rect 33518 8430 33570 8482
rect 33570 8430 33572 8482
rect 33516 8428 33572 8430
rect 33404 8204 33460 8260
rect 32620 7644 32676 7700
rect 32732 7084 32788 7140
rect 31724 6636 31780 6692
rect 31388 5404 31444 5460
rect 31276 5292 31332 5348
rect 31500 5292 31556 5348
rect 30044 2828 30100 2884
rect 30380 4060 30436 4116
rect 31500 4060 31556 4116
rect 31500 3612 31556 3668
rect 30940 3052 30996 3108
rect 29708 2156 29764 2212
rect 29596 1874 29652 1876
rect 29596 1822 29598 1874
rect 29598 1822 29650 1874
rect 29650 1822 29652 1874
rect 29596 1820 29652 1822
rect 29484 1372 29540 1428
rect 29596 1484 29652 1540
rect 28476 1148 28532 1204
rect 27804 140 27860 196
rect 30156 2210 30212 2212
rect 30156 2158 30158 2210
rect 30158 2158 30210 2210
rect 30210 2158 30212 2210
rect 30156 2156 30212 2158
rect 30492 2210 30548 2212
rect 30492 2158 30494 2210
rect 30494 2158 30546 2210
rect 30546 2158 30548 2210
rect 30492 2156 30548 2158
rect 30156 1820 30212 1876
rect 29932 812 29988 868
rect 30044 1708 30100 1764
rect 30156 700 30212 756
rect 30044 364 30100 420
rect 31836 6076 31892 6132
rect 32284 6636 32340 6692
rect 32060 5794 32116 5796
rect 32060 5742 32062 5794
rect 32062 5742 32114 5794
rect 32114 5742 32116 5794
rect 32060 5740 32116 5742
rect 31836 5516 31892 5572
rect 32060 5516 32116 5572
rect 31948 5404 32004 5460
rect 31836 4172 31892 4228
rect 31836 3612 31892 3668
rect 32620 6130 32676 6132
rect 32620 6078 32622 6130
rect 32622 6078 32674 6130
rect 32674 6078 32676 6130
rect 32620 6076 32676 6078
rect 32396 5852 32452 5908
rect 32620 5852 32676 5908
rect 32508 3052 32564 3108
rect 31836 2268 31892 2324
rect 32732 5628 32788 5684
rect 32732 4844 32788 4900
rect 33068 6860 33124 6916
rect 32956 6636 33012 6692
rect 33628 6524 33684 6580
rect 33628 6076 33684 6132
rect 34972 10610 35028 10612
rect 34972 10558 34974 10610
rect 34974 10558 35026 10610
rect 35026 10558 35028 10610
rect 34972 10556 35028 10558
rect 34524 9772 34580 9828
rect 34412 9324 34468 9380
rect 34076 8146 34132 8148
rect 34076 8094 34078 8146
rect 34078 8094 34130 8146
rect 34130 8094 34132 8146
rect 34076 8092 34132 8094
rect 34300 7586 34356 7588
rect 34300 7534 34302 7586
rect 34302 7534 34354 7586
rect 34354 7534 34356 7586
rect 34300 7532 34356 7534
rect 33964 6300 34020 6356
rect 33180 5794 33236 5796
rect 33180 5742 33182 5794
rect 33182 5742 33234 5794
rect 33234 5742 33236 5794
rect 33180 5740 33236 5742
rect 33628 5516 33684 5572
rect 34188 5516 34244 5572
rect 33628 5234 33684 5236
rect 33628 5182 33630 5234
rect 33630 5182 33682 5234
rect 33682 5182 33684 5234
rect 33628 5180 33684 5182
rect 34076 5180 34132 5236
rect 33068 4844 33124 4900
rect 33516 4956 33572 5012
rect 33516 3164 33572 3220
rect 33628 3836 33684 3892
rect 33068 2658 33124 2660
rect 33068 2606 33070 2658
rect 33070 2606 33122 2658
rect 33122 2606 33124 2658
rect 33068 2604 33124 2606
rect 32732 2492 32788 2548
rect 33292 2156 33348 2212
rect 32620 1932 32676 1988
rect 32844 1932 32900 1988
rect 33628 700 33684 756
rect 33740 2380 33796 2436
rect 32844 588 32900 644
rect 33964 2044 34020 2100
rect 33852 1708 33908 1764
rect 33852 1484 33908 1540
rect 33964 476 34020 532
rect 33740 364 33796 420
rect 33628 140 33684 196
rect 34524 7980 34580 8036
rect 34524 5234 34580 5236
rect 34524 5182 34526 5234
rect 34526 5182 34578 5234
rect 34578 5182 34580 5234
rect 34524 5180 34580 5182
rect 34972 8818 35028 8820
rect 34972 8766 34974 8818
rect 34974 8766 35026 8818
rect 35026 8766 35028 8818
rect 34972 8764 35028 8766
rect 35308 13692 35364 13748
rect 36092 13916 36148 13972
rect 35644 13132 35700 13188
rect 35308 13020 35364 13076
rect 36204 12796 36260 12852
rect 35308 12236 35364 12292
rect 35868 11788 35924 11844
rect 35308 11004 35364 11060
rect 35532 11004 35588 11060
rect 35084 8370 35140 8372
rect 35084 8318 35086 8370
rect 35086 8318 35138 8370
rect 35138 8318 35140 8370
rect 35084 8316 35140 8318
rect 35420 7980 35476 8036
rect 35308 7756 35364 7812
rect 34972 7586 35028 7588
rect 34972 7534 34974 7586
rect 34974 7534 35026 7586
rect 35026 7534 35028 7586
rect 34972 7532 35028 7534
rect 35196 7644 35252 7700
rect 34860 5852 34916 5908
rect 34748 5292 34804 5348
rect 34636 4620 34692 4676
rect 34860 5180 34916 5236
rect 35308 5068 35364 5124
rect 35196 4284 35252 4340
rect 34860 4172 34916 4228
rect 34972 4060 35028 4116
rect 35308 4172 35364 4228
rect 35420 3724 35476 3780
rect 35196 3276 35252 3332
rect 35756 10220 35812 10276
rect 35756 8370 35812 8372
rect 35756 8318 35758 8370
rect 35758 8318 35810 8370
rect 35810 8318 35812 8370
rect 35756 8316 35812 8318
rect 35980 10892 36036 10948
rect 35980 10220 36036 10276
rect 35980 8652 36036 8708
rect 36092 7868 36148 7924
rect 35756 7644 35812 7700
rect 35644 7586 35700 7588
rect 35644 7534 35646 7586
rect 35646 7534 35698 7586
rect 35698 7534 35700 7586
rect 35644 7532 35700 7534
rect 35868 7308 35924 7364
rect 35756 6300 35812 6356
rect 35644 5516 35700 5572
rect 36092 7196 36148 7252
rect 35980 5516 36036 5572
rect 35756 5068 35812 5124
rect 35756 4732 35812 4788
rect 36316 12236 36372 12292
rect 36988 13244 37044 13300
rect 36876 13020 36932 13076
rect 36988 12348 37044 12404
rect 36540 11340 36596 11396
rect 36764 11676 36820 11732
rect 36540 10892 36596 10948
rect 36316 9042 36372 9044
rect 36316 8990 36318 9042
rect 36318 8990 36370 9042
rect 36370 8990 36372 9042
rect 36316 8988 36372 8990
rect 36428 8204 36484 8260
rect 36316 7532 36372 7588
rect 36316 7362 36372 7364
rect 36316 7310 36318 7362
rect 36318 7310 36370 7362
rect 36370 7310 36372 7362
rect 36316 7308 36372 7310
rect 36652 8988 36708 9044
rect 36652 7308 36708 7364
rect 36428 7196 36484 7252
rect 36876 8316 36932 8372
rect 37324 11788 37380 11844
rect 38332 13580 38388 13636
rect 38780 12908 38836 12964
rect 37884 12290 37940 12292
rect 37884 12238 37886 12290
rect 37886 12238 37938 12290
rect 37938 12238 37940 12290
rect 37884 12236 37940 12238
rect 37884 11340 37940 11396
rect 37324 10332 37380 10388
rect 37436 8258 37492 8260
rect 37436 8206 37438 8258
rect 37438 8206 37490 8258
rect 37490 8206 37492 8258
rect 37436 8204 37492 8206
rect 36764 6636 36820 6692
rect 37212 7980 37268 8036
rect 37100 7532 37156 7588
rect 37772 8204 37828 8260
rect 37772 7980 37828 8036
rect 37548 7196 37604 7252
rect 37772 6636 37828 6692
rect 37772 6300 37828 6356
rect 38220 11788 38276 11844
rect 37996 11228 38052 11284
rect 38332 11340 38388 11396
rect 38108 9212 38164 9268
rect 38220 9100 38276 9156
rect 37996 8370 38052 8372
rect 37996 8318 37998 8370
rect 37998 8318 38050 8370
rect 38050 8318 38052 8370
rect 37996 8316 38052 8318
rect 37996 7980 38052 8036
rect 37996 6300 38052 6356
rect 36876 5180 36932 5236
rect 37100 5180 37156 5236
rect 39004 9772 39060 9828
rect 38332 7756 38388 7812
rect 38444 7868 38500 7924
rect 39004 8482 39060 8484
rect 39004 8430 39006 8482
rect 39006 8430 39058 8482
rect 39058 8430 39060 8482
rect 39004 8428 39060 8430
rect 38556 8204 38612 8260
rect 38780 8204 38836 8260
rect 38780 7868 38836 7924
rect 39900 12236 39956 12292
rect 39900 11676 39956 11732
rect 39676 11004 39732 11060
rect 40012 10668 40068 10724
rect 40124 13468 40180 13524
rect 39452 9996 39508 10052
rect 39900 9996 39956 10052
rect 39452 9042 39508 9044
rect 39452 8990 39454 9042
rect 39454 8990 39506 9042
rect 39506 8990 39508 9042
rect 39452 8988 39508 8990
rect 39676 8930 39732 8932
rect 39676 8878 39678 8930
rect 39678 8878 39730 8930
rect 39730 8878 39732 8930
rect 39676 8876 39732 8878
rect 40012 8764 40068 8820
rect 39564 8540 39620 8596
rect 39228 7868 39284 7924
rect 39340 7980 39396 8036
rect 37436 5516 37492 5572
rect 37436 4620 37492 4676
rect 36204 3948 36260 4004
rect 37660 3724 37716 3780
rect 36092 3276 36148 3332
rect 37324 3330 37380 3332
rect 37324 3278 37326 3330
rect 37326 3278 37378 3330
rect 37378 3278 37380 3330
rect 37324 3276 37380 3278
rect 36764 3052 36820 3108
rect 36764 2716 36820 2772
rect 36204 2268 36260 2324
rect 37100 2044 37156 2100
rect 37100 1596 37156 1652
rect 34412 140 34468 196
rect 35644 1484 35700 1540
rect 38220 5180 38276 5236
rect 38668 6860 38724 6916
rect 38556 6188 38612 6244
rect 38444 5906 38500 5908
rect 38444 5854 38446 5906
rect 38446 5854 38498 5906
rect 38498 5854 38500 5906
rect 38444 5852 38500 5854
rect 39452 6636 39508 6692
rect 38668 5740 38724 5796
rect 39228 5906 39284 5908
rect 39228 5854 39230 5906
rect 39230 5854 39282 5906
rect 39282 5854 39284 5906
rect 39228 5852 39284 5854
rect 41020 13804 41076 13860
rect 41356 12572 41412 12628
rect 40572 11340 40628 11396
rect 41244 12124 41300 12180
rect 41804 13132 41860 13188
rect 41804 12178 41860 12180
rect 41804 12126 41806 12178
rect 41806 12126 41858 12178
rect 41858 12126 41860 12178
rect 41804 12124 41860 12126
rect 42140 13186 42196 13188
rect 42140 13134 42142 13186
rect 42142 13134 42194 13186
rect 42194 13134 42196 13186
rect 42140 13132 42196 13134
rect 42252 12684 42308 12740
rect 42812 13356 42868 13412
rect 42588 13132 42644 13188
rect 42364 12348 42420 12404
rect 42476 12908 42532 12964
rect 42028 12124 42084 12180
rect 41468 11564 41524 11620
rect 41916 11452 41972 11508
rect 40460 10386 40516 10388
rect 40460 10334 40462 10386
rect 40462 10334 40514 10386
rect 40514 10334 40516 10386
rect 40460 10332 40516 10334
rect 40124 8316 40180 8372
rect 40236 9436 40292 9492
rect 40124 7644 40180 7700
rect 39788 6188 39844 6244
rect 38668 5234 38724 5236
rect 38668 5182 38670 5234
rect 38670 5182 38722 5234
rect 38722 5182 38724 5234
rect 38668 5180 38724 5182
rect 38332 3276 38388 3332
rect 38444 4284 38500 4340
rect 39676 5234 39732 5236
rect 39676 5182 39678 5234
rect 39678 5182 39730 5234
rect 39730 5182 39732 5234
rect 39676 5180 39732 5182
rect 40684 9996 40740 10052
rect 40908 10220 40964 10276
rect 40684 8764 40740 8820
rect 40572 8540 40628 8596
rect 40684 8316 40740 8372
rect 41580 9996 41636 10052
rect 41132 8988 41188 9044
rect 41468 8930 41524 8932
rect 41468 8878 41470 8930
rect 41470 8878 41522 8930
rect 41522 8878 41524 8930
rect 41468 8876 41524 8878
rect 41244 8316 41300 8372
rect 40908 7980 40964 8036
rect 40684 7084 40740 7140
rect 40796 7868 40852 7924
rect 40236 6636 40292 6692
rect 40684 6748 40740 6804
rect 40460 6300 40516 6356
rect 40124 5964 40180 6020
rect 40572 5852 40628 5908
rect 40348 3836 40404 3892
rect 39004 3164 39060 3220
rect 38892 2156 38948 2212
rect 38780 1932 38836 1988
rect 38332 1708 38388 1764
rect 38668 1708 38724 1764
rect 37660 1260 37716 1316
rect 37884 1260 37940 1316
rect 37212 812 37268 868
rect 38780 924 38836 980
rect 38892 588 38948 644
rect 39004 364 39060 420
rect 40684 5740 40740 5796
rect 40684 4844 40740 4900
rect 40684 4620 40740 4676
rect 40684 2828 40740 2884
rect 40348 2716 40404 2772
rect 40348 1820 40404 1876
rect 39788 1484 39844 1540
rect 40236 1708 40292 1764
rect 41020 7868 41076 7924
rect 42252 10332 42308 10388
rect 42140 10050 42196 10052
rect 42140 9998 42142 10050
rect 42142 9998 42194 10050
rect 42194 9998 42196 10050
rect 42140 9996 42196 9998
rect 42364 10220 42420 10276
rect 43708 13132 43764 13188
rect 43260 12460 43316 12516
rect 43484 12908 43540 12964
rect 43260 12236 43316 12292
rect 42700 12178 42756 12180
rect 42700 12126 42702 12178
rect 42702 12126 42754 12178
rect 42754 12126 42756 12178
rect 42700 12124 42756 12126
rect 43148 11004 43204 11060
rect 42476 10108 42532 10164
rect 42588 9996 42644 10052
rect 42364 9212 42420 9268
rect 42028 8818 42084 8820
rect 42028 8766 42030 8818
rect 42030 8766 42082 8818
rect 42082 8766 42084 8818
rect 42028 8764 42084 8766
rect 42252 8428 42308 8484
rect 41692 7868 41748 7924
rect 41356 6860 41412 6916
rect 42140 7868 42196 7924
rect 41804 7308 41860 7364
rect 42028 6802 42084 6804
rect 42028 6750 42030 6802
rect 42030 6750 42082 6802
rect 42082 6750 42084 6802
rect 42028 6748 42084 6750
rect 41468 6636 41524 6692
rect 41468 6300 41524 6356
rect 42252 7250 42308 7252
rect 42252 7198 42254 7250
rect 42254 7198 42306 7250
rect 42306 7198 42308 7250
rect 42252 7196 42308 7198
rect 43148 9212 43204 9268
rect 43148 9042 43204 9044
rect 43148 8990 43150 9042
rect 43150 8990 43202 9042
rect 43202 8990 43204 9042
rect 43148 8988 43204 8990
rect 43260 8876 43316 8932
rect 43372 10220 43428 10276
rect 43372 8204 43428 8260
rect 42364 6748 42420 6804
rect 42252 6300 42308 6356
rect 41804 6018 41860 6020
rect 41804 5966 41806 6018
rect 41806 5966 41858 6018
rect 41858 5966 41860 6018
rect 41804 5964 41860 5966
rect 42140 5404 42196 5460
rect 41244 5292 41300 5348
rect 41132 5180 41188 5236
rect 42028 5068 42084 5124
rect 41916 4956 41972 5012
rect 41692 3836 41748 3892
rect 41580 2882 41636 2884
rect 41580 2830 41582 2882
rect 41582 2830 41634 2882
rect 41634 2830 41636 2882
rect 41580 2828 41636 2830
rect 40908 2210 40964 2212
rect 40908 2158 40910 2210
rect 40910 2158 40962 2210
rect 40962 2158 40964 2210
rect 40908 2156 40964 2158
rect 41132 2210 41188 2212
rect 41132 2158 41134 2210
rect 41134 2158 41186 2210
rect 41186 2158 41188 2210
rect 41132 2156 41188 2158
rect 42700 7196 42756 7252
rect 43148 7250 43204 7252
rect 43148 7198 43150 7250
rect 43150 7198 43202 7250
rect 43202 7198 43204 7250
rect 43148 7196 43204 7198
rect 42812 6860 42868 6916
rect 43148 6300 43204 6356
rect 42588 4620 42644 4676
rect 42700 4956 42756 5012
rect 42028 4284 42084 4340
rect 42476 3948 42532 4004
rect 42476 3500 42532 3556
rect 41916 1820 41972 1876
rect 40796 1484 40852 1540
rect 40348 924 40404 980
rect 41916 1372 41972 1428
rect 40236 700 40292 756
rect 41692 140 41748 196
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 44156 12124 44212 12180
rect 44268 12066 44324 12068
rect 44268 12014 44270 12066
rect 44270 12014 44322 12066
rect 44322 12014 44324 12066
rect 44268 12012 44324 12014
rect 44940 12796 44996 12852
rect 45052 12236 45108 12292
rect 45052 12066 45108 12068
rect 45052 12014 45054 12066
rect 45054 12014 45106 12066
rect 45106 12014 45108 12066
rect 45052 12012 45108 12014
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44828 11788 44884 11844
rect 44672 11732 44728 11734
rect 45388 11228 45444 11284
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 44828 10668 44884 10724
rect 43596 10332 43652 10388
rect 44464 10218 44520 10220
rect 44156 10108 44212 10164
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 43708 7196 43764 7252
rect 43820 7084 43876 7140
rect 43820 6860 43876 6916
rect 43596 6300 43652 6356
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 43596 6076 43652 6132
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 43596 4508 43652 4564
rect 44828 10108 44884 10164
rect 44268 8876 44324 8932
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 44268 8092 44324 8148
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44268 5852 44324 5908
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 44268 4844 44324 4900
rect 44940 4508 44996 4564
rect 44464 3946 44520 3948
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 45388 10668 45444 10724
rect 45836 13580 45892 13636
rect 45500 9660 45556 9716
rect 45612 11452 45668 11508
rect 45276 8428 45332 8484
rect 45724 11282 45780 11284
rect 45724 11230 45726 11282
rect 45726 11230 45778 11282
rect 45778 11230 45780 11282
rect 45724 11228 45780 11230
rect 45724 9548 45780 9604
rect 45612 8316 45668 8372
rect 45388 7756 45444 7812
rect 45388 6748 45444 6804
rect 45948 13244 46004 13300
rect 45948 12460 46004 12516
rect 46060 11900 46116 11956
rect 46396 11228 46452 11284
rect 46620 10386 46676 10388
rect 46620 10334 46622 10386
rect 46622 10334 46674 10386
rect 46674 10334 46676 10386
rect 46620 10332 46676 10334
rect 46620 10108 46676 10164
rect 46060 9548 46116 9604
rect 46396 9548 46452 9604
rect 46060 9042 46116 9044
rect 46060 8990 46062 9042
rect 46062 8990 46114 9042
rect 46114 8990 46116 9042
rect 46060 8988 46116 8990
rect 45948 8428 46004 8484
rect 46396 8204 46452 8260
rect 45724 5292 45780 5348
rect 45500 3836 45556 3892
rect 43804 3162 43860 3164
rect 43372 2828 43428 2884
rect 43596 3052 43652 3108
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 43596 2828 43652 2884
rect 43932 2604 43988 2660
rect 43708 2268 43764 2324
rect 43708 1932 43764 1988
rect 44156 2604 44212 2660
rect 45052 2604 45108 2660
rect 44156 2380 44212 2436
rect 44464 2378 44520 2380
rect 44268 2268 44324 2324
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 44828 2268 44884 2324
rect 43932 1932 43988 1988
rect 43596 1596 43652 1652
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 42588 812 42644 868
rect 42476 364 42532 420
rect 41916 140 41972 196
rect 45724 2940 45780 2996
rect 46844 12962 46900 12964
rect 46844 12910 46846 12962
rect 46846 12910 46898 12962
rect 46898 12910 46900 12962
rect 46844 12908 46900 12910
rect 47180 12012 47236 12068
rect 46844 10780 46900 10836
rect 46844 10332 46900 10388
rect 47068 10386 47124 10388
rect 47068 10334 47070 10386
rect 47070 10334 47122 10386
rect 47122 10334 47124 10386
rect 47068 10332 47124 10334
rect 46956 10108 47012 10164
rect 46956 8540 47012 8596
rect 46956 7644 47012 7700
rect 46732 5964 46788 6020
rect 46396 4956 46452 5012
rect 46620 5180 46676 5236
rect 46732 4508 46788 4564
rect 47852 13356 47908 13412
rect 48188 13132 48244 13188
rect 48412 13074 48468 13076
rect 48412 13022 48414 13074
rect 48414 13022 48466 13074
rect 48466 13022 48468 13074
rect 48412 13020 48468 13022
rect 47964 12908 48020 12964
rect 49084 13580 49140 13636
rect 48972 13186 49028 13188
rect 48972 13134 48974 13186
rect 48974 13134 49026 13186
rect 49026 13134 49028 13186
rect 48972 13132 49028 13134
rect 48076 12236 48132 12292
rect 47740 11788 47796 11844
rect 47516 11282 47572 11284
rect 47516 11230 47518 11282
rect 47518 11230 47570 11282
rect 47570 11230 47572 11282
rect 47516 11228 47572 11230
rect 49420 12124 49476 12180
rect 48972 11506 49028 11508
rect 48972 11454 48974 11506
rect 48974 11454 49026 11506
rect 49026 11454 49028 11506
rect 48972 11452 49028 11454
rect 48524 11340 48580 11396
rect 48188 10556 48244 10612
rect 48748 11116 48804 11172
rect 48972 11004 49028 11060
rect 48300 10498 48356 10500
rect 48300 10446 48302 10498
rect 48302 10446 48354 10498
rect 48354 10446 48356 10498
rect 48300 10444 48356 10446
rect 48860 10332 48916 10388
rect 48188 9938 48244 9940
rect 48188 9886 48190 9938
rect 48190 9886 48242 9938
rect 48242 9886 48244 9938
rect 48188 9884 48244 9886
rect 48524 9938 48580 9940
rect 48524 9886 48526 9938
rect 48526 9886 48578 9938
rect 48578 9886 48580 9938
rect 48524 9884 48580 9886
rect 48524 8988 48580 9044
rect 47292 7868 47348 7924
rect 47964 8428 48020 8484
rect 47404 4732 47460 4788
rect 47068 2940 47124 2996
rect 46620 2828 46676 2884
rect 46284 2716 46340 2772
rect 46732 1372 46788 1428
rect 47068 1484 47124 1540
rect 45500 924 45556 980
rect 45724 924 45780 980
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 10780 28 10836 84
rect 48300 7756 48356 7812
rect 48076 6748 48132 6804
rect 48076 3164 48132 3220
rect 47964 2716 48020 2772
rect 47516 2156 47572 2212
rect 48748 7532 48804 7588
rect 48748 6524 48804 6580
rect 48636 6018 48692 6020
rect 48636 5966 48638 6018
rect 48638 5966 48690 6018
rect 48690 5966 48692 6018
rect 48636 5964 48692 5966
rect 49084 9996 49140 10052
rect 49532 11564 49588 11620
rect 49868 13244 49924 13300
rect 49644 11004 49700 11060
rect 49756 10108 49812 10164
rect 49420 9826 49476 9828
rect 49420 9774 49422 9826
rect 49422 9774 49474 9826
rect 49474 9774 49476 9826
rect 49420 9772 49476 9774
rect 49084 8540 49140 8596
rect 49420 8146 49476 8148
rect 49420 8094 49422 8146
rect 49422 8094 49474 8146
rect 49474 8094 49476 8146
rect 49420 8092 49476 8094
rect 49420 6972 49476 7028
rect 48972 5964 49028 6020
rect 49980 13020 50036 13076
rect 50428 12348 50484 12404
rect 50204 11900 50260 11956
rect 50428 11954 50484 11956
rect 50428 11902 50430 11954
rect 50430 11902 50482 11954
rect 50482 11902 50484 11954
rect 50428 11900 50484 11902
rect 50316 11618 50372 11620
rect 50316 11566 50318 11618
rect 50318 11566 50370 11618
rect 50370 11566 50372 11618
rect 50316 11564 50372 11566
rect 50540 10668 50596 10724
rect 49980 9884 50036 9940
rect 50204 10220 50260 10276
rect 49868 9772 49924 9828
rect 50428 9212 50484 9268
rect 49756 8092 49812 8148
rect 49644 7868 49700 7924
rect 50204 8930 50260 8932
rect 50204 8878 50206 8930
rect 50206 8878 50258 8930
rect 50258 8878 50260 8930
rect 50204 8876 50260 8878
rect 50316 8370 50372 8372
rect 50316 8318 50318 8370
rect 50318 8318 50370 8370
rect 50370 8318 50372 8370
rect 50316 8316 50372 8318
rect 50204 6690 50260 6692
rect 50204 6638 50206 6690
rect 50206 6638 50258 6690
rect 50258 6638 50260 6690
rect 50204 6636 50260 6638
rect 49532 5794 49588 5796
rect 49532 5742 49534 5794
rect 49534 5742 49586 5794
rect 49586 5742 49588 5794
rect 49532 5740 49588 5742
rect 51100 13580 51156 13636
rect 50876 11564 50932 11620
rect 50876 11116 50932 11172
rect 50764 9436 50820 9492
rect 50988 8764 51044 8820
rect 50988 8258 51044 8260
rect 50988 8206 50990 8258
rect 50990 8206 51042 8258
rect 51042 8206 51044 8258
rect 50988 8204 51044 8206
rect 50540 7474 50596 7476
rect 50540 7422 50542 7474
rect 50542 7422 50594 7474
rect 50594 7422 50596 7474
rect 50540 7420 50596 7422
rect 50652 6972 50708 7028
rect 50540 6690 50596 6692
rect 50540 6638 50542 6690
rect 50542 6638 50594 6690
rect 50594 6638 50596 6690
rect 50540 6636 50596 6638
rect 50540 6300 50596 6356
rect 50540 4844 50596 4900
rect 50316 3836 50372 3892
rect 50204 3276 50260 3332
rect 50428 3276 50484 3332
rect 52220 13132 52276 13188
rect 51772 12684 51828 12740
rect 51324 11676 51380 11732
rect 51996 12572 52052 12628
rect 51884 11618 51940 11620
rect 51884 11566 51886 11618
rect 51886 11566 51938 11618
rect 51938 11566 51940 11618
rect 51884 11564 51940 11566
rect 51324 10892 51380 10948
rect 51548 9772 51604 9828
rect 51212 9324 51268 9380
rect 51436 7362 51492 7364
rect 51436 7310 51438 7362
rect 51438 7310 51490 7362
rect 51490 7310 51492 7362
rect 51436 7308 51492 7310
rect 51100 6860 51156 6916
rect 51100 6690 51156 6692
rect 51100 6638 51102 6690
rect 51102 6638 51154 6690
rect 51154 6638 51156 6690
rect 51100 6636 51156 6638
rect 50652 4060 50708 4116
rect 48300 1932 48356 1988
rect 48748 1874 48804 1876
rect 48748 1822 48750 1874
rect 48750 1822 48802 1874
rect 48802 1822 48804 1874
rect 48748 1820 48804 1822
rect 49308 1820 49364 1876
rect 47628 1484 47684 1540
rect 47404 1372 47460 1428
rect 50652 1596 50708 1652
rect 50428 1314 50484 1316
rect 50428 1262 50430 1314
rect 50430 1262 50482 1314
rect 50482 1262 50484 1314
rect 50428 1260 50484 1262
rect 50764 1260 50820 1316
rect 50988 1202 51044 1204
rect 50988 1150 50990 1202
rect 50990 1150 51042 1202
rect 51042 1150 51044 1202
rect 50988 1148 51044 1150
rect 52108 10780 52164 10836
rect 51996 9602 52052 9604
rect 51996 9550 51998 9602
rect 51998 9550 52050 9602
rect 52050 9550 52052 9602
rect 51996 9548 52052 9550
rect 51884 9436 51940 9492
rect 52108 9100 52164 9156
rect 53116 13244 53172 13300
rect 52892 13074 52948 13076
rect 52892 13022 52894 13074
rect 52894 13022 52946 13074
rect 52946 13022 52948 13074
rect 52892 13020 52948 13022
rect 52556 12402 52612 12404
rect 52556 12350 52558 12402
rect 52558 12350 52610 12402
rect 52610 12350 52612 12402
rect 52556 12348 52612 12350
rect 52556 11676 52612 11732
rect 53788 13020 53844 13076
rect 52332 9996 52388 10052
rect 52556 8988 52612 9044
rect 52220 8316 52276 8372
rect 51996 6972 52052 7028
rect 52444 6860 52500 6916
rect 52556 6748 52612 6804
rect 51660 5122 51716 5124
rect 51660 5070 51662 5122
rect 51662 5070 51714 5122
rect 51714 5070 51716 5122
rect 51660 5068 51716 5070
rect 52108 5292 52164 5348
rect 51996 5122 52052 5124
rect 51996 5070 51998 5122
rect 51998 5070 52050 5122
rect 52050 5070 52052 5122
rect 51996 5068 52052 5070
rect 52332 4508 52388 4564
rect 52220 4396 52276 4452
rect 51884 3276 51940 3332
rect 51324 3164 51380 3220
rect 52108 2770 52164 2772
rect 52108 2718 52110 2770
rect 52110 2718 52162 2770
rect 52162 2718 52164 2770
rect 52108 2716 52164 2718
rect 51436 2044 51492 2100
rect 52220 2098 52276 2100
rect 52220 2046 52222 2098
rect 52222 2046 52274 2098
rect 52274 2046 52276 2098
rect 52220 2044 52276 2046
rect 51660 1596 51716 1652
rect 51100 924 51156 980
rect 51772 1372 51828 1428
rect 49532 588 49588 644
rect 49756 700 49812 756
rect 47740 364 47796 420
rect 52668 5852 52724 5908
rect 52668 4508 52724 4564
rect 53788 11004 53844 11060
rect 53788 10780 53844 10836
rect 53228 10444 53284 10500
rect 53116 9660 53172 9716
rect 53004 9266 53060 9268
rect 53004 9214 53006 9266
rect 53006 9214 53058 9266
rect 53058 9214 53060 9266
rect 53004 9212 53060 9214
rect 53004 7868 53060 7924
rect 52892 6636 52948 6692
rect 53004 6130 53060 6132
rect 53004 6078 53006 6130
rect 53006 6078 53058 6130
rect 53058 6078 53060 6130
rect 53004 6076 53060 6078
rect 53788 9548 53844 9604
rect 54124 12684 54180 12740
rect 54684 13468 54740 13524
rect 54236 11452 54292 11508
rect 54012 9212 54068 9268
rect 53340 8370 53396 8372
rect 53340 8318 53342 8370
rect 53342 8318 53394 8370
rect 53394 8318 53396 8370
rect 53340 8316 53396 8318
rect 53228 4226 53284 4228
rect 53228 4174 53230 4226
rect 53230 4174 53282 4226
rect 53282 4174 53284 4226
rect 53228 4172 53284 4174
rect 52780 3164 52836 3220
rect 52556 2828 52612 2884
rect 52780 2658 52836 2660
rect 52780 2606 52782 2658
rect 52782 2606 52834 2658
rect 52834 2606 52836 2658
rect 52780 2604 52836 2606
rect 53564 7196 53620 7252
rect 53564 6524 53620 6580
rect 54460 11394 54516 11396
rect 54460 11342 54462 11394
rect 54462 11342 54514 11394
rect 54514 11342 54516 11394
rect 54460 11340 54516 11342
rect 54348 11116 54404 11172
rect 54236 9324 54292 9380
rect 54124 8652 54180 8708
rect 54348 8540 54404 8596
rect 54908 13356 54964 13412
rect 54908 13186 54964 13188
rect 54908 13134 54910 13186
rect 54910 13134 54962 13186
rect 54962 13134 54964 13186
rect 54908 13132 54964 13134
rect 55356 12908 55412 12964
rect 55692 13244 55748 13300
rect 54684 10220 54740 10276
rect 54572 10108 54628 10164
rect 54124 7756 54180 7812
rect 54572 7196 54628 7252
rect 53900 6188 53956 6244
rect 54124 5628 54180 5684
rect 54572 5852 54628 5908
rect 54236 5180 54292 5236
rect 53564 4956 53620 5012
rect 53564 3724 53620 3780
rect 54572 4562 54628 4564
rect 54572 4510 54574 4562
rect 54574 4510 54626 4562
rect 54626 4510 54628 4562
rect 54572 4508 54628 4510
rect 53676 3612 53732 3668
rect 54124 3554 54180 3556
rect 54124 3502 54126 3554
rect 54126 3502 54178 3554
rect 54178 3502 54180 3554
rect 54124 3500 54180 3502
rect 53564 3442 53620 3444
rect 53564 3390 53566 3442
rect 53566 3390 53618 3442
rect 53618 3390 53620 3442
rect 53564 3388 53620 3390
rect 54572 3164 54628 3220
rect 53564 3052 53620 3108
rect 53452 2268 53508 2324
rect 54124 2492 54180 2548
rect 53564 1874 53620 1876
rect 53564 1822 53566 1874
rect 53566 1822 53618 1874
rect 53618 1822 53620 1874
rect 53564 1820 53620 1822
rect 53564 1426 53620 1428
rect 53564 1374 53566 1426
rect 53566 1374 53618 1426
rect 53618 1374 53620 1426
rect 53564 1372 53620 1374
rect 51996 924 52052 980
rect 53788 812 53844 868
rect 55356 11228 55412 11284
rect 55580 11228 55636 11284
rect 55468 10332 55524 10388
rect 55132 9436 55188 9492
rect 55020 8428 55076 8484
rect 56252 12460 56308 12516
rect 55804 10444 55860 10500
rect 56140 8988 56196 9044
rect 55580 8316 55636 8372
rect 55916 8092 55972 8148
rect 55132 7644 55188 7700
rect 56140 7698 56196 7700
rect 56140 7646 56142 7698
rect 56142 7646 56194 7698
rect 56194 7646 56196 7698
rect 56140 7644 56196 7646
rect 54908 7084 54964 7140
rect 56140 6748 56196 6804
rect 55132 6300 55188 6356
rect 57036 13916 57092 13972
rect 57036 11452 57092 11508
rect 57260 12124 57316 12180
rect 57260 7868 57316 7924
rect 56700 6076 56756 6132
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 55132 4844 55188 4900
rect 56140 5404 56196 5460
rect 55132 4338 55188 4340
rect 55132 4286 55134 4338
rect 55134 4286 55186 4338
rect 55186 4286 55188 4338
rect 55132 4284 55188 4286
rect 56140 4060 56196 4116
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 55132 2940 55188 2996
rect 56700 3388 56756 3444
rect 56140 2716 56196 2772
rect 54908 2268 54964 2324
rect 56476 2604 56532 2660
rect 55132 1090 55188 1092
rect 55132 1038 55134 1090
rect 55134 1038 55186 1090
rect 55186 1038 55188 1090
rect 55132 1036 55188 1038
rect 54796 700 54852 756
rect 56476 476 56532 532
rect 55804 140 55860 196
rect 47068 28 47124 84
rect 56700 28 56756 84
<< metal3 >>
rect 17042 14140 17052 14196
rect 17108 14140 30044 14196
rect 30100 14140 30110 14196
rect 12908 14028 24276 14084
rect 25330 14028 25340 14084
rect 25396 14028 25900 14084
rect 25956 14028 25966 14084
rect 26450 14028 26460 14084
rect 26516 14028 32508 14084
rect 32564 14028 32574 14084
rect 0 13972 112 14000
rect 12908 13972 12964 14028
rect 24220 13972 24276 14028
rect 57344 13972 57456 14000
rect 0 13916 476 13972
rect 532 13916 542 13972
rect 9762 13916 9772 13972
rect 9828 13916 11900 13972
rect 11956 13916 11966 13972
rect 12898 13916 12908 13972
rect 12964 13916 12974 13972
rect 20626 13916 20636 13972
rect 20692 13916 24164 13972
rect 24220 13916 26572 13972
rect 26628 13916 26638 13972
rect 26786 13916 26796 13972
rect 26852 13916 36092 13972
rect 36148 13916 36158 13972
rect 57026 13916 57036 13972
rect 57092 13916 57456 13972
rect 0 13888 112 13916
rect 24108 13860 24164 13916
rect 57344 13888 57456 13916
rect 14802 13804 14812 13860
rect 14868 13804 23884 13860
rect 23940 13804 23950 13860
rect 24108 13804 28028 13860
rect 28084 13804 28094 13860
rect 30034 13804 30044 13860
rect 30100 13804 30156 13860
rect 30212 13804 30222 13860
rect 30930 13804 30940 13860
rect 30996 13804 41020 13860
rect 41076 13804 41086 13860
rect 11890 13692 11900 13748
rect 11956 13692 25732 13748
rect 26674 13692 26684 13748
rect 26740 13692 27356 13748
rect 27412 13692 27422 13748
rect 35298 13692 35308 13748
rect 35364 13692 44156 13748
rect 44212 13692 44222 13748
rect 2258 13580 2268 13636
rect 2324 13580 3388 13636
rect 3444 13580 3454 13636
rect 14354 13580 14364 13636
rect 14420 13580 25228 13636
rect 25284 13580 25294 13636
rect 0 13524 112 13552
rect 25676 13524 25732 13692
rect 25890 13580 25900 13636
rect 25956 13580 31612 13636
rect 31668 13580 31678 13636
rect 38322 13580 38332 13636
rect 38388 13580 45836 13636
rect 45892 13580 45902 13636
rect 49074 13580 49084 13636
rect 49140 13580 51100 13636
rect 51156 13580 51166 13636
rect 57344 13524 57456 13552
rect 0 13468 140 13524
rect 196 13468 206 13524
rect 3602 13468 3612 13524
rect 3668 13468 4732 13524
rect 4788 13468 4798 13524
rect 23986 13468 23996 13524
rect 24052 13468 25452 13524
rect 25508 13468 25518 13524
rect 25676 13468 26796 13524
rect 26852 13468 26862 13524
rect 27682 13468 27692 13524
rect 27748 13468 40124 13524
rect 40180 13468 40190 13524
rect 54674 13468 54684 13524
rect 54740 13468 57456 13524
rect 0 13440 112 13468
rect 57344 13440 57456 13468
rect 13794 13356 13804 13412
rect 13860 13356 21868 13412
rect 21924 13356 21934 13412
rect 22092 13356 24388 13412
rect 25218 13356 25228 13412
rect 25284 13356 28924 13412
rect 28980 13356 28990 13412
rect 30818 13356 30828 13412
rect 30884 13356 42812 13412
rect 42868 13356 42878 13412
rect 47842 13356 47852 13412
rect 47908 13356 54908 13412
rect 54964 13356 54974 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 22092 13300 22148 13356
rect 2146 13244 2156 13300
rect 2212 13244 4284 13300
rect 4340 13244 4350 13300
rect 7522 13244 7532 13300
rect 7588 13244 9660 13300
rect 9716 13244 9726 13300
rect 13346 13244 13356 13300
rect 13412 13244 15036 13300
rect 15092 13244 15102 13300
rect 15810 13244 15820 13300
rect 15876 13244 22148 13300
rect 24332 13188 24388 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 24892 13244 25900 13300
rect 25956 13244 25966 13300
rect 26786 13244 26796 13300
rect 26852 13244 26862 13300
rect 35634 13244 35644 13300
rect 35700 13244 36988 13300
rect 37044 13244 37054 13300
rect 45938 13244 45948 13300
rect 46004 13244 49868 13300
rect 49924 13244 49934 13300
rect 53106 13244 53116 13300
rect 53172 13244 55692 13300
rect 55748 13244 55758 13300
rect 24892 13188 24948 13244
rect 26796 13188 26852 13244
rect 3714 13132 3724 13188
rect 3780 13132 5628 13188
rect 5684 13132 5694 13188
rect 5954 13132 5964 13188
rect 6020 13132 7420 13188
rect 7476 13132 7486 13188
rect 11330 13132 11340 13188
rect 11396 13132 13244 13188
rect 13300 13132 13310 13188
rect 17378 13132 17388 13188
rect 17444 13132 18620 13188
rect 18676 13132 18686 13188
rect 18946 13132 18956 13188
rect 19012 13132 19964 13188
rect 20020 13132 20030 13188
rect 22530 13132 22540 13188
rect 22596 13132 24108 13188
rect 24164 13132 24174 13188
rect 24332 13132 24948 13188
rect 25442 13132 25452 13188
rect 25508 13132 26852 13188
rect 28242 13132 28252 13188
rect 28308 13132 35644 13188
rect 35700 13132 35710 13188
rect 41794 13132 41804 13188
rect 41860 13132 42140 13188
rect 42196 13132 42588 13188
rect 42644 13132 43708 13188
rect 43764 13132 43774 13188
rect 48178 13132 48188 13188
rect 48244 13132 48972 13188
rect 49028 13132 49038 13188
rect 52210 13132 52220 13188
rect 52276 13132 54908 13188
rect 54964 13132 54974 13188
rect 0 13076 112 13104
rect 57344 13076 57456 13104
rect 0 13020 1484 13076
rect 1540 13020 1550 13076
rect 6066 13020 6076 13076
rect 6132 13020 6142 13076
rect 8194 13020 8204 13076
rect 8260 13020 10108 13076
rect 10164 13020 10174 13076
rect 14914 13020 14924 13076
rect 14980 13020 16828 13076
rect 16884 13020 16894 13076
rect 17154 13020 17164 13076
rect 17220 13020 35308 13076
rect 35364 13020 35374 13076
rect 36866 13020 36876 13076
rect 36932 13020 48412 13076
rect 48468 13020 48478 13076
rect 49970 13020 49980 13076
rect 50036 13020 52892 13076
rect 52948 13020 52958 13076
rect 53778 13020 53788 13076
rect 53844 13020 57456 13076
rect 0 12992 112 13020
rect 6076 12964 6132 13020
rect 57344 12992 57456 13020
rect 4274 12908 4284 12964
rect 4340 12908 5852 12964
rect 5908 12908 5918 12964
rect 6076 12908 6524 12964
rect 6580 12908 6590 12964
rect 16594 12908 16604 12964
rect 16660 12908 21420 12964
rect 21476 12908 21486 12964
rect 22194 12908 22204 12964
rect 22260 12908 38668 12964
rect 38770 12908 38780 12964
rect 38836 12908 42476 12964
rect 42532 12908 42542 12964
rect 43474 12908 43484 12964
rect 43540 12908 46844 12964
rect 46900 12908 46910 12964
rect 47954 12908 47964 12964
rect 48020 12908 55356 12964
rect 55412 12908 55422 12964
rect 38612 12852 38668 12908
rect 14466 12796 14476 12852
rect 14532 12796 20524 12852
rect 20580 12796 20590 12852
rect 20748 12796 31388 12852
rect 31444 12796 31724 12852
rect 31780 12796 31790 12852
rect 32274 12796 32284 12852
rect 32340 12796 36204 12852
rect 36260 12796 36270 12852
rect 38612 12796 40572 12852
rect 40628 12796 40638 12852
rect 40786 12796 40796 12852
rect 40852 12796 44940 12852
rect 44996 12796 45006 12852
rect 20748 12740 20804 12796
rect 9314 12684 9324 12740
rect 9380 12684 15596 12740
rect 15652 12684 15662 12740
rect 19282 12684 19292 12740
rect 19348 12684 20804 12740
rect 21298 12684 21308 12740
rect 21364 12684 21980 12740
rect 22036 12684 22046 12740
rect 22978 12684 22988 12740
rect 23044 12684 42252 12740
rect 42308 12684 42318 12740
rect 42476 12684 45500 12740
rect 45556 12684 45566 12740
rect 51762 12684 51772 12740
rect 51828 12684 54124 12740
rect 54180 12684 54190 12740
rect 0 12628 112 12656
rect 42476 12628 42532 12684
rect 57344 12628 57456 12656
rect 0 12572 364 12628
rect 420 12572 430 12628
rect 15250 12572 15260 12628
rect 15316 12572 20972 12628
rect 21028 12572 21038 12628
rect 24210 12572 24220 12628
rect 24276 12572 26236 12628
rect 26292 12572 26302 12628
rect 27458 12572 27468 12628
rect 27524 12572 41356 12628
rect 41412 12572 41422 12628
rect 42130 12572 42140 12628
rect 42196 12572 42532 12628
rect 51986 12572 51996 12628
rect 52052 12572 57456 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 57344 12544 57456 12572
rect 13458 12460 13468 12516
rect 13524 12460 16604 12516
rect 16660 12460 16670 12516
rect 16818 12460 16828 12516
rect 16884 12460 17556 12516
rect 20850 12460 20860 12516
rect 20916 12460 21868 12516
rect 21924 12460 21934 12516
rect 24210 12460 24220 12516
rect 24276 12460 25452 12516
rect 25508 12460 25518 12516
rect 25778 12460 25788 12516
rect 25844 12460 27244 12516
rect 27300 12460 27310 12516
rect 28690 12460 28700 12516
rect 28756 12460 30716 12516
rect 30772 12460 30782 12516
rect 32498 12460 32508 12516
rect 32564 12460 43260 12516
rect 43316 12460 43326 12516
rect 45938 12460 45948 12516
rect 46004 12460 56252 12516
rect 56308 12460 56318 12516
rect 17500 12404 17556 12460
rect 2818 12348 2828 12404
rect 2884 12348 3388 12404
rect 6962 12348 6972 12404
rect 7028 12348 8316 12404
rect 8372 12348 8382 12404
rect 10098 12348 10108 12404
rect 10164 12348 11004 12404
rect 11060 12348 11070 12404
rect 12002 12348 12012 12404
rect 12068 12348 12796 12404
rect 12852 12348 12862 12404
rect 14802 12348 14812 12404
rect 14868 12348 15932 12404
rect 15988 12348 15998 12404
rect 16370 12348 16380 12404
rect 16436 12348 17276 12404
rect 17332 12348 17342 12404
rect 17500 12348 21140 12404
rect 23090 12348 23100 12404
rect 23156 12348 23548 12404
rect 23604 12348 23614 12404
rect 23772 12348 30156 12404
rect 30212 12348 30222 12404
rect 36978 12348 36988 12404
rect 37044 12348 42364 12404
rect 42420 12348 42430 12404
rect 50418 12348 50428 12404
rect 50484 12348 52556 12404
rect 52612 12348 52622 12404
rect 3332 12292 3388 12348
rect 21084 12292 21140 12348
rect 23772 12292 23828 12348
rect 3332 12236 20860 12292
rect 20916 12236 20926 12292
rect 21084 12236 23828 12292
rect 23986 12236 23996 12292
rect 24052 12236 24444 12292
rect 24500 12236 24510 12292
rect 25442 12236 25452 12292
rect 25508 12236 27132 12292
rect 27188 12236 27198 12292
rect 29362 12236 29372 12292
rect 29428 12236 31052 12292
rect 31108 12236 32284 12292
rect 32340 12236 32350 12292
rect 35298 12236 35308 12292
rect 35364 12236 36316 12292
rect 36372 12236 37884 12292
rect 37940 12236 37950 12292
rect 38612 12236 39900 12292
rect 39956 12236 39966 12292
rect 40562 12236 40572 12292
rect 40628 12236 43260 12292
rect 43316 12236 43326 12292
rect 45042 12236 45052 12292
rect 45108 12236 48076 12292
rect 48132 12236 48142 12292
rect 0 12180 112 12208
rect 38612 12180 38668 12236
rect 57344 12180 57456 12208
rect 0 12124 588 12180
rect 644 12124 654 12180
rect 5058 12124 5068 12180
rect 5124 12124 11004 12180
rect 11060 12124 11070 12180
rect 11554 12124 11564 12180
rect 11620 12124 14084 12180
rect 14242 12124 14252 12180
rect 14308 12124 15148 12180
rect 15204 12124 15214 12180
rect 15362 12124 15372 12180
rect 15428 12124 18396 12180
rect 18452 12124 18462 12180
rect 20626 12124 20636 12180
rect 20692 12124 21420 12180
rect 21476 12124 28476 12180
rect 28532 12124 28542 12180
rect 29474 12124 29484 12180
rect 29540 12124 38668 12180
rect 41234 12124 41244 12180
rect 41300 12124 41804 12180
rect 41860 12124 41870 12180
rect 42018 12124 42028 12180
rect 42084 12124 42700 12180
rect 42756 12124 42766 12180
rect 44146 12124 44156 12180
rect 44212 12124 49420 12180
rect 49476 12124 49486 12180
rect 57250 12124 57260 12180
rect 57316 12124 57456 12180
rect 0 12096 112 12124
rect 14028 12068 14084 12124
rect 57344 12096 57456 12124
rect 1922 12012 1932 12068
rect 1988 12012 9436 12068
rect 9492 12012 9502 12068
rect 10658 12012 10668 12068
rect 10724 12012 13580 12068
rect 13636 12012 13646 12068
rect 14028 12012 15148 12068
rect 15092 11956 15148 12012
rect 16716 12012 19964 12068
rect 20020 12012 20030 12068
rect 20962 12012 20972 12068
rect 21028 12012 25676 12068
rect 25732 12012 25742 12068
rect 25890 12012 25900 12068
rect 25956 12012 27804 12068
rect 27860 12012 27870 12068
rect 34850 12012 34860 12068
rect 34916 12012 38668 12068
rect 40338 12012 40348 12068
rect 40404 12012 44268 12068
rect 44324 12012 44334 12068
rect 45042 12012 45052 12068
rect 45108 12012 47180 12068
rect 47236 12012 47246 12068
rect 16716 11956 16772 12012
rect 38612 11956 38668 12012
rect 8418 11900 8428 11956
rect 8484 11900 14252 11956
rect 14308 11900 14318 11956
rect 15092 11900 16772 11956
rect 18162 11900 18172 11956
rect 18228 11900 23548 11956
rect 23604 11900 23614 11956
rect 24546 11900 24556 11956
rect 24612 11900 25956 11956
rect 26338 11900 26348 11956
rect 26404 11900 29820 11956
rect 29876 11900 29886 11956
rect 35186 11900 35196 11956
rect 35252 11900 38500 11956
rect 38612 11900 42140 11956
rect 42196 11900 42206 11956
rect 42354 11900 42364 11956
rect 42420 11900 46060 11956
rect 46116 11900 46126 11956
rect 46386 11900 46396 11956
rect 46452 11900 50204 11956
rect 50260 11900 50428 11956
rect 50484 11900 50494 11956
rect 1138 11788 1148 11844
rect 1204 11788 2268 11844
rect 2324 11788 2334 11844
rect 5730 11788 5740 11844
rect 5796 11788 8596 11844
rect 10098 11788 10108 11844
rect 10164 11788 19348 11844
rect 19506 11788 19516 11844
rect 19572 11788 20636 11844
rect 20692 11788 20702 11844
rect 21186 11788 21196 11844
rect 21252 11788 23324 11844
rect 23380 11788 23390 11844
rect 24994 11788 25004 11844
rect 25060 11788 25340 11844
rect 25396 11788 25406 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 8540 11732 8596 11788
rect 19292 11732 19348 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 25900 11732 25956 11900
rect 38444 11844 38500 11900
rect 27570 11788 27580 11844
rect 27636 11788 29260 11844
rect 29316 11788 29326 11844
rect 31378 11788 31388 11844
rect 31444 11788 35868 11844
rect 35924 11788 35934 11844
rect 37314 11788 37324 11844
rect 37380 11788 38220 11844
rect 38276 11788 38286 11844
rect 38444 11788 42476 11844
rect 42532 11788 42542 11844
rect 44818 11788 44828 11844
rect 44884 11788 47740 11844
rect 47796 11788 47806 11844
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 57344 11732 57456 11760
rect 0 11676 3556 11732
rect 8540 11676 16940 11732
rect 16996 11676 17006 11732
rect 18246 11676 18284 11732
rect 18340 11676 18350 11732
rect 19292 11676 21084 11732
rect 21140 11676 21150 11732
rect 21298 11676 21308 11732
rect 21364 11676 24220 11732
rect 24276 11676 24286 11732
rect 25900 11676 28924 11732
rect 28980 11676 28990 11732
rect 32610 11676 32620 11732
rect 32676 11676 34132 11732
rect 34738 11676 34748 11732
rect 34804 11676 36764 11732
rect 36820 11676 36830 11732
rect 39890 11676 39900 11732
rect 39956 11676 42364 11732
rect 42420 11676 42430 11732
rect 51314 11676 51324 11732
rect 51380 11676 52556 11732
rect 52612 11676 52622 11732
rect 55412 11676 57456 11732
rect 0 11648 112 11676
rect 1474 11564 1484 11620
rect 1540 11564 2940 11620
rect 2996 11564 3006 11620
rect 3500 11396 3556 11676
rect 34076 11620 34132 11676
rect 55412 11620 55468 11676
rect 57344 11648 57456 11676
rect 4610 11564 4620 11620
rect 4676 11564 5180 11620
rect 5236 11564 5246 11620
rect 6178 11564 6188 11620
rect 6244 11564 6860 11620
rect 6916 11564 6926 11620
rect 7746 11564 7756 11620
rect 7812 11564 8764 11620
rect 8820 11564 8830 11620
rect 15698 11564 15708 11620
rect 15764 11564 21308 11620
rect 21364 11564 21374 11620
rect 23426 11564 23436 11620
rect 23492 11564 27468 11620
rect 27524 11564 27534 11620
rect 30482 11564 30492 11620
rect 30548 11564 33852 11620
rect 33908 11564 33918 11620
rect 34076 11564 41468 11620
rect 41524 11564 41534 11620
rect 49522 11564 49532 11620
rect 49588 11564 50316 11620
rect 50372 11564 50382 11620
rect 50866 11564 50876 11620
rect 50932 11564 51884 11620
rect 51940 11564 51950 11620
rect 52108 11564 55468 11620
rect 52108 11508 52164 11564
rect 15138 11452 15148 11508
rect 15204 11452 19516 11508
rect 19572 11452 19582 11508
rect 19954 11452 19964 11508
rect 20020 11452 25564 11508
rect 25620 11452 25630 11508
rect 25778 11452 25788 11508
rect 25844 11452 41916 11508
rect 41972 11452 41982 11508
rect 42466 11452 42476 11508
rect 42532 11452 45612 11508
rect 45668 11452 45678 11508
rect 48962 11452 48972 11508
rect 49028 11452 52164 11508
rect 54226 11452 54236 11508
rect 54292 11452 57036 11508
rect 57092 11452 57102 11508
rect 578 11340 588 11396
rect 644 11340 3388 11396
rect 3500 11340 14588 11396
rect 14644 11340 14654 11396
rect 18050 11340 18060 11396
rect 18116 11340 21756 11396
rect 21812 11340 21822 11396
rect 23538 11340 23548 11396
rect 23604 11340 26684 11396
rect 26740 11340 26750 11396
rect 27010 11340 27020 11396
rect 27076 11340 35196 11396
rect 35252 11340 35262 11396
rect 36530 11340 36540 11396
rect 36596 11340 37884 11396
rect 37940 11340 37950 11396
rect 38322 11340 38332 11396
rect 38388 11340 40572 11396
rect 40628 11340 40638 11396
rect 48514 11340 48524 11396
rect 48580 11340 54460 11396
rect 54516 11340 54526 11396
rect 0 11284 112 11312
rect 3332 11284 3388 11340
rect 57344 11284 57456 11312
rect 0 11228 252 11284
rect 308 11228 318 11284
rect 3332 11228 9324 11284
rect 9380 11228 9390 11284
rect 18386 11228 18396 11284
rect 18452 11228 22428 11284
rect 22484 11228 22494 11284
rect 23986 11228 23996 11284
rect 24052 11228 26460 11284
rect 26516 11228 26526 11284
rect 26684 11228 34300 11284
rect 34356 11228 34366 11284
rect 37986 11228 37996 11284
rect 38052 11228 45388 11284
rect 45444 11228 45454 11284
rect 45714 11228 45724 11284
rect 45780 11228 46396 11284
rect 46452 11228 46462 11284
rect 47506 11228 47516 11284
rect 47572 11228 55356 11284
rect 55412 11228 55422 11284
rect 55570 11228 55580 11284
rect 55636 11228 57456 11284
rect 0 11200 112 11228
rect 26684 11172 26740 11228
rect 57344 11200 57456 11228
rect 466 11116 476 11172
rect 532 11116 10108 11172
rect 10164 11116 10174 11172
rect 16146 11116 16156 11172
rect 16212 11116 18172 11172
rect 18228 11116 18238 11172
rect 20066 11116 20076 11172
rect 20132 11116 25060 11172
rect 26002 11116 26012 11172
rect 26068 11116 26740 11172
rect 27010 11116 27020 11172
rect 27076 11116 27972 11172
rect 28130 11116 28140 11172
rect 28196 11116 38220 11172
rect 38276 11116 38286 11172
rect 38994 11116 39004 11172
rect 39060 11116 48748 11172
rect 48804 11116 48814 11172
rect 50866 11116 50876 11172
rect 50932 11116 54348 11172
rect 54404 11116 54414 11172
rect 25004 11060 25060 11116
rect 27916 11060 27972 11116
rect 13570 11004 13580 11060
rect 13636 11004 22428 11060
rect 22484 11004 22494 11060
rect 24210 11004 24220 11060
rect 24276 11004 24556 11060
rect 24612 11004 24622 11060
rect 25004 11004 27692 11060
rect 27748 11004 27758 11060
rect 27916 11004 31836 11060
rect 31892 11004 31902 11060
rect 32162 11004 32172 11060
rect 32228 11004 33124 11060
rect 33618 11004 33628 11060
rect 33684 11004 34412 11060
rect 34468 11004 35308 11060
rect 35364 11004 35374 11060
rect 35522 11004 35532 11060
rect 35588 11004 38780 11060
rect 38836 11004 38846 11060
rect 39666 11004 39676 11060
rect 39732 11004 43148 11060
rect 43204 11004 43214 11060
rect 45948 11004 48972 11060
rect 49028 11004 49038 11060
rect 49634 11004 49644 11060
rect 49700 11004 53788 11060
rect 53844 11004 53854 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 9426 10892 9436 10948
rect 9492 10892 20076 10948
rect 20132 10892 20142 10948
rect 20402 10892 20412 10948
rect 20468 10892 21308 10948
rect 21364 10892 21374 10948
rect 24882 10892 24892 10948
rect 24948 10892 25676 10948
rect 25732 10892 25742 10948
rect 25890 10892 25900 10948
rect 25956 10892 26012 10948
rect 26068 10892 26078 10948
rect 26562 10892 26572 10948
rect 26628 10892 27020 10948
rect 27076 10892 27086 10948
rect 27234 10892 27244 10948
rect 27300 10892 29596 10948
rect 29652 10892 29662 10948
rect 29810 10892 29820 10948
rect 29876 10892 32844 10948
rect 32900 10892 32910 10948
rect 0 10836 112 10864
rect 33068 10836 33124 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 33282 10892 33292 10948
rect 33348 10892 35084 10948
rect 35140 10892 35150 10948
rect 35970 10892 35980 10948
rect 36036 10892 36540 10948
rect 36596 10892 36606 10948
rect 45948 10836 46004 11004
rect 46162 10892 46172 10948
rect 46228 10892 51324 10948
rect 51380 10892 51390 10948
rect 57344 10836 57456 10864
rect 0 10780 4956 10836
rect 5012 10780 5022 10836
rect 5282 10780 5292 10836
rect 5348 10780 19516 10836
rect 19572 10780 19582 10836
rect 20300 10780 32508 10836
rect 32564 10780 32574 10836
rect 33068 10780 46004 10836
rect 46834 10780 46844 10836
rect 46900 10780 52108 10836
rect 52164 10780 52174 10836
rect 53778 10780 53788 10836
rect 53844 10780 57456 10836
rect 0 10752 112 10780
rect 20300 10724 20356 10780
rect 57344 10752 57456 10780
rect 8978 10668 8988 10724
rect 9044 10668 18060 10724
rect 18116 10668 18126 10724
rect 18274 10668 18284 10724
rect 18340 10668 19180 10724
rect 19236 10668 19404 10724
rect 19460 10668 20356 10724
rect 21298 10668 21308 10724
rect 21364 10668 25004 10724
rect 25060 10668 25070 10724
rect 25218 10668 25228 10724
rect 25284 10668 28700 10724
rect 28756 10668 28766 10724
rect 30146 10668 30156 10724
rect 30212 10668 33516 10724
rect 33572 10668 33582 10724
rect 34850 10668 34860 10724
rect 34916 10668 37772 10724
rect 37828 10668 37838 10724
rect 40002 10668 40012 10724
rect 40068 10668 44828 10724
rect 44884 10668 44894 10724
rect 45378 10668 45388 10724
rect 45444 10668 50540 10724
rect 50596 10668 50606 10724
rect 3332 10556 10164 10612
rect 11330 10556 11340 10612
rect 11396 10556 11676 10612
rect 11732 10556 12572 10612
rect 12628 10556 12638 10612
rect 16594 10556 16604 10612
rect 16660 10556 19292 10612
rect 19348 10556 19358 10612
rect 20178 10556 20188 10612
rect 20244 10556 32788 10612
rect 34962 10556 34972 10612
rect 35028 10556 48188 10612
rect 48244 10556 48254 10612
rect 3266 10444 3276 10500
rect 3332 10444 3388 10556
rect 10108 10500 10164 10556
rect 32732 10500 32788 10556
rect 8866 10444 8876 10500
rect 8932 10444 9884 10500
rect 9940 10444 9950 10500
rect 10108 10444 11900 10500
rect 11956 10444 11966 10500
rect 12114 10444 12124 10500
rect 12180 10444 14252 10500
rect 14308 10444 14318 10500
rect 16482 10444 16492 10500
rect 16548 10444 17164 10500
rect 17220 10444 17230 10500
rect 18722 10444 18732 10500
rect 18788 10444 21084 10500
rect 21140 10444 21150 10500
rect 21410 10444 21420 10500
rect 21476 10444 25340 10500
rect 25396 10444 25406 10500
rect 25666 10444 25676 10500
rect 25732 10444 26572 10500
rect 26628 10444 27580 10500
rect 27636 10444 28364 10500
rect 28420 10444 28430 10500
rect 29362 10444 29372 10500
rect 29428 10444 30940 10500
rect 30996 10444 31006 10500
rect 32732 10444 48300 10500
rect 48356 10444 48366 10500
rect 53218 10444 53228 10500
rect 53284 10444 55804 10500
rect 55860 10444 55870 10500
rect 0 10388 112 10416
rect 57344 10388 57456 10416
rect 0 10332 1372 10388
rect 1428 10332 1438 10388
rect 4386 10332 4396 10388
rect 4452 10332 16548 10388
rect 20066 10332 20076 10388
rect 20132 10332 20524 10388
rect 20580 10332 20590 10388
rect 21858 10332 21868 10388
rect 21924 10332 37324 10388
rect 37380 10332 37390 10388
rect 37548 10332 40292 10388
rect 40450 10332 40460 10388
rect 40516 10332 42252 10388
rect 42308 10332 42318 10388
rect 43586 10332 43596 10388
rect 43652 10332 46620 10388
rect 46676 10332 46844 10388
rect 46900 10332 46910 10388
rect 47058 10332 47068 10388
rect 47124 10332 48860 10388
rect 48916 10332 48926 10388
rect 55458 10332 55468 10388
rect 55524 10332 57456 10388
rect 0 10304 112 10332
rect 7410 10220 7420 10276
rect 7476 10220 16436 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 11106 10108 11116 10164
rect 11172 10108 11900 10164
rect 11956 10108 11966 10164
rect 12338 10108 12348 10164
rect 12404 10108 13132 10164
rect 13188 10108 13198 10164
rect 13346 10108 13356 10164
rect 13412 10108 15820 10164
rect 15876 10108 15886 10164
rect 4946 9996 4956 10052
rect 5012 9996 8316 10052
rect 8372 9996 8382 10052
rect 10322 9996 10332 10052
rect 10388 9996 12908 10052
rect 12964 9996 12974 10052
rect 14242 9996 14252 10052
rect 14308 9996 16156 10052
rect 16212 9996 16222 10052
rect 0 9940 112 9968
rect 16380 9940 16436 10220
rect 16492 10052 16548 10332
rect 37548 10276 37604 10332
rect 40236 10276 40292 10332
rect 57344 10304 57456 10332
rect 18050 10220 18060 10276
rect 18116 10220 22204 10276
rect 22260 10220 22270 10276
rect 23314 10220 23324 10276
rect 23380 10220 24220 10276
rect 24276 10220 24286 10276
rect 26114 10220 26124 10276
rect 26180 10220 26236 10276
rect 26292 10220 26460 10276
rect 26516 10220 26526 10276
rect 26898 10220 26908 10276
rect 26964 10220 28364 10276
rect 28420 10220 28430 10276
rect 28578 10220 28588 10276
rect 28644 10220 29708 10276
rect 29764 10220 30044 10276
rect 30100 10220 30380 10276
rect 30436 10220 30446 10276
rect 31154 10220 31164 10276
rect 31220 10220 35756 10276
rect 35812 10220 35822 10276
rect 35970 10220 35980 10276
rect 36036 10220 37604 10276
rect 37762 10220 37772 10276
rect 37828 10220 40180 10276
rect 40236 10220 40908 10276
rect 40964 10220 40974 10276
rect 42354 10220 42364 10276
rect 42420 10220 43372 10276
rect 43428 10220 43438 10276
rect 50194 10220 50204 10276
rect 50260 10220 54684 10276
rect 54740 10220 54750 10276
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 40124 10164 40180 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 17826 10108 17836 10164
rect 17892 10108 19964 10164
rect 20020 10108 20030 10164
rect 20188 10108 22092 10164
rect 22148 10108 22158 10164
rect 25218 10108 25228 10164
rect 25284 10108 28476 10164
rect 28532 10108 28542 10164
rect 28700 10108 39228 10164
rect 39284 10108 39294 10164
rect 40124 10108 42252 10164
rect 42308 10108 42318 10164
rect 42466 10108 42476 10164
rect 42532 10108 44156 10164
rect 44212 10108 44222 10164
rect 44818 10108 44828 10164
rect 44884 10108 46620 10164
rect 46676 10108 46686 10164
rect 46946 10108 46956 10164
rect 47012 10108 49756 10164
rect 49812 10108 49822 10164
rect 54562 10108 54572 10164
rect 54628 10108 55468 10164
rect 20188 10052 20244 10108
rect 28700 10052 28756 10108
rect 16492 9996 18060 10052
rect 18116 9996 18126 10052
rect 18834 9996 18844 10052
rect 18900 9996 20244 10052
rect 21858 9996 21868 10052
rect 21924 9996 24220 10052
rect 24276 9996 24286 10052
rect 25330 9996 25340 10052
rect 25396 9996 28756 10052
rect 31266 9996 31276 10052
rect 31332 9996 39116 10052
rect 39172 9996 39182 10052
rect 39442 9996 39452 10052
rect 39508 9996 39900 10052
rect 39956 9996 40684 10052
rect 40740 9996 41580 10052
rect 41636 9996 41646 10052
rect 42130 9996 42140 10052
rect 42196 9996 42588 10052
rect 42644 9996 42654 10052
rect 44146 9996 44156 10052
rect 44212 9996 46060 10052
rect 46116 9996 46126 10052
rect 49074 9996 49084 10052
rect 49140 9996 52332 10052
rect 52388 9996 52398 10052
rect 55412 9940 55468 10108
rect 57344 9940 57456 9968
rect 0 9884 1036 9940
rect 1092 9884 1102 9940
rect 9538 9884 9548 9940
rect 9604 9884 16044 9940
rect 16100 9884 16110 9940
rect 16380 9884 21532 9940
rect 21588 9884 21598 9940
rect 22082 9884 22092 9940
rect 22148 9884 22316 9940
rect 22372 9884 22382 9940
rect 23202 9884 23212 9940
rect 23268 9884 23996 9940
rect 24052 9884 24444 9940
rect 24500 9884 25452 9940
rect 25508 9884 25518 9940
rect 26114 9884 26124 9940
rect 26180 9884 29932 9940
rect 29988 9884 29998 9940
rect 30146 9884 30156 9940
rect 30212 9884 48188 9940
rect 48244 9884 48524 9940
rect 48580 9884 48590 9940
rect 49970 9884 49980 9940
rect 50036 9884 52220 9940
rect 52276 9884 52286 9940
rect 55412 9884 57456 9940
rect 0 9856 112 9884
rect 57344 9856 57456 9884
rect 3332 9772 16716 9828
rect 16772 9772 16782 9828
rect 17378 9772 17388 9828
rect 17444 9772 18732 9828
rect 18788 9772 18798 9828
rect 20290 9772 20300 9828
rect 20356 9772 21084 9828
rect 21140 9772 24780 9828
rect 24836 9772 24846 9828
rect 25106 9772 25116 9828
rect 25172 9772 28252 9828
rect 28308 9772 28318 9828
rect 29250 9772 29260 9828
rect 29316 9772 34524 9828
rect 34580 9772 34590 9828
rect 38994 9772 39004 9828
rect 39060 9772 49420 9828
rect 49476 9772 49486 9828
rect 49858 9772 49868 9828
rect 49924 9772 51548 9828
rect 51604 9772 51614 9828
rect 3332 9716 3388 9772
rect 2706 9660 2716 9716
rect 2772 9660 3388 9716
rect 10210 9660 10220 9716
rect 10276 9660 11676 9716
rect 11732 9660 11742 9716
rect 13234 9660 13244 9716
rect 13300 9660 23100 9716
rect 23156 9660 23166 9716
rect 24546 9660 24556 9716
rect 24612 9660 26012 9716
rect 26068 9660 27580 9716
rect 27636 9660 27646 9716
rect 28354 9660 28364 9716
rect 28420 9660 30268 9716
rect 30324 9660 30334 9716
rect 30594 9660 30604 9716
rect 30660 9660 37324 9716
rect 37380 9660 37390 9716
rect 38210 9660 38220 9716
rect 38276 9660 44156 9716
rect 44212 9660 44222 9716
rect 45490 9660 45500 9716
rect 45556 9660 53116 9716
rect 53172 9660 53182 9716
rect 7298 9548 7308 9604
rect 7364 9548 11564 9604
rect 11620 9548 11630 9604
rect 16034 9548 16044 9604
rect 16100 9548 17500 9604
rect 17556 9548 19292 9604
rect 19348 9548 21308 9604
rect 21364 9548 21374 9604
rect 21746 9548 21756 9604
rect 21812 9548 25732 9604
rect 26198 9548 26236 9604
rect 26292 9548 27020 9604
rect 27076 9548 30940 9604
rect 30996 9548 31724 9604
rect 31780 9548 31790 9604
rect 32498 9548 32508 9604
rect 32564 9548 45724 9604
rect 45780 9548 45790 9604
rect 46050 9548 46060 9604
rect 46116 9548 46396 9604
rect 46452 9548 46462 9604
rect 51986 9548 51996 9604
rect 52052 9548 53788 9604
rect 53844 9548 53854 9604
rect 0 9492 112 9520
rect 0 9436 1932 9492
rect 1988 9436 1998 9492
rect 17714 9436 17724 9492
rect 17780 9436 18284 9492
rect 18340 9436 18956 9492
rect 19012 9436 19180 9492
rect 19236 9436 22876 9492
rect 22932 9436 22942 9492
rect 24210 9436 24220 9492
rect 24276 9436 24948 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 24892 9380 24948 9436
rect 14802 9324 14812 9380
rect 14868 9324 20860 9380
rect 20916 9324 20926 9380
rect 24882 9324 24892 9380
rect 24948 9324 24958 9380
rect 25676 9268 25732 9548
rect 46060 9492 46116 9548
rect 57344 9492 57456 9520
rect 27234 9436 27244 9492
rect 27300 9436 30716 9492
rect 30772 9436 30782 9492
rect 32274 9436 32284 9492
rect 32340 9436 40236 9492
rect 40292 9436 40302 9492
rect 45266 9436 45276 9492
rect 45332 9436 46116 9492
rect 50754 9436 50764 9492
rect 50820 9436 51884 9492
rect 51940 9436 51950 9492
rect 55122 9436 55132 9492
rect 55188 9436 57456 9492
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 57344 9408 57456 9436
rect 27346 9324 27356 9380
rect 27412 9324 28140 9380
rect 28196 9324 28206 9380
rect 28802 9324 28812 9380
rect 28868 9324 30380 9380
rect 30436 9324 30828 9380
rect 30884 9324 30894 9380
rect 31052 9324 33628 9380
rect 33684 9324 33694 9380
rect 34402 9324 34412 9380
rect 34468 9324 38388 9380
rect 38546 9324 38556 9380
rect 38612 9324 40908 9380
rect 40964 9324 40974 9380
rect 44258 9324 44268 9380
rect 44324 9324 46396 9380
rect 46452 9324 46462 9380
rect 51202 9324 51212 9380
rect 51268 9324 54236 9380
rect 54292 9324 54302 9380
rect 31052 9268 31108 9324
rect 38332 9268 38388 9324
rect 130 9212 140 9268
rect 196 9212 308 9268
rect 1586 9212 1596 9268
rect 1652 9212 15260 9268
rect 15316 9212 15326 9268
rect 15586 9212 15596 9268
rect 15652 9212 18284 9268
rect 18340 9212 18350 9268
rect 18834 9212 18844 9268
rect 18900 9212 21420 9268
rect 21476 9212 21486 9268
rect 21634 9212 21644 9268
rect 21700 9212 25004 9268
rect 25060 9212 25070 9268
rect 25218 9212 25228 9268
rect 25284 9212 25452 9268
rect 25508 9212 25518 9268
rect 25676 9212 29484 9268
rect 29540 9212 29550 9268
rect 30258 9212 30268 9268
rect 30324 9212 31108 9268
rect 31266 9212 31276 9268
rect 31332 9212 33068 9268
rect 33124 9212 33134 9268
rect 33506 9212 33516 9268
rect 33572 9212 38108 9268
rect 38164 9212 38174 9268
rect 38332 9212 42364 9268
rect 42420 9212 42430 9268
rect 43138 9212 43148 9268
rect 43204 9212 50428 9268
rect 50484 9212 50494 9268
rect 52994 9212 53004 9268
rect 53060 9212 54012 9268
rect 54068 9212 54078 9268
rect 252 9156 308 9212
rect 252 9100 10220 9156
rect 10276 9100 10286 9156
rect 10434 9100 10444 9156
rect 10500 9100 11788 9156
rect 11844 9100 11854 9156
rect 12898 9100 12908 9156
rect 12964 9100 14364 9156
rect 14420 9100 14430 9156
rect 20178 9100 20188 9156
rect 20244 9100 32844 9156
rect 32900 9100 32910 9156
rect 33618 9100 33628 9156
rect 33684 9100 37996 9156
rect 38052 9100 38062 9156
rect 38210 9100 38220 9156
rect 38276 9100 52108 9156
rect 52164 9100 52174 9156
rect 0 9044 112 9072
rect 57344 9044 57456 9072
rect 0 8988 3276 9044
rect 3332 8988 3342 9044
rect 12002 8988 12012 9044
rect 12068 8988 15484 9044
rect 15540 8988 15550 9044
rect 20290 8988 20300 9044
rect 20356 8988 21532 9044
rect 21588 8988 21598 9044
rect 21746 8988 21756 9044
rect 21812 8988 22316 9044
rect 22372 8988 25004 9044
rect 25060 8988 26572 9044
rect 26628 8988 26638 9044
rect 26786 8988 26796 9044
rect 26852 8988 29820 9044
rect 29876 8988 29886 9044
rect 30706 8988 30716 9044
rect 30772 8988 32284 9044
rect 32340 8988 33516 9044
rect 33572 8988 33582 9044
rect 33740 8988 36316 9044
rect 36372 8988 36382 9044
rect 36642 8988 36652 9044
rect 36708 8988 39452 9044
rect 39508 8988 39518 9044
rect 41122 8988 41132 9044
rect 41188 8988 43148 9044
rect 43204 8988 43214 9044
rect 43372 8988 45052 9044
rect 45108 8988 45118 9044
rect 46050 8988 46060 9044
rect 46116 8988 46172 9044
rect 46228 8988 46238 9044
rect 48514 8988 48524 9044
rect 48580 8988 52556 9044
rect 52612 8988 52622 9044
rect 56130 8988 56140 9044
rect 56196 8988 57456 9044
rect 0 8960 112 8988
rect 33740 8932 33796 8988
rect 43372 8932 43428 8988
rect 57344 8960 57456 8988
rect 4162 8876 4172 8932
rect 4228 8876 7476 8932
rect 7634 8876 7644 8932
rect 7700 8876 20524 8932
rect 20580 8876 20590 8932
rect 22418 8876 22428 8932
rect 22484 8876 24892 8932
rect 24948 8876 24958 8932
rect 25218 8876 25228 8932
rect 25284 8876 25452 8932
rect 25508 8876 25518 8932
rect 26114 8876 26124 8932
rect 26180 8876 31276 8932
rect 31332 8876 31342 8932
rect 31612 8876 33796 8932
rect 39666 8876 39676 8932
rect 39732 8876 41468 8932
rect 41524 8876 41534 8932
rect 43250 8876 43260 8932
rect 43316 8876 43428 8932
rect 44258 8876 44268 8932
rect 44324 8876 50204 8932
rect 50260 8876 50270 8932
rect 1698 8764 1708 8820
rect 1764 8764 4508 8820
rect 4564 8764 4956 8820
rect 5012 8764 5022 8820
rect 7420 8708 7476 8876
rect 31612 8820 31668 8876
rect 10210 8764 10220 8820
rect 10276 8764 16716 8820
rect 16772 8764 16782 8820
rect 19954 8764 19964 8820
rect 20020 8764 21980 8820
rect 22036 8764 22046 8820
rect 22194 8764 22204 8820
rect 22260 8764 31668 8820
rect 31724 8764 32508 8820
rect 32564 8764 32574 8820
rect 34962 8764 34972 8820
rect 35028 8764 40012 8820
rect 40068 8764 40684 8820
rect 40740 8764 40750 8820
rect 41990 8764 42028 8820
rect 42084 8764 42094 8820
rect 42252 8764 44884 8820
rect 45042 8764 45052 8820
rect 45108 8764 50988 8820
rect 51044 8764 51054 8820
rect 7420 8652 23548 8708
rect 23604 8652 23614 8708
rect 24882 8652 24892 8708
rect 24948 8652 28700 8708
rect 28756 8652 28766 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 31724 8596 31780 8764
rect 42252 8708 42308 8764
rect 32050 8652 32060 8708
rect 32116 8652 35980 8708
rect 36036 8652 36046 8708
rect 0 8540 3276 8596
rect 3332 8540 3342 8596
rect 14690 8540 14700 8596
rect 14756 8540 18620 8596
rect 18676 8540 18686 8596
rect 18956 8540 20468 8596
rect 24882 8540 24892 8596
rect 24948 8540 27020 8596
rect 27076 8540 31276 8596
rect 31332 8540 31342 8596
rect 31490 8540 31500 8596
rect 31556 8540 31780 8596
rect 32274 8540 32284 8596
rect 32340 8540 38444 8596
rect 38500 8540 38510 8596
rect 0 8512 112 8540
rect 18956 8484 19012 8540
rect 2594 8428 2604 8484
rect 2660 8428 9268 8484
rect 12114 8428 12124 8484
rect 12180 8428 12460 8484
rect 12516 8428 13020 8484
rect 13076 8428 14028 8484
rect 14084 8428 15148 8484
rect 16146 8428 16156 8484
rect 16212 8428 17836 8484
rect 17892 8428 17902 8484
rect 18274 8428 18284 8484
rect 18340 8428 19012 8484
rect 20178 8428 20188 8484
rect 20244 8428 20254 8484
rect 9212 8260 9268 8428
rect 15092 8372 15148 8428
rect 20188 8372 20244 8428
rect 11890 8316 11900 8372
rect 11956 8316 12908 8372
rect 12964 8316 13468 8372
rect 13524 8316 13534 8372
rect 13906 8316 13916 8372
rect 13972 8316 14364 8372
rect 14420 8316 14430 8372
rect 15092 8316 20244 8372
rect 20412 8372 20468 8540
rect 38612 8484 38668 8708
rect 38724 8652 38734 8708
rect 39106 8652 39116 8708
rect 39172 8652 42308 8708
rect 44828 8708 44884 8764
rect 44828 8652 54124 8708
rect 54180 8652 54190 8708
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 57344 8596 57456 8624
rect 39554 8540 39564 8596
rect 39620 8540 40572 8596
rect 40628 8540 40638 8596
rect 41122 8540 41132 8596
rect 41188 8540 44268 8596
rect 44324 8540 44334 8596
rect 46946 8540 46956 8596
rect 47012 8540 49084 8596
rect 49140 8540 49150 8596
rect 54338 8540 54348 8596
rect 54404 8540 57456 8596
rect 57344 8512 57456 8540
rect 21858 8428 21868 8484
rect 21924 8428 27244 8484
rect 27300 8428 27310 8484
rect 28476 8428 32956 8484
rect 33012 8428 33292 8484
rect 33348 8428 33516 8484
rect 33572 8428 33582 8484
rect 33842 8428 33852 8484
rect 33908 8428 38668 8484
rect 38994 8428 39004 8484
rect 39060 8428 42252 8484
rect 42308 8428 42318 8484
rect 43596 8428 45276 8484
rect 45332 8428 45342 8484
rect 45938 8428 45948 8484
rect 46004 8428 47964 8484
rect 48020 8428 48030 8484
rect 48188 8428 55020 8484
rect 55076 8428 55086 8484
rect 28476 8372 28532 8428
rect 43596 8372 43652 8428
rect 48188 8372 48244 8428
rect 20412 8316 21924 8372
rect 22754 8316 22764 8372
rect 22820 8316 28028 8372
rect 28084 8316 28094 8372
rect 28466 8316 28476 8372
rect 28532 8316 28542 8372
rect 35046 8316 35084 8372
rect 35140 8316 35150 8372
rect 35746 8316 35756 8372
rect 35812 8316 36876 8372
rect 36932 8316 36942 8372
rect 37436 8316 37996 8372
rect 38052 8316 38062 8372
rect 40114 8316 40124 8372
rect 40180 8316 40684 8372
rect 40740 8316 40750 8372
rect 41234 8316 41244 8372
rect 41300 8316 43652 8372
rect 45602 8316 45612 8372
rect 45668 8316 48244 8372
rect 50306 8316 50316 8372
rect 50372 8316 52220 8372
rect 52276 8316 52286 8372
rect 53330 8316 53340 8372
rect 53396 8316 55580 8372
rect 55636 8316 55646 8372
rect 21868 8260 21924 8316
rect 37436 8260 37492 8316
rect 6262 8204 6300 8260
rect 6356 8204 6366 8260
rect 9212 8204 15148 8260
rect 16706 8204 16716 8260
rect 16772 8204 21644 8260
rect 21700 8204 21710 8260
rect 21868 8204 23212 8260
rect 23268 8204 23278 8260
rect 23538 8204 23548 8260
rect 23604 8204 24220 8260
rect 24276 8204 24286 8260
rect 25218 8204 25228 8260
rect 25284 8204 32620 8260
rect 32676 8204 32686 8260
rect 33394 8204 33404 8260
rect 33460 8204 36428 8260
rect 36484 8204 37436 8260
rect 37492 8204 37502 8260
rect 37762 8204 37772 8260
rect 37828 8204 38556 8260
rect 38612 8204 38622 8260
rect 38770 8204 38780 8260
rect 38836 8204 43372 8260
rect 43428 8204 43438 8260
rect 46386 8204 46396 8260
rect 46452 8204 50988 8260
rect 51044 8204 51054 8260
rect 0 8148 112 8176
rect 15092 8148 15148 8204
rect 57344 8148 57456 8176
rect 0 8092 7420 8148
rect 7476 8092 7756 8148
rect 7812 8092 7822 8148
rect 9762 8092 9772 8148
rect 9828 8092 12348 8148
rect 12404 8092 12414 8148
rect 13132 8092 14700 8148
rect 14756 8092 14766 8148
rect 15092 8092 21868 8148
rect 21924 8092 21934 8148
rect 22082 8092 22092 8148
rect 22148 8092 26012 8148
rect 26068 8092 26078 8148
rect 26674 8092 26684 8148
rect 26740 8092 27020 8148
rect 27076 8092 27086 8148
rect 27356 8092 31164 8148
rect 31220 8092 31230 8148
rect 34066 8092 34076 8148
rect 34132 8092 44268 8148
rect 44324 8092 44334 8148
rect 49410 8092 49420 8148
rect 49476 8092 49756 8148
rect 49812 8092 49822 8148
rect 55906 8092 55916 8148
rect 55972 8092 57456 8148
rect 0 8064 112 8092
rect 13132 8036 13188 8092
rect 27356 8036 27412 8092
rect 57344 8064 57456 8092
rect 8418 7980 8428 8036
rect 8484 7980 9324 8036
rect 9380 7980 13188 8036
rect 13346 7980 13356 8036
rect 13412 7980 16604 8036
rect 16660 7980 16670 8036
rect 18498 7980 18508 8036
rect 18564 7980 19180 8036
rect 19236 7980 22652 8036
rect 22708 7980 22718 8036
rect 22866 7980 22876 8036
rect 22932 7980 24444 8036
rect 24500 7980 24510 8036
rect 24658 7980 24668 8036
rect 24724 7980 26460 8036
rect 26516 7980 26526 8036
rect 26898 7980 26908 8036
rect 26964 7980 27412 8036
rect 28578 7980 28588 8036
rect 28644 7980 30492 8036
rect 30548 7980 30558 8036
rect 34514 7980 34524 8036
rect 34580 7980 35420 8036
rect 35476 7980 37212 8036
rect 37268 7980 37772 8036
rect 37828 7980 37838 8036
rect 37986 7980 37996 8036
rect 38052 7980 39340 8036
rect 39396 7980 39406 8036
rect 40898 7980 40908 8036
rect 40964 7980 44828 8036
rect 44884 7980 44894 8036
rect 8306 7868 8316 7924
rect 8372 7868 16380 7924
rect 16436 7868 16446 7924
rect 16604 7868 23548 7924
rect 23604 7868 23614 7924
rect 24210 7868 24220 7924
rect 24276 7868 26684 7924
rect 26740 7868 26750 7924
rect 27682 7868 27692 7924
rect 27748 7868 27916 7924
rect 27972 7868 27982 7924
rect 29586 7868 29596 7924
rect 29652 7868 35868 7924
rect 35924 7868 35934 7924
rect 36082 7868 36092 7924
rect 36148 7868 38444 7924
rect 38500 7868 38780 7924
rect 38836 7868 38846 7924
rect 39218 7868 39228 7924
rect 39284 7868 40796 7924
rect 40852 7868 40862 7924
rect 41010 7868 41020 7924
rect 41076 7868 41692 7924
rect 41748 7868 42140 7924
rect 42196 7868 42206 7924
rect 44146 7868 44156 7924
rect 44212 7868 46844 7924
rect 46900 7868 46910 7924
rect 47282 7868 47292 7924
rect 47348 7868 49644 7924
rect 49700 7868 49710 7924
rect 52994 7868 53004 7924
rect 53060 7868 57260 7924
rect 57316 7868 57326 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 16604 7812 16660 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 12226 7756 12236 7812
rect 12292 7756 12796 7812
rect 12852 7756 12862 7812
rect 14018 7756 14028 7812
rect 14084 7756 14476 7812
rect 14532 7756 14542 7812
rect 14690 7756 14700 7812
rect 14756 7756 15820 7812
rect 15876 7756 15886 7812
rect 16034 7756 16044 7812
rect 16100 7756 16660 7812
rect 19618 7756 19628 7812
rect 19684 7756 20748 7812
rect 20804 7756 20814 7812
rect 20962 7756 20972 7812
rect 21028 7756 22204 7812
rect 22260 7756 22270 7812
rect 24220 7756 29596 7812
rect 29652 7756 29662 7812
rect 30146 7756 30156 7812
rect 30212 7756 33292 7812
rect 33348 7756 33358 7812
rect 35298 7756 35308 7812
rect 35364 7756 38332 7812
rect 38388 7756 38398 7812
rect 45378 7756 45388 7812
rect 45444 7756 47236 7812
rect 48290 7756 48300 7812
rect 48356 7756 54124 7812
rect 54180 7756 54190 7812
rect 0 7700 112 7728
rect 24220 7700 24276 7756
rect 47180 7700 47236 7756
rect 57344 7700 57456 7728
rect 0 7644 8876 7700
rect 8932 7644 8942 7700
rect 11330 7644 11340 7700
rect 11396 7644 18732 7700
rect 18788 7644 18798 7700
rect 19394 7644 19404 7700
rect 19460 7644 19796 7700
rect 20066 7644 20076 7700
rect 20132 7644 24276 7700
rect 24434 7644 24444 7700
rect 24500 7644 32620 7700
rect 32676 7644 32686 7700
rect 35186 7644 35196 7700
rect 35252 7644 35756 7700
rect 35812 7644 35822 7700
rect 35970 7644 35980 7700
rect 36036 7644 40124 7700
rect 40180 7644 40190 7700
rect 41906 7644 41916 7700
rect 41972 7644 46956 7700
rect 47012 7644 47022 7700
rect 47180 7644 55132 7700
rect 55188 7644 55198 7700
rect 56130 7644 56140 7700
rect 56196 7644 57456 7700
rect 0 7616 112 7644
rect 19740 7588 19796 7644
rect 57344 7616 57456 7644
rect 1474 7532 1484 7588
rect 1540 7532 7980 7588
rect 8036 7532 8046 7588
rect 12114 7532 12124 7588
rect 12180 7532 15148 7588
rect 15810 7532 15820 7588
rect 15876 7532 16156 7588
rect 16212 7532 16222 7588
rect 18274 7532 18284 7588
rect 18340 7532 19516 7588
rect 19572 7532 19582 7588
rect 19740 7532 20636 7588
rect 20692 7532 20702 7588
rect 20850 7532 20860 7588
rect 20916 7532 27132 7588
rect 27188 7532 27198 7588
rect 28018 7532 28028 7588
rect 28084 7532 32060 7588
rect 32116 7532 32126 7588
rect 34290 7532 34300 7588
rect 34356 7532 34972 7588
rect 35028 7532 35644 7588
rect 35700 7532 36316 7588
rect 36372 7532 37100 7588
rect 37156 7532 37166 7588
rect 37314 7532 37324 7588
rect 37380 7532 48748 7588
rect 48804 7532 48814 7588
rect 15092 7476 15148 7532
rect 1026 7420 1036 7476
rect 1092 7420 3388 7476
rect 6850 7420 6860 7476
rect 6916 7420 12796 7476
rect 12852 7420 12862 7476
rect 13122 7420 13132 7476
rect 13188 7420 13580 7476
rect 13636 7420 14476 7476
rect 14532 7420 14700 7476
rect 14756 7420 14766 7476
rect 15092 7420 23996 7476
rect 24052 7420 24062 7476
rect 25778 7420 25788 7476
rect 25844 7420 28812 7476
rect 28868 7420 28878 7476
rect 29036 7420 32172 7476
rect 32228 7420 32238 7476
rect 32610 7420 32620 7476
rect 32676 7420 50540 7476
rect 50596 7420 50606 7476
rect 3332 7364 3388 7420
rect 29036 7364 29092 7420
rect 3332 7308 7308 7364
rect 7364 7308 7374 7364
rect 7746 7308 7756 7364
rect 7812 7308 8652 7364
rect 8708 7308 8718 7364
rect 8876 7308 15372 7364
rect 15428 7308 15438 7364
rect 17714 7308 17724 7364
rect 17780 7308 18284 7364
rect 18340 7308 18350 7364
rect 19282 7308 19292 7364
rect 19348 7308 19740 7364
rect 19796 7308 19806 7364
rect 19954 7308 19964 7364
rect 20020 7308 29092 7364
rect 29250 7308 29260 7364
rect 29316 7308 30492 7364
rect 30548 7308 30558 7364
rect 31602 7308 31612 7364
rect 31668 7308 35644 7364
rect 35700 7308 35710 7364
rect 35858 7308 35868 7364
rect 35924 7308 36316 7364
rect 36372 7308 36382 7364
rect 36642 7308 36652 7364
rect 36708 7308 41804 7364
rect 41860 7308 41870 7364
rect 42242 7308 42252 7364
rect 42308 7308 44940 7364
rect 44996 7308 45006 7364
rect 45378 7308 45388 7364
rect 45444 7308 51436 7364
rect 51492 7308 51502 7364
rect 0 7252 112 7280
rect 0 7196 1596 7252
rect 1652 7196 1662 7252
rect 2930 7196 2940 7252
rect 2996 7196 5236 7252
rect 0 7168 112 7196
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 5180 7028 5236 7196
rect 8876 7140 8932 7308
rect 57344 7252 57456 7280
rect 9874 7196 9884 7252
rect 9940 7196 10556 7252
rect 10612 7196 12124 7252
rect 12180 7196 13916 7252
rect 13972 7196 13982 7252
rect 14354 7196 14364 7252
rect 14420 7196 14430 7252
rect 14578 7196 14588 7252
rect 14644 7196 21644 7252
rect 21700 7196 21710 7252
rect 21858 7196 21868 7252
rect 21924 7196 30156 7252
rect 30212 7196 30222 7252
rect 31826 7196 31836 7252
rect 31892 7196 33068 7252
rect 33124 7196 33134 7252
rect 36082 7196 36092 7252
rect 36148 7196 36428 7252
rect 36484 7196 36494 7252
rect 37538 7196 37548 7252
rect 37604 7196 41916 7252
rect 41972 7196 41982 7252
rect 42242 7196 42252 7252
rect 42308 7196 42700 7252
rect 42756 7196 43148 7252
rect 43204 7196 43708 7252
rect 43764 7196 43774 7252
rect 44268 7196 53564 7252
rect 53620 7196 53630 7252
rect 54562 7196 54572 7252
rect 54628 7196 57456 7252
rect 14364 7140 14420 7196
rect 6066 7084 6076 7140
rect 6132 7084 8932 7140
rect 12674 7084 12684 7140
rect 12740 7084 13132 7140
rect 13188 7084 13198 7140
rect 14364 7084 15148 7140
rect 15204 7084 21420 7140
rect 21476 7084 21486 7140
rect 22194 7084 22204 7140
rect 22260 7084 24332 7140
rect 24388 7084 24398 7140
rect 24994 7084 25004 7140
rect 25060 7084 25452 7140
rect 25508 7084 25518 7140
rect 26450 7084 26460 7140
rect 26516 7084 32732 7140
rect 32788 7084 32798 7140
rect 36978 7084 36988 7140
rect 37044 7084 40348 7140
rect 40404 7084 40414 7140
rect 40674 7084 40684 7140
rect 40740 7084 43820 7140
rect 43876 7084 43886 7140
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 44268 7028 44324 7196
rect 57344 7168 57456 7196
rect 44818 7084 44828 7140
rect 44884 7084 54908 7140
rect 54964 7084 54974 7140
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 5180 6972 15148 7028
rect 15250 6972 15260 7028
rect 15316 6972 20916 7028
rect 21634 6972 21644 7028
rect 21700 6972 24220 7028
rect 24276 6972 24286 7028
rect 24892 6972 28476 7028
rect 28532 6972 28542 7028
rect 31378 6972 31388 7028
rect 31444 6972 44324 7028
rect 44828 6972 49420 7028
rect 49476 6972 49486 7028
rect 50642 6972 50652 7028
rect 50708 6972 51996 7028
rect 52052 6972 52062 7028
rect 15092 6916 15148 6972
rect 20860 6916 20916 6972
rect 24892 6916 24948 6972
rect 44828 6916 44884 6972
rect 1922 6860 1932 6916
rect 1988 6860 10108 6916
rect 10164 6860 10174 6916
rect 15092 6860 20076 6916
rect 20132 6860 20142 6916
rect 20850 6860 20860 6916
rect 20916 6860 20926 6916
rect 21186 6860 21196 6916
rect 21252 6860 24948 6916
rect 25106 6860 25116 6916
rect 25172 6860 28028 6916
rect 28084 6860 28094 6916
rect 28242 6860 28252 6916
rect 28308 6860 30044 6916
rect 30100 6860 30110 6916
rect 33058 6860 33068 6916
rect 33124 6860 34860 6916
rect 34916 6860 34926 6916
rect 38658 6860 38668 6916
rect 38724 6860 41132 6916
rect 41188 6860 41198 6916
rect 41346 6860 41356 6916
rect 41412 6860 42812 6916
rect 42868 6860 42878 6916
rect 43810 6860 43820 6916
rect 43876 6860 44884 6916
rect 45164 6860 46452 6916
rect 51090 6860 51100 6916
rect 51156 6860 52444 6916
rect 52500 6860 52510 6916
rect 0 6804 112 6832
rect 45164 6804 45220 6860
rect 0 6748 6860 6804
rect 6916 6748 6926 6804
rect 7084 6748 12068 6804
rect 13010 6748 13020 6804
rect 13076 6748 13356 6804
rect 13412 6748 13422 6804
rect 16370 6748 16380 6804
rect 16436 6748 17332 6804
rect 17714 6748 17724 6804
rect 17780 6748 23884 6804
rect 23940 6748 23950 6804
rect 24322 6748 24332 6804
rect 24388 6748 25228 6804
rect 25284 6748 25294 6804
rect 25442 6748 25452 6804
rect 25508 6748 26684 6804
rect 26740 6748 26750 6804
rect 26852 6748 28364 6804
rect 28420 6748 28430 6804
rect 28578 6748 28588 6804
rect 28644 6748 28924 6804
rect 28980 6748 28990 6804
rect 30268 6748 35476 6804
rect 0 6720 112 6748
rect 7084 6580 7140 6748
rect 12012 6692 12068 6748
rect 11106 6636 11116 6692
rect 11172 6636 11788 6692
rect 11844 6636 11854 6692
rect 12012 6636 17052 6692
rect 17108 6636 17118 6692
rect 17276 6580 17332 6748
rect 26852 6692 26908 6748
rect 30268 6692 30324 6748
rect 18386 6636 18396 6692
rect 18452 6636 18844 6692
rect 18900 6636 18910 6692
rect 20514 6636 20524 6692
rect 20580 6636 26908 6692
rect 27010 6636 27020 6692
rect 27076 6636 28252 6692
rect 28308 6636 28318 6692
rect 28466 6636 28476 6692
rect 28532 6636 30324 6692
rect 31714 6636 31724 6692
rect 31780 6636 32284 6692
rect 32340 6636 32956 6692
rect 33012 6636 33022 6692
rect 35420 6580 35476 6748
rect 37548 6748 40684 6804
rect 40740 6748 42028 6804
rect 42084 6748 42094 6804
rect 42354 6748 42364 6804
rect 42420 6748 45220 6804
rect 45378 6748 45388 6804
rect 45444 6748 45454 6804
rect 37548 6692 37604 6748
rect 45388 6692 45444 6748
rect 36754 6636 36764 6692
rect 36820 6636 37604 6692
rect 37762 6636 37772 6692
rect 37828 6636 39452 6692
rect 39508 6636 39518 6692
rect 40226 6636 40236 6692
rect 40292 6636 41468 6692
rect 41524 6636 41534 6692
rect 41682 6636 41692 6692
rect 41748 6636 45444 6692
rect 46396 6692 46452 6860
rect 57344 6804 57456 6832
rect 48066 6748 48076 6804
rect 48132 6748 52556 6804
rect 52612 6748 52622 6804
rect 56130 6748 56140 6804
rect 56196 6748 57456 6804
rect 57344 6720 57456 6748
rect 46396 6636 50204 6692
rect 50260 6636 50540 6692
rect 50596 6636 50606 6692
rect 51090 6636 51100 6692
rect 51156 6636 52892 6692
rect 52948 6636 52958 6692
rect 1138 6524 1148 6580
rect 1204 6524 7140 6580
rect 7970 6524 7980 6580
rect 8036 6524 16492 6580
rect 16548 6524 16558 6580
rect 17276 6524 21868 6580
rect 21924 6524 21934 6580
rect 22642 6524 22652 6580
rect 22708 6524 26236 6580
rect 26292 6524 26302 6580
rect 26450 6524 26460 6580
rect 26516 6524 33628 6580
rect 33684 6524 33694 6580
rect 35420 6524 45388 6580
rect 45444 6524 45454 6580
rect 48738 6524 48748 6580
rect 48804 6524 53564 6580
rect 53620 6524 53630 6580
rect 242 6412 252 6468
rect 308 6412 15596 6468
rect 15652 6412 16268 6468
rect 16324 6412 16334 6468
rect 16706 6412 16716 6468
rect 16772 6412 28476 6468
rect 28532 6412 28542 6468
rect 28690 6412 28700 6468
rect 28756 6412 32676 6468
rect 32946 6412 32956 6468
rect 33012 6412 46956 6468
rect 47012 6412 47022 6468
rect 0 6356 112 6384
rect 0 6300 1036 6356
rect 1092 6300 1102 6356
rect 14130 6300 14140 6356
rect 14196 6300 23660 6356
rect 23716 6300 23726 6356
rect 24210 6300 24220 6356
rect 24276 6300 32396 6356
rect 32452 6300 32462 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 32620 6244 32676 6412
rect 57344 6356 57456 6384
rect 32834 6300 32844 6356
rect 32900 6300 33964 6356
rect 34020 6300 34030 6356
rect 35746 6300 35756 6356
rect 35812 6300 37772 6356
rect 37828 6300 37838 6356
rect 37986 6300 37996 6356
rect 38052 6300 40460 6356
rect 40516 6300 41468 6356
rect 41524 6300 42252 6356
rect 42308 6300 43148 6356
rect 43204 6300 43214 6356
rect 43586 6300 43596 6356
rect 43652 6300 43662 6356
rect 47068 6300 50540 6356
rect 50596 6300 50606 6356
rect 55122 6300 55132 6356
rect 55188 6300 57456 6356
rect 43596 6244 43652 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 47068 6244 47124 6300
rect 57344 6272 57456 6300
rect 7858 6188 7868 6244
rect 7924 6188 8316 6244
rect 8372 6188 9324 6244
rect 9380 6188 9390 6244
rect 11778 6188 11788 6244
rect 11844 6188 16716 6244
rect 16772 6188 16782 6244
rect 18284 6188 19404 6244
rect 19460 6188 19470 6244
rect 20738 6188 20748 6244
rect 20804 6188 21308 6244
rect 21364 6188 21644 6244
rect 21700 6188 21710 6244
rect 23202 6188 23212 6244
rect 23268 6188 23548 6244
rect 23604 6188 23614 6244
rect 24210 6188 24220 6244
rect 24276 6188 27188 6244
rect 27458 6188 27468 6244
rect 27524 6188 31948 6244
rect 32004 6188 32014 6244
rect 32620 6188 38556 6244
rect 38612 6188 38622 6244
rect 39778 6188 39788 6244
rect 39844 6188 43652 6244
rect 45490 6188 45500 6244
rect 45556 6188 47124 6244
rect 50372 6188 53900 6244
rect 53956 6188 53966 6244
rect 18284 6132 18340 6188
rect 27132 6132 27188 6188
rect 50372 6132 50428 6188
rect 6514 6076 6524 6132
rect 6580 6076 12012 6132
rect 12068 6076 12078 6132
rect 12450 6076 12460 6132
rect 12516 6076 15932 6132
rect 15988 6076 18340 6132
rect 18498 6076 18508 6132
rect 18564 6076 26796 6132
rect 26852 6076 26862 6132
rect 27132 6076 31612 6132
rect 31668 6076 31678 6132
rect 31826 6076 31836 6132
rect 31892 6076 32620 6132
rect 32676 6076 32686 6132
rect 32844 6076 32956 6132
rect 33012 6076 33022 6132
rect 33618 6076 33628 6132
rect 33684 6076 43596 6132
rect 43652 6076 43662 6132
rect 44044 6076 50428 6132
rect 52994 6076 53004 6132
rect 53060 6076 56700 6132
rect 56756 6076 56766 6132
rect 32844 6020 32900 6076
rect 1362 5964 1372 6020
rect 1428 5964 6412 6020
rect 6468 5964 6748 6020
rect 6804 5964 7420 6020
rect 7476 5964 8316 6020
rect 8372 5964 8382 6020
rect 8988 5964 16044 6020
rect 16100 5964 16110 6020
rect 17602 5964 17612 6020
rect 17668 5964 21756 6020
rect 21812 5964 21822 6020
rect 22166 5964 22204 6020
rect 22260 5964 22270 6020
rect 22418 5964 22428 6020
rect 22484 5964 26460 6020
rect 26516 5964 26526 6020
rect 26674 5964 26684 6020
rect 26740 5964 32900 6020
rect 33058 5964 33068 6020
rect 33124 5964 35140 6020
rect 40114 5964 40124 6020
rect 40180 5964 41804 6020
rect 41860 5964 41870 6020
rect 0 5908 112 5936
rect 8988 5908 9044 5964
rect 0 5852 1148 5908
rect 1204 5852 1214 5908
rect 6962 5852 6972 5908
rect 7028 5852 9044 5908
rect 14242 5852 14252 5908
rect 14308 5852 15708 5908
rect 15764 5852 16268 5908
rect 16324 5852 16334 5908
rect 19394 5852 19404 5908
rect 19460 5852 26012 5908
rect 26068 5852 26078 5908
rect 26226 5852 26236 5908
rect 26292 5852 26572 5908
rect 26628 5852 27356 5908
rect 27412 5852 27580 5908
rect 27636 5852 27646 5908
rect 27804 5852 29148 5908
rect 29204 5852 29214 5908
rect 29810 5852 29820 5908
rect 29876 5852 30268 5908
rect 30324 5852 32396 5908
rect 32452 5852 32462 5908
rect 32610 5852 32620 5908
rect 32676 5852 34860 5908
rect 34916 5852 34926 5908
rect 0 5824 112 5852
rect 27804 5796 27860 5852
rect 35084 5796 35140 5964
rect 44044 5908 44100 6076
rect 46722 5964 46732 6020
rect 46788 5964 48636 6020
rect 48692 5964 48972 6020
rect 49028 5964 49038 6020
rect 57344 5908 57456 5936
rect 38434 5852 38444 5908
rect 38500 5852 39228 5908
rect 39284 5852 39294 5908
rect 40562 5852 40572 5908
rect 40628 5852 44100 5908
rect 44258 5852 44268 5908
rect 44324 5852 52668 5908
rect 52724 5852 52734 5908
rect 54562 5852 54572 5908
rect 54628 5852 57456 5908
rect 57344 5824 57456 5852
rect 2818 5740 2828 5796
rect 2884 5740 3388 5796
rect 14578 5740 14588 5796
rect 14644 5740 25676 5796
rect 25732 5740 25742 5796
rect 26338 5740 26348 5796
rect 26404 5740 27132 5796
rect 27188 5740 27860 5796
rect 27916 5740 28252 5796
rect 28308 5740 29036 5796
rect 29092 5740 29260 5796
rect 29316 5740 29326 5796
rect 29698 5740 29708 5796
rect 29764 5740 31892 5796
rect 32050 5740 32060 5796
rect 32116 5740 33180 5796
rect 33236 5740 33246 5796
rect 35084 5740 38668 5796
rect 38724 5740 38734 5796
rect 40674 5740 40684 5796
rect 40740 5740 49532 5796
rect 49588 5740 49598 5796
rect 3332 5684 3388 5740
rect 27916 5684 27972 5740
rect 3332 5628 15148 5684
rect 16930 5628 16940 5684
rect 16996 5628 21028 5684
rect 21410 5628 21420 5684
rect 21476 5628 21486 5684
rect 21746 5628 21756 5684
rect 21812 5628 22540 5684
rect 22596 5628 22606 5684
rect 23426 5628 23436 5684
rect 23492 5628 26572 5684
rect 26628 5628 26638 5684
rect 26786 5628 26796 5684
rect 26852 5628 27468 5684
rect 27524 5628 27534 5684
rect 27682 5628 27692 5684
rect 27748 5628 27972 5684
rect 28130 5628 28140 5684
rect 28196 5628 28364 5684
rect 28420 5628 28430 5684
rect 28802 5628 28812 5684
rect 28868 5628 29932 5684
rect 29988 5628 30716 5684
rect 30772 5628 30782 5684
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 15092 5460 15148 5628
rect 16034 5516 16044 5572
rect 16100 5516 20636 5572
rect 20692 5516 20702 5572
rect 20972 5460 21028 5628
rect 21420 5572 21476 5628
rect 31836 5572 31892 5740
rect 32722 5628 32732 5684
rect 32788 5628 54124 5684
rect 54180 5628 54190 5684
rect 21420 5516 23324 5572
rect 23380 5516 23390 5572
rect 23650 5516 23660 5572
rect 23716 5516 24332 5572
rect 24388 5516 24398 5572
rect 25666 5516 25676 5572
rect 25732 5516 26124 5572
rect 26180 5516 30380 5572
rect 30436 5516 30446 5572
rect 31798 5516 31836 5572
rect 31892 5516 32060 5572
rect 32116 5516 33628 5572
rect 33684 5516 33694 5572
rect 34178 5516 34188 5572
rect 34244 5516 35644 5572
rect 35700 5516 35710 5572
rect 35970 5516 35980 5572
rect 36036 5516 37436 5572
rect 37492 5516 37502 5572
rect 38658 5516 38668 5572
rect 38724 5516 41972 5572
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 0 5404 3388 5460
rect 15092 5404 20748 5460
rect 20804 5404 20814 5460
rect 20972 5404 24220 5460
rect 24276 5404 24286 5460
rect 27020 5404 31388 5460
rect 31444 5404 31454 5460
rect 31938 5404 31948 5460
rect 32004 5404 41692 5460
rect 41748 5404 41758 5460
rect 0 5376 112 5404
rect 3332 5348 3388 5404
rect 27020 5348 27076 5404
rect 3332 5292 9772 5348
rect 9828 5292 9838 5348
rect 15474 5292 15484 5348
rect 15540 5292 16044 5348
rect 16100 5292 16110 5348
rect 16594 5292 16604 5348
rect 16660 5292 20748 5348
rect 20804 5292 20814 5348
rect 20962 5292 20972 5348
rect 21028 5292 22652 5348
rect 22708 5292 22718 5348
rect 23986 5292 23996 5348
rect 24052 5292 25956 5348
rect 26226 5292 26236 5348
rect 26292 5292 27076 5348
rect 27234 5292 27244 5348
rect 27300 5292 31276 5348
rect 31332 5292 31342 5348
rect 31490 5292 31500 5348
rect 31556 5292 34748 5348
rect 34804 5292 34814 5348
rect 38770 5292 38780 5348
rect 38836 5292 41244 5348
rect 41300 5292 41310 5348
rect 25900 5236 25956 5292
rect 41916 5236 41972 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 57344 5460 57456 5488
rect 42130 5404 42140 5460
rect 42196 5404 44268 5460
rect 44324 5404 44334 5460
rect 56130 5404 56140 5460
rect 56196 5404 57456 5460
rect 57344 5376 57456 5404
rect 42690 5292 42700 5348
rect 42756 5292 45276 5348
rect 45332 5292 45342 5348
rect 45714 5292 45724 5348
rect 45780 5292 52108 5348
rect 52164 5292 52174 5348
rect 2258 5180 2268 5236
rect 2324 5180 4956 5236
rect 5012 5180 5022 5236
rect 6850 5180 6860 5236
rect 6916 5180 14532 5236
rect 14690 5180 14700 5236
rect 14756 5180 16380 5236
rect 16436 5180 16446 5236
rect 17042 5180 17052 5236
rect 17108 5180 22428 5236
rect 22484 5180 22494 5236
rect 23650 5180 23660 5236
rect 23716 5180 25676 5236
rect 25732 5180 25742 5236
rect 25900 5180 33628 5236
rect 33684 5180 34076 5236
rect 34132 5180 34524 5236
rect 34580 5180 34590 5236
rect 34850 5180 34860 5236
rect 34916 5180 36876 5236
rect 36932 5180 36942 5236
rect 37090 5180 37100 5236
rect 37156 5180 38220 5236
rect 38276 5180 38668 5236
rect 38724 5180 38734 5236
rect 39666 5180 39676 5236
rect 39732 5180 41132 5236
rect 41188 5180 41198 5236
rect 41916 5180 46620 5236
rect 46676 5180 46686 5236
rect 46834 5180 46844 5236
rect 46900 5180 54236 5236
rect 54292 5180 54302 5236
rect 10882 5068 10892 5124
rect 10948 5068 11788 5124
rect 11844 5068 11854 5124
rect 12226 5068 12236 5124
rect 12292 5068 12460 5124
rect 12516 5068 12526 5124
rect 13346 5068 13356 5124
rect 13412 5068 14252 5124
rect 14308 5068 14318 5124
rect 0 5012 112 5040
rect 14476 5012 14532 5180
rect 15810 5068 15820 5124
rect 15876 5068 18396 5124
rect 18452 5068 18462 5124
rect 18834 5068 18844 5124
rect 18900 5068 19404 5124
rect 19460 5068 19470 5124
rect 19852 5068 20972 5124
rect 21028 5068 21038 5124
rect 21196 5068 21308 5124
rect 21364 5068 21374 5124
rect 21858 5068 21868 5124
rect 21924 5068 22316 5124
rect 22372 5068 22382 5124
rect 22530 5068 22540 5124
rect 22596 5068 26460 5124
rect 26516 5068 26526 5124
rect 26674 5068 26684 5124
rect 26740 5068 27580 5124
rect 27636 5068 27646 5124
rect 27794 5068 27804 5124
rect 27860 5068 27916 5124
rect 27972 5068 27982 5124
rect 28252 5068 28476 5124
rect 28532 5068 28542 5124
rect 28690 5068 28700 5124
rect 28756 5068 29708 5124
rect 29764 5068 29774 5124
rect 30146 5068 30156 5124
rect 30212 5068 35308 5124
rect 35364 5068 35374 5124
rect 35746 5068 35756 5124
rect 35812 5068 42028 5124
rect 42084 5068 42094 5124
rect 42252 5068 51660 5124
rect 51716 5068 51996 5124
rect 52052 5068 52062 5124
rect 54898 5068 54908 5124
rect 54964 5068 55468 5124
rect 0 4956 924 5012
rect 980 4956 990 5012
rect 1148 4956 11676 5012
rect 11732 4956 11742 5012
rect 12114 4956 12124 5012
rect 12180 4956 13468 5012
rect 13524 4956 13534 5012
rect 14476 4956 15148 5012
rect 15250 4956 15260 5012
rect 15316 4956 17724 5012
rect 17780 4956 17790 5012
rect 18274 4956 18284 5012
rect 18340 4956 19628 5012
rect 19684 4956 19694 5012
rect 0 4928 112 4956
rect 1148 4900 1204 4956
rect 15092 4900 15148 4956
rect 19852 4900 19908 5068
rect 21196 5012 21252 5068
rect 28252 5012 28308 5068
rect 20738 4956 20748 5012
rect 20804 4956 21252 5012
rect 21410 4956 21420 5012
rect 21476 4956 23212 5012
rect 23268 4956 23278 5012
rect 23538 4956 23548 5012
rect 23604 4956 25340 5012
rect 25396 4956 25406 5012
rect 25554 4956 25564 5012
rect 25620 4956 26908 5012
rect 26964 4956 26974 5012
rect 27458 4956 27468 5012
rect 27524 4956 28308 5012
rect 28466 4956 28476 5012
rect 28532 4956 28924 5012
rect 28980 4956 28990 5012
rect 29138 4956 29148 5012
rect 29204 4956 29932 5012
rect 29988 4956 29998 5012
rect 30146 4956 30156 5012
rect 30212 4956 33516 5012
rect 33572 4956 33582 5012
rect 39218 4956 39228 5012
rect 39284 4956 41916 5012
rect 41972 4956 41982 5012
rect 42252 4900 42308 5068
rect 55412 5012 55468 5068
rect 57344 5012 57456 5040
rect 42690 4956 42700 5012
rect 42756 4956 46396 5012
rect 46452 4956 46462 5012
rect 50372 4956 53564 5012
rect 53620 4956 53630 5012
rect 55412 4956 57456 5012
rect 50372 4900 50428 4956
rect 57344 4928 57456 4956
rect 354 4844 364 4900
rect 420 4844 1204 4900
rect 3266 4844 3276 4900
rect 3332 4844 8764 4900
rect 8820 4844 8830 4900
rect 9884 4844 13244 4900
rect 13300 4844 13310 4900
rect 15092 4844 19908 4900
rect 20066 4844 20076 4900
rect 20132 4844 23436 4900
rect 23492 4844 23502 4900
rect 24658 4844 24668 4900
rect 24724 4844 26908 4900
rect 26964 4844 26974 4900
rect 27122 4844 27132 4900
rect 27188 4844 31612 4900
rect 31668 4844 31678 4900
rect 32722 4844 32732 4900
rect 32788 4844 33068 4900
rect 33124 4844 33134 4900
rect 33282 4844 33292 4900
rect 33348 4844 40684 4900
rect 40740 4844 40750 4900
rect 41916 4844 42308 4900
rect 42812 4844 44268 4900
rect 44324 4844 44334 4900
rect 44930 4844 44940 4900
rect 44996 4844 50428 4900
rect 50530 4844 50540 4900
rect 50596 4844 55132 4900
rect 55188 4844 55198 4900
rect 9884 4788 9940 4844
rect 41916 4788 41972 4844
rect 5842 4732 5852 4788
rect 5908 4732 9940 4788
rect 10098 4732 10108 4788
rect 10164 4732 20188 4788
rect 20244 4732 20254 4788
rect 21410 4732 21420 4788
rect 21476 4732 23660 4788
rect 23716 4732 23726 4788
rect 24322 4732 24332 4788
rect 24388 4732 35756 4788
rect 35812 4732 35822 4788
rect 37986 4732 37996 4788
rect 38052 4732 41972 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 6290 4620 6300 4676
rect 6356 4620 13468 4676
rect 13524 4620 13534 4676
rect 15092 4620 15260 4676
rect 15316 4620 15326 4676
rect 15474 4620 15484 4676
rect 15540 4620 18508 4676
rect 18564 4620 18574 4676
rect 19618 4620 19628 4676
rect 19684 4620 20412 4676
rect 20468 4620 20478 4676
rect 21522 4620 21532 4676
rect 21588 4620 23660 4676
rect 23716 4620 23726 4676
rect 24220 4620 34636 4676
rect 34692 4620 34702 4676
rect 37426 4620 37436 4676
rect 37492 4620 40516 4676
rect 40674 4620 40684 4676
rect 40740 4620 42588 4676
rect 42644 4620 42654 4676
rect 0 4564 112 4592
rect 0 4508 14924 4564
rect 14980 4508 14990 4564
rect 0 4480 112 4508
rect 15092 4452 15148 4620
rect 24220 4564 24276 4620
rect 40460 4564 40516 4620
rect 42812 4564 42868 4844
rect 44258 4732 44268 4788
rect 44324 4732 47404 4788
rect 47460 4732 47470 4788
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 57344 4564 57456 4592
rect 15250 4508 15260 4564
rect 15316 4508 24276 4564
rect 24434 4508 24444 4564
rect 24500 4508 30156 4564
rect 30212 4508 30222 4564
rect 30370 4508 30380 4564
rect 30436 4508 31724 4564
rect 31780 4508 31790 4564
rect 31938 4508 31948 4564
rect 32004 4508 38556 4564
rect 38612 4508 38622 4564
rect 40460 4508 42868 4564
rect 43586 4508 43596 4564
rect 43652 4508 44940 4564
rect 44996 4508 45006 4564
rect 46722 4508 46732 4564
rect 46788 4508 52332 4564
rect 52388 4508 52668 4564
rect 52724 4508 52734 4564
rect 54562 4508 54572 4564
rect 54628 4508 57456 4564
rect 57344 4480 57456 4508
rect 1586 4396 1596 4452
rect 1652 4396 15148 4452
rect 15362 4396 15372 4452
rect 15428 4396 25564 4452
rect 25620 4396 25630 4452
rect 25778 4396 25788 4452
rect 25844 4396 52220 4452
rect 52276 4396 52286 4452
rect 5170 4284 5180 4340
rect 5236 4284 10276 4340
rect 15026 4284 15036 4340
rect 15092 4284 17948 4340
rect 18004 4284 18014 4340
rect 18386 4284 18396 4340
rect 18452 4284 21308 4340
rect 21364 4284 21374 4340
rect 21858 4284 21868 4340
rect 21924 4284 22540 4340
rect 22596 4284 22606 4340
rect 23426 4284 23436 4340
rect 23492 4284 28812 4340
rect 28868 4284 28878 4340
rect 29586 4284 29596 4340
rect 29652 4284 35196 4340
rect 35252 4284 35262 4340
rect 38434 4284 38444 4340
rect 38500 4284 38780 4340
rect 38836 4284 38846 4340
rect 42018 4284 42028 4340
rect 42084 4284 55132 4340
rect 55188 4284 55198 4340
rect 3052 4172 5068 4228
rect 5124 4172 5134 4228
rect 9090 4172 9100 4228
rect 9156 4172 9772 4228
rect 9828 4172 9838 4228
rect 0 4116 112 4144
rect 3052 4116 3108 4172
rect 10220 4116 10276 4284
rect 13794 4172 13804 4228
rect 13860 4172 24220 4228
rect 24276 4172 24286 4228
rect 26562 4172 26572 4228
rect 26628 4172 27244 4228
rect 27300 4172 27310 4228
rect 27794 4172 27804 4228
rect 27860 4172 31836 4228
rect 31892 4172 31902 4228
rect 32162 4172 32172 4228
rect 32228 4172 34860 4228
rect 34916 4172 34926 4228
rect 35298 4172 35308 4228
rect 35364 4172 44828 4228
rect 44884 4172 44894 4228
rect 45378 4172 45388 4228
rect 45444 4172 53228 4228
rect 53284 4172 53294 4228
rect 57344 4116 57456 4144
rect 0 4060 3108 4116
rect 3266 4060 3276 4116
rect 3332 4060 9268 4116
rect 10220 4060 18956 4116
rect 19012 4060 19022 4116
rect 19170 4060 19180 4116
rect 19236 4060 27132 4116
rect 27188 4060 27198 4116
rect 27346 4060 27356 4116
rect 27412 4060 28588 4116
rect 28644 4060 30380 4116
rect 30436 4060 30446 4116
rect 31490 4060 31500 4116
rect 31556 4060 33852 4116
rect 33908 4060 33918 4116
rect 34962 4060 34972 4116
rect 35028 4060 50652 4116
rect 50708 4060 50718 4116
rect 56130 4060 56140 4116
rect 56196 4060 57456 4116
rect 0 4032 112 4060
rect 9212 4004 9268 4060
rect 57344 4032 57456 4060
rect 9212 3948 18564 4004
rect 18722 3948 18732 4004
rect 18788 3948 24332 4004
rect 24388 3948 24398 4004
rect 24892 3948 35308 4004
rect 35364 3948 35374 4004
rect 36194 3948 36204 4004
rect 36260 3948 42476 4004
rect 42532 3948 42542 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 18508 3892 18564 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 6738 3836 6748 3892
rect 6804 3836 13020 3892
rect 13076 3836 13086 3892
rect 13234 3836 13244 3892
rect 13300 3836 15148 3892
rect 15204 3836 15214 3892
rect 18508 3836 23324 3892
rect 23380 3836 23390 3892
rect 24892 3780 24948 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 26002 3836 26012 3892
rect 26068 3836 33628 3892
rect 33684 3836 33694 3892
rect 33852 3836 40348 3892
rect 40404 3836 40414 3892
rect 41682 3836 41692 3892
rect 41748 3836 42980 3892
rect 45490 3836 45500 3892
rect 45556 3836 50316 3892
rect 50372 3836 50382 3892
rect 33852 3780 33908 3836
rect 42924 3780 42980 3836
rect 10210 3724 10220 3780
rect 10276 3724 15036 3780
rect 15092 3724 15102 3780
rect 18274 3724 18284 3780
rect 18340 3724 21476 3780
rect 21634 3724 21644 3780
rect 21700 3724 24948 3780
rect 27122 3724 27132 3780
rect 27188 3724 27580 3780
rect 27636 3724 27646 3780
rect 27794 3724 27804 3780
rect 27860 3724 33908 3780
rect 34962 3724 34972 3780
rect 35028 3724 35420 3780
rect 35476 3724 35486 3780
rect 37650 3724 37660 3780
rect 37716 3724 42700 3780
rect 42756 3724 42766 3780
rect 42924 3724 53564 3780
rect 53620 3724 53630 3780
rect 0 3668 112 3696
rect 21420 3668 21476 3724
rect 57344 3668 57456 3696
rect 0 3612 3332 3668
rect 3602 3612 3612 3668
rect 3668 3612 13356 3668
rect 13412 3612 13422 3668
rect 17826 3612 17836 3668
rect 17892 3612 19068 3668
rect 19124 3612 19134 3668
rect 21420 3612 23492 3668
rect 23650 3612 23660 3668
rect 23716 3612 27244 3668
rect 27300 3612 27310 3668
rect 27458 3612 27468 3668
rect 27524 3612 28700 3668
rect 28756 3612 28766 3668
rect 28914 3612 28924 3668
rect 28980 3612 31500 3668
rect 31556 3612 31566 3668
rect 31826 3612 31836 3668
rect 31892 3612 40180 3668
rect 40338 3612 40348 3668
rect 40404 3612 42308 3668
rect 44818 3612 44828 3668
rect 44884 3612 53676 3668
rect 53732 3612 53742 3668
rect 54898 3612 54908 3668
rect 54964 3612 57456 3668
rect 0 3584 112 3612
rect 3276 3332 3332 3612
rect 23436 3556 23492 3612
rect 8418 3500 8428 3556
rect 8484 3500 18396 3556
rect 18452 3500 18462 3556
rect 19516 3500 21756 3556
rect 21812 3500 21822 3556
rect 23436 3500 25788 3556
rect 25844 3500 25854 3556
rect 26338 3500 26348 3556
rect 26404 3500 26796 3556
rect 26852 3500 29708 3556
rect 29764 3500 29774 3556
rect 29932 3500 36876 3556
rect 36932 3500 36942 3556
rect 19516 3444 19572 3500
rect 29932 3444 29988 3500
rect 40124 3444 40180 3612
rect 42252 3444 42308 3612
rect 57344 3584 57456 3612
rect 42466 3500 42476 3556
rect 42532 3500 54124 3556
rect 54180 3500 54190 3556
rect 12786 3388 12796 3444
rect 12852 3388 15764 3444
rect 18610 3388 18620 3444
rect 18676 3388 19572 3444
rect 20626 3388 20636 3444
rect 20692 3388 23100 3444
rect 23156 3388 23166 3444
rect 23314 3388 23324 3444
rect 23380 3388 26684 3444
rect 26740 3388 26750 3444
rect 27234 3388 27244 3444
rect 27300 3388 29988 3444
rect 30146 3388 30156 3444
rect 30212 3388 38668 3444
rect 38724 3388 38734 3444
rect 40124 3388 41860 3444
rect 42252 3388 45388 3444
rect 45444 3388 45454 3444
rect 53554 3388 53564 3444
rect 53620 3388 56700 3444
rect 56756 3388 56766 3444
rect 15708 3332 15764 3388
rect 41804 3332 42084 3388
rect 3276 3276 6748 3332
rect 6804 3276 6814 3332
rect 13346 3276 13356 3332
rect 13412 3276 15484 3332
rect 15540 3276 15550 3332
rect 15708 3276 23436 3332
rect 23492 3276 23502 3332
rect 23660 3276 26012 3332
rect 26068 3276 26078 3332
rect 27020 3276 34972 3332
rect 35028 3276 35038 3332
rect 35186 3276 35196 3332
rect 35252 3276 36092 3332
rect 36148 3276 36158 3332
rect 37314 3276 37324 3332
rect 37380 3276 38332 3332
rect 38388 3276 38398 3332
rect 38612 3276 40348 3332
rect 40404 3276 40414 3332
rect 42028 3276 50204 3332
rect 50260 3276 50270 3332
rect 50418 3276 50428 3332
rect 50484 3276 51884 3332
rect 51940 3276 51950 3332
rect 0 3220 112 3248
rect 23660 3220 23716 3276
rect 27020 3220 27076 3276
rect 38612 3220 38668 3276
rect 57344 3220 57456 3248
rect 0 3164 3668 3220
rect 10434 3164 10444 3220
rect 10500 3164 19180 3220
rect 19236 3164 19246 3220
rect 20178 3164 20188 3220
rect 20244 3164 21756 3220
rect 21812 3164 21822 3220
rect 22978 3164 22988 3220
rect 23044 3164 23716 3220
rect 24210 3164 24220 3220
rect 24276 3164 26908 3220
rect 27010 3164 27020 3220
rect 27076 3164 27086 3220
rect 27346 3164 27356 3220
rect 27412 3164 32788 3220
rect 33506 3164 33516 3220
rect 33572 3164 38668 3220
rect 38994 3164 39004 3220
rect 39060 3164 42028 3220
rect 42084 3164 42094 3220
rect 45948 3164 48076 3220
rect 48132 3164 48142 3220
rect 51314 3164 51324 3220
rect 51380 3164 52780 3220
rect 52836 3164 52846 3220
rect 54562 3164 54572 3220
rect 54628 3164 57456 3220
rect 0 3136 112 3164
rect 3612 2996 3668 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 26852 3108 26908 3164
rect 32732 3108 32788 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 18722 3052 18732 3108
rect 18788 3052 23660 3108
rect 23716 3052 23726 3108
rect 24210 3052 24220 3108
rect 24276 3052 26236 3108
rect 26292 3052 26302 3108
rect 26852 3052 27972 3108
rect 28354 3052 28364 3108
rect 28420 3052 30940 3108
rect 30996 3052 32508 3108
rect 32564 3052 32574 3108
rect 32732 3052 36764 3108
rect 36820 3052 36830 3108
rect 36978 3052 36988 3108
rect 37044 3052 43596 3108
rect 43652 3052 43662 3108
rect 27916 2996 27972 3052
rect 3612 2940 10332 2996
rect 10388 2940 10398 2996
rect 15026 2940 15036 2996
rect 15092 2940 27692 2996
rect 27748 2940 27758 2996
rect 27916 2940 29484 2996
rect 29540 2940 29550 2996
rect 30258 2940 30268 2996
rect 30324 2940 45724 2996
rect 45780 2940 45790 2996
rect 45948 2884 46004 3164
rect 57344 3136 57456 3164
rect 46946 3052 46956 3108
rect 47012 3052 53564 3108
rect 53620 3052 53630 3108
rect 47058 2940 47068 2996
rect 47124 2940 55132 2996
rect 55188 2940 55198 2996
rect 1138 2828 1148 2884
rect 1204 2828 5628 2884
rect 5684 2828 5694 2884
rect 8194 2828 8204 2884
rect 8260 2828 14252 2884
rect 14308 2828 14318 2884
rect 14914 2828 14924 2884
rect 14980 2828 20188 2884
rect 21746 2828 21756 2884
rect 21812 2828 24780 2884
rect 24836 2828 25676 2884
rect 25732 2828 25742 2884
rect 26002 2828 26012 2884
rect 26068 2828 26908 2884
rect 28914 2828 28924 2884
rect 28980 2828 29820 2884
rect 29876 2828 29886 2884
rect 30034 2828 30044 2884
rect 30100 2828 36596 2884
rect 36866 2828 36876 2884
rect 36932 2828 40684 2884
rect 40740 2828 40750 2884
rect 41570 2828 41580 2884
rect 41636 2828 43372 2884
rect 43428 2828 43438 2884
rect 43586 2828 43596 2884
rect 43652 2828 46004 2884
rect 46610 2828 46620 2884
rect 46676 2828 52556 2884
rect 52612 2828 52622 2884
rect 0 2772 112 2800
rect 20132 2772 20188 2828
rect 26852 2772 26908 2828
rect 0 2716 1596 2772
rect 1652 2716 1662 2772
rect 7298 2716 7308 2772
rect 7364 2716 18620 2772
rect 18676 2716 18686 2772
rect 20132 2716 25116 2772
rect 25172 2716 25182 2772
rect 26852 2716 36484 2772
rect 0 2688 112 2716
rect 5282 2604 5292 2660
rect 5348 2604 33068 2660
rect 33124 2604 33134 2660
rect 12338 2492 12348 2548
rect 12404 2492 15540 2548
rect 18498 2492 18508 2548
rect 18564 2492 25508 2548
rect 26002 2492 26012 2548
rect 26068 2492 32732 2548
rect 32788 2492 32798 2548
rect 15484 2436 15540 2492
rect 25452 2436 25508 2492
rect 7522 2380 7532 2436
rect 7588 2380 15260 2436
rect 15316 2380 15326 2436
rect 15484 2380 20188 2436
rect 22082 2380 22092 2436
rect 22148 2380 24220 2436
rect 24276 2380 24286 2436
rect 25452 2380 28812 2436
rect 28868 2380 28878 2436
rect 32050 2380 32060 2436
rect 32116 2380 33740 2436
rect 33796 2380 33806 2436
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 20132 2324 20188 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 36428 2324 36484 2716
rect 36540 2548 36596 2828
rect 57344 2772 57456 2800
rect 36754 2716 36764 2772
rect 36820 2716 40124 2772
rect 40180 2716 40190 2772
rect 40338 2716 40348 2772
rect 40404 2716 46284 2772
rect 46340 2716 46350 2772
rect 47954 2716 47964 2772
rect 48020 2716 52108 2772
rect 52164 2716 52174 2772
rect 56130 2716 56140 2772
rect 56196 2716 57456 2772
rect 57344 2688 57456 2716
rect 38546 2604 38556 2660
rect 38612 2604 43932 2660
rect 43988 2604 43998 2660
rect 44146 2604 44156 2660
rect 44212 2604 45052 2660
rect 45108 2604 45118 2660
rect 52770 2604 52780 2660
rect 52836 2604 56476 2660
rect 56532 2604 56542 2660
rect 36540 2492 54124 2548
rect 54180 2492 54190 2548
rect 38658 2380 38668 2436
rect 38724 2380 44156 2436
rect 44212 2380 44222 2436
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 57344 2324 57456 2352
rect 0 2268 3276 2324
rect 3332 2268 3342 2324
rect 10770 2268 10780 2324
rect 10836 2268 19964 2324
rect 20020 2268 20030 2324
rect 20132 2268 23324 2324
rect 23380 2268 23390 2324
rect 25554 2268 25564 2324
rect 25620 2268 31836 2324
rect 31892 2268 31902 2324
rect 35298 2268 35308 2324
rect 35364 2268 36204 2324
rect 36260 2268 36270 2324
rect 36428 2268 42084 2324
rect 43698 2268 43708 2324
rect 43764 2268 44268 2324
rect 44324 2268 44334 2324
rect 44818 2268 44828 2324
rect 44884 2268 53452 2324
rect 53508 2268 53518 2324
rect 54898 2268 54908 2324
rect 54964 2268 57456 2324
rect 0 2240 112 2268
rect 42028 2212 42084 2268
rect 57344 2240 57456 2268
rect 4946 2156 4956 2212
rect 5012 2156 15372 2212
rect 15428 2156 15438 2212
rect 18386 2156 18396 2212
rect 18452 2156 20524 2212
rect 20580 2156 20590 2212
rect 22418 2156 22428 2212
rect 22484 2156 23100 2212
rect 23156 2156 23436 2212
rect 23492 2156 24332 2212
rect 24388 2156 25116 2212
rect 25172 2156 25182 2212
rect 29698 2156 29708 2212
rect 29764 2156 30156 2212
rect 30212 2156 30492 2212
rect 30548 2156 33292 2212
rect 33348 2156 33358 2212
rect 33628 2156 38892 2212
rect 38948 2156 38958 2212
rect 40870 2156 40908 2212
rect 40964 2156 41132 2212
rect 41188 2156 41198 2212
rect 42028 2156 47516 2212
rect 47572 2156 47582 2212
rect 33628 2100 33684 2156
rect 6626 2044 6636 2100
rect 6692 2044 14252 2100
rect 14308 2044 14318 2100
rect 18498 2044 18508 2100
rect 18564 2044 26012 2100
rect 26068 2044 26078 2100
rect 26786 2044 26796 2100
rect 26852 2044 33684 2100
rect 33954 2044 33964 2100
rect 34020 2044 36876 2100
rect 36932 2044 36942 2100
rect 37090 2044 37100 2100
rect 37156 2044 51436 2100
rect 51492 2044 51502 2100
rect 52182 2044 52220 2100
rect 52276 2044 52286 2100
rect 8082 1932 8092 1988
rect 8148 1932 28140 1988
rect 28196 1932 28206 1988
rect 28466 1932 28476 1988
rect 28532 1932 32620 1988
rect 32676 1932 32686 1988
rect 32834 1932 32844 1988
rect 32900 1932 36988 1988
rect 37044 1932 37054 1988
rect 38770 1932 38780 1988
rect 38836 1932 43708 1988
rect 43764 1932 43774 1988
rect 43922 1932 43932 1988
rect 43988 1932 48300 1988
rect 48356 1932 48366 1988
rect 0 1876 112 1904
rect 57344 1876 57456 1904
rect 0 1820 9772 1876
rect 9828 1820 9838 1876
rect 14242 1820 14252 1876
rect 14308 1820 29596 1876
rect 29652 1820 29662 1876
rect 30146 1820 30156 1876
rect 30212 1820 40348 1876
rect 40404 1820 40414 1876
rect 41906 1820 41916 1876
rect 41972 1820 48748 1876
rect 48804 1820 49308 1876
rect 49364 1820 49374 1876
rect 53554 1820 53564 1876
rect 53620 1820 57456 1876
rect 0 1792 112 1820
rect 57344 1792 57456 1820
rect 1708 1708 6972 1764
rect 7028 1708 7038 1764
rect 15474 1708 15484 1764
rect 15540 1708 23436 1764
rect 23492 1708 23502 1764
rect 23660 1708 24276 1764
rect 25778 1708 25788 1764
rect 25844 1708 29820 1764
rect 29876 1708 29886 1764
rect 30034 1708 30044 1764
rect 30100 1708 33684 1764
rect 33842 1708 33852 1764
rect 33908 1708 38332 1764
rect 38388 1708 38398 1764
rect 38658 1708 38668 1764
rect 38724 1708 38734 1764
rect 40226 1708 40236 1764
rect 40292 1708 47012 1764
rect 1708 1540 1764 1708
rect 9874 1596 9884 1652
rect 9940 1596 18508 1652
rect 18564 1596 18574 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23660 1540 23716 1708
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 24220 1540 24276 1708
rect 33628 1652 33684 1708
rect 38668 1652 38724 1708
rect 46956 1652 47012 1708
rect 25218 1596 25228 1652
rect 25284 1596 32284 1652
rect 32340 1596 32350 1652
rect 33628 1596 37100 1652
rect 37156 1596 37166 1652
rect 38668 1596 43596 1652
rect 43652 1596 43662 1652
rect 46956 1596 50652 1652
rect 50708 1596 51660 1652
rect 51716 1596 51726 1652
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 1148 1484 1764 1540
rect 5506 1484 5516 1540
rect 5572 1484 8428 1540
rect 15586 1484 15596 1540
rect 15652 1484 23716 1540
rect 24220 1484 26012 1540
rect 26068 1484 26078 1540
rect 29586 1484 29596 1540
rect 29652 1484 33852 1540
rect 33908 1484 33918 1540
rect 35634 1484 35644 1540
rect 35700 1484 39788 1540
rect 39844 1484 39854 1540
rect 40786 1484 40796 1540
rect 40852 1484 43708 1540
rect 47058 1484 47068 1540
rect 47124 1484 47628 1540
rect 47684 1484 47694 1540
rect 0 1428 112 1456
rect 1148 1428 1204 1484
rect 0 1372 1204 1428
rect 1362 1372 1372 1428
rect 1428 1372 6860 1428
rect 6916 1372 6926 1428
rect 0 1344 112 1372
rect 8372 1316 8428 1484
rect 43652 1428 43708 1484
rect 57344 1428 57456 1456
rect 11666 1372 11676 1428
rect 11732 1372 21644 1428
rect 21700 1372 21710 1428
rect 23538 1372 23548 1428
rect 23604 1372 25788 1428
rect 25844 1372 25854 1428
rect 29474 1372 29484 1428
rect 29540 1372 41916 1428
rect 41972 1372 41982 1428
rect 43652 1372 46732 1428
rect 46788 1372 46798 1428
rect 47394 1372 47404 1428
rect 47460 1372 51772 1428
rect 51828 1372 51838 1428
rect 53554 1372 53564 1428
rect 53620 1372 57456 1428
rect 57344 1344 57456 1372
rect 3378 1260 3388 1316
rect 3444 1260 5964 1316
rect 6020 1260 6030 1316
rect 8372 1260 28756 1316
rect 29810 1260 29820 1316
rect 29876 1260 37660 1316
rect 37716 1260 37726 1316
rect 37874 1260 37884 1316
rect 37940 1260 50428 1316
rect 50484 1260 50764 1316
rect 50820 1260 50830 1316
rect 28700 1204 28756 1260
rect 11554 1148 11564 1204
rect 11620 1148 21084 1204
rect 21140 1148 21150 1204
rect 21308 1148 22988 1204
rect 23044 1148 23054 1204
rect 23314 1148 23324 1204
rect 23380 1148 28476 1204
rect 28532 1148 28542 1204
rect 28700 1148 50988 1204
rect 51044 1148 51054 1204
rect 21308 1092 21364 1148
rect 19506 1036 19516 1092
rect 19572 1036 21364 1092
rect 21522 1036 21532 1092
rect 21588 1036 26796 1092
rect 26852 1036 26862 1092
rect 27458 1036 27468 1092
rect 27524 1036 55132 1092
rect 55188 1036 55198 1092
rect 0 980 112 1008
rect 57344 980 57456 1008
rect 0 924 1484 980
rect 1540 924 1550 980
rect 3042 924 3052 980
rect 3108 924 23996 980
rect 24052 924 24062 980
rect 24210 924 24220 980
rect 24276 924 38780 980
rect 38836 924 38846 980
rect 40338 924 40348 980
rect 40404 924 45500 980
rect 45556 924 45566 980
rect 45714 924 45724 980
rect 45780 924 51100 980
rect 51156 924 51166 980
rect 51986 924 51996 980
rect 52052 924 57456 980
rect 0 896 112 924
rect 57344 896 57456 924
rect 5058 812 5068 868
rect 5124 812 18732 868
rect 18788 812 18798 868
rect 25554 812 25564 868
rect 25620 812 29932 868
rect 29988 812 29998 868
rect 37202 812 37212 868
rect 37268 812 42588 868
rect 42644 812 42654 868
rect 46050 812 46060 868
rect 46116 812 53788 868
rect 53844 812 53854 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 5618 700 5628 756
rect 5684 700 18396 756
rect 18452 700 18462 756
rect 23202 700 23212 756
rect 23268 700 24332 756
rect 24388 700 24398 756
rect 24882 700 24892 756
rect 24948 700 30156 756
rect 30212 700 30222 756
rect 33618 700 33628 756
rect 33684 700 40236 756
rect 40292 700 40302 756
rect 49746 700 49756 756
rect 49812 700 54796 756
rect 54852 700 54862 756
rect 914 588 924 644
rect 980 588 13244 644
rect 13300 588 13310 644
rect 17266 588 17276 644
rect 17332 588 32844 644
rect 32900 588 32910 644
rect 38882 588 38892 644
rect 38948 588 49532 644
rect 49588 588 49598 644
rect 0 532 112 560
rect 57344 532 57456 560
rect 0 476 5180 532
rect 5236 476 5246 532
rect 14354 476 14364 532
rect 14420 476 33964 532
rect 34020 476 34030 532
rect 56466 476 56476 532
rect 56532 476 57456 532
rect 0 448 112 476
rect 57344 448 57456 476
rect 8530 364 8540 420
rect 8596 364 30044 420
rect 30100 364 30110 420
rect 33730 364 33740 420
rect 33796 364 39004 420
rect 39060 364 39070 420
rect 42466 364 42476 420
rect 42532 364 47740 420
rect 47796 364 47806 420
rect 23986 252 23996 308
rect 24052 252 26572 308
rect 26628 252 26638 308
rect 9426 140 9436 196
rect 9492 140 9884 196
rect 9940 140 9950 196
rect 11442 140 11452 196
rect 11508 140 11900 196
rect 11956 140 11966 196
rect 13458 140 13468 196
rect 13524 140 13916 196
rect 13972 140 13982 196
rect 18946 140 18956 196
rect 19012 140 20188 196
rect 21074 140 21084 196
rect 21140 140 27804 196
rect 27860 140 27870 196
rect 33618 140 33628 196
rect 33684 140 34412 196
rect 34468 140 34478 196
rect 41682 140 41692 196
rect 41748 140 41758 196
rect 41906 140 41916 196
rect 41972 140 55804 196
rect 55860 140 55870 196
rect 0 84 112 112
rect 20132 84 20188 140
rect 41692 84 41748 140
rect 57344 84 57456 112
rect 0 28 10780 84
rect 10836 28 10846 84
rect 20132 28 30156 84
rect 30212 28 30222 84
rect 41692 28 47068 84
rect 47124 28 47134 84
rect 56690 28 56700 84
rect 56756 28 57456 84
rect 0 0 112 28
rect 57344 0 57456 28
<< via3 >>
rect 25900 14028 25956 14084
rect 30156 13804 30212 13860
rect 44156 13692 44212 13748
rect 25228 13580 25284 13636
rect 26796 13468 26852 13524
rect 21868 13356 21924 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 35644 13244 35700 13300
rect 25452 13132 25508 13188
rect 16604 12908 16660 12964
rect 22204 12908 22260 12964
rect 40572 12796 40628 12852
rect 40796 12796 40852 12852
rect 45500 12684 45556 12740
rect 20972 12572 21028 12628
rect 42140 12572 42196 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 16604 12460 16660 12516
rect 24220 12460 24276 12516
rect 25452 12460 25508 12516
rect 40572 12236 40628 12292
rect 20972 12012 21028 12068
rect 25676 12012 25732 12068
rect 27804 12012 27860 12068
rect 40348 12012 40404 12068
rect 35196 11900 35252 11956
rect 42140 11900 42196 11956
rect 42364 11900 42420 11956
rect 46396 11900 46452 11956
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 42476 11788 42532 11844
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 18284 11676 18340 11732
rect 24220 11676 24276 11732
rect 42364 11676 42420 11732
rect 21308 11564 21364 11620
rect 25788 11452 25844 11508
rect 42476 11452 42532 11508
rect 14588 11340 14644 11396
rect 26684 11340 26740 11396
rect 27020 11340 27076 11396
rect 35196 11340 35252 11396
rect 26460 11228 26516 11284
rect 16156 11116 16212 11172
rect 20076 11116 20132 11172
rect 26012 11116 26068 11172
rect 38220 11116 38276 11172
rect 39004 11116 39060 11172
rect 22428 11004 22484 11060
rect 27692 11004 27748 11060
rect 31836 11004 31892 11060
rect 38780 11004 38836 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 20076 10892 20132 10948
rect 25900 10892 25956 10948
rect 26572 10892 26628 10948
rect 27244 10892 27300 10948
rect 29596 10892 29652 10948
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 35084 10892 35140 10948
rect 46172 10892 46228 10948
rect 18060 10668 18116 10724
rect 21308 10668 21364 10724
rect 25004 10668 25060 10724
rect 33516 10668 33572 10724
rect 34860 10668 34916 10724
rect 37772 10668 37828 10724
rect 16492 10444 16548 10500
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 14252 9996 14308 10052
rect 16156 9996 16212 10052
rect 18060 10220 18116 10276
rect 26124 10220 26180 10276
rect 26908 10220 26964 10276
rect 28364 10220 28420 10276
rect 37772 10220 37828 10276
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 25228 10108 25284 10164
rect 28476 10108 28532 10164
rect 39228 10108 39284 10164
rect 42252 10108 42308 10164
rect 21868 9996 21924 10052
rect 39116 9996 39172 10052
rect 44156 9996 44212 10052
rect 46060 9996 46116 10052
rect 26124 9884 26180 9940
rect 52220 9884 52276 9940
rect 28364 9660 28420 9716
rect 30268 9660 30324 9716
rect 37324 9660 37380 9716
rect 38220 9660 38276 9716
rect 44156 9660 44212 9716
rect 26236 9548 26292 9604
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 45276 9436 45332 9492
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 28140 9324 28196 9380
rect 38556 9324 38612 9380
rect 40908 9324 40964 9380
rect 44268 9324 44324 9380
rect 46396 9324 46452 9380
rect 30268 9212 30324 9268
rect 31276 9212 31332 9268
rect 33516 9212 33572 9268
rect 37996 9100 38052 9156
rect 45052 8988 45108 9044
rect 46172 8988 46228 9044
rect 24892 8876 24948 8932
rect 42028 8764 42084 8820
rect 45052 8764 45108 8820
rect 24892 8652 24948 8708
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 32060 8652 32116 8708
rect 31276 8540 31332 8596
rect 32284 8540 32340 8596
rect 38444 8540 38500 8596
rect 38668 8652 38724 8708
rect 39116 8652 39172 8708
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 41132 8540 41188 8596
rect 44268 8540 44324 8596
rect 21868 8428 21924 8484
rect 33852 8428 33908 8484
rect 35084 8316 35140 8372
rect 6300 8204 6356 8260
rect 25228 8204 25284 8260
rect 32620 8204 32676 8260
rect 14700 8092 14756 8148
rect 21868 8092 21924 8148
rect 26684 8092 26740 8148
rect 27020 8092 27076 8148
rect 26908 7980 26964 8036
rect 28588 7980 28644 8036
rect 30492 7980 30548 8036
rect 44828 7980 44884 8036
rect 26684 7868 26740 7924
rect 27916 7868 27972 7924
rect 29596 7868 29652 7924
rect 35868 7868 35924 7924
rect 44156 7868 44212 7924
rect 46844 7868 46900 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 14700 7756 14756 7812
rect 20972 7756 21028 7812
rect 30156 7756 30212 7812
rect 33292 7756 33348 7812
rect 35980 7644 36036 7700
rect 41916 7644 41972 7700
rect 20636 7532 20692 7588
rect 27132 7532 27188 7588
rect 28028 7532 28084 7588
rect 32060 7532 32116 7588
rect 37324 7532 37380 7588
rect 32620 7420 32676 7476
rect 31612 7308 31668 7364
rect 35644 7308 35700 7364
rect 42252 7308 42308 7364
rect 44940 7308 44996 7364
rect 45388 7308 45444 7364
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 14588 7196 14644 7252
rect 30156 7196 30212 7252
rect 31836 7196 31892 7252
rect 33068 7196 33124 7252
rect 41916 7196 41972 7252
rect 21420 7084 21476 7140
rect 25452 7084 25508 7140
rect 26460 7084 26516 7140
rect 36988 7084 37044 7140
rect 40348 7084 40404 7140
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44828 7084 44884 7140
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 24220 6972 24276 7028
rect 28028 6860 28084 6916
rect 34860 6860 34916 6916
rect 41132 6860 41188 6916
rect 25452 6748 25508 6804
rect 26684 6748 26740 6804
rect 28252 6636 28308 6692
rect 41692 6636 41748 6692
rect 16492 6524 16548 6580
rect 26236 6524 26292 6580
rect 45388 6524 45444 6580
rect 28700 6412 28756 6468
rect 32956 6412 33012 6468
rect 46956 6412 47012 6468
rect 23660 6300 23716 6356
rect 24220 6300 24276 6356
rect 32396 6300 32452 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 32844 6300 32900 6356
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 27468 6188 27524 6244
rect 31948 6188 32004 6244
rect 45500 6188 45556 6244
rect 31612 6076 31668 6132
rect 32956 6076 33012 6132
rect 22204 5964 22260 6020
rect 22428 5964 22484 6020
rect 26684 5964 26740 6020
rect 33068 5964 33124 6020
rect 26012 5852 26068 5908
rect 21420 5628 21476 5684
rect 21756 5628 21812 5684
rect 23436 5628 23492 5684
rect 26572 5628 26628 5684
rect 26796 5628 26852 5684
rect 27468 5628 27524 5684
rect 28140 5628 28196 5684
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 20636 5516 20692 5572
rect 23324 5516 23380 5572
rect 23660 5516 23716 5572
rect 26124 5516 26180 5572
rect 38668 5516 38724 5572
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 41692 5404 41748 5460
rect 20748 5292 20804 5348
rect 27244 5292 27300 5348
rect 38780 5292 38836 5348
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 44268 5404 44324 5460
rect 42700 5292 42756 5348
rect 45276 5292 45332 5348
rect 23660 5180 23716 5236
rect 46844 5180 46900 5236
rect 26460 5068 26516 5124
rect 27916 5068 27972 5124
rect 28476 5068 28532 5124
rect 15260 4956 15316 5012
rect 21420 4956 21476 5012
rect 25564 4956 25620 5012
rect 26908 4956 26964 5012
rect 29148 4956 29204 5012
rect 29932 4956 29988 5012
rect 30156 4956 30212 5012
rect 39228 4956 39284 5012
rect 13244 4844 13300 4900
rect 23436 4844 23492 4900
rect 27132 4844 27188 4900
rect 31612 4844 31668 4900
rect 33292 4844 33348 4900
rect 44940 4844 44996 4900
rect 23660 4732 23716 4788
rect 37996 4732 38052 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 6300 4620 6356 4676
rect 15260 4620 15316 4676
rect 44268 4732 44324 4788
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 30380 4508 30436 4564
rect 31724 4508 31780 4564
rect 31948 4508 32004 4564
rect 38556 4508 38612 4564
rect 25564 4396 25620 4452
rect 25788 4396 25844 4452
rect 38780 4284 38836 4340
rect 27244 4172 27300 4228
rect 32172 4172 32228 4228
rect 44828 4172 44884 4228
rect 45388 4172 45444 4228
rect 27132 4060 27188 4116
rect 33852 4060 33908 4116
rect 35308 3948 35364 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 13244 3836 13300 3892
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 18284 3724 18340 3780
rect 27132 3724 27188 3780
rect 27580 3724 27636 3780
rect 34972 3724 35028 3780
rect 42700 3724 42756 3780
rect 27244 3612 27300 3668
rect 28924 3612 28980 3668
rect 40348 3612 40404 3668
rect 44828 3612 44884 3668
rect 25788 3500 25844 3556
rect 36876 3500 36932 3556
rect 23100 3388 23156 3444
rect 23324 3388 23380 3444
rect 27244 3388 27300 3444
rect 30156 3388 30212 3444
rect 38668 3388 38724 3444
rect 45388 3388 45444 3444
rect 34972 3276 35028 3332
rect 40348 3276 40404 3332
rect 27356 3164 27412 3220
rect 42028 3164 42084 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 24220 3052 24276 3108
rect 36988 3052 37044 3108
rect 30268 2940 30324 2996
rect 46956 3052 47012 3108
rect 14252 2828 14308 2884
rect 36876 2828 36932 2884
rect 26012 2492 26068 2548
rect 24220 2380 24276 2436
rect 32060 2380 32116 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 40124 2716 40180 2772
rect 38556 2604 38612 2660
rect 38668 2380 38724 2436
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 35308 2268 35364 2324
rect 40908 2156 40964 2212
rect 14252 2044 14308 2100
rect 26012 2044 26068 2100
rect 36876 2044 36932 2100
rect 52220 2044 52276 2100
rect 36988 1932 37044 1988
rect 14252 1820 14308 1876
rect 29820 1708 29876 1764
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 32284 1596 32340 1652
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 29820 1260 29876 1316
rect 21084 1148 21140 1204
rect 27468 1036 27524 1092
rect 46060 812 46116 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 23212 700 23268 756
rect 21084 140 21140 196
rect 30156 28 30212 84
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14224
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 21868 13412 21924 13422
rect 16604 12964 16660 12974
rect 16604 12516 16660 12908
rect 16604 12450 16660 12460
rect 20972 12628 21028 12638
rect 20972 12068 21028 12572
rect 20972 12002 21028 12012
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 18284 11732 18340 11742
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 14588 11396 14644 11406
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 14252 10052 14308 10062
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 6300 8260 6356 8270
rect 6300 4676 6356 8204
rect 6300 4610 6356 4620
rect 13244 4900 13300 4910
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 13244 3892 13300 4844
rect 13244 3826 13300 3836
rect 14252 2884 14308 9996
rect 14588 7252 14644 11340
rect 16156 11172 16212 11182
rect 16156 10052 16212 11116
rect 18060 10724 18116 10734
rect 16156 9986 16212 9996
rect 16492 10500 16548 10510
rect 14700 8148 14756 8158
rect 14700 7812 14756 8092
rect 14700 7746 14756 7756
rect 14588 7186 14644 7196
rect 16492 6580 16548 10444
rect 18060 10276 18116 10668
rect 18060 10210 18116 10220
rect 16492 6514 16548 6524
rect 15260 5012 15316 5022
rect 15260 4676 15316 4956
rect 15260 4610 15316 4620
rect 18284 3780 18340 11676
rect 21308 11620 21364 11630
rect 20076 11172 20132 11182
rect 20076 10948 20132 11116
rect 20076 10882 20132 10892
rect 21308 10724 21364 11564
rect 21308 10658 21364 10668
rect 21868 10052 21924 13356
rect 21868 9986 21924 9996
rect 22204 12964 22260 12974
rect 21868 8484 21924 8494
rect 21868 8148 21924 8428
rect 21868 8082 21924 8092
rect 20972 7812 21028 7822
rect 20972 7678 21028 7756
rect 20636 7622 21028 7678
rect 20636 7588 20692 7622
rect 20636 7522 20692 7532
rect 21420 7140 21476 7150
rect 21420 5684 21476 7084
rect 22204 6020 22260 12908
rect 23776 12572 24096 14224
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 24436 13356 24756 14224
rect 25900 14084 25956 14094
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 22204 5954 22260 5964
rect 22428 11060 22484 11070
rect 22428 6020 22484 11004
rect 23776 11004 24096 12516
rect 24220 12516 24276 12526
rect 24220 11732 24276 12460
rect 24220 11666 24276 11676
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 22428 5954 22484 5964
rect 23660 6356 23716 6366
rect 21420 5618 21476 5628
rect 21756 5684 21812 5694
rect 20636 5572 20692 5582
rect 21756 5518 21812 5628
rect 23436 5684 23492 5694
rect 20636 5158 20692 5516
rect 20748 5462 21812 5518
rect 23324 5572 23380 5582
rect 20748 5348 20804 5462
rect 20748 5282 20804 5292
rect 20636 5102 21476 5158
rect 21420 5012 21476 5102
rect 21420 4946 21476 4956
rect 18284 3714 18340 3724
rect 23100 3482 23268 3538
rect 23100 3444 23156 3482
rect 23100 3378 23156 3388
rect 14252 2818 14308 2828
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 14252 2100 14308 2110
rect 14252 1876 14308 2044
rect 14252 1810 14308 1820
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 21084 1204 21140 1214
rect 21084 196 21140 1148
rect 23212 756 23268 3482
rect 23324 3444 23380 5516
rect 23436 4900 23492 5628
rect 23660 5572 23716 6300
rect 23660 5506 23716 5516
rect 23776 6300 24096 7812
rect 24436 10220 24756 11732
rect 25228 13636 25284 13646
rect 25004 10724 25060 10734
rect 25004 10558 25060 10668
rect 25004 10502 25172 10558
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 25116 10018 25172 10502
rect 25228 10164 25284 13580
rect 25452 13188 25508 13198
rect 25452 12516 25508 13132
rect 25452 12450 25508 12460
rect 25676 12068 25732 12078
rect 25676 11998 25732 12012
rect 25676 11942 25844 11998
rect 25788 11508 25844 11942
rect 25788 11442 25844 11452
rect 25900 10948 25956 14028
rect 30156 13860 30212 13870
rect 26796 13524 26852 13534
rect 26796 12898 26852 13468
rect 26796 12842 27076 12898
rect 27020 12538 27076 12842
rect 27020 12482 27300 12538
rect 26684 11396 26740 11406
rect 26460 11284 26516 11294
rect 25900 10882 25956 10892
rect 26012 11172 26068 11182
rect 25228 10098 25284 10108
rect 25116 9962 25284 10018
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24892 8932 24948 8942
rect 24892 8708 24948 8876
rect 24892 8642 24948 8652
rect 24436 7084 24756 8596
rect 25228 8260 25284 9962
rect 25228 8194 25284 8204
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 24220 7028 24276 7038
rect 24220 6356 24276 6972
rect 24220 6290 24276 6300
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 23436 4834 23492 4844
rect 23660 5236 23716 5246
rect 23660 4788 23716 5180
rect 23660 4722 23716 4732
rect 23776 4732 24096 6244
rect 23324 3378 23380 3388
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23212 690 23268 700
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 24436 5516 24756 7028
rect 25452 7140 25508 7150
rect 25452 6804 25508 7084
rect 25452 6738 25508 6748
rect 26012 5908 26068 11116
rect 26012 5842 26068 5852
rect 26124 10276 26180 10286
rect 26124 9940 26180 10220
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 26124 5572 26180 9884
rect 26236 9604 26292 9614
rect 26236 6580 26292 9548
rect 26460 7140 26516 11228
rect 26460 7074 26516 7084
rect 26572 10948 26628 10958
rect 26236 6514 26292 6524
rect 26572 5684 26628 10892
rect 26684 8148 26740 11340
rect 27020 11396 27076 11406
rect 26684 8082 26740 8092
rect 26796 11222 26964 11278
rect 26684 7924 26740 7934
rect 26684 7858 26740 7868
rect 26796 7858 26852 11222
rect 26908 10276 26964 11222
rect 26908 10210 26964 10220
rect 27020 8148 27076 11340
rect 27244 10948 27300 12482
rect 27804 12068 27860 12078
rect 27244 10882 27300 10892
rect 27692 11060 27748 11070
rect 27020 8082 27076 8092
rect 26684 7802 26852 7858
rect 26908 8036 26964 8046
rect 26684 6804 26740 6814
rect 26684 6020 26740 6748
rect 26684 5954 26740 5964
rect 26572 5618 26628 5628
rect 26796 5684 26852 5694
rect 26124 5506 26180 5516
rect 24436 3948 24756 5460
rect 26796 5158 26852 5628
rect 26460 5124 26852 5158
rect 26516 5102 26852 5124
rect 26460 5058 26516 5068
rect 25564 5012 25620 5022
rect 25564 4452 25620 4956
rect 26908 5012 26964 7980
rect 26908 4946 26964 4956
rect 27132 7588 27188 7598
rect 27132 4900 27188 7532
rect 27468 6244 27524 6254
rect 27468 5684 27524 6188
rect 27468 5618 27524 5628
rect 27692 5518 27748 11004
rect 27356 5462 27748 5518
rect 27132 4834 27188 4844
rect 27244 5348 27300 5358
rect 25564 4386 25620 4396
rect 25788 4452 25844 4462
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 23776 1596 24096 3108
rect 24220 3108 24276 3118
rect 24220 2436 24276 3052
rect 24220 2370 24276 2380
rect 24436 2380 24756 3892
rect 25788 3556 25844 4396
rect 27244 4228 27300 5292
rect 27244 4162 27300 4172
rect 27132 4116 27188 4126
rect 27132 3780 27188 4060
rect 27132 3714 27188 3724
rect 25788 3490 25844 3500
rect 27244 3668 27300 3678
rect 27244 3444 27300 3612
rect 27244 3378 27300 3388
rect 27356 3220 27412 5462
rect 27804 5338 27860 12012
rect 29596 10948 29652 10958
rect 28364 10276 28420 10286
rect 28364 9716 28420 10220
rect 28476 10164 28644 10198
rect 28532 10142 28644 10164
rect 28476 10098 28532 10108
rect 28364 9650 28420 9660
rect 28140 9380 28196 9390
rect 27356 3154 27412 3164
rect 27468 5282 27860 5338
rect 27916 7924 27972 7934
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 21084 130 21140 140
rect 23776 0 24096 1540
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 26012 2548 26068 2558
rect 26012 2100 26068 2492
rect 26012 2034 26068 2044
rect 27468 1092 27524 5282
rect 27916 5124 27972 7868
rect 28028 7588 28084 7598
rect 28028 6916 28084 7532
rect 28028 6850 28084 6860
rect 28140 5684 28196 9324
rect 28588 8036 28644 10142
rect 28588 7970 28644 7980
rect 29596 7924 29652 10892
rect 29596 7858 29652 7868
rect 30156 7812 30212 13804
rect 35644 13300 35700 13310
rect 35196 11956 35252 11966
rect 35196 11396 35252 11900
rect 35196 11330 35252 11340
rect 31836 11060 31892 11070
rect 30268 9716 30324 9726
rect 30268 9268 30324 9660
rect 30268 9202 30324 9212
rect 31276 9268 31332 9278
rect 31276 8596 31332 9212
rect 31276 8530 31332 8540
rect 30156 7746 30212 7756
rect 30492 8036 30548 8046
rect 30156 7252 30212 7262
rect 28252 6692 28308 6702
rect 28252 6598 28308 6636
rect 28252 6542 28756 6598
rect 28700 6468 28756 6542
rect 28700 6402 28756 6412
rect 28140 5618 28196 5628
rect 27916 5058 27972 5068
rect 28476 5124 29204 5158
rect 28532 5102 29204 5124
rect 28476 5058 28532 5068
rect 29148 5012 29204 5102
rect 29148 4946 29204 4956
rect 29932 5012 29988 5022
rect 29932 4618 29988 4956
rect 30156 5012 30212 7196
rect 30156 4946 30212 4956
rect 29932 4564 30436 4618
rect 29932 4562 30380 4564
rect 30380 4498 30436 4508
rect 30492 4438 30548 7980
rect 31612 7364 31668 7374
rect 31612 6132 31668 7308
rect 31836 7252 31892 11004
rect 35084 10948 35140 10958
rect 33516 10724 33572 10734
rect 33516 9268 33572 10668
rect 33516 9202 33572 9212
rect 34860 10724 34916 10734
rect 32060 8708 32116 8718
rect 32060 7588 32116 8652
rect 32060 7522 32116 7532
rect 32284 8596 32340 8606
rect 31836 7186 31892 7196
rect 31612 6066 31668 6076
rect 31948 6244 32004 6254
rect 30268 4382 30548 4438
rect 31612 4900 31668 4910
rect 27580 3780 27636 3790
rect 27580 3718 27636 3724
rect 27580 3668 28980 3718
rect 27580 3662 28924 3668
rect 28924 3602 28980 3612
rect 30156 3444 30212 3454
rect 29820 1764 29876 1774
rect 29820 1316 29876 1708
rect 29820 1250 29876 1260
rect 27468 1026 27524 1036
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 30156 84 30212 3388
rect 30268 2996 30324 4382
rect 31612 4078 31668 4844
rect 31724 4564 31780 4574
rect 31724 4258 31780 4508
rect 31948 4564 32004 6188
rect 31948 4498 32004 4508
rect 31724 4228 32228 4258
rect 31724 4202 32172 4228
rect 32172 4162 32228 4172
rect 31612 4022 32116 4078
rect 30268 2930 30324 2940
rect 32060 2436 32116 4022
rect 32060 2370 32116 2380
rect 32284 1652 32340 8540
rect 33852 8484 33908 8494
rect 32620 8260 32676 8270
rect 32620 7476 32676 8204
rect 32620 7410 32676 7420
rect 33292 7812 33348 7822
rect 33068 7252 33124 7262
rect 32956 6468 33012 6478
rect 32396 6362 32900 6418
rect 32396 6356 32452 6362
rect 32396 6290 32452 6300
rect 32844 6356 32900 6362
rect 32844 6290 32900 6300
rect 32956 6132 33012 6412
rect 32956 6066 33012 6076
rect 33068 6020 33124 7196
rect 33068 5954 33124 5964
rect 33292 4900 33348 7756
rect 33292 4834 33348 4844
rect 33852 4116 33908 8428
rect 34860 6916 34916 10668
rect 35084 8372 35140 10892
rect 35084 8306 35140 8316
rect 35644 7364 35700 13244
rect 40572 12852 40628 12862
rect 40572 12292 40628 12796
rect 40572 12226 40628 12236
rect 40796 12852 40852 12862
rect 40348 12068 40404 12078
rect 38220 11172 38276 11182
rect 37772 10724 37828 10734
rect 37772 10276 37828 10668
rect 37772 10210 37828 10220
rect 37324 9716 37380 9726
rect 35868 7924 35924 7934
rect 35868 7858 35924 7868
rect 35868 7802 36036 7858
rect 35980 7700 36036 7802
rect 35980 7634 36036 7644
rect 37324 7588 37380 9660
rect 38220 9716 38276 11116
rect 39004 11172 39060 11182
rect 39004 11098 39060 11116
rect 38780 11060 39060 11098
rect 38836 11042 39060 11060
rect 38780 10994 38836 11004
rect 39228 10164 39284 10174
rect 38220 9650 38276 9660
rect 39116 10052 39172 10062
rect 38556 9380 38612 9390
rect 37324 7522 37380 7532
rect 37996 9156 38052 9166
rect 35644 7298 35700 7308
rect 34860 6850 34916 6860
rect 36988 7140 37044 7150
rect 36988 5158 37044 7084
rect 33852 4050 33908 4060
rect 36876 5102 37044 5158
rect 35308 4004 35364 4014
rect 34972 3780 35028 3790
rect 34972 3332 35028 3724
rect 34972 3266 35028 3276
rect 35308 2324 35364 3948
rect 36876 3556 36932 5102
rect 37996 4788 38052 9100
rect 38556 8758 38612 9324
rect 38444 8702 38612 8758
rect 38668 8708 38724 8718
rect 38444 8596 38500 8702
rect 38444 8530 38500 8540
rect 38668 5572 38724 8652
rect 39116 8708 39172 9996
rect 39116 8642 39172 8652
rect 38668 5506 38724 5516
rect 37996 4722 38052 4732
rect 38780 5348 38836 5358
rect 36876 3490 36932 3500
rect 38556 4564 38612 4574
rect 36988 3108 37044 3118
rect 35308 2258 35364 2268
rect 36876 2884 36932 2894
rect 36876 2100 36932 2828
rect 36876 2034 36932 2044
rect 36988 1988 37044 3052
rect 38556 2660 38612 4508
rect 38780 4340 38836 5292
rect 39228 5012 39284 10108
rect 40348 7140 40404 12012
rect 40348 7074 40404 7084
rect 39228 4946 39284 4956
rect 38780 4274 38836 4284
rect 40348 3668 40404 3678
rect 38556 2594 38612 2604
rect 38668 3444 38724 3454
rect 38668 2436 38724 3388
rect 40348 3332 40404 3612
rect 40348 3266 40404 3276
rect 40796 2818 40852 12796
rect 42140 12628 42196 12638
rect 42140 11956 42196 12572
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 42140 11890 42196 11900
rect 42364 11956 42420 11966
rect 42364 11732 42420 11900
rect 42364 11666 42420 11676
rect 42476 11844 42532 11854
rect 42476 11508 42532 11788
rect 42476 11442 42532 11452
rect 43776 11004 44096 12516
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 42252 10164 42308 10174
rect 40124 2772 40852 2818
rect 40180 2762 40852 2772
rect 40908 9380 40964 9390
rect 40124 2706 40180 2716
rect 38668 2370 38724 2380
rect 40908 2212 40964 9324
rect 42028 8820 42084 8830
rect 41132 8596 41188 8606
rect 41132 6916 41188 8540
rect 41916 7700 41972 7710
rect 41916 7252 41972 7644
rect 41916 7186 41972 7196
rect 41132 6850 41188 6860
rect 41692 6692 41748 6702
rect 41692 5460 41748 6636
rect 41692 5394 41748 5404
rect 42028 3220 42084 8764
rect 42252 7364 42308 10108
rect 42252 7298 42308 7308
rect 43776 9436 44096 10948
rect 44156 13748 44212 13758
rect 44156 10052 44212 13692
rect 44156 9986 44212 9996
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 44156 9716 44212 9726
rect 44156 7924 44212 9660
rect 44268 9380 44324 9390
rect 44268 8596 44324 9324
rect 44268 8530 44324 8540
rect 44436 8652 44756 10164
rect 45500 12740 45556 12750
rect 45276 9492 45332 9502
rect 45052 9044 45108 9054
rect 45052 8820 45108 8988
rect 45052 8754 45108 8764
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44156 7858 44212 7868
rect 43776 6300 44096 7812
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 42700 5348 42756 5358
rect 42700 3780 42756 5292
rect 42700 3714 42756 3724
rect 43776 4732 44096 6244
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44828 8036 44884 8046
rect 44828 7140 44884 7980
rect 44828 7074 44884 7084
rect 44940 7364 44996 7374
rect 44436 5516 44756 7028
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 44268 5460 44324 5470
rect 44268 4788 44324 5404
rect 44268 4722 44324 4732
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 42028 3154 42084 3164
rect 43776 3164 44096 4676
rect 40908 2146 40964 2156
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 36988 1922 37044 1932
rect 32284 1586 32340 1596
rect 43776 1596 44096 3108
rect 30156 18 30212 28
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 43776 0 44096 1540
rect 44436 3948 44756 5460
rect 44940 4900 44996 7308
rect 45276 5348 45332 9436
rect 45388 7364 45444 7374
rect 45388 6580 45444 7308
rect 45388 6514 45444 6524
rect 45500 6244 45556 12684
rect 46396 11956 46452 11966
rect 46172 10948 46228 10958
rect 45500 6178 45556 6188
rect 46060 10052 46116 10062
rect 45276 5282 45332 5292
rect 44940 4834 44996 4844
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 44828 4228 44884 4238
rect 44828 3668 44884 4172
rect 44828 3602 44884 3612
rect 45388 4228 45444 4238
rect 45388 3444 45444 4172
rect 45388 3378 45444 3388
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 46060 868 46116 9996
rect 46172 9044 46228 10892
rect 46396 9380 46452 11900
rect 46396 9314 46452 9324
rect 52220 9940 52276 9950
rect 46172 8978 46228 8988
rect 46844 7924 46900 7934
rect 46844 5236 46900 7868
rect 46844 5170 46900 5180
rect 46956 6468 47012 6478
rect 46956 3108 47012 6412
rect 46956 3042 47012 3052
rect 52220 2100 52276 9884
rect 52220 2034 52276 2044
rect 46060 802 46116 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _043_
timestamp 1486834041
transform 1 0 41440 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _044_
timestamp 1486834041
transform 1 0 40544 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _045_
timestamp 1486834041
transform -1 0 42784 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _046_
timestamp 1486834041
transform -1 0 39760 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _047_
timestamp 1486834041
transform 1 0 38528 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _048_
timestamp 1486834041
transform -1 0 19264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _049_
timestamp 1486834041
transform 1 0 18144 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _050_
timestamp 1486834041
transform -1 0 27552 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _051_
timestamp 1486834041
transform 1 0 26656 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _052_
timestamp 1486834041
transform 1 0 10416 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _053_
timestamp 1486834041
transform -1 0 11872 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _054_
timestamp 1486834041
transform -1 0 39312 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _055_
timestamp 1486834041
transform -1 0 42448 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _056_
timestamp 1486834041
transform -1 0 36960 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _057_
timestamp 1486834041
transform 1 0 39424 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _058_
timestamp 1486834041
transform 1 0 42560 0 -1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _059_
timestamp 1486834041
transform 1 0 40992 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _060_
timestamp 1486834041
transform -1 0 40992 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _061_
timestamp 1486834041
transform -1 0 41440 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _062_
timestamp 1486834041
transform -1 0 43792 0 1 8624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _063_
timestamp 1486834041
transform 1 0 40880 0 -1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _064_
timestamp 1486834041
transform 1 0 40656 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _065_
timestamp 1486834041
transform -1 0 39760 0 1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _066_
timestamp 1486834041
transform -1 0 39872 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _067_
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _068_
timestamp 1486834041
transform -1 0 37520 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _069_
timestamp 1486834041
transform -1 0 38864 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _070_
timestamp 1486834041
transform 1 0 17696 0 1 3920
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _071_
timestamp 1486834041
transform -1 0 18928 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _072_
timestamp 1486834041
transform 1 0 18256 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_
timestamp 1486834041
transform 1 0 18256 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _074_
timestamp 1486834041
transform 1 0 20832 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _075_
timestamp 1486834041
transform -1 0 20160 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _076_
timestamp 1486834041
transform 1 0 18592 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _077_
timestamp 1486834041
transform 1 0 26432 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _078_
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _079_
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _080_
timestamp 1486834041
transform -1 0 27776 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _081_
timestamp 1486834041
transform 1 0 28784 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _082_
timestamp 1486834041
transform -1 0 30128 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _083_
timestamp 1486834041
transform 1 0 28560 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _084_
timestamp 1486834041
transform 1 0 10752 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _085_
timestamp 1486834041
transform 1 0 12544 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _086_
timestamp 1486834041
transform -1 0 12432 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _087_
timestamp 1486834041
transform 1 0 10864 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _088_
timestamp 1486834041
transform 1 0 12320 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _089_
timestamp 1486834041
transform -1 0 12320 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _090_
timestamp 1486834041
transform 1 0 11760 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _091_
timestamp 1486834041
transform 1 0 22064 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _092_
timestamp 1486834041
transform 1 0 32368 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _093_
timestamp 1486834041
transform 1 0 26432 0 -1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _094_
timestamp 1486834041
transform 1 0 31136 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _095_
timestamp 1486834041
transform 1 0 29680 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _096_
timestamp 1486834041
transform 1 0 25872 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _097_
timestamp 1486834041
transform 1 0 30128 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _098_
timestamp 1486834041
transform 1 0 21056 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _099_
timestamp 1486834041
transform 1 0 9184 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _100_
timestamp 1486834041
transform 1 0 7952 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _101_
timestamp 1486834041
transform 1 0 8960 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _102_
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _103_
timestamp 1486834041
transform 1 0 24976 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _104_
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _105_
timestamp 1486834041
transform 1 0 7504 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _106_
timestamp 1486834041
transform 1 0 20944 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _107_
timestamp 1486834041
transform 1 0 15792 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _108_
timestamp 1486834041
transform 1 0 34048 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _109_
timestamp 1486834041
transform 1 0 33824 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _110_
timestamp 1486834041
transform 1 0 36288 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _111_
timestamp 1486834041
transform 1 0 35392 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _112_
timestamp 1486834041
transform 1 0 37520 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _113_
timestamp 1486834041
transform 1 0 33040 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _115_
timestamp 1486834041
transform 1 0 50288 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _116_
timestamp 1486834041
transform 1 0 45248 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _117_
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _118_
timestamp 1486834041
transform 1 0 51856 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _119_
timestamp 1486834041
transform 1 0 9744 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _120_
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _121_
timestamp 1486834041
transform 1 0 25200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _122_
timestamp 1486834041
transform 1 0 13104 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _123_
timestamp 1486834041
transform 1 0 31584 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _124_
timestamp 1486834041
transform 1 0 44352 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _125_
timestamp 1486834041
transform 1 0 40992 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _126_
timestamp 1486834041
transform 1 0 23296 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _127_
timestamp 1486834041
transform 1 0 13216 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _128_
timestamp 1486834041
transform 1 0 29904 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _129_
timestamp 1486834041
transform 1 0 27440 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _130_
timestamp 1486834041
transform 1 0 30800 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _131_
timestamp 1486834041
transform 1 0 21392 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _132_
timestamp 1486834041
transform 1 0 9072 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _133_
timestamp 1486834041
transform 1 0 7616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _134_
timestamp 1486834041
transform 1 0 9184 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _135_
timestamp 1486834041
transform 1 0 24528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _136_
timestamp 1486834041
transform 1 0 25424 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _137_
timestamp 1486834041
transform 1 0 23296 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _138_
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _139_
timestamp 1486834041
transform 1 0 21504 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _140_
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _141_
timestamp 1486834041
transform 1 0 34272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _142_
timestamp 1486834041
transform 1 0 34272 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _143_
timestamp 1486834041
transform 1 0 36512 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _144_
timestamp 1486834041
transform 1 0 35056 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _145_
timestamp 1486834041
transform 1 0 38304 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _146_
timestamp 1486834041
transform 1 0 33376 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _147_
timestamp 1486834041
transform 1 0 36176 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _148_
timestamp 1486834041
transform 1 0 51520 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _149_
timestamp 1486834041
transform 1 0 49728 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _150_
timestamp 1486834041
transform 1 0 46256 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _151_
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _152_
timestamp 1486834041
transform 1 0 49616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _153_
timestamp 1486834041
transform 1 0 45360 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _154_
timestamp 1486834041
transform 1 0 46256 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _155_
timestamp 1486834041
transform 1 0 50400 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _156_
timestamp 1486834041
transform 1 0 39872 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _157_
timestamp 1486834041
transform 1 0 50624 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _158_
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _159_
timestamp 1486834041
transform 1 0 47712 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _160_
timestamp 1486834041
transform -1 0 38640 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _161_
timestamp 1486834041
transform 1 0 51296 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _162_
timestamp 1486834041
transform -1 0 42336 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _163_
timestamp 1486834041
transform -1 0 55216 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _164_
timestamp 1486834041
transform -1 0 32144 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _165_
timestamp 1486834041
transform 1 0 1344 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _166_
timestamp 1486834041
transform -1 0 13664 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _167_
timestamp 1486834041
transform -1 0 31920 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _168_
timestamp 1486834041
transform 1 0 26544 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _169_
timestamp 1486834041
transform -1 0 32032 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _170_
timestamp 1486834041
transform -1 0 22064 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _171_
timestamp 1486834041
transform 1 0 32144 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _172_
timestamp 1486834041
transform -1 0 18816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _173_
timestamp 1486834041
transform -1 0 21616 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _174_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _175_
timestamp 1486834041
transform -1 0 38864 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _176_
timestamp 1486834041
transform -1 0 24192 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _177_
timestamp 1486834041
transform 1 0 32368 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _178_
timestamp 1486834041
transform -1 0 15904 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _179_
timestamp 1486834041
transform -1 0 35280 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _180_
timestamp 1486834041
transform -1 0 22288 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _181_
timestamp 1486834041
transform -1 0 30352 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _182_
timestamp 1486834041
transform -1 0 14224 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _183_
timestamp 1486834041
transform -1 0 37072 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _184_
timestamp 1486834041
transform -1 0 21280 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _185_
timestamp 1486834041
transform -1 0 28896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _186_
timestamp 1486834041
transform -1 0 12432 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _187_
timestamp 1486834041
transform 1 0 52528 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _188_
timestamp 1486834041
transform 1 0 50736 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _189_
timestamp 1486834041
transform 1 0 46816 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _190_
timestamp 1486834041
transform 1 0 44352 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _191_
timestamp 1486834041
transform 1 0 45696 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _192_
timestamp 1486834041
transform 1 0 50736 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _193_
timestamp 1486834041
transform 1 0 49168 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _194_
timestamp 1486834041
transform -1 0 5712 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _195_
timestamp 1486834041
transform -1 0 42560 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _196_
timestamp 1486834041
transform -1 0 18704 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _197_
timestamp 1486834041
transform -1 0 26432 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _198_
timestamp 1486834041
transform 1 0 11424 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _199_
timestamp 1486834041
transform -1 0 43344 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _200_
timestamp 1486834041
transform -1 0 19824 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _201_
timestamp 1486834041
transform -1 0 29232 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _202_
timestamp 1486834041
transform 1 0 12768 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _203_
timestamp 1486834041
transform 1 0 49840 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _204_
timestamp 1486834041
transform 1 0 48832 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _205_
timestamp 1486834041
transform -1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _206_
timestamp 1486834041
transform 1 0 51520 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _207_
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _208_
timestamp 1486834041
transform 1 0 48272 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _209_
timestamp 1486834041
transform 1 0 47600 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _210_
timestamp 1486834041
transform 1 0 49728 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _211_
timestamp 1486834041
transform -1 0 42112 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _212_
timestamp 1486834041
transform -1 0 18144 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _213_
timestamp 1486834041
transform -1 0 28784 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _214_
timestamp 1486834041
transform 1 0 13328 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _215_
timestamp 1486834041
transform -1 0 43008 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _216_
timestamp 1486834041
transform 1 0 18144 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _217_
timestamp 1486834041
transform -1 0 29680 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _218_
timestamp 1486834041
transform 1 0 14224 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _219_
timestamp 1486834041
transform -1 0 49616 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1486834041
transform 1 0 42112 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I0
timestamp 1486834041
transform 1 0 37408 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I1
timestamp 1486834041
transform 1 0 37184 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I0
timestamp 1486834041
transform -1 0 35280 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I1
timestamp 1486834041
transform -1 0 35056 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I0
timestamp 1486834041
transform -1 0 42784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I1
timestamp 1486834041
transform 1 0 42000 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I0
timestamp 1486834041
transform 1 0 42672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I1
timestamp 1486834041
transform -1 0 43120 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I0
timestamp 1486834041
transform 1 0 40656 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I1
timestamp 1486834041
transform 1 0 40432 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I0
timestamp 1486834041
transform 1 0 42336 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I1
timestamp 1486834041
transform 1 0 42560 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I0
timestamp 1486834041
transform -1 0 36176 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I1
timestamp 1486834041
transform -1 0 35504 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I2
timestamp 1486834041
transform -1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I3
timestamp 1486834041
transform -1 0 35728 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I0
timestamp 1486834041
transform 1 0 19376 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I1
timestamp 1486834041
transform 1 0 19600 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I0
timestamp 1486834041
transform 1 0 18928 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I1
timestamp 1486834041
transform 1 0 19152 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I0
timestamp 1486834041
transform -1 0 24640 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I1
timestamp 1486834041
transform -1 0 25312 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I2
timestamp 1486834041
transform -1 0 24864 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I3
timestamp 1486834041
transform -1 0 25088 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I0
timestamp 1486834041
transform -1 0 28336 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I1
timestamp 1486834041
transform -1 0 28560 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I0
timestamp 1486834041
transform 1 0 30016 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I1
timestamp 1486834041
transform -1 0 30464 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I0
timestamp 1486834041
transform -1 0 28784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I1
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I2
timestamp 1486834041
transform 1 0 32368 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I3
timestamp 1486834041
transform 1 0 33264 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I0
timestamp 1486834041
transform -1 0 12544 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I1
timestamp 1486834041
transform 1 0 12544 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I0
timestamp 1486834041
transform -1 0 14448 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I1
timestamp 1486834041
transform 1 0 14448 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I0
timestamp 1486834041
transform -1 0 16128 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I1
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I2
timestamp 1486834041
transform 1 0 15904 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I3
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I0
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I1
timestamp 1486834041
transform 1 0 20944 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I0
timestamp 1486834041
transform 1 0 31808 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I1
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I0
timestamp 1486834041
transform 1 0 25984 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I1
timestamp 1486834041
transform -1 0 26432 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I0
timestamp 1486834041
transform 1 0 30688 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I1
timestamp 1486834041
transform 1 0 30912 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__D
timestamp 1486834041
transform -1 0 29680 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__D
timestamp 1486834041
transform 1 0 25648 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__D
timestamp 1486834041
transform 1 0 29904 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__D
timestamp 1486834041
transform 1 0 20832 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__D
timestamp 1486834041
transform 1 0 8848 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__D
timestamp 1486834041
transform 1 0 7728 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__D
timestamp 1486834041
transform 1 0 8736 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__D
timestamp 1486834041
transform 1 0 23968 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__D
timestamp 1486834041
transform 1 0 24752 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__D
timestamp 1486834041
transform -1 0 24416 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__D
timestamp 1486834041
transform -1 0 7504 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__D
timestamp 1486834041
transform 1 0 20720 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__D
timestamp 1486834041
transform 1 0 15568 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__D
timestamp 1486834041
transform 1 0 33824 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__D
timestamp 1486834041
transform 1 0 33600 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__D
timestamp 1486834041
transform -1 0 36288 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__D
timestamp 1486834041
transform 1 0 35168 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__D
timestamp 1486834041
transform 1 0 37296 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__D
timestamp 1486834041
transform 1 0 32816 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I
timestamp 1486834041
transform -1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__I
timestamp 1486834041
transform 1 0 45024 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1486834041
transform -1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__I
timestamp 1486834041
transform 1 0 51632 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1486834041
transform -1 0 9744 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1486834041
transform 1 0 24192 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1486834041
transform -1 0 25200 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1486834041
transform -1 0 13104 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1486834041
transform -1 0 44352 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1486834041
transform -1 0 40992 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1486834041
transform 1 0 23072 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1486834041
transform -1 0 13216 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1486834041
transform 1 0 29680 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1486834041
transform 1 0 28336 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1486834041
transform -1 0 30800 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1486834041
transform 1 0 21168 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1486834041
transform 1 0 8848 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1486834041
transform 1 0 7392 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1486834041
transform -1 0 9184 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1486834041
transform 1 0 24304 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1486834041
transform 1 0 25200 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__I
timestamp 1486834041
transform 1 0 23072 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1486834041
transform 1 0 6384 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I
timestamp 1486834041
transform 1 0 21280 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1486834041
transform -1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I
timestamp 1486834041
transform 1 0 34048 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__I
timestamp 1486834041
transform 1 0 34048 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I
timestamp 1486834041
transform -1 0 36512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1486834041
transform 1 0 34832 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I
timestamp 1486834041
transform -1 0 38304 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1486834041
transform -1 0 33376 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I
timestamp 1486834041
transform 1 0 50624 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1486834041
transform 1 0 49504 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I
timestamp 1486834041
transform 1 0 46032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1486834041
transform 1 0 48160 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I
timestamp 1486834041
transform 1 0 49392 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__I
timestamp 1486834041
transform -1 0 45360 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1486834041
transform 1 0 45696 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1486834041
transform 1 0 50176 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1486834041
transform -1 0 39872 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__I
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1486834041
transform 1 0 46592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1486834041
transform -1 0 47712 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1486834041
transform 1 0 38640 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1486834041
transform 1 0 51072 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1486834041
transform -1 0 42560 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1486834041
transform 1 0 55216 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__I
timestamp 1486834041
transform -1 0 1344 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1486834041
transform -1 0 13888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1486834041
transform 1 0 31024 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1486834041
transform 1 0 18816 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1486834041
transform -1 0 20720 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1486834041
transform 1 0 37744 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1486834041
transform -1 0 32480 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1486834041
transform 1 0 16128 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1486834041
transform -1 0 34384 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1486834041
transform 1 0 22288 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1486834041
transform -1 0 30576 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1486834041
transform 1 0 14224 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1486834041
transform 1 0 35728 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1486834041
transform -1 0 20384 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1486834041
transform -1 0 29120 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1486834041
transform 1 0 52304 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1486834041
transform 1 0 50512 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1486834041
transform -1 0 46816 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1486834041
transform 1 0 44128 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1486834041
transform -1 0 45696 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1486834041
transform 1 0 50512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I
timestamp 1486834041
transform -1 0 49168 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1486834041
transform 1 0 5712 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1486834041
transform 1 0 41440 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1486834041
transform -1 0 18928 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1486834041
transform -1 0 26656 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__I
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1486834041
transform 1 0 42224 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1486834041
transform -1 0 20048 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I
timestamp 1486834041
transform 1 0 29232 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1486834041
transform 1 0 13888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1486834041
transform 1 0 49616 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I
timestamp 1486834041
transform 1 0 48608 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I
timestamp 1486834041
transform -1 0 46592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I
timestamp 1486834041
transform -1 0 51520 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__I
timestamp 1486834041
transform -1 0 53088 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__I
timestamp 1486834041
transform 1 0 48048 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1486834041
transform -1 0 47600 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__I
timestamp 1486834041
transform 1 0 49504 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__I
timestamp 1486834041
transform 1 0 42112 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__I
timestamp 1486834041
transform -1 0 19488 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__I
timestamp 1486834041
transform 1 0 28784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I
timestamp 1486834041
transform 1 0 14672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1486834041
transform 1 0 41888 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1486834041
transform -1 0 19264 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__I
timestamp 1486834041
transform 1 0 29680 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__I
timestamp 1486834041
transform 1 0 15120 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__I
timestamp 1486834041
transform 1 0 48720 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout5_I
timestamp 1486834041
transform 1 0 25648 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout6_I
timestamp 1486834041
transform -1 0 26096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout5
timestamp 1486834041
transform 1 0 25872 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout6
timestamp 1486834041
transform 1 0 26096 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78
timestamp 1486834041
transform 1 0 9408 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93
timestamp 1486834041
transform 1 0 11088 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1486834041
transform 1 0 11984 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1486834041
transform 1 0 13216 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114
timestamp 1486834041
transform 1 0 13440 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129
timestamp 1486834041
transform 1 0 15120 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133
timestamp 1486834041
transform 1 0 15568 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135
timestamp 1486834041
transform 1 0 15792 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_212
timestamp 1486834041
transform 1 0 24416 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_216
timestamp 1486834041
transform 1 0 24864 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_218
timestamp 1486834041
transform 1 0 25088 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_229
timestamp 1486834041
transform 1 0 26320 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_237
timestamp 1486834041
transform 1 0 27216 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_426
timestamp 1486834041
transform 1 0 48384 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_434
timestamp 1486834041
transform 1 0 49280 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_438
timestamp 1486834041
transform 1 0 49728 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 54656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 54880 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_88
timestamp 1486834041
transform 1 0 10528 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_96
timestamp 1486834041
transform 1 0 11424 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_111
timestamp 1486834041
transform 1 0 13104 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_127
timestamp 1486834041
transform 1 0 14896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1486834041
transform 1 0 15792 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_174
timestamp 1486834041
transform 1 0 20160 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_190
timestamp 1486834041
transform 1 0 21952 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_198
timestamp 1486834041
transform 1 0 22848 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_232
timestamp 1486834041
transform 1 0 26656 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_240
timestamp 1486834041
transform 1 0 27552 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_254
timestamp 1486834041
transform 1 0 29120 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_256
timestamp 1486834041
transform 1 0 29344 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_267
timestamp 1486834041
transform 1 0 30576 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_275
timestamp 1486834041
transform 1 0 31472 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_279
timestamp 1486834041
transform 1 0 31920 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_284
timestamp 1486834041
transform 1 0 32480 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_328
timestamp 1486834041
transform 1 0 37408 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_330
timestamp 1486834041
transform 1 0 37632 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_341
timestamp 1486834041
transform 1 0 38864 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_349
timestamp 1486834041
transform 1 0 39760 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_356
timestamp 1486834041
transform 1 0 40544 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_368
timestamp 1486834041
transform 1 0 41888 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_400
timestamp 1486834041
transform 1 0 45472 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_408
timestamp 1486834041
transform 1 0 46368 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_426
timestamp 1486834041
transform 1 0 48384 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1486834041
transform 1 0 48608 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_437
timestamp 1486834041
transform 1 0 49616 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 55776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 56224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_181
timestamp 1486834041
transform 1 0 20944 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_193
timestamp 1486834041
transform 1 0 22288 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_213
timestamp 1486834041
transform 1 0 24528 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_237
timestamp 1486834041
transform 1 0 27216 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_293
timestamp 1486834041
transform 1 0 33488 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_301
timestamp 1486834041
transform 1 0 34384 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_338
timestamp 1486834041
transform 1 0 38528 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_346
timestamp 1486834041
transform 1 0 39424 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_358
timestamp 1486834041
transform 1 0 40768 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_362
timestamp 1486834041
transform 1 0 41216 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_374
timestamp 1486834041
transform 1 0 42560 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_382
timestamp 1486834041
transform 1 0 43456 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_384
timestamp 1486834041
transform 1 0 43680 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_403
timestamp 1486834041
transform 1 0 45808 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_411
timestamp 1486834041
transform 1 0 46704 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_415
timestamp 1486834041
transform 1 0 47152 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_417
timestamp 1486834041
transform 1 0 47376 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_428
timestamp 1486834041
transform 1 0 48608 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_444
timestamp 1486834041
transform 1 0 50400 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_84
timestamp 1486834041
transform 1 0 10080 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_116
timestamp 1486834041
transform 1 0 13664 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_132
timestamp 1486834041
transform 1 0 15456 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_150
timestamp 1486834041
transform 1 0 17472 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_152
timestamp 1486834041
transform 1 0 17696 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_173
timestamp 1486834041
transform 1 0 20048 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_205
timestamp 1486834041
transform 1 0 23632 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_228
timestamp 1486834041
transform 1 0 26208 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_240
timestamp 1486834041
transform 1 0 27552 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_248
timestamp 1486834041
transform 1 0 28448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_263
timestamp 1486834041
transform 1 0 30128 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1486834041
transform 1 0 31920 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_282
timestamp 1486834041
transform 1 0 32256 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_285
timestamp 1486834041
transform 1 0 32592 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_301
timestamp 1486834041
transform 1 0 34384 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_305
timestamp 1486834041
transform 1 0 34832 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_307
timestamp 1486834041
transform 1 0 35056 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_330
timestamp 1486834041
transform 1 0 37632 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_346
timestamp 1486834041
transform 1 0 39424 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 47264 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_438
timestamp 1486834041
transform 1 0 49728 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_446
timestamp 1486834041
transform 1 0 50624 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_450
timestamp 1486834041
transform 1 0 51072 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 56224 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 56448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_71
timestamp 1486834041
transform 1 0 8624 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_94
timestamp 1486834041
transform 1 0 11200 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_96
timestamp 1486834041
transform 1 0 11424 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_109
timestamp 1486834041
transform 1 0 12880 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_123
timestamp 1486834041
transform 1 0 14448 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_127
timestamp 1486834041
transform 1 0 14896 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_140
timestamp 1486834041
transform 1 0 16352 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_148
timestamp 1486834041
transform 1 0 17248 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1486834041
transform 1 0 20720 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_202
timestamp 1486834041
transform 1 0 23296 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_242
timestamp 1486834041
transform 1 0 27776 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_244
timestamp 1486834041
transform 1 0 28000 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_252
timestamp 1486834041
transform 1 0 28896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_284
timestamp 1486834041
transform 1 0 32480 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_292
timestamp 1486834041
transform 1 0 33376 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_296
timestamp 1486834041
transform 1 0 33824 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_308
timestamp 1486834041
transform 1 0 35168 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_312
timestamp 1486834041
transform 1 0 35616 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_314
timestamp 1486834041
transform 1 0 35840 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_317
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_333
timestamp 1486834041
transform 1 0 37968 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_341
timestamp 1486834041
transform 1 0 38864 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_349
timestamp 1486834041
transform 1 0 39760 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_381
timestamp 1486834041
transform 1 0 43344 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_387
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_398
timestamp 1486834041
transform 1 0 45248 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_430
timestamp 1486834041
transform 1 0 48832 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_434
timestamp 1486834041
transform 1 0 49280 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_446
timestamp 1486834041
transform 1 0 50624 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_454
timestamp 1486834041
transform 1 0 51520 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_457
timestamp 1486834041
transform 1 0 51856 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_34
timestamp 1486834041
transform 1 0 4480 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_50
timestamp 1486834041
transform 1 0 6272 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_58
timestamp 1486834041
transform 1 0 7168 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_61
timestamp 1486834041
transform 1 0 7504 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_69
timestamp 1486834041
transform 1 0 8400 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_88
timestamp 1486834041
transform 1 0 10528 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_96
timestamp 1486834041
transform 1 0 11424 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_144
timestamp 1486834041
transform 1 0 16800 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_176
timestamp 1486834041
transform 1 0 20384 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_180
timestamp 1486834041
transform 1 0 20832 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_208
timestamp 1486834041
transform 1 0 23968 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_232
timestamp 1486834041
transform 1 0 26656 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_240
timestamp 1486834041
transform 1 0 27552 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_244
timestamp 1486834041
transform 1 0 28000 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_249
timestamp 1486834041
transform 1 0 28560 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_265
timestamp 1486834041
transform 1 0 30352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_277
timestamp 1486834041
transform 1 0 31696 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_284
timestamp 1486834041
transform 1 0 32480 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_292
timestamp 1486834041
transform 1 0 33376 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_316
timestamp 1486834041
transform 1 0 36064 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_332
timestamp 1486834041
transform 1 0 37856 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_336
timestamp 1486834041
transform 1 0 38304 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 47264 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_454
timestamp 1486834041
transform 1 0 51520 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_465
timestamp 1486834041
transform 1 0 52752 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 55776 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 56224 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_45
timestamp 1486834041
transform 1 0 5712 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_49
timestamp 1486834041
transform 1 0 6160 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_81
timestamp 1486834041
transform 1 0 9744 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_89
timestamp 1486834041
transform 1 0 10640 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_93
timestamp 1486834041
transform 1 0 11088 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_95
timestamp 1486834041
transform 1 0 11312 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_100
timestamp 1486834041
transform 1 0 11872 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_181
timestamp 1486834041
transform 1 0 20944 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_183
timestamp 1486834041
transform 1 0 21168 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_194
timestamp 1486834041
transform 1 0 22400 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_210
timestamp 1486834041
transform 1 0 24192 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_221
timestamp 1486834041
transform 1 0 25424 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_257
timestamp 1486834041
transform 1 0 29456 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_298
timestamp 1486834041
transform 1 0 34048 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 35840 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_321
timestamp 1486834041
transform 1 0 36624 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_329
timestamp 1486834041
transform 1 0 37520 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_341
timestamp 1486834041
transform 1 0 38864 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_343
timestamp 1486834041
transform 1 0 39088 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_349
timestamp 1486834041
transform 1 0 39760 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_357
timestamp 1486834041
transform 1 0 40656 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_361
timestamp 1486834041
transform 1 0 41104 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_363
timestamp 1486834041
transform 1 0 41328 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_376
timestamp 1486834041
transform 1 0 42784 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 43680 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_419
timestamp 1486834041
transform 1 0 47600 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_427
timestamp 1486834041
transform 1 0 48496 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_438
timestamp 1486834041
transform 1 0 49728 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_446
timestamp 1486834041
transform 1 0 50624 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_452
timestamp 1486834041
transform 1 0 51296 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1486834041
transform 1 0 51520 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 8064 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_80
timestamp 1486834041
transform 1 0 9632 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_84
timestamp 1486834041
transform 1 0 10080 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_86
timestamp 1486834041
transform 1 0 10304 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_107
timestamp 1486834041
transform 1 0 12656 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_123
timestamp 1486834041
transform 1 0 14448 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_131
timestamp 1486834041
transform 1 0 15344 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_135
timestamp 1486834041
transform 1 0 15792 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_137
timestamp 1486834041
transform 1 0 16016 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_150
timestamp 1486834041
transform 1 0 17472 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_154
timestamp 1486834041
transform 1 0 17920 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_156
timestamp 1486834041
transform 1 0 18144 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_165
timestamp 1486834041
transform 1 0 19152 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_173
timestamp 1486834041
transform 1 0 20048 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_177
timestamp 1486834041
transform 1 0 20496 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_201
timestamp 1486834041
transform 1 0 23184 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_205
timestamp 1486834041
transform 1 0 23632 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_207
timestamp 1486834041
transform 1 0 23856 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_232
timestamp 1486834041
transform 1 0 26656 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_264
timestamp 1486834041
transform 1 0 30240 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_314
timestamp 1486834041
transform 1 0 35840 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_317
timestamp 1486834041
transform 1 0 36176 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_349
timestamp 1486834041
transform 1 0 39760 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1486834041
transform 1 0 40320 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_389
timestamp 1486834041
transform 1 0 44240 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_397
timestamp 1486834041
transform 1 0 45136 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_399
timestamp 1486834041
transform 1 0 45360 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_410
timestamp 1486834041
transform 1 0 46592 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_418
timestamp 1486834041
transform 1 0 47488 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_438
timestamp 1486834041
transform 1 0 49728 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_460
timestamp 1486834041
transform 1 0 52192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 55776 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 56224 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_53
timestamp 1486834041
transform 1 0 6608 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_61
timestamp 1486834041
transform 1 0 7504 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_85
timestamp 1486834041
transform 1 0 10192 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_93
timestamp 1486834041
transform 1 0 11088 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_97
timestamp 1486834041
transform 1 0 11536 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_99
timestamp 1486834041
transform 1 0 11760 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_111
timestamp 1486834041
transform 1 0 13104 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_127
timestamp 1486834041
transform 1 0 14896 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_131
timestamp 1486834041
transform 1 0 15344 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 20160 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_266
timestamp 1486834041
transform 1 0 30464 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_298
timestamp 1486834041
transform 1 0 34048 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_301
timestamp 1486834041
transform 1 0 34384 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_349
timestamp 1486834041
transform 1 0 39760 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_365
timestamp 1486834041
transform 1 0 41552 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_435
timestamp 1486834041
transform 1 0 49392 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_16
timestamp 1486834041
transform 1 0 2464 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_48
timestamp 1486834041
transform 1 0 6048 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_56
timestamp 1486834041
transform 1 0 6944 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_131
timestamp 1486834041
transform 1 0 15344 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_139
timestamp 1486834041
transform 1 0 16240 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_150
timestamp 1486834041
transform 1 0 17472 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_156
timestamp 1486834041
transform 1 0 18144 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_198
timestamp 1486834041
transform 1 0 22848 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 23744 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_228
timestamp 1486834041
transform 1 0 26208 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_236
timestamp 1486834041
transform 1 0 27104 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_240
timestamp 1486834041
transform 1 0 27552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_242
timestamp 1486834041
transform 1 0 27776 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_261
timestamp 1486834041
transform 1 0 29904 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_269
timestamp 1486834041
transform 1 0 30800 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 31920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_282
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_300
timestamp 1486834041
transform 1 0 34272 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_324
timestamp 1486834041
transform 1 0 36960 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_345
timestamp 1486834041
transform 1 0 39312 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_349
timestamp 1486834041
transform 1 0 39760 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_373
timestamp 1486834041
transform 1 0 42448 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1486834041
transform 1 0 46032 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1486834041
transform 1 0 46928 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1486834041
transform 1 0 47376 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1486834041
transform 1 0 47600 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_430
timestamp 1486834041
transform 1 0 48832 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_433
timestamp 1486834041
transform 1 0 49168 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_447
timestamp 1486834041
transform 1 0 50736 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 56224 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 56448 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1486834041
transform 1 0 1120 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_19
timestamp 1486834041
transform 1 0 2800 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_27
timestamp 1486834041
transform 1 0 3696 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_31
timestamp 1486834041
transform 1 0 4144 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_45
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_77
timestamp 1486834041
transform 1 0 9296 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_89
timestamp 1486834041
transform 1 0 10640 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_120
timestamp 1486834041
transform 1 0 14112 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_152
timestamp 1486834041
transform 1 0 17696 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_164
timestamp 1486834041
transform 1 0 19040 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_172
timestamp 1486834041
transform 1 0 19936 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1486834041
transform 1 0 20160 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1486834041
transform 1 0 20720 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_220
timestamp 1486834041
transform 1 0 25312 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_228
timestamp 1486834041
transform 1 0 26208 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_230
timestamp 1486834041
transform 1 0 26432 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_239
timestamp 1486834041
transform 1 0 27440 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_243
timestamp 1486834041
transform 1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_253
timestamp 1486834041
transform 1 0 29008 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_261
timestamp 1486834041
transform 1 0 29904 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_265
timestamp 1486834041
transform 1 0 30352 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_267
timestamp 1486834041
transform 1 0 30576 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_309
timestamp 1486834041
transform 1 0 35280 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_325
timestamp 1486834041
transform 1 0 37072 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_329
timestamp 1486834041
transform 1 0 37520 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_341
timestamp 1486834041
transform 1 0 38864 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_345
timestamp 1486834041
transform 1 0 39312 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_354
timestamp 1486834041
transform 1 0 40320 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_360
timestamp 1486834041
transform 1 0 40992 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_395
timestamp 1486834041
transform 1 0 44912 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_407
timestamp 1486834041
transform 1 0 46256 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_6
timestamp 1486834041
transform 1 0 1344 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_8
timestamp 1486834041
transform 1 0 1568 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_23
timestamp 1486834041
transform 1 0 3248 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_27
timestamp 1486834041
transform 1 0 3696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_47
timestamp 1486834041
transform 1 0 5936 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_63
timestamp 1486834041
transform 1 0 7728 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1486834041
transform 1 0 8176 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1486834041
transform 1 0 8400 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_103
timestamp 1486834041
transform 1 0 12208 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_105
timestamp 1486834041
transform 1 0 12432 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_116
timestamp 1486834041
transform 1 0 13664 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 15344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_146
timestamp 1486834041
transform 1 0 17024 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_168
timestamp 1486834041
transform 1 0 19488 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_172
timestamp 1486834041
transform 1 0 19936 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_184
timestamp 1486834041
transform 1 0 21280 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_195
timestamp 1486834041
transform 1 0 22512 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_199
timestamp 1486834041
transform 1 0 22960 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_214
timestamp 1486834041
transform 1 0 24640 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_222
timestamp 1486834041
transform 1 0 25536 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_245
timestamp 1486834041
transform 1 0 28112 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_253
timestamp 1486834041
transform 1 0 29008 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_257
timestamp 1486834041
transform 1 0 29456 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_269
timestamp 1486834041
transform 1 0 30800 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_277
timestamp 1486834041
transform 1 0 31696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 39424 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_368
timestamp 1486834041
transform 1 0 41888 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_376
timestamp 1486834041
transform 1 0 42784 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_392
timestamp 1486834041
transform 1 0 44576 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_400
timestamp 1486834041
transform 1 0 45472 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_404
timestamp 1486834041
transform 1 0 45920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_415
timestamp 1486834041
transform 1 0 47152 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 56224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 56448 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_45
timestamp 1486834041
transform 1 0 5712 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_47
timestamp 1486834041
transform 1 0 5936 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1486834041
transform 1 0 12320 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_109
timestamp 1486834041
transform 1 0 12880 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_179
timestamp 1486834041
transform 1 0 20720 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_195
timestamp 1486834041
transform 1 0 22512 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_203
timestamp 1486834041
transform 1 0 23408 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_207
timestamp 1486834041
transform 1 0 23856 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_209
timestamp 1486834041
transform 1 0 24080 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_212
timestamp 1486834041
transform 1 0 24416 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_220
timestamp 1486834041
transform 1 0 25312 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_222
timestamp 1486834041
transform 1 0 25536 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_255
timestamp 1486834041
transform 1 0 29232 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_279
timestamp 1486834041
transform 1 0 31920 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_295
timestamp 1486834041
transform 1 0 33712 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_297
timestamp 1486834041
transform 1 0 33936 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_308
timestamp 1486834041
transform 1 0 35168 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_312
timestamp 1486834041
transform 1 0 35616 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_314
timestamp 1486834041
transform 1 0 35840 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_349
timestamp 1486834041
transform 1 0 39760 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_353
timestamp 1486834041
transform 1 0 40208 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_379
timestamp 1486834041
transform 1 0 43120 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_383
timestamp 1486834041
transform 1 0 43568 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_403
timestamp 1486834041
transform 1 0 45808 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_407
timestamp 1486834041
transform 1 0 46256 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_412
timestamp 1486834041
transform 1 0 46816 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_83
timestamp 1486834041
transform 1 0 9968 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_222
timestamp 1486834041
transform 1 0 25536 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_249
timestamp 1486834041
transform 1 0 28560 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_265
timestamp 1486834041
transform 1 0 30352 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_273
timestamp 1486834041
transform 1 0 31248 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_277
timestamp 1486834041
transform 1 0 31696 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 31920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_284
timestamp 1486834041
transform 1 0 32480 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_292
timestamp 1486834041
transform 1 0 33376 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_318
timestamp 1486834041
transform 1 0 36288 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_344
timestamp 1486834041
transform 1 0 39200 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_348
timestamp 1486834041
transform 1 0 39648 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_356
timestamp 1486834041
transform 1 0 40544 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_376
timestamp 1486834041
transform 1 0 42784 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_392
timestamp 1486834041
transform 1 0 44576 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_398
timestamp 1486834041
transform 1 0 45248 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 55440 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 56224 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 56448 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_47
timestamp 1486834041
transform 1 0 5936 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_107
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_215
timestamp 1486834041
transform 1 0 24752 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1486834041
transform 1 0 27664 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_247
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_263
timestamp 1486834041
transform 1 0 30128 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_289
timestamp 1486834041
transform 1 0 33040 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_305
timestamp 1486834041
transform 1 0 34832 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 35728 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_325
timestamp 1486834041
transform 1 0 37072 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_349
timestamp 1486834041
transform 1 0 39760 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_357
timestamp 1486834041
transform 1 0 40656 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_361
timestamp 1486834041
transform 1 0 41104 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_378
timestamp 1486834041
transform 1 0 43008 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_382
timestamp 1486834041
transform 1 0 43456 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_384
timestamp 1486834041
transform 1 0 43680 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_406
timestamp 1486834041
transform 1 0 46144 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 51184 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_224
timestamp 1486834041
transform 1 0 25760 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_227
timestamp 1486834041
transform 1 0 26096 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_235
timestamp 1486834041
transform 1 0 26992 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_237
timestamp 1486834041
transform 1 0 27216 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_284
timestamp 1486834041
transform 1 0 32480 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_300
timestamp 1486834041
transform 1 0 34272 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_304
timestamp 1486834041
transform 1 0 34720 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_342
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_358
timestamp 1486834041
transform 1 0 40768 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_366
timestamp 1486834041
transform 1 0 41664 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_372
timestamp 1486834041
transform 1 0 42336 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_376
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_392
timestamp 1486834041
transform 1 0 44576 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_439
timestamp 1486834041
transform 1 0 49840 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_472
timestamp 1486834041
transform 1 0 53536 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1486834041
transform 1 0 55776 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_496
timestamp 1486834041
transform 1 0 56224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_498
timestamp 1486834041
transform 1 0 56448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform -1 0 15120 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 52416 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 53424 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 53984 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 54992 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 53424 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 53984 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 54992 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 53424 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 54992 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 54992 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 53424 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 54992 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 53984 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 53424 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 53984 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 50848 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 52416 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 48048 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 50848 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 50848 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 49280 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 52416 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 52416 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 53984 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 54992 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 53424 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 53984 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 48272 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 52752 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 54992 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 52416 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 51632 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 46704 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 52416 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 44800 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 50288 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 49616 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 51968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 51184 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 51856 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 53424 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 54208 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 2800 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 3248 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 3024 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 3808 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 4592 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 3024 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 2912 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 4592 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 4480 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 7728 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 7616 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 6720 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 9184 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 7728 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 8512 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 10640 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 8288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 14112 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 14336 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 16352 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 15680 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 9296 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 12208 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 15344 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 22960 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 20384 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform -1 0 23184 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 24752 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform -1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 18256 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform -1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform -1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 19824 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 20272 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform -1 0 19712 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 21392 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output105
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output106
timestamp 1486834041
transform -1 0 6720 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output107
timestamp 1486834041
transform -1 0 8288 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output108
timestamp 1486834041
transform -1 0 11088 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output109
timestamp 1486834041
transform -1 0 13104 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output110
timestamp 1486834041
transform 1 0 46928 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  S_WARMBOOT_111
timestamp 1486834041
transform -1 0 25760 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 53984 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal2 s 13440 0 13552 112 0 FreeSans 448 0 0 0 BOOT_top
port 0 nsew signal output
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 CONFIGURED_top
port 1 nsew signal input
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 Co
port 2 nsew signal output
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 3 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 4 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 5 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 6 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 7 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 8 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 9 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 10 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 11 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 12 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 13 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 14 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 15 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 16 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 17 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 18 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 19 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 20 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 21 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 22 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 23 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 24 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 25 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 26 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 27 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 28 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 29 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 30 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 31 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 32 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 33 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 34 nsew signal input
flabel metal3 s 57344 0 57456 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 35 nsew signal output
flabel metal3 s 57344 4480 57456 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 36 nsew signal output
flabel metal3 s 57344 4928 57456 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 37 nsew signal output
flabel metal3 s 57344 5376 57456 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 38 nsew signal output
flabel metal3 s 57344 5824 57456 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 39 nsew signal output
flabel metal3 s 57344 6272 57456 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 40 nsew signal output
flabel metal3 s 57344 6720 57456 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 41 nsew signal output
flabel metal3 s 57344 7168 57456 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 42 nsew signal output
flabel metal3 s 57344 7616 57456 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 43 nsew signal output
flabel metal3 s 57344 8064 57456 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 44 nsew signal output
flabel metal3 s 57344 8512 57456 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 45 nsew signal output
flabel metal3 s 57344 448 57456 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 46 nsew signal output
flabel metal3 s 57344 8960 57456 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 47 nsew signal output
flabel metal3 s 57344 9408 57456 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 48 nsew signal output
flabel metal3 s 57344 9856 57456 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 49 nsew signal output
flabel metal3 s 57344 10304 57456 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 50 nsew signal output
flabel metal3 s 57344 10752 57456 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 51 nsew signal output
flabel metal3 s 57344 11200 57456 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 52 nsew signal output
flabel metal3 s 57344 11648 57456 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 53 nsew signal output
flabel metal3 s 57344 12096 57456 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 54 nsew signal output
flabel metal3 s 57344 12544 57456 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 55 nsew signal output
flabel metal3 s 57344 12992 57456 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 56 nsew signal output
flabel metal3 s 57344 896 57456 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 57 nsew signal output
flabel metal3 s 57344 13440 57456 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 58 nsew signal output
flabel metal3 s 57344 13888 57456 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 59 nsew signal output
flabel metal3 s 57344 1344 57456 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 60 nsew signal output
flabel metal3 s 57344 1792 57456 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 61 nsew signal output
flabel metal3 s 57344 2240 57456 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 62 nsew signal output
flabel metal3 s 57344 2688 57456 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 63 nsew signal output
flabel metal3 s 57344 3136 57456 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 64 nsew signal output
flabel metal3 s 57344 3584 57456 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 65 nsew signal output
flabel metal3 s 57344 4032 57456 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 66 nsew signal output
flabel metal2 s 17472 0 17584 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 67 nsew signal input
flabel metal2 s 37632 0 37744 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 68 nsew signal input
flabel metal2 s 39648 0 39760 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 69 nsew signal input
flabel metal2 s 41664 0 41776 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 70 nsew signal input
flabel metal2 s 43680 0 43792 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 71 nsew signal input
flabel metal2 s 45696 0 45808 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 72 nsew signal input
flabel metal2 s 47712 0 47824 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 73 nsew signal input
flabel metal2 s 49728 0 49840 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 74 nsew signal input
flabel metal2 s 51744 0 51856 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 75 nsew signal input
flabel metal2 s 53760 0 53872 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 76 nsew signal input
flabel metal2 s 55776 0 55888 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 77 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 78 nsew signal input
flabel metal2 s 21504 0 21616 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 79 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 80 nsew signal input
flabel metal2 s 25536 0 25648 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 81 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 82 nsew signal input
flabel metal2 s 29568 0 29680 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 83 nsew signal input
flabel metal2 s 31584 0 31696 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 84 nsew signal input
flabel metal2 s 33600 0 33712 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 85 nsew signal input
flabel metal2 s 35616 0 35728 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 86 nsew signal input
flabel metal2 s 48160 14112 48272 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 87 nsew signal output
flabel metal2 s 52640 14112 52752 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 88 nsew signal output
flabel metal2 s 53088 14112 53200 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 89 nsew signal output
flabel metal2 s 53536 14112 53648 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 90 nsew signal output
flabel metal2 s 53984 14112 54096 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 91 nsew signal output
flabel metal2 s 54432 14112 54544 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 92 nsew signal output
flabel metal2 s 54880 14112 54992 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 93 nsew signal output
flabel metal2 s 55328 14112 55440 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 94 nsew signal output
flabel metal2 s 55776 14112 55888 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 95 nsew signal output
flabel metal2 s 56224 14112 56336 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 96 nsew signal output
flabel metal2 s 56672 14112 56784 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 97 nsew signal output
flabel metal2 s 48608 14112 48720 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 98 nsew signal output
flabel metal2 s 49056 14112 49168 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 99 nsew signal output
flabel metal2 s 49504 14112 49616 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 100 nsew signal output
flabel metal2 s 49952 14112 50064 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 101 nsew signal output
flabel metal2 s 50400 14112 50512 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 102 nsew signal output
flabel metal2 s 50848 14112 50960 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 103 nsew signal output
flabel metal2 s 51296 14112 51408 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 104 nsew signal output
flabel metal2 s 51744 14112 51856 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 105 nsew signal output
flabel metal2 s 52192 14112 52304 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 106 nsew signal output
flabel metal2 s 672 14112 784 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 107 nsew signal output
flabel metal2 s 1120 14112 1232 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 108 nsew signal output
flabel metal2 s 1568 14112 1680 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 109 nsew signal output
flabel metal2 s 2016 14112 2128 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 110 nsew signal output
flabel metal2 s 2464 14112 2576 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 111 nsew signal output
flabel metal2 s 2912 14112 3024 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 112 nsew signal output
flabel metal2 s 3360 14112 3472 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 113 nsew signal output
flabel metal2 s 3808 14112 3920 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 114 nsew signal output
flabel metal2 s 4256 14112 4368 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 115 nsew signal output
flabel metal2 s 4704 14112 4816 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 116 nsew signal output
flabel metal2 s 5152 14112 5264 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 117 nsew signal output
flabel metal2 s 5600 14112 5712 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 118 nsew signal output
flabel metal2 s 6048 14112 6160 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 119 nsew signal output
flabel metal2 s 6496 14112 6608 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 120 nsew signal output
flabel metal2 s 6944 14112 7056 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 121 nsew signal output
flabel metal2 s 7392 14112 7504 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 122 nsew signal output
flabel metal2 s 7840 14112 7952 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 123 nsew signal output
flabel metal2 s 8288 14112 8400 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 124 nsew signal output
flabel metal2 s 8736 14112 8848 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 125 nsew signal output
flabel metal2 s 9184 14112 9296 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 126 nsew signal output
flabel metal2 s 9632 14112 9744 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 127 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 128 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 129 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 130 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 131 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 132 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 133 nsew signal output
flabel metal2 s 10080 14112 10192 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 134 nsew signal output
flabel metal2 s 10528 14112 10640 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 135 nsew signal output
flabel metal2 s 10976 14112 11088 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 136 nsew signal output
flabel metal2 s 11424 14112 11536 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 137 nsew signal output
flabel metal2 s 11872 14112 11984 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 138 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 139 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 140 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 141 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 142 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 143 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 144 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 145 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 146 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 147 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 148 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 149 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 150 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 151 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 152 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 153 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 154 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 155 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 156 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 157 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 158 nsew signal output
flabel metal2 s 1344 0 1456 112 0 FreeSans 448 0 0 0 RESET_top
port 159 nsew signal input
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[0]
port 160 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S1END[1]
port 161 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S1END[2]
port 162 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S1END[3]
port 163 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S2END[0]
port 164 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S2END[1]
port 165 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S2END[2]
port 166 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S2END[3]
port 167 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S2END[4]
port 168 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 S2END[5]
port 169 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 S2END[6]
port 170 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 S2END[7]
port 171 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 172 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 173 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 174 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 175 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 176 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 177 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 178 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 179 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 S4END[0]
port 180 nsew signal input
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 S4END[10]
port 181 nsew signal input
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 S4END[11]
port 182 nsew signal input
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 S4END[12]
port 183 nsew signal input
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 S4END[13]
port 184 nsew signal input
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 S4END[14]
port 185 nsew signal input
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 S4END[15]
port 186 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 S4END[1]
port 187 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 S4END[2]
port 188 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 S4END[3]
port 189 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 S4END[4]
port 190 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 S4END[5]
port 191 nsew signal input
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 S4END[6]
port 192 nsew signal input
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 S4END[7]
port 193 nsew signal input
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 S4END[8]
port 194 nsew signal input
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 S4END[9]
port 195 nsew signal input
flabel metal2 s 5376 0 5488 112 0 FreeSans 448 0 0 0 SLOT_top0
port 196 nsew signal output
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 SLOT_top1
port 197 nsew signal output
flabel metal2 s 9408 0 9520 112 0 FreeSans 448 0 0 0 SLOT_top2
port 198 nsew signal output
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 SLOT_top3
port 199 nsew signal output
flabel metal2 s 40544 14112 40656 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 200 nsew signal input
flabel metal2 s 45024 14112 45136 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 201 nsew signal input
flabel metal2 s 45472 14112 45584 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 202 nsew signal input
flabel metal2 s 45920 14112 46032 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 203 nsew signal input
flabel metal2 s 46368 14112 46480 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 204 nsew signal input
flabel metal2 s 46816 14112 46928 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 205 nsew signal input
flabel metal2 s 47264 14112 47376 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 206 nsew signal input
flabel metal2 s 40992 14112 41104 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 207 nsew signal input
flabel metal2 s 41440 14112 41552 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 208 nsew signal input
flabel metal2 s 41888 14112 42000 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 209 nsew signal input
flabel metal2 s 42336 14112 42448 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 210 nsew signal input
flabel metal2 s 42784 14112 42896 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 211 nsew signal input
flabel metal2 s 43232 14112 43344 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 212 nsew signal input
flabel metal2 s 43680 14112 43792 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 213 nsew signal input
flabel metal2 s 44128 14112 44240 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 214 nsew signal input
flabel metal2 s 44576 14112 44688 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 215 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 UserCLK
port 216 nsew signal input
flabel metal2 s 47712 14112 47824 14224 0 FreeSans 448 0 0 0 UserCLKo
port 217 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
rlabel metal1 28728 12544 28728 12544 0 VDD
rlabel metal1 28728 13328 28728 13328 0 VSS
rlabel metal2 13496 126 13496 126 0 BOOT_top
rlabel metal2 3416 686 3416 686 0 CONFIGURED_top
rlabel metal2 10808 1176 10808 1176 0 FrameData[0]
rlabel metal2 25144 2632 25144 2632 0 FrameData[10]
rlabel metal3 518 4984 518 4984 0 FrameData[11]
rlabel metal3 1722 5432 1722 5432 0 FrameData[12]
rlabel metal3 630 5880 630 5880 0 FrameData[13]
rlabel metal3 574 6328 574 6328 0 FrameData[14]
rlabel metal3 19600 3304 19600 3304 0 FrameData[15]
rlabel metal3 854 7224 854 7224 0 FrameData[16]
rlabel metal2 8904 8680 8904 8680 0 FrameData[17]
rlabel metal2 7784 8176 7784 8176 0 FrameData[18]
rlabel metal3 1694 8568 1694 8568 0 FrameData[19]
rlabel metal3 2646 504 2646 504 0 FrameData[1]
rlabel metal3 1694 9016 1694 9016 0 FrameData[20]
rlabel metal3 23296 2856 23296 2856 0 FrameData[21]
rlabel metal2 1120 7672 1120 7672 0 FrameData[22]
rlabel metal3 742 10360 742 10360 0 FrameData[23]
rlabel metal2 20776 7336 20776 7336 0 FrameData[24]
rlabel metal3 182 11256 182 11256 0 FrameData[25]
rlabel metal4 24248 6664 24248 6664 0 FrameData[26]
rlabel metal3 350 12152 350 12152 0 FrameData[27]
rlabel metal3 784 4872 784 4872 0 FrameData[28]
rlabel metal3 798 13048 798 13048 0 FrameData[29]
rlabel metal3 798 952 798 952 0 FrameData[2]
rlabel metal3 126 13496 126 13496 0 FrameData[30]
rlabel metal3 294 13944 294 13944 0 FrameData[31]
rlabel metal3 630 1400 630 1400 0 FrameData[3]
rlabel metal3 4942 1848 4942 1848 0 FrameData[4]
rlabel metal3 1694 2296 1694 2296 0 FrameData[5]
rlabel metal3 854 2744 854 2744 0 FrameData[6]
rlabel metal3 1862 3192 1862 3192 0 FrameData[7]
rlabel metal3 1694 3640 1694 3640 0 FrameData[8]
rlabel metal3 1582 4088 1582 4088 0 FrameData[9]
rlabel metal3 57050 56 57050 56 0 FrameData_O[0]
rlabel metal3 55986 4536 55986 4536 0 FrameData_O[10]
rlabel metal3 55188 5096 55188 5096 0 FrameData_O[11]
rlabel metal2 56168 4984 56168 4984 0 FrameData_O[12]
rlabel metal2 54600 5936 54600 5936 0 FrameData_O[13]
rlabel metal2 55160 6384 55160 6384 0 FrameData_O[14]
rlabel metal2 56168 6440 56168 6440 0 FrameData_O[15]
rlabel metal2 54600 7392 54600 7392 0 FrameData_O[16]
rlabel metal3 56770 7672 56770 7672 0 FrameData_O[17]
rlabel metal3 56658 8120 56658 8120 0 FrameData_O[18]
rlabel metal2 54376 8736 54376 8736 0 FrameData_O[19]
rlabel metal3 56938 504 56938 504 0 FrameData_O[1]
rlabel metal3 56770 9016 56770 9016 0 FrameData_O[20]
rlabel metal2 55160 9520 55160 9520 0 FrameData_O[21]
rlabel metal2 54600 10416 54600 10416 0 FrameData_O[22]
rlabel metal2 55160 8232 55160 8232 0 FrameData_O[23]
rlabel metal3 52920 9576 52920 9576 0 FrameData_O[24]
rlabel metal3 54488 8344 54488 8344 0 FrameData_O[25]
rlabel metal3 52136 11536 52136 11536 0 FrameData_O[26]
rlabel metal2 53032 7784 53032 7784 0 FrameData_O[27]
rlabel metal2 51912 9800 51912 9800 0 FrameData_O[28]
rlabel metal2 53816 12040 53816 12040 0 FrameData_O[29]
rlabel metal2 52024 1120 52024 1120 0 FrameData_O[2]
rlabel metal2 54712 11872 54712 11872 0 FrameData_O[30]
rlabel metal2 51240 9296 51240 9296 0 FrameData_O[31]
rlabel metal3 55482 1400 55482 1400 0 FrameData_O[3]
rlabel metal3 55482 1848 55482 1848 0 FrameData_O[4]
rlabel metal2 54936 2184 54936 2184 0 FrameData_O[5]
rlabel metal2 56168 2072 56168 2072 0 FrameData_O[6]
rlabel metal2 54600 3080 54600 3080 0 FrameData_O[7]
rlabel metal3 56154 3640 56154 3640 0 FrameData_O[8]
rlabel metal2 56168 3528 56168 3528 0 FrameData_O[9]
rlabel metal2 17528 1470 17528 1470 0 FrameStrobe[0]
rlabel metal2 50792 1624 50792 1624 0 FrameStrobe[10]
rlabel metal2 39704 1722 39704 1722 0 FrameStrobe[11]
rlabel metal2 47656 2016 47656 2016 0 FrameStrobe[12]
rlabel metal2 43736 742 43736 742 0 FrameStrobe[13]
rlabel metal2 51128 3304 51128 3304 0 FrameStrobe[14]
rlabel metal2 47768 238 47768 238 0 FrameStrobe[15]
rlabel metal2 49784 406 49784 406 0 FrameStrobe[16]
rlabel metal2 51800 742 51800 742 0 FrameStrobe[17]
rlabel metal2 53816 462 53816 462 0 FrameStrobe[18]
rlabel metal2 41944 784 41944 784 0 FrameStrobe[19]
rlabel metal3 21336 1120 21336 1120 0 FrameStrobe[1]
rlabel metal2 21560 574 21560 574 0 FrameStrobe[2]
rlabel metal2 23576 742 23576 742 0 FrameStrobe[3]
rlabel metal2 25592 462 25592 462 0 FrameStrobe[4]
rlabel metal2 49448 7560 49448 7560 0 FrameStrobe[5]
rlabel metal2 45304 8624 45304 8624 0 FrameStrobe[6]
rlabel metal2 45752 10416 45752 10416 0 FrameStrobe[7]
rlabel metal3 46424 6776 46424 6776 0 FrameStrobe[8]
rlabel metal2 39816 2016 39816 2016 0 FrameStrobe[9]
rlabel metal2 48216 13650 48216 13650 0 FrameStrobe_O[0]
rlabel metal2 52696 13538 52696 13538 0 FrameStrobe_O[10]
rlabel metal2 53144 13706 53144 13706 0 FrameStrobe_O[11]
rlabel metal2 53480 10192 53480 10192 0 FrameStrobe_O[12]
rlabel metal3 53536 9240 53536 9240 0 FrameStrobe_O[13]
rlabel metal2 54488 13202 54488 13202 0 FrameStrobe_O[14]
rlabel metal2 54936 13762 54936 13762 0 FrameStrobe_O[15]
rlabel metal2 55384 13538 55384 13538 0 FrameStrobe_O[16]
rlabel metal2 53256 8512 53256 8512 0 FrameStrobe_O[17]
rlabel metal2 56280 13314 56280 13314 0 FrameStrobe_O[18]
rlabel metal3 54880 6104 54880 6104 0 FrameStrobe_O[19]
rlabel metal2 49112 12656 49112 12656 0 FrameStrobe_O[1]
rlabel metal2 51128 13384 51128 13384 0 FrameStrobe_O[2]
rlabel metal3 49952 11592 49952 11592 0 FrameStrobe_O[3]
rlabel metal2 50008 13594 50008 13594 0 FrameStrobe_O[4]
rlabel metal2 50456 13258 50456 13258 0 FrameStrobe_O[5]
rlabel metal2 50904 12866 50904 12866 0 FrameStrobe_O[6]
rlabel metal2 51352 12922 51352 12922 0 FrameStrobe_O[7]
rlabel metal2 51800 13426 51800 13426 0 FrameStrobe_O[8]
rlabel metal2 52248 13650 52248 13650 0 FrameStrobe_O[9]
rlabel metal2 31920 8904 31920 8904 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 27832 10080 27832 10080 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 32648 5768 32648 5768 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 23016 4872 23016 4872 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 11928 9576 11928 9576 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 13048 7224 13048 7224 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 11368 5096 11368 5096 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 26376 6104 26376 6104 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 26936 3164 26936 3164 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 26600 3528 26600 3528 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 17528 10080 17528 10080 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 22680 7952 22680 7952 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 18032 7336 18032 7336 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 41832 7560 41832 7560 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 39480 6216 39480 6216 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 37128 5432 37128 5432 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 42392 10416 42392 10416 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 40712 10192 40712 10192 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 40040 8904 40040 8904 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 31640 8512 31640 8512 0 Inst_S_WARMBOOT_switch_matrix.N1BEG0
rlabel metal2 26712 9296 26712 9296 0 Inst_S_WARMBOOT_switch_matrix.N1BEG1
rlabel metal3 32256 6104 32256 6104 0 Inst_S_WARMBOOT_switch_matrix.N1BEG2
rlabel metal3 22120 5096 22120 5096 0 Inst_S_WARMBOOT_switch_matrix.N1BEG3
rlabel metal2 1288 8260 1288 8260 0 N1BEG[0]
rlabel metal2 2072 9352 2072 9352 0 N1BEG[1]
rlabel metal2 1624 13034 1624 13034 0 N1BEG[2]
rlabel metal2 2184 11144 2184 11144 0 N1BEG[3]
rlabel metal2 2520 12698 2520 12698 0 N2BEG[0]
rlabel metal2 2968 13202 2968 13202 0 N2BEG[1]
rlabel metal2 2296 12992 2296 12992 0 N2BEG[2]
rlabel metal2 3864 13426 3864 13426 0 N2BEG[3]
rlabel metal2 2184 13216 2184 13216 0 N2BEG[4]
rlabel metal2 4760 13818 4760 13818 0 N2BEG[5]
rlabel metal3 4928 11592 4928 11592 0 N2BEG[6]
rlabel metal2 5656 13650 5656 13650 0 N2BEG[7]
rlabel metal2 6104 13594 6104 13594 0 N2BEGb[0]
rlabel metal2 6440 11984 6440 11984 0 N2BEGb[1]
rlabel metal3 6552 11592 6552 11592 0 N2BEGb[2]
rlabel metal3 6720 13160 6720 13160 0 N2BEGb[3]
rlabel metal2 7952 10808 7952 10808 0 N2BEGb[4]
rlabel metal2 8344 13258 8344 13258 0 N2BEGb[5]
rlabel metal3 8288 11592 8288 11592 0 N2BEGb[6]
rlabel metal2 9240 13538 9240 13538 0 N2BEGb[7]
rlabel metal2 7560 13216 7560 13216 0 N4BEG[0]
rlabel metal2 14056 12376 14056 12376 0 N4BEG[10]
rlabel metal2 14616 13202 14616 13202 0 N4BEG[11]
rlabel metal2 13384 13160 13384 13160 0 N4BEG[12]
rlabel metal2 15512 12698 15512 12698 0 N4BEG[13]
rlabel metal2 15960 13258 15960 13258 0 N4BEG[14]
rlabel metal2 16408 13930 16408 13930 0 N4BEG[15]
rlabel metal2 10136 13594 10136 13594 0 N4BEG[1]
rlabel metal2 10584 11914 10584 11914 0 N4BEG[2]
rlabel metal2 11032 13258 11032 13258 0 N4BEG[3]
rlabel metal2 10920 11760 10920 11760 0 N4BEG[4]
rlabel metal2 9800 13552 9800 13552 0 N4BEG[5]
rlabel metal2 12376 12698 12376 12698 0 N4BEG[6]
rlabel metal3 12432 12376 12432 12376 0 N4BEG[7]
rlabel metal3 12320 13160 12320 13160 0 N4BEG[8]
rlabel metal2 13720 13034 13720 13034 0 N4BEG[9]
rlabel metal2 16856 13594 16856 13594 0 NN4BEG[0]
rlabel metal2 21336 13426 21336 13426 0 NN4BEG[10]
rlabel via1 21560 12847 21560 12847 0 NN4BEG[11]
rlabel metal2 22232 13202 22232 13202 0 NN4BEG[12]
rlabel metal2 22680 13650 22680 13650 0 NN4BEG[13]
rlabel metal3 23352 12376 23352 12376 0 NN4BEG[14]
rlabel metal2 23576 13818 23576 13818 0 NN4BEG[15]
rlabel metal2 17304 13258 17304 13258 0 NN4BEG[1]
rlabel metal2 17528 12096 17528 12096 0 NN4BEG[2]
rlabel metal2 18200 13258 18200 13258 0 NN4BEG[3]
rlabel metal3 18032 13160 18032 13160 0 NN4BEG[4]
rlabel metal2 19096 12866 19096 12866 0 NN4BEG[5]
rlabel metal2 19544 13650 19544 13650 0 NN4BEG[6]
rlabel metal3 19488 13160 19488 13160 0 NN4BEG[7]
rlabel metal2 20440 12810 20440 12810 0 NN4BEG[8]
rlabel metal2 20888 13314 20888 13314 0 NN4BEG[9]
rlabel metal2 1400 742 1400 742 0 RESET_top
rlabel metal2 23688 7840 23688 7840 0 S1END[0]
rlabel metal2 24920 12530 24920 12530 0 S1END[1]
rlabel metal2 27608 9800 27608 9800 0 S1END[2]
rlabel metal2 25816 13314 25816 13314 0 S1END[3]
rlabel metal3 18312 6160 18312 6160 0 S2END[0]
rlabel metal3 29400 2856 29400 2856 0 S2END[1]
rlabel metal2 24808 9352 24808 9352 0 S2END[2]
rlabel metal2 35784 9688 35784 9688 0 S2END[3]
rlabel metal2 15736 8288 15736 8288 0 S2END[4]
rlabel metal3 31920 2184 31920 2184 0 S2END[5]
rlabel metal2 22344 9352 22344 9352 0 S2END[6]
rlabel metal2 36344 7784 36344 7784 0 S2END[7]
rlabel metal3 18704 5320 18704 5320 0 S2MID[0]
rlabel metal2 28392 4256 28392 4256 0 S2MID[1]
rlabel metal2 23240 9464 23240 9464 0 S2MID[2]
rlabel metal2 35448 7784 35448 7784 0 S2MID[3]
rlabel metal2 20552 11536 20552 11536 0 S2MID[4]
rlabel metal3 21056 12152 21056 12152 0 S2MID[5]
rlabel metal2 18872 9184 18872 9184 0 S2MID[6]
rlabel metal3 30240 12264 30240 12264 0 S2MID[7]
rlabel metal3 20216 8400 20216 8400 0 S4END[0]
rlabel metal2 50624 8120 50624 8120 0 S4END[10]
rlabel metal2 45864 10136 45864 10136 0 S4END[11]
rlabel metal2 44184 7280 44184 7280 0 S4END[12]
rlabel metal2 46760 1624 46760 1624 0 S4END[13]
rlabel metal2 50568 3640 50568 3640 0 S4END[14]
rlabel metal2 52360 4480 52360 4480 0 S4END[15]
rlabel metal2 29288 6664 29288 6664 0 S4END[1]
rlabel metal2 19432 5152 19432 5152 0 S4END[2]
rlabel metal2 40712 6720 40712 6720 0 S4END[3]
rlabel metal2 23352 1736 23352 1736 0 S4END[4]
rlabel metal3 31976 13160 31976 13160 0 S4END[5]
rlabel metal2 19656 4536 19656 4536 0 S4END[6]
rlabel metal2 40488 6440 40488 6440 0 S4END[7]
rlabel metal2 24248 5824 24248 5824 0 S4END[8]
rlabel metal2 49112 8512 49112 8512 0 S4END[9]
rlabel metal2 5432 686 5432 686 0 SLOT_top0
rlabel metal2 7448 686 7448 686 0 SLOT_top1
rlabel metal2 9464 126 9464 126 0 SLOT_top2
rlabel metal2 11480 126 11480 126 0 SLOT_top3
rlabel metal2 26712 3080 26712 3080 0 SS4END[0]
rlabel metal2 48104 10696 48104 10696 0 SS4END[10]
rlabel metal2 53088 5320 53088 5320 0 SS4END[11]
rlabel metal2 51520 3752 51520 3752 0 SS4END[12]
rlabel metal2 46536 11760 46536 11760 0 SS4END[13]
rlabel metal3 47712 5992 47712 5992 0 SS4END[14]
rlabel metal2 49672 7728 49672 7728 0 SS4END[15]
rlabel metal2 41048 13986 41048 13986 0 SS4END[1]
rlabel metal2 19208 9576 19208 9576 0 SS4END[2]
rlabel metal2 41944 13650 41944 13650 0 SS4END[3]
rlabel metal2 18648 8176 18648 8176 0 SS4END[4]
rlabel metal2 42840 13762 42840 13762 0 SS4END[5]
rlabel metal3 19768 10696 19768 10696 0 SS4END[6]
rlabel metal3 42952 13160 42952 13160 0 SS4END[7]
rlabel metal2 49616 4424 49616 4424 0 SS4END[8]
rlabel metal2 47768 11200 47768 11200 0 SS4END[9]
rlabel metal2 23520 1736 23520 1736 0 UserCLK
rlabel metal2 47432 11368 47432 11368 0 UserCLKo
rlabel metal3 28112 3640 28112 3640 0 _000_
rlabel metal2 29960 2968 29960 2968 0 _001_
rlabel metal2 29288 3472 29288 3472 0 _002_
rlabel metal2 11032 7728 11032 7728 0 _003_
rlabel metal2 12264 7616 12264 7616 0 _004_
rlabel metal2 12152 6720 12152 6720 0 _005_
rlabel metal3 11480 6664 11480 6664 0 _006_
rlabel metal3 12824 4984 12824 4984 0 _007_
rlabel metal2 12040 5544 12040 5544 0 _008_
rlabel metal2 41720 7952 41720 7952 0 _009_
rlabel metal2 40824 8512 40824 8512 0 _010_
rlabel metal2 42504 9240 42504 9240 0 _011_
rlabel metal2 39480 4816 39480 4816 0 _012_
rlabel metal2 38976 5096 38976 5096 0 _013_
rlabel metal2 18760 6888 18760 6888 0 _014_
rlabel metal3 18648 6664 18648 6664 0 _015_
rlabel metal2 27272 3976 27272 3976 0 _016_
rlabel metal2 26992 3752 26992 3752 0 _017_
rlabel metal2 11256 6552 11256 6552 0 _018_
rlabel metal2 11592 6384 11592 6384 0 _019_
rlabel metal2 42280 8400 42280 8400 0 _020_
rlabel metal2 41888 8456 41888 8456 0 _021_
rlabel metal2 36680 8680 36680 8680 0 _022_
rlabel metal3 40600 8904 40600 8904 0 _023_
rlabel metal2 42840 6776 42840 6776 0 _024_
rlabel metal2 41048 10472 41048 10472 0 _025_
rlabel metal3 41384 10360 41384 10360 0 _026_
rlabel metal2 41160 8680 41160 8680 0 _027_
rlabel metal3 40432 5208 40432 5208 0 _028_
rlabel metal2 39592 7224 39592 7224 0 _029_
rlabel metal3 38864 5880 38864 5880 0 _030_
rlabel metal2 39480 5376 39480 5376 0 _031_
rlabel metal2 37352 6664 37352 6664 0 _032_
rlabel metal2 37688 5768 37688 5768 0 _033_
rlabel metal2 17976 5600 17976 5600 0 _034_
rlabel metal2 18424 9352 18424 9352 0 _035_
rlabel metal2 18928 7448 18928 7448 0 _036_
rlabel metal2 18648 7168 18648 7168 0 _037_
rlabel metal2 19992 8232 19992 8232 0 _038_
rlabel metal2 19768 7448 19768 7448 0 _039_
rlabel metal2 27608 4704 27608 4704 0 _040_
rlabel metal2 28504 4648 28504 4648 0 _041_
rlabel metal2 28952 3808 28952 3808 0 _042_
rlabel metal2 39032 1792 39032 1792 0 net1
rlabel metal2 50568 5600 50568 5600 0 net10
rlabel metal3 25704 9408 25704 9408 0 net100
rlabel metal2 52248 4032 52248 4032 0 net101
rlabel metal2 53704 4312 53704 4312 0 net102
rlabel metal2 19992 7392 19992 7392 0 net103
rlabel metal2 20216 11312 20216 11312 0 net104
rlabel metal3 23800 728 23800 728 0 net105
rlabel metal2 23408 11592 23408 11592 0 net106
rlabel metal3 18088 9800 18088 9800 0 net107
rlabel metal3 9296 6104 9296 6104 0 net108
rlabel metal3 25480 2464 25480 2464 0 net109
rlabel metal2 22120 2520 22120 2520 0 net11
rlabel metal2 18760 7448 18760 7448 0 net110
rlabel metal3 24248 14000 24248 14000 0 net111
rlabel metal2 49000 2184 49000 2184 0 net112
rlabel metal2 25480 13328 25480 13328 0 net113
rlabel metal2 55160 7560 55160 7560 0 net12
rlabel metal2 55048 8680 55048 8680 0 net13
rlabel metal4 26040 2296 26040 2296 0 net14
rlabel metal3 50064 2744 50064 2744 0 net15
rlabel metal2 55048 10472 55048 10472 0 net16
rlabel metal2 54152 9240 54152 9240 0 net17
rlabel metal2 24248 1400 24248 1400 0 net18
rlabel metal2 43960 2296 43960 2296 0 net19
rlabel metal3 51800 6888 51800 6888 0 net2
rlabel metal2 51016 9296 51016 9296 0 net20
rlabel metal3 45976 3024 45976 3024 0 net21
rlabel metal2 48216 10976 48216 10976 0 net22
rlabel metal2 50680 5544 50680 5544 0 net23
rlabel metal2 42616 2100 42616 2100 0 net24
rlabel via3 38808 11051 38808 11051 0 net25
rlabel metal3 6972 1512 6972 1512 0 net26
rlabel metal2 39032 10528 39032 10528 0 net27
rlabel metal2 44296 8512 44296 8512 0 net28
rlabel metal2 52528 1176 52528 1176 0 net29
rlabel metal2 53592 3976 53592 3976 0 net3
rlabel metal3 49616 2856 49616 2856 0 net30
rlabel metal2 54152 2296 54152 2296 0 net31
rlabel metal3 41328 1064 41328 1064 0 net32
rlabel metal3 50288 3080 50288 3080 0 net33
rlabel metal3 34272 12824 34272 12824 0 net34
rlabel metal3 51128 2968 51128 2968 0 net35
rlabel metal2 36904 12656 36904 12656 0 net36
rlabel metal3 52080 3192 52080 3192 0 net37
rlabel metal2 55384 11704 55384 11704 0 net38
rlabel metal2 48496 2856 48496 2856 0 net39
rlabel metal2 54152 5432 54152 5432 0 net4
rlabel metal2 52136 9072 52136 9072 0 net40
rlabel metal2 51800 6552 51800 6552 0 net41
rlabel metal3 42504 2856 42504 2856 0 net42
rlabel metal2 48552 11704 48552 11704 0 net43
rlabel metal2 52696 6272 52696 6272 0 net44
rlabel metal2 1960 11648 1960 11648 0 net45
rlabel metal2 52136 5600 52136 5600 0 net46
rlabel metal4 52248 5992 52248 5992 0 net47
rlabel metal2 51968 6776 51968 6776 0 net48
rlabel metal2 46984 10024 46984 10024 0 net49
rlabel metal3 16016 7560 16016 7560 0 net5
rlabel metal2 52360 11480 52360 11480 0 net50
rlabel metal2 52248 10248 52248 10248 0 net51
rlabel metal2 51352 11144 51352 11144 0 net52
rlabel metal2 52136 10696 52136 10696 0 net53
rlabel metal3 52024 6664 52024 6664 0 net54
rlabel metal2 53928 7308 53928 7308 0 net55
rlabel metal2 2296 6720 2296 6720 0 net56
rlabel metal2 2632 8680 2632 8680 0 net57
rlabel metal2 24024 616 24024 616 0 net58
rlabel metal2 2856 8120 2856 8120 0 net59
rlabel metal2 25256 3024 25256 3024 0 net6
rlabel metal3 14448 3304 14448 3304 0 net60
rlabel metal2 18088 9576 18088 9576 0 net61
rlabel metal2 2856 12264 2856 12264 0 net62
rlabel metal2 19544 10752 19544 10752 0 net63
rlabel metal2 2744 11312 2744 11312 0 net64
rlabel metal2 23576 9184 23576 9184 0 net65
rlabel metal3 19208 2632 19208 2632 0 net66
rlabel metal2 15176 4032 15176 4032 0 net67
rlabel metal3 11424 2408 11424 2408 0 net68
rlabel metal3 16408 10080 16408 10080 0 net69
rlabel metal4 23688 5936 23688 5936 0 net7
rlabel metal4 14280 1960 14280 1960 0 net70
rlabel metal2 13496 4536 13496 4536 0 net71
rlabel metal4 18088 10472 18088 10472 0 net72
rlabel metal2 20552 9296 20552 9296 0 net73
rlabel metal3 18144 1960 18144 1960 0 net74
rlabel metal2 11872 4424 11872 4424 0 net75
rlabel metal2 16408 7336 16408 7336 0 net76
rlabel metal2 14616 8568 14616 8568 0 net77
rlabel metal3 13216 10472 13216 10472 0 net78
rlabel metal3 41664 4648 41664 4648 0 net79
rlabel metal2 53592 6216 53592 6216 0 net8
rlabel metal3 18480 3640 18480 3640 0 net80
rlabel metal4 24920 8792 24920 8792 0 net81
rlabel metal2 15848 10304 15848 10304 0 net82
rlabel metal2 51464 2352 51464 2352 0 net83
rlabel metal3 23688 1624 23688 1624 0 net84
rlabel metal4 22456 8512 22456 8512 0 net85
rlabel metal4 21112 672 21112 672 0 net86
rlabel metal2 16744 6328 16744 6328 0 net87
rlabel metal3 46144 3304 46144 3304 0 net88
rlabel metal2 5096 12208 5096 12208 0 net89
rlabel metal2 54264 5936 54264 5936 0 net9
rlabel metal3 25704 13608 25704 13608 0 net90
rlabel metal2 17976 3976 17976 3976 0 net91
rlabel metal4 25256 9111 25256 9111 0 net92
rlabel metal2 22792 9856 22792 9856 0 net93
rlabel metal2 20552 12880 20552 12880 0 net94
rlabel metal2 23016 12432 23016 12432 0 net95
rlabel metal2 18872 9968 18872 9968 0 net96
rlabel metal2 28952 10024 28952 10024 0 net97
rlabel metal2 23912 13440 23912 13440 0 net98
rlabel metal2 17080 13160 17080 13160 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 14224
<< end >>
