module S_term_single2 (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 gf180mcu_fd_sc_mcu7t5v0__buf_2 _000_ (.I(FrameData[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _001_ (.I(FrameData[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _002_ (.I(FrameData[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _003_ (.I(FrameData[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _004_ (.I(FrameData[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _005_ (.I(FrameData[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _006_ (.I(FrameData[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _007_ (.I(FrameData[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _008_ (.I(FrameData[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _009_ (.I(FrameData[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _010_ (.I(FrameData[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _011_ (.I(FrameData[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _012_ (.I(FrameData[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _013_ (.I(FrameData[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _014_ (.I(FrameData[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _015_ (.I(FrameData[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _016_ (.I(FrameData[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _017_ (.I(FrameData[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _018_ (.I(FrameData[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _019_ (.I(FrameData[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _020_ (.I(FrameData[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _021_ (.I(FrameData[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _022_ (.I(FrameData[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _023_ (.I(FrameData[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _024_ (.I(FrameData[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _025_ (.I(FrameData[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _026_ (.I(FrameData[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _027_ (.I(FrameData[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _028_ (.I(FrameData[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _029_ (.I(FrameData[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _030_ (.I(FrameData[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _031_ (.I(FrameData[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _032_ (.I(FrameStrobe[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _033_ (.I(FrameStrobe[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _034_ (.I(FrameStrobe[2]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _035_ (.I(FrameStrobe[3]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _036_ (.I(FrameStrobe[4]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _037_ (.I(FrameStrobe[5]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _038_ (.I(FrameStrobe[6]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _039_ (.I(FrameStrobe[7]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _040_ (.I(FrameStrobe[8]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _041_ (.I(FrameStrobe[9]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _042_ (.I(FrameStrobe[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _043_ (.I(FrameStrobe[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _044_ (.I(FrameStrobe[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _045_ (.I(FrameStrobe[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _046_ (.I(FrameStrobe[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _047_ (.I(FrameStrobe[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _048_ (.I(FrameStrobe[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _049_ (.I(FrameStrobe[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _050_ (.I(FrameStrobe[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _051_ (.I(FrameStrobe[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _052_ (.I(S1END[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _053_ (.I(S1END[2]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _054_ (.I(S1END[1]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _055_ (.I(S1END[0]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _056_ (.I(S2MID[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _057_ (.I(S2MID[6]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _058_ (.I(S2MID[5]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _059_ (.I(S2MID[4]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _060_ (.I(S2MID[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _061_ (.I(S2MID[2]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _062_ (.I(S2MID[1]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _063_ (.I(S2MID[0]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _064_ (.I(S2END[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _065_ (.I(S2END[6]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _066_ (.I(S2END[5]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _067_ (.I(S2END[4]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _068_ (.I(S2END[3]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _069_ (.I(S2END[2]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _070_ (.I(S2END[1]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _071_ (.I(S2END[0]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _072_ (.I(S4END[15]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _073_ (.I(S4END[14]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _074_ (.I(S4END[13]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _075_ (.I(S4END[12]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _076_ (.I(S4END[11]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _077_ (.I(S4END[10]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _078_ (.I(S4END[9]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _079_ (.I(S4END[8]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _080_ (.I(S4END[7]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _081_ (.I(S4END[6]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _082_ (.I(S4END[5]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _083_ (.I(S4END[4]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _084_ (.I(S4END[3]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _085_ (.I(S4END[2]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _086_ (.I(S4END[1]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _087_ (.I(S4END[0]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _088_ (.I(SS4END[15]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _089_ (.I(SS4END[14]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _090_ (.I(SS4END[13]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _091_ (.I(SS4END[12]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _092_ (.I(SS4END[11]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _093_ (.I(SS4END[10]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _094_ (.I(SS4END[9]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _095_ (.I(SS4END[8]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _096_ (.I(SS4END[7]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _097_ (.I(SS4END[6]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _098_ (.I(SS4END[5]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _099_ (.I(SS4END[4]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _100_ (.I(SS4END[3]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _101_ (.I(SS4END[2]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _102_ (.I(SS4END[1]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _103_ (.I(SS4END[0]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _104_ (.I(UserCLK),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_175 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output1 (.I(net1),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output2 (.I(net2),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output3 (.I(net3),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output4 (.I(net4),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output5 (.I(net5),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output6 (.I(net6),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output7 (.I(net7),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output8 (.I(net8),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output9 (.I(net9),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output10 (.I(net10),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output11 (.I(net11),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output12 (.I(net12),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output13 (.I(net13),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output14 (.I(net14),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output15 (.I(net15),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output16 (.I(net16),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output17 (.I(net17),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output18 (.I(net18),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output19 (.I(net19),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output20 (.I(net20),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output21 (.I(net21),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output22 (.I(net22),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output23 (.I(net23),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output24 (.I(net24),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output25 (.I(net25),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output26 (.I(net26),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output27 (.I(net27),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output28 (.I(net28),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output29 (.I(net29),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output30 (.I(net30),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output31 (.I(net31),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output32 (.I(net32),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output33 (.I(net33),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output34 (.I(net34),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output35 (.I(net35),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output36 (.I(net36),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output37 (.I(net37),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output38 (.I(net38),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output39 (.I(net39),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output40 (.I(net40),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output41 (.I(net41),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output42 (.I(net42),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output43 (.I(net43),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output44 (.I(net44),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output45 (.I(net45),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output46 (.I(net46),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output47 (.I(net47),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output48 (.I(net48),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output49 (.I(net49),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output50 (.I(net50),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output51 (.I(net51),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output52 (.I(net52),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output53 (.I(net53),
    .Z(N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output54 (.I(net54),
    .Z(N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output55 (.I(net55),
    .Z(N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output56 (.I(net56),
    .Z(N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output57 (.I(net57),
    .Z(N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output58 (.I(net58),
    .Z(N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output59 (.I(net59),
    .Z(N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output60 (.I(net60),
    .Z(N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output61 (.I(net61),
    .Z(N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output62 (.I(net62),
    .Z(N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output63 (.I(net63),
    .Z(N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output64 (.I(net64),
    .Z(N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output65 (.I(net65),
    .Z(N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output66 (.I(net66),
    .Z(N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output67 (.I(net67),
    .Z(N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output68 (.I(net68),
    .Z(N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output69 (.I(net69),
    .Z(N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output70 (.I(net70),
    .Z(N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output71 (.I(net71),
    .Z(N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output72 (.I(net72),
    .Z(N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output73 (.I(net73),
    .Z(N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output74 (.I(net74),
    .Z(N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output75 (.I(net75),
    .Z(N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output76 (.I(net76),
    .Z(N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output77 (.I(net77),
    .Z(N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output78 (.I(net78),
    .Z(N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output79 (.I(net79),
    .Z(N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output80 (.I(net80),
    .Z(N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output81 (.I(net81),
    .Z(N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output82 (.I(net82),
    .Z(N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output83 (.I(net83),
    .Z(N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output84 (.I(net84),
    .Z(N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output85 (.I(net85),
    .Z(N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output86 (.I(net86),
    .Z(N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output87 (.I(net87),
    .Z(N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output88 (.I(net88),
    .Z(N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output89 (.I(net89),
    .Z(NN4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output90 (.I(net90),
    .Z(NN4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output91 (.I(net91),
    .Z(NN4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output92 (.I(net92),
    .Z(NN4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output93 (.I(net93),
    .Z(NN4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output94 (.I(net94),
    .Z(NN4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output95 (.I(net95),
    .Z(NN4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output96 (.I(net96),
    .Z(NN4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output97 (.I(net97),
    .Z(NN4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output98 (.I(net98),
    .Z(NN4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output99 (.I(net99),
    .Z(NN4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output100 (.I(net100),
    .Z(NN4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output101 (.I(net101),
    .Z(NN4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output102 (.I(net102),
    .Z(NN4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output103 (.I(net103),
    .Z(NN4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output104 (.I(net104),
    .Z(NN4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_560 ();
endmodule
