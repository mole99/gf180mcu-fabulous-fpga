magic
tech gf180mcuD
magscale 1 5
timestamp 1764323744
<< metal1 >>
rect 336 6677 31864 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 22233 6677
rect 22259 6651 22285 6677
rect 22311 6651 22337 6677
rect 22363 6651 31864 6677
rect 336 6634 31864 6651
rect 1863 6593 1889 6599
rect 1863 6561 1889 6567
rect 2983 6593 3009 6599
rect 2983 6561 3009 6567
rect 3767 6593 3793 6599
rect 3767 6561 3793 6567
rect 4887 6593 4913 6599
rect 4887 6561 4913 6567
rect 5671 6593 5697 6599
rect 5671 6561 5697 6567
rect 8695 6593 8721 6599
rect 8695 6561 8721 6567
rect 9479 6593 9505 6599
rect 9479 6561 9505 6567
rect 10599 6593 10625 6599
rect 10599 6561 10625 6567
rect 11383 6593 11409 6599
rect 11383 6561 11409 6567
rect 12503 6593 12529 6599
rect 12503 6561 12529 6567
rect 13287 6593 13313 6599
rect 26055 6593 26081 6599
rect 25433 6567 25439 6593
rect 25465 6567 25471 6593
rect 13287 6561 13313 6567
rect 26055 6561 26081 6567
rect 27455 6593 27481 6599
rect 27455 6561 27481 6567
rect 28239 6593 28265 6599
rect 28239 6561 28265 6567
rect 31263 6593 31289 6599
rect 31263 6561 31289 6567
rect 30249 6511 30255 6537
rect 30281 6511 30287 6537
rect 25607 6481 25633 6487
rect 849 6455 855 6481
rect 881 6455 887 6481
rect 2137 6455 2143 6481
rect 2169 6455 2175 6481
rect 3257 6455 3263 6481
rect 3289 6455 3295 6481
rect 4041 6455 4047 6481
rect 4073 6455 4079 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 5945 6455 5951 6481
rect 5977 6455 5983 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 7849 6455 7855 6481
rect 7881 6455 7887 6481
rect 8913 6455 8919 6481
rect 8945 6455 8951 6481
rect 9753 6455 9759 6481
rect 9785 6455 9791 6481
rect 10817 6455 10823 6481
rect 10849 6455 10855 6481
rect 11657 6455 11663 6481
rect 11689 6455 11695 6481
rect 12777 6455 12783 6481
rect 12809 6455 12815 6481
rect 13561 6455 13567 6481
rect 13593 6455 13599 6481
rect 14457 6455 14463 6481
rect 14489 6455 14495 6481
rect 25769 6455 25775 6481
rect 25801 6455 25807 6481
rect 27169 6455 27175 6481
rect 27201 6455 27207 6481
rect 27953 6455 27959 6481
rect 27985 6455 27991 6481
rect 29073 6455 29079 6481
rect 29105 6455 29111 6481
rect 29857 6455 29863 6481
rect 29889 6455 29895 6481
rect 30977 6455 30983 6481
rect 31009 6455 31015 6481
rect 25607 6449 25633 6455
rect 1247 6425 1273 6431
rect 1247 6393 1273 6399
rect 6959 6425 6985 6431
rect 13959 6425 13985 6431
rect 7401 6399 7407 6425
rect 7433 6399 7439 6425
rect 29409 6399 29415 6425
rect 29441 6399 29447 6425
rect 6959 6393 6985 6399
rect 13959 6393 13985 6399
rect 336 6285 31864 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 21903 6285
rect 21929 6259 21955 6285
rect 21981 6259 22007 6285
rect 22033 6259 31864 6285
rect 336 6242 31864 6259
rect 3487 6201 3513 6207
rect 3487 6169 3513 6175
rect 4271 6201 4297 6207
rect 4271 6169 4297 6175
rect 5839 6201 5865 6207
rect 5839 6169 5865 6175
rect 8191 6201 8217 6207
rect 8191 6169 8217 6175
rect 8975 6201 9001 6207
rect 8975 6169 9001 6175
rect 9927 6201 9953 6207
rect 9927 6169 9953 6175
rect 11215 6201 11241 6207
rect 11215 6169 11241 6175
rect 11999 6201 12025 6207
rect 11999 6169 12025 6175
rect 12559 6201 12585 6207
rect 12559 6169 12585 6175
rect 26279 6201 26305 6207
rect 26279 6169 26305 6175
rect 27063 6201 27089 6207
rect 27063 6169 27089 6175
rect 27847 6201 27873 6207
rect 27847 6169 27873 6175
rect 28631 6201 28657 6207
rect 28631 6169 28657 6175
rect 14911 6145 14937 6151
rect 1801 6119 1807 6145
rect 1833 6119 1839 6145
rect 4993 6119 4999 6145
rect 5025 6119 5031 6145
rect 7457 6119 7463 6145
rect 7489 6119 7495 6145
rect 13449 6119 13455 6145
rect 13481 6119 13487 6145
rect 14911 6113 14937 6119
rect 15191 6145 15217 6151
rect 30305 6119 30311 6145
rect 30337 6119 30343 6145
rect 31089 6119 31095 6145
rect 31121 6119 31127 6145
rect 15191 6113 15217 6119
rect 15471 6089 15497 6095
rect 20679 6089 20705 6095
rect 5329 6063 5335 6089
rect 5361 6063 5367 6089
rect 9193 6063 9199 6089
rect 9225 6063 9231 6089
rect 9417 6063 9423 6089
rect 9449 6063 9455 6089
rect 12161 6063 12167 6089
rect 12193 6063 12199 6089
rect 14681 6063 14687 6089
rect 14713 6063 14719 6089
rect 17649 6063 17655 6089
rect 17681 6063 17687 6089
rect 26049 6063 26055 6089
rect 26081 6063 26087 6089
rect 26777 6063 26783 6089
rect 26809 6063 26815 6089
rect 15471 6057 15497 6063
rect 20679 6057 20705 6063
rect 17879 6033 17905 6039
rect 2193 6007 2199 6033
rect 2225 6007 2231 6033
rect 3761 6007 3767 6033
rect 3793 6007 3799 6033
rect 4545 6007 4551 6033
rect 4577 6007 4583 6033
rect 6113 6007 6119 6033
rect 6145 6007 6151 6033
rect 7065 6007 7071 6033
rect 7097 6007 7103 6033
rect 8465 6007 8471 6033
rect 8497 6007 8503 6033
rect 11489 6007 11495 6033
rect 11521 6007 11527 6033
rect 13057 6007 13063 6033
rect 13089 6007 13095 6033
rect 13841 6007 13847 6033
rect 13873 6007 13879 6033
rect 17879 6001 17905 6007
rect 21799 6033 21825 6039
rect 29583 6033 29609 6039
rect 27561 6007 27567 6033
rect 27593 6007 27599 6033
rect 28345 6007 28351 6033
rect 28377 6007 28383 6033
rect 29913 6007 29919 6033
rect 29945 6007 29951 6033
rect 30697 6007 30703 6033
rect 30729 6007 30735 6033
rect 21799 6001 21825 6007
rect 29583 6001 29609 6007
rect 20399 5977 20425 5983
rect 20399 5945 20425 5951
rect 21519 5977 21545 5983
rect 21519 5945 21545 5951
rect 29303 5977 29329 5983
rect 29303 5945 29329 5951
rect 336 5893 31864 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 22233 5893
rect 22259 5867 22285 5893
rect 22311 5867 22337 5893
rect 22363 5867 31864 5893
rect 336 5850 31864 5867
rect 2311 5809 2337 5815
rect 2311 5777 2337 5783
rect 3879 5809 3905 5815
rect 3879 5777 3905 5783
rect 5447 5809 5473 5815
rect 5447 5777 5473 5783
rect 9311 5809 9337 5815
rect 9311 5777 9337 5783
rect 10151 5809 10177 5815
rect 10151 5777 10177 5783
rect 14015 5809 14041 5815
rect 14015 5777 14041 5783
rect 26503 5809 26529 5815
rect 26503 5777 26529 5783
rect 27287 5809 27313 5815
rect 27287 5777 27313 5783
rect 28239 5809 28265 5815
rect 28239 5777 28265 5783
rect 29023 5809 29049 5815
rect 29023 5777 29049 5783
rect 29807 5809 29833 5815
rect 29807 5777 29833 5783
rect 30591 5809 30617 5815
rect 30591 5777 30617 5783
rect 23367 5697 23393 5703
rect 31095 5697 31121 5703
rect 1129 5671 1135 5697
rect 1161 5671 1167 5697
rect 2585 5671 2591 5697
rect 2617 5671 2623 5697
rect 3313 5671 3319 5697
rect 3345 5671 3351 5697
rect 4153 5671 4159 5697
rect 4185 5671 4191 5697
rect 5721 5671 5727 5697
rect 5753 5671 5759 5697
rect 6505 5671 6511 5697
rect 6537 5671 6543 5697
rect 6729 5671 6735 5697
rect 6761 5671 6767 5697
rect 7457 5671 7463 5697
rect 7489 5671 7495 5697
rect 9025 5671 9031 5697
rect 9057 5671 9063 5697
rect 10313 5671 10319 5697
rect 10345 5671 10351 5697
rect 11209 5671 11215 5697
rect 11241 5671 11247 5697
rect 11993 5671 11999 5697
rect 12025 5671 12031 5697
rect 13617 5671 13623 5697
rect 13649 5671 13655 5697
rect 26217 5671 26223 5697
rect 26249 5671 26255 5697
rect 27001 5671 27007 5697
rect 27033 5671 27039 5697
rect 28009 5671 28015 5697
rect 28041 5671 28047 5697
rect 28737 5671 28743 5697
rect 28769 5671 28775 5697
rect 29521 5671 29527 5697
rect 29553 5671 29559 5697
rect 30361 5671 30367 5697
rect 30393 5671 30399 5697
rect 23367 5665 23393 5671
rect 31095 5665 31121 5671
rect 7183 5641 7209 5647
rect 961 5615 967 5641
rect 993 5615 999 5641
rect 3033 5615 3039 5641
rect 3065 5615 3071 5641
rect 6169 5615 6175 5641
rect 6201 5615 6207 5641
rect 7183 5609 7209 5615
rect 7967 5641 7993 5647
rect 7967 5609 7993 5615
rect 10711 5641 10737 5647
rect 13119 5641 13145 5647
rect 11545 5615 11551 5641
rect 11577 5615 11583 5641
rect 14233 5615 14239 5641
rect 14265 5615 14271 5641
rect 23137 5615 23143 5641
rect 23169 5615 23175 5641
rect 31313 5615 31319 5641
rect 31345 5615 31351 5641
rect 10711 5609 10737 5615
rect 13119 5609 13145 5615
rect 336 5501 31864 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 21903 5501
rect 21929 5475 21955 5501
rect 21981 5475 22007 5501
rect 22033 5475 31864 5501
rect 336 5458 31864 5475
rect 4831 5417 4857 5423
rect 4831 5385 4857 5391
rect 5615 5417 5641 5423
rect 5615 5385 5641 5391
rect 7183 5417 7209 5423
rect 7183 5385 7209 5391
rect 8135 5417 8161 5423
rect 8135 5385 8161 5391
rect 8919 5417 8945 5423
rect 8919 5385 8945 5391
rect 9535 5417 9561 5423
rect 9535 5385 9561 5391
rect 11103 5417 11129 5423
rect 11103 5385 11129 5391
rect 11999 5417 12025 5423
rect 11999 5385 12025 5391
rect 30759 5361 30785 5367
rect 3369 5335 3375 5361
rect 3401 5335 3407 5361
rect 4097 5335 4103 5361
rect 4129 5335 4135 5361
rect 28569 5335 28575 5361
rect 28601 5335 28607 5361
rect 29409 5335 29415 5361
rect 29441 5335 29447 5361
rect 30759 5329 30785 5335
rect 8633 5279 8639 5305
rect 8665 5279 8671 5305
rect 9977 5279 9983 5305
rect 10009 5279 10015 5305
rect 11601 5279 11607 5305
rect 11633 5279 11639 5305
rect 27673 5279 27679 5305
rect 27705 5279 27711 5305
rect 29017 5279 29023 5305
rect 29049 5279 29055 5305
rect 30305 5279 30311 5305
rect 30337 5279 30343 5305
rect 31089 5279 31095 5305
rect 31121 5279 31127 5305
rect 6791 5249 6817 5255
rect 10767 5249 10793 5255
rect 21799 5249 21825 5255
rect 3761 5223 3767 5249
rect 3793 5223 3799 5249
rect 4545 5223 4551 5249
rect 4577 5223 4583 5249
rect 5329 5223 5335 5249
rect 5361 5223 5367 5249
rect 6113 5223 6119 5249
rect 6145 5223 6151 5249
rect 7681 5223 7687 5249
rect 7713 5223 7719 5249
rect 7849 5223 7855 5249
rect 7881 5223 7887 5249
rect 12497 5223 12503 5249
rect 12529 5223 12535 5249
rect 28065 5223 28071 5249
rect 28097 5223 28103 5249
rect 28233 5223 28239 5249
rect 28265 5223 28271 5249
rect 31425 5223 31431 5249
rect 31457 5223 31463 5249
rect 6791 5217 6817 5223
rect 10767 5217 10793 5223
rect 21799 5217 21825 5223
rect 6511 5193 6537 5199
rect 6511 5161 6537 5167
rect 10487 5193 10513 5199
rect 10487 5161 10513 5167
rect 21519 5193 21545 5199
rect 21519 5161 21545 5167
rect 336 5109 31864 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 22233 5109
rect 22259 5083 22285 5109
rect 22311 5083 22337 5109
rect 22363 5083 31864 5109
rect 336 5066 31864 5083
rect 3879 5025 3905 5031
rect 3879 4993 3905 4999
rect 28961 4943 28967 4969
rect 28993 4943 28999 4969
rect 27959 4913 27985 4919
rect 5777 4887 5783 4913
rect 5809 4887 5815 4913
rect 7513 4887 7519 4913
rect 7545 4887 7551 4913
rect 28681 4887 28687 4913
rect 28713 4887 28719 4913
rect 29409 4887 29415 4913
rect 29441 4887 29447 4913
rect 29745 4887 29751 4913
rect 29777 4887 29783 4913
rect 30137 4887 30143 4913
rect 30169 4887 30175 4913
rect 30977 4887 30983 4913
rect 31009 4887 31015 4913
rect 27959 4881 27985 4887
rect 4159 4857 4185 4863
rect 4159 4825 4185 4831
rect 5279 4857 5305 4863
rect 5279 4825 5305 4831
rect 7071 4857 7097 4863
rect 7071 4825 7097 4831
rect 28239 4857 28265 4863
rect 28239 4825 28265 4831
rect 30647 4857 30673 4863
rect 31369 4831 31375 4857
rect 31401 4831 31407 4857
rect 30647 4825 30673 4831
rect 336 4717 31864 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 21903 4717
rect 21929 4691 21955 4717
rect 21981 4691 22007 4717
rect 22033 4691 31864 4717
rect 336 4674 31864 4691
rect 29359 4633 29385 4639
rect 29359 4601 29385 4607
rect 30759 4633 30785 4639
rect 30759 4601 30785 4607
rect 2759 4577 2785 4583
rect 1409 4551 1415 4577
rect 1441 4551 1447 4577
rect 2759 4545 2785 4551
rect 24095 4577 24121 4583
rect 26609 4551 26615 4577
rect 26641 4551 26647 4577
rect 28345 4551 28351 4577
rect 28377 4551 28383 4577
rect 28793 4551 28799 4577
rect 28825 4551 28831 4577
rect 24095 4545 24121 4551
rect 1639 4521 1665 4527
rect 14799 4521 14825 4527
rect 2529 4495 2535 4521
rect 2561 4495 2567 4521
rect 1639 4489 1665 4495
rect 14799 4489 14825 4495
rect 20511 4521 20537 4527
rect 20511 4489 20537 4495
rect 26391 4521 26417 4527
rect 26391 4489 26417 4495
rect 28127 4521 28153 4527
rect 29577 4495 29583 4521
rect 29609 4495 29615 4521
rect 31145 4495 31151 4521
rect 31177 4495 31183 4521
rect 28127 4489 28153 4495
rect 8919 4465 8945 4471
rect 8919 4433 8945 4439
rect 10823 4465 10849 4471
rect 10823 4433 10849 4439
rect 11103 4465 11129 4471
rect 11103 4433 11129 4439
rect 14519 4465 14545 4471
rect 14519 4433 14545 4439
rect 20231 4465 20257 4471
rect 30249 4439 30255 4465
rect 30281 4439 30287 4465
rect 31425 4439 31431 4465
rect 31457 4439 31463 4465
rect 20231 4433 20257 4439
rect 8639 4409 8665 4415
rect 8639 4377 8665 4383
rect 23815 4409 23841 4415
rect 23815 4377 23841 4383
rect 28575 4409 28601 4415
rect 28575 4377 28601 4383
rect 336 4325 31864 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 22233 4325
rect 22259 4299 22285 4325
rect 22311 4299 22337 4325
rect 22363 4299 31864 4325
rect 336 4282 31864 4299
rect 2367 4241 2393 4247
rect 2367 4209 2393 4215
rect 28463 4241 28489 4247
rect 28463 4209 28489 4215
rect 28239 4185 28265 4191
rect 28239 4153 28265 4159
rect 28743 4185 28769 4191
rect 28743 4153 28769 4159
rect 28911 4185 28937 4191
rect 30529 4159 30535 4185
rect 30561 4159 30567 4185
rect 28911 4153 28937 4159
rect 2647 4129 2673 4135
rect 2647 4097 2673 4103
rect 6231 4129 6257 4135
rect 6231 4097 6257 4103
rect 21967 4129 21993 4135
rect 21967 4097 21993 4103
rect 27959 4129 27985 4135
rect 27959 4097 27985 4103
rect 29191 4129 29217 4135
rect 29353 4103 29359 4129
rect 29385 4103 29391 4129
rect 30193 4103 30199 4129
rect 30225 4103 30231 4129
rect 30921 4103 30927 4129
rect 30953 4103 30959 4129
rect 29191 4097 29217 4103
rect 6511 4073 6537 4079
rect 29863 4073 29889 4079
rect 21737 4047 21743 4073
rect 21769 4047 21775 4073
rect 6511 4041 6537 4047
rect 29863 4041 29889 4047
rect 31431 4017 31457 4023
rect 31431 3985 31457 3991
rect 336 3933 31864 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 21903 3933
rect 21929 3907 21955 3933
rect 21981 3907 22007 3933
rect 22033 3907 31864 3933
rect 336 3890 31864 3907
rect 31543 3849 31569 3855
rect 31543 3817 31569 3823
rect 20847 3793 20873 3799
rect 30759 3793 30785 3799
rect 7401 3767 7407 3793
rect 7433 3767 7439 3793
rect 29577 3767 29583 3793
rect 29609 3767 29615 3793
rect 20847 3761 20873 3767
rect 30759 3761 30785 3767
rect 7631 3737 7657 3743
rect 7631 3705 7657 3711
rect 17431 3737 17457 3743
rect 17431 3705 17457 3711
rect 21127 3737 21153 3743
rect 21127 3705 21153 3711
rect 28911 3737 28937 3743
rect 29409 3711 29415 3737
rect 29441 3711 29447 3737
rect 30249 3711 30255 3737
rect 30281 3711 30287 3737
rect 31145 3711 31151 3737
rect 31177 3711 31183 3737
rect 28911 3705 28937 3711
rect 17711 3681 17737 3687
rect 17711 3649 17737 3655
rect 29191 3681 29217 3687
rect 29191 3649 29217 3655
rect 336 3541 31864 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 22233 3541
rect 22259 3515 22285 3541
rect 22311 3515 22337 3541
rect 22363 3515 31864 3541
rect 336 3498 31864 3515
rect 15359 3457 15385 3463
rect 15359 3425 15385 3431
rect 8751 3345 8777 3351
rect 18439 3345 18465 3351
rect 25215 3345 25241 3351
rect 8969 3319 8975 3345
rect 9001 3319 9007 3345
rect 23529 3319 23535 3345
rect 23561 3319 23567 3345
rect 8751 3313 8777 3319
rect 18439 3313 18465 3319
rect 25215 3313 25241 3319
rect 25495 3345 25521 3351
rect 25495 3313 25521 3319
rect 29247 3345 29273 3351
rect 29247 3313 29273 3319
rect 29695 3345 29721 3351
rect 29695 3313 29721 3319
rect 29975 3345 30001 3351
rect 30137 3319 30143 3345
rect 30169 3319 30175 3345
rect 31033 3319 31039 3345
rect 31065 3319 31071 3345
rect 29975 3313 30001 3319
rect 18159 3289 18185 3295
rect 31431 3289 31457 3295
rect 15129 3263 15135 3289
rect 15161 3263 15167 3289
rect 23697 3263 23703 3289
rect 23729 3263 23735 3289
rect 29465 3263 29471 3289
rect 29497 3263 29503 3289
rect 18159 3257 18185 3263
rect 31431 3257 31457 3263
rect 30647 3233 30673 3239
rect 30647 3201 30673 3207
rect 336 3149 31864 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 21903 3149
rect 21929 3123 21955 3149
rect 21981 3123 22007 3149
rect 22033 3123 31864 3149
rect 336 3106 31864 3123
rect 30759 3065 30785 3071
rect 30759 3033 30785 3039
rect 31543 3065 31569 3071
rect 31543 3033 31569 3039
rect 4047 3009 4073 3015
rect 1017 2983 1023 3009
rect 1049 2983 1055 3009
rect 4047 2977 4073 2983
rect 13287 3009 13313 3015
rect 13287 2977 13313 2983
rect 14799 3009 14825 3015
rect 14799 2977 14825 2983
rect 28967 3009 28993 3015
rect 28967 2977 28993 2983
rect 29639 3009 29665 3015
rect 29639 2977 29665 2983
rect 4327 2953 4353 2959
rect 4327 2921 4353 2927
rect 13567 2953 13593 2959
rect 29409 2927 29415 2953
rect 29441 2927 29447 2953
rect 30249 2927 30255 2953
rect 30281 2927 30287 2953
rect 31089 2927 31095 2953
rect 31121 2927 31127 2953
rect 13567 2921 13593 2927
rect 15079 2897 15105 2903
rect 15079 2865 15105 2871
rect 22079 2897 22105 2903
rect 22079 2865 22105 2871
rect 22359 2897 22385 2903
rect 22359 2865 22385 2871
rect 1247 2841 1273 2847
rect 1247 2809 1273 2815
rect 28687 2841 28713 2847
rect 28687 2809 28713 2815
rect 336 2757 31864 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 22233 2757
rect 22259 2731 22285 2757
rect 22311 2731 22337 2757
rect 22363 2731 31864 2757
rect 336 2714 31864 2731
rect 1247 2673 1273 2679
rect 1247 2641 1273 2647
rect 8639 2673 8665 2679
rect 8639 2641 8665 2647
rect 10935 2673 10961 2679
rect 10935 2641 10961 2647
rect 12559 2673 12585 2679
rect 12559 2641 12585 2647
rect 20175 2673 20201 2679
rect 20175 2641 20201 2647
rect 21183 2673 21209 2679
rect 21183 2641 21209 2647
rect 29695 2673 29721 2679
rect 29695 2641 29721 2647
rect 967 2617 993 2623
rect 967 2585 993 2591
rect 9367 2617 9393 2623
rect 9367 2585 9393 2591
rect 9647 2617 9673 2623
rect 9647 2585 9673 2591
rect 10655 2617 10681 2623
rect 10655 2585 10681 2591
rect 12279 2617 12305 2623
rect 12279 2585 12305 2591
rect 14519 2617 14545 2623
rect 14519 2585 14545 2591
rect 20455 2617 20481 2623
rect 20455 2585 20481 2591
rect 20903 2617 20929 2623
rect 20903 2585 20929 2591
rect 21743 2617 21769 2623
rect 21743 2585 21769 2591
rect 25439 2617 25465 2623
rect 25439 2585 25465 2591
rect 28631 2617 28657 2623
rect 28631 2585 28657 2591
rect 29191 2617 29217 2623
rect 30137 2591 30143 2617
rect 30169 2591 30175 2617
rect 30529 2591 30535 2617
rect 30561 2591 30567 2617
rect 31313 2591 31319 2617
rect 31345 2591 31351 2617
rect 29191 2585 29217 2591
rect 14799 2561 14825 2567
rect 14799 2529 14825 2535
rect 21463 2561 21489 2567
rect 28351 2561 28377 2567
rect 25209 2535 25215 2561
rect 25241 2535 25247 2561
rect 21463 2529 21489 2535
rect 28351 2529 28377 2535
rect 28911 2561 28937 2567
rect 28911 2529 28937 2535
rect 29975 2561 30001 2567
rect 30921 2535 30927 2561
rect 30953 2535 30959 2561
rect 29975 2529 30001 2535
rect 8409 2479 8415 2505
rect 8441 2479 8447 2505
rect 336 2365 31864 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 21903 2365
rect 21929 2339 21955 2365
rect 21981 2339 22007 2365
rect 22033 2339 31864 2365
rect 336 2322 31864 2339
rect 31543 2281 31569 2287
rect 31543 2249 31569 2255
rect 8247 2225 8273 2231
rect 961 2199 967 2225
rect 993 2199 999 2225
rect 27841 2199 27847 2225
rect 27873 2199 27879 2225
rect 8247 2193 8273 2199
rect 21295 2169 21321 2175
rect 21295 2137 21321 2143
rect 24543 2169 24569 2175
rect 31089 2143 31095 2169
rect 31121 2143 31127 2169
rect 24543 2137 24569 2143
rect 21015 2113 21041 2119
rect 21015 2081 21041 2087
rect 24263 2113 24289 2119
rect 30249 2087 30255 2113
rect 30281 2087 30287 2113
rect 30641 2087 30647 2113
rect 30673 2087 30679 2113
rect 24263 2081 24289 2087
rect 1191 2057 1217 2063
rect 1191 2025 1217 2031
rect 8527 2057 8553 2063
rect 8527 2025 8553 2031
rect 28071 2057 28097 2063
rect 28071 2025 28097 2031
rect 336 1973 31864 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 22233 1973
rect 22259 1947 22285 1973
rect 22311 1947 22337 1973
rect 22363 1947 31864 1973
rect 336 1930 31864 1947
rect 2591 1889 2617 1895
rect 2591 1857 2617 1863
rect 11999 1889 12025 1895
rect 11999 1857 12025 1863
rect 20399 1889 20425 1895
rect 20399 1857 20425 1863
rect 25271 1889 25297 1895
rect 25271 1857 25297 1863
rect 2871 1833 2897 1839
rect 2871 1801 2897 1807
rect 22191 1833 22217 1839
rect 22191 1801 22217 1807
rect 22471 1833 22497 1839
rect 22471 1801 22497 1807
rect 23255 1833 23281 1839
rect 23255 1801 23281 1807
rect 24991 1833 25017 1839
rect 24991 1801 25017 1807
rect 1303 1777 1329 1783
rect 29695 1777 29721 1783
rect 8577 1751 8583 1777
rect 8609 1751 8615 1777
rect 23473 1751 23479 1777
rect 23505 1751 23511 1777
rect 1303 1745 1329 1751
rect 29695 1745 29721 1751
rect 29975 1777 30001 1783
rect 30137 1751 30143 1777
rect 30169 1751 30175 1777
rect 30921 1751 30927 1777
rect 30953 1751 30959 1777
rect 29975 1745 30001 1751
rect 30647 1721 30673 1727
rect 1073 1695 1079 1721
rect 1105 1695 1111 1721
rect 8409 1695 8415 1721
rect 8441 1695 8447 1721
rect 11769 1695 11775 1721
rect 11801 1695 11807 1721
rect 20169 1695 20175 1721
rect 20201 1695 20207 1721
rect 30647 1689 30673 1695
rect 31431 1721 31457 1727
rect 31431 1689 31457 1695
rect 336 1581 31864 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 21903 1581
rect 21929 1555 21955 1581
rect 21981 1555 22007 1581
rect 22033 1555 31864 1581
rect 336 1538 31864 1555
rect 31543 1497 31569 1503
rect 31543 1465 31569 1471
rect 26049 1415 26055 1441
rect 26081 1415 26087 1441
rect 29639 1385 29665 1391
rect 29409 1359 29415 1385
rect 29441 1359 29447 1385
rect 31089 1359 31095 1385
rect 31121 1359 31127 1385
rect 29639 1353 29665 1359
rect 29191 1329 29217 1335
rect 30249 1303 30255 1329
rect 30281 1303 30287 1329
rect 30641 1303 30647 1329
rect 30673 1303 30679 1329
rect 29191 1297 29217 1303
rect 26279 1273 26305 1279
rect 26279 1241 26305 1247
rect 28911 1273 28937 1279
rect 28911 1241 28937 1247
rect 336 1189 31864 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 22233 1189
rect 22259 1163 22285 1189
rect 22311 1163 22337 1189
rect 22363 1163 31864 1189
rect 336 1146 31864 1163
rect 6231 1105 6257 1111
rect 6231 1073 6257 1079
rect 7631 1105 7657 1111
rect 7631 1073 7657 1079
rect 8079 1105 8105 1111
rect 8079 1073 8105 1079
rect 11439 1105 11465 1111
rect 16479 1105 16505 1111
rect 15409 1079 15415 1105
rect 15441 1079 15447 1105
rect 11439 1073 11465 1079
rect 16479 1073 16505 1079
rect 17935 1105 17961 1111
rect 17935 1073 17961 1079
rect 18439 1105 18465 1111
rect 18439 1073 18465 1079
rect 19727 1105 19753 1111
rect 19727 1073 19753 1079
rect 20903 1105 20929 1111
rect 20903 1073 20929 1079
rect 21351 1105 21377 1111
rect 21351 1073 21377 1079
rect 21799 1105 21825 1111
rect 21799 1073 21825 1079
rect 22919 1105 22945 1111
rect 22919 1073 22945 1079
rect 29695 1105 29721 1111
rect 29695 1073 29721 1079
rect 967 1049 993 1055
rect 967 1017 993 1023
rect 4831 1049 4857 1055
rect 4831 1017 4857 1023
rect 7351 1049 7377 1055
rect 7351 1017 7377 1023
rect 7799 1049 7825 1055
rect 7799 1017 7825 1023
rect 17655 1049 17681 1055
rect 17655 1017 17681 1023
rect 18159 1049 18185 1055
rect 18159 1017 18185 1023
rect 18775 1049 18801 1055
rect 18775 1017 18801 1023
rect 19447 1049 19473 1055
rect 19447 1017 19473 1023
rect 20623 1049 20649 1055
rect 20623 1017 20649 1023
rect 21071 1049 21097 1055
rect 21071 1017 21097 1023
rect 21519 1049 21545 1055
rect 21519 1017 21545 1023
rect 24319 1049 24345 1055
rect 24319 1017 24345 1023
rect 24879 1049 24905 1055
rect 24879 1017 24905 1023
rect 25439 1049 25465 1055
rect 25439 1017 25465 1023
rect 28799 1049 28825 1055
rect 28799 1017 28825 1023
rect 29247 1049 29273 1055
rect 30137 1023 30143 1049
rect 30169 1023 30175 1049
rect 29247 1017 29273 1023
rect 1247 993 1273 999
rect 1247 961 1273 967
rect 4551 993 4577 999
rect 15247 993 15273 999
rect 5049 967 5055 993
rect 5081 967 5087 993
rect 4551 961 4577 967
rect 15247 961 15273 967
rect 19055 993 19081 999
rect 19055 961 19081 967
rect 24039 993 24065 999
rect 24039 961 24065 967
rect 24599 993 24625 999
rect 28967 993 28993 999
rect 25209 967 25215 993
rect 25241 967 25247 993
rect 28569 967 28575 993
rect 28601 967 28607 993
rect 24599 961 24625 967
rect 28967 961 28993 967
rect 29975 993 30001 999
rect 30921 967 30927 993
rect 30953 967 30959 993
rect 29975 961 30001 967
rect 5279 937 5305 943
rect 5279 905 5305 911
rect 6511 937 6537 943
rect 6511 905 6537 911
rect 11159 937 11185 943
rect 11159 905 11185 911
rect 16199 937 16225 943
rect 31431 937 31457 943
rect 22689 911 22695 937
rect 22721 911 22727 937
rect 16199 905 16225 911
rect 31431 905 31457 911
rect 30647 881 30673 887
rect 30647 849 30673 855
rect 336 797 31864 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 21903 797
rect 21929 771 21955 797
rect 21981 771 22007 797
rect 22033 771 31864 797
rect 336 754 31864 771
rect 31543 713 31569 719
rect 31543 681 31569 687
rect 911 657 937 663
rect 911 625 937 631
rect 29807 657 29833 663
rect 29807 625 29833 631
rect 30591 657 30617 663
rect 30591 625 30617 631
rect 5049 575 5055 601
rect 5081 575 5087 601
rect 30081 575 30087 601
rect 30113 575 30119 601
rect 31089 575 31095 601
rect 31121 575 31127 601
rect 5279 545 5305 551
rect 29297 519 29303 545
rect 29329 519 29335 545
rect 5279 513 5305 519
rect 1191 489 1217 495
rect 1191 457 1217 463
rect 336 405 31864 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 22233 405
rect 22259 379 22285 405
rect 22311 379 22337 405
rect 22363 379 31864 405
rect 336 362 31864 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 22233 6651 22259 6677
rect 22285 6651 22311 6677
rect 22337 6651 22363 6677
rect 1863 6567 1889 6593
rect 2983 6567 3009 6593
rect 3767 6567 3793 6593
rect 4887 6567 4913 6593
rect 5671 6567 5697 6593
rect 8695 6567 8721 6593
rect 9479 6567 9505 6593
rect 10599 6567 10625 6593
rect 11383 6567 11409 6593
rect 12503 6567 12529 6593
rect 13287 6567 13313 6593
rect 25439 6567 25465 6593
rect 26055 6567 26081 6593
rect 27455 6567 27481 6593
rect 28239 6567 28265 6593
rect 31263 6567 31289 6593
rect 30255 6511 30281 6537
rect 855 6455 881 6481
rect 2143 6455 2169 6481
rect 3263 6455 3289 6481
rect 4047 6455 4073 6481
rect 5167 6455 5193 6481
rect 5951 6455 5977 6481
rect 6455 6455 6481 6481
rect 7855 6455 7881 6481
rect 8919 6455 8945 6481
rect 9759 6455 9785 6481
rect 10823 6455 10849 6481
rect 11663 6455 11689 6481
rect 12783 6455 12809 6481
rect 13567 6455 13593 6481
rect 14463 6455 14489 6481
rect 25607 6455 25633 6481
rect 25775 6455 25801 6481
rect 27175 6455 27201 6481
rect 27959 6455 27985 6481
rect 29079 6455 29105 6481
rect 29863 6455 29889 6481
rect 30983 6455 31009 6481
rect 1247 6399 1273 6425
rect 6959 6399 6985 6425
rect 7407 6399 7433 6425
rect 13959 6399 13985 6425
rect 29415 6399 29441 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 21903 6259 21929 6285
rect 21955 6259 21981 6285
rect 22007 6259 22033 6285
rect 3487 6175 3513 6201
rect 4271 6175 4297 6201
rect 5839 6175 5865 6201
rect 8191 6175 8217 6201
rect 8975 6175 9001 6201
rect 9927 6175 9953 6201
rect 11215 6175 11241 6201
rect 11999 6175 12025 6201
rect 12559 6175 12585 6201
rect 26279 6175 26305 6201
rect 27063 6175 27089 6201
rect 27847 6175 27873 6201
rect 28631 6175 28657 6201
rect 1807 6119 1833 6145
rect 4999 6119 5025 6145
rect 7463 6119 7489 6145
rect 13455 6119 13481 6145
rect 14911 6119 14937 6145
rect 15191 6119 15217 6145
rect 30311 6119 30337 6145
rect 31095 6119 31121 6145
rect 5335 6063 5361 6089
rect 9199 6063 9225 6089
rect 9423 6063 9449 6089
rect 12167 6063 12193 6089
rect 14687 6063 14713 6089
rect 15471 6063 15497 6089
rect 17655 6063 17681 6089
rect 20679 6063 20705 6089
rect 26055 6063 26081 6089
rect 26783 6063 26809 6089
rect 2199 6007 2225 6033
rect 3767 6007 3793 6033
rect 4551 6007 4577 6033
rect 6119 6007 6145 6033
rect 7071 6007 7097 6033
rect 8471 6007 8497 6033
rect 11495 6007 11521 6033
rect 13063 6007 13089 6033
rect 13847 6007 13873 6033
rect 17879 6007 17905 6033
rect 21799 6007 21825 6033
rect 27567 6007 27593 6033
rect 28351 6007 28377 6033
rect 29583 6007 29609 6033
rect 29919 6007 29945 6033
rect 30703 6007 30729 6033
rect 20399 5951 20425 5977
rect 21519 5951 21545 5977
rect 29303 5951 29329 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 22233 5867 22259 5893
rect 22285 5867 22311 5893
rect 22337 5867 22363 5893
rect 2311 5783 2337 5809
rect 3879 5783 3905 5809
rect 5447 5783 5473 5809
rect 9311 5783 9337 5809
rect 10151 5783 10177 5809
rect 14015 5783 14041 5809
rect 26503 5783 26529 5809
rect 27287 5783 27313 5809
rect 28239 5783 28265 5809
rect 29023 5783 29049 5809
rect 29807 5783 29833 5809
rect 30591 5783 30617 5809
rect 1135 5671 1161 5697
rect 2591 5671 2617 5697
rect 3319 5671 3345 5697
rect 4159 5671 4185 5697
rect 5727 5671 5753 5697
rect 6511 5671 6537 5697
rect 6735 5671 6761 5697
rect 7463 5671 7489 5697
rect 9031 5671 9057 5697
rect 10319 5671 10345 5697
rect 11215 5671 11241 5697
rect 11999 5671 12025 5697
rect 13623 5671 13649 5697
rect 23367 5671 23393 5697
rect 26223 5671 26249 5697
rect 27007 5671 27033 5697
rect 28015 5671 28041 5697
rect 28743 5671 28769 5697
rect 29527 5671 29553 5697
rect 30367 5671 30393 5697
rect 31095 5671 31121 5697
rect 967 5615 993 5641
rect 3039 5615 3065 5641
rect 6175 5615 6201 5641
rect 7183 5615 7209 5641
rect 7967 5615 7993 5641
rect 10711 5615 10737 5641
rect 11551 5615 11577 5641
rect 13119 5615 13145 5641
rect 14239 5615 14265 5641
rect 23143 5615 23169 5641
rect 31319 5615 31345 5641
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 21903 5475 21929 5501
rect 21955 5475 21981 5501
rect 22007 5475 22033 5501
rect 4831 5391 4857 5417
rect 5615 5391 5641 5417
rect 7183 5391 7209 5417
rect 8135 5391 8161 5417
rect 8919 5391 8945 5417
rect 9535 5391 9561 5417
rect 11103 5391 11129 5417
rect 11999 5391 12025 5417
rect 3375 5335 3401 5361
rect 4103 5335 4129 5361
rect 28575 5335 28601 5361
rect 29415 5335 29441 5361
rect 30759 5335 30785 5361
rect 8639 5279 8665 5305
rect 9983 5279 10009 5305
rect 11607 5279 11633 5305
rect 27679 5279 27705 5305
rect 29023 5279 29049 5305
rect 30311 5279 30337 5305
rect 31095 5279 31121 5305
rect 3767 5223 3793 5249
rect 4551 5223 4577 5249
rect 5335 5223 5361 5249
rect 6119 5223 6145 5249
rect 6791 5223 6817 5249
rect 7687 5223 7713 5249
rect 7855 5223 7881 5249
rect 10767 5223 10793 5249
rect 12503 5223 12529 5249
rect 21799 5223 21825 5249
rect 28071 5223 28097 5249
rect 28239 5223 28265 5249
rect 31431 5223 31457 5249
rect 6511 5167 6537 5193
rect 10487 5167 10513 5193
rect 21519 5167 21545 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 22233 5083 22259 5109
rect 22285 5083 22311 5109
rect 22337 5083 22363 5109
rect 3879 4999 3905 5025
rect 28967 4943 28993 4969
rect 5783 4887 5809 4913
rect 7519 4887 7545 4913
rect 27959 4887 27985 4913
rect 28687 4887 28713 4913
rect 29415 4887 29441 4913
rect 29751 4887 29777 4913
rect 30143 4887 30169 4913
rect 30983 4887 31009 4913
rect 4159 4831 4185 4857
rect 5279 4831 5305 4857
rect 7071 4831 7097 4857
rect 28239 4831 28265 4857
rect 30647 4831 30673 4857
rect 31375 4831 31401 4857
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 21903 4691 21929 4717
rect 21955 4691 21981 4717
rect 22007 4691 22033 4717
rect 29359 4607 29385 4633
rect 30759 4607 30785 4633
rect 1415 4551 1441 4577
rect 2759 4551 2785 4577
rect 24095 4551 24121 4577
rect 26615 4551 26641 4577
rect 28351 4551 28377 4577
rect 28799 4551 28825 4577
rect 1639 4495 1665 4521
rect 2535 4495 2561 4521
rect 14799 4495 14825 4521
rect 20511 4495 20537 4521
rect 26391 4495 26417 4521
rect 28127 4495 28153 4521
rect 29583 4495 29609 4521
rect 31151 4495 31177 4521
rect 8919 4439 8945 4465
rect 10823 4439 10849 4465
rect 11103 4439 11129 4465
rect 14519 4439 14545 4465
rect 20231 4439 20257 4465
rect 30255 4439 30281 4465
rect 31431 4439 31457 4465
rect 8639 4383 8665 4409
rect 23815 4383 23841 4409
rect 28575 4383 28601 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 22233 4299 22259 4325
rect 22285 4299 22311 4325
rect 22337 4299 22363 4325
rect 2367 4215 2393 4241
rect 28463 4215 28489 4241
rect 28239 4159 28265 4185
rect 28743 4159 28769 4185
rect 28911 4159 28937 4185
rect 30535 4159 30561 4185
rect 2647 4103 2673 4129
rect 6231 4103 6257 4129
rect 21967 4103 21993 4129
rect 27959 4103 27985 4129
rect 29191 4103 29217 4129
rect 29359 4103 29385 4129
rect 30199 4103 30225 4129
rect 30927 4103 30953 4129
rect 6511 4047 6537 4073
rect 21743 4047 21769 4073
rect 29863 4047 29889 4073
rect 31431 3991 31457 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 21903 3907 21929 3933
rect 21955 3907 21981 3933
rect 22007 3907 22033 3933
rect 31543 3823 31569 3849
rect 7407 3767 7433 3793
rect 20847 3767 20873 3793
rect 29583 3767 29609 3793
rect 30759 3767 30785 3793
rect 7631 3711 7657 3737
rect 17431 3711 17457 3737
rect 21127 3711 21153 3737
rect 28911 3711 28937 3737
rect 29415 3711 29441 3737
rect 30255 3711 30281 3737
rect 31151 3711 31177 3737
rect 17711 3655 17737 3681
rect 29191 3655 29217 3681
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 22233 3515 22259 3541
rect 22285 3515 22311 3541
rect 22337 3515 22363 3541
rect 15359 3431 15385 3457
rect 8751 3319 8777 3345
rect 8975 3319 9001 3345
rect 18439 3319 18465 3345
rect 23535 3319 23561 3345
rect 25215 3319 25241 3345
rect 25495 3319 25521 3345
rect 29247 3319 29273 3345
rect 29695 3319 29721 3345
rect 29975 3319 30001 3345
rect 30143 3319 30169 3345
rect 31039 3319 31065 3345
rect 15135 3263 15161 3289
rect 18159 3263 18185 3289
rect 23703 3263 23729 3289
rect 29471 3263 29497 3289
rect 31431 3263 31457 3289
rect 30647 3207 30673 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 21903 3123 21929 3149
rect 21955 3123 21981 3149
rect 22007 3123 22033 3149
rect 30759 3039 30785 3065
rect 31543 3039 31569 3065
rect 1023 2983 1049 3009
rect 4047 2983 4073 3009
rect 13287 2983 13313 3009
rect 14799 2983 14825 3009
rect 28967 2983 28993 3009
rect 29639 2983 29665 3009
rect 4327 2927 4353 2953
rect 13567 2927 13593 2953
rect 29415 2927 29441 2953
rect 30255 2927 30281 2953
rect 31095 2927 31121 2953
rect 15079 2871 15105 2897
rect 22079 2871 22105 2897
rect 22359 2871 22385 2897
rect 1247 2815 1273 2841
rect 28687 2815 28713 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 22233 2731 22259 2757
rect 22285 2731 22311 2757
rect 22337 2731 22363 2757
rect 1247 2647 1273 2673
rect 8639 2647 8665 2673
rect 10935 2647 10961 2673
rect 12559 2647 12585 2673
rect 20175 2647 20201 2673
rect 21183 2647 21209 2673
rect 29695 2647 29721 2673
rect 967 2591 993 2617
rect 9367 2591 9393 2617
rect 9647 2591 9673 2617
rect 10655 2591 10681 2617
rect 12279 2591 12305 2617
rect 14519 2591 14545 2617
rect 20455 2591 20481 2617
rect 20903 2591 20929 2617
rect 21743 2591 21769 2617
rect 25439 2591 25465 2617
rect 28631 2591 28657 2617
rect 29191 2591 29217 2617
rect 30143 2591 30169 2617
rect 30535 2591 30561 2617
rect 31319 2591 31345 2617
rect 14799 2535 14825 2561
rect 21463 2535 21489 2561
rect 25215 2535 25241 2561
rect 28351 2535 28377 2561
rect 28911 2535 28937 2561
rect 29975 2535 30001 2561
rect 30927 2535 30953 2561
rect 8415 2479 8441 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 21903 2339 21929 2365
rect 21955 2339 21981 2365
rect 22007 2339 22033 2365
rect 31543 2255 31569 2281
rect 967 2199 993 2225
rect 8247 2199 8273 2225
rect 27847 2199 27873 2225
rect 21295 2143 21321 2169
rect 24543 2143 24569 2169
rect 31095 2143 31121 2169
rect 21015 2087 21041 2113
rect 24263 2087 24289 2113
rect 30255 2087 30281 2113
rect 30647 2087 30673 2113
rect 1191 2031 1217 2057
rect 8527 2031 8553 2057
rect 28071 2031 28097 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 22233 1947 22259 1973
rect 22285 1947 22311 1973
rect 22337 1947 22363 1973
rect 2591 1863 2617 1889
rect 11999 1863 12025 1889
rect 20399 1863 20425 1889
rect 25271 1863 25297 1889
rect 2871 1807 2897 1833
rect 22191 1807 22217 1833
rect 22471 1807 22497 1833
rect 23255 1807 23281 1833
rect 24991 1807 25017 1833
rect 1303 1751 1329 1777
rect 8583 1751 8609 1777
rect 23479 1751 23505 1777
rect 29695 1751 29721 1777
rect 29975 1751 30001 1777
rect 30143 1751 30169 1777
rect 30927 1751 30953 1777
rect 1079 1695 1105 1721
rect 8415 1695 8441 1721
rect 11775 1695 11801 1721
rect 20175 1695 20201 1721
rect 30647 1695 30673 1721
rect 31431 1695 31457 1721
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 21903 1555 21929 1581
rect 21955 1555 21981 1581
rect 22007 1555 22033 1581
rect 31543 1471 31569 1497
rect 26055 1415 26081 1441
rect 29415 1359 29441 1385
rect 29639 1359 29665 1385
rect 31095 1359 31121 1385
rect 29191 1303 29217 1329
rect 30255 1303 30281 1329
rect 30647 1303 30673 1329
rect 26279 1247 26305 1273
rect 28911 1247 28937 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 22233 1163 22259 1189
rect 22285 1163 22311 1189
rect 22337 1163 22363 1189
rect 6231 1079 6257 1105
rect 7631 1079 7657 1105
rect 8079 1079 8105 1105
rect 11439 1079 11465 1105
rect 15415 1079 15441 1105
rect 16479 1079 16505 1105
rect 17935 1079 17961 1105
rect 18439 1079 18465 1105
rect 19727 1079 19753 1105
rect 20903 1079 20929 1105
rect 21351 1079 21377 1105
rect 21799 1079 21825 1105
rect 22919 1079 22945 1105
rect 29695 1079 29721 1105
rect 967 1023 993 1049
rect 4831 1023 4857 1049
rect 7351 1023 7377 1049
rect 7799 1023 7825 1049
rect 17655 1023 17681 1049
rect 18159 1023 18185 1049
rect 18775 1023 18801 1049
rect 19447 1023 19473 1049
rect 20623 1023 20649 1049
rect 21071 1023 21097 1049
rect 21519 1023 21545 1049
rect 24319 1023 24345 1049
rect 24879 1023 24905 1049
rect 25439 1023 25465 1049
rect 28799 1023 28825 1049
rect 29247 1023 29273 1049
rect 30143 1023 30169 1049
rect 1247 967 1273 993
rect 4551 967 4577 993
rect 5055 967 5081 993
rect 15247 967 15273 993
rect 19055 967 19081 993
rect 24039 967 24065 993
rect 24599 967 24625 993
rect 25215 967 25241 993
rect 28575 967 28601 993
rect 28967 967 28993 993
rect 29975 967 30001 993
rect 30927 967 30953 993
rect 5279 911 5305 937
rect 6511 911 6537 937
rect 11159 911 11185 937
rect 16199 911 16225 937
rect 22695 911 22721 937
rect 31431 911 31457 937
rect 30647 855 30673 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 21903 771 21929 797
rect 21955 771 21981 797
rect 22007 771 22033 797
rect 31543 687 31569 713
rect 911 631 937 657
rect 29807 631 29833 657
rect 30591 631 30617 657
rect 5055 575 5081 601
rect 30087 575 30113 601
rect 31095 575 31121 601
rect 5279 519 5305 545
rect 29303 519 29329 545
rect 1191 463 1217 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
rect 22233 379 22259 405
rect 22285 379 22311 405
rect 22337 379 22363 405
<< metal2 >>
rect 2128 7056 2184 7112
rect 2352 7056 2408 7112
rect 2576 7056 2632 7112
rect 2800 7056 2856 7112
rect 3024 7056 3080 7112
rect 3248 7056 3304 7112
rect 3472 7056 3528 7112
rect 3696 7056 3752 7112
rect 3920 7056 3976 7112
rect 4144 7056 4200 7112
rect 4368 7056 4424 7112
rect 4592 7056 4648 7112
rect 4816 7056 4872 7112
rect 5040 7056 5096 7112
rect 5264 7056 5320 7112
rect 5488 7056 5544 7112
rect 5712 7056 5768 7112
rect 5936 7056 5992 7112
rect 6160 7056 6216 7112
rect 6384 7056 6440 7112
rect 6608 7056 6664 7112
rect 6832 7056 6888 7112
rect 7056 7056 7112 7112
rect 7280 7056 7336 7112
rect 7504 7056 7560 7112
rect 7728 7056 7784 7112
rect 7952 7056 8008 7112
rect 8176 7056 8232 7112
rect 8400 7056 8456 7112
rect 8624 7056 8680 7112
rect 8848 7056 8904 7112
rect 9072 7056 9128 7112
rect 9296 7056 9352 7112
rect 9520 7056 9576 7112
rect 9744 7056 9800 7112
rect 9968 7056 10024 7112
rect 10192 7056 10248 7112
rect 10416 7056 10472 7112
rect 10640 7056 10696 7112
rect 10864 7056 10920 7112
rect 11088 7056 11144 7112
rect 11312 7056 11368 7112
rect 11536 7056 11592 7112
rect 11760 7056 11816 7112
rect 11984 7056 12040 7112
rect 12208 7056 12264 7112
rect 12432 7056 12488 7112
rect 12656 7056 12712 7112
rect 12880 7056 12936 7112
rect 13104 7056 13160 7112
rect 13328 7056 13384 7112
rect 13552 7056 13608 7112
rect 13776 7056 13832 7112
rect 14000 7056 14056 7112
rect 14224 7056 14280 7112
rect 14448 7056 14504 7112
rect 14672 7056 14728 7112
rect 14896 7056 14952 7112
rect 15120 7056 15176 7112
rect 15344 7056 15400 7112
rect 15568 7056 15624 7112
rect 15792 7056 15848 7112
rect 16016 7056 16072 7112
rect 16240 7056 16296 7112
rect 16464 7056 16520 7112
rect 16688 7056 16744 7112
rect 16912 7056 16968 7112
rect 17136 7056 17192 7112
rect 17360 7056 17416 7112
rect 17584 7056 17640 7112
rect 17808 7056 17864 7112
rect 18032 7056 18088 7112
rect 18256 7056 18312 7112
rect 18480 7056 18536 7112
rect 18704 7056 18760 7112
rect 18928 7056 18984 7112
rect 19152 7056 19208 7112
rect 19376 7056 19432 7112
rect 19600 7056 19656 7112
rect 19824 7056 19880 7112
rect 20048 7056 20104 7112
rect 20272 7056 20328 7112
rect 20496 7056 20552 7112
rect 20720 7056 20776 7112
rect 20944 7056 21000 7112
rect 21168 7056 21224 7112
rect 21392 7056 21448 7112
rect 21616 7056 21672 7112
rect 21840 7056 21896 7112
rect 22064 7056 22120 7112
rect 22288 7056 22344 7112
rect 22512 7056 22568 7112
rect 22736 7056 22792 7112
rect 22960 7056 23016 7112
rect 23184 7056 23240 7112
rect 23408 7056 23464 7112
rect 23632 7056 23688 7112
rect 23856 7056 23912 7112
rect 24080 7056 24136 7112
rect 24304 7056 24360 7112
rect 24528 7056 24584 7112
rect 24752 7056 24808 7112
rect 24976 7056 25032 7112
rect 25200 7056 25256 7112
rect 25424 7056 25480 7112
rect 25648 7056 25704 7112
rect 25872 7056 25928 7112
rect 26096 7056 26152 7112
rect 26320 7056 26376 7112
rect 26544 7056 26600 7112
rect 26768 7056 26824 7112
rect 26992 7056 27048 7112
rect 27216 7056 27272 7112
rect 27440 7056 27496 7112
rect 27664 7056 27720 7112
rect 27888 7056 27944 7112
rect 28112 7056 28168 7112
rect 28336 7056 28392 7112
rect 28560 7056 28616 7112
rect 28784 7056 28840 7112
rect 29008 7056 29064 7112
rect 29232 7056 29288 7112
rect 29456 7056 29512 7112
rect 29680 7056 29736 7112
rect 29904 7056 29960 7112
rect 126 6986 154 6991
rect 126 3458 154 6958
rect 1862 6818 1890 6823
rect 1806 6762 1834 6767
rect 1246 6594 1274 6599
rect 798 6538 826 6543
rect 462 6314 490 6319
rect 462 5250 490 6286
rect 462 5217 490 5222
rect 798 5026 826 6510
rect 798 4993 826 4998
rect 854 6481 882 6487
rect 854 6455 855 6481
rect 881 6455 882 6481
rect 854 4214 882 6455
rect 1078 6482 1106 6487
rect 966 5642 994 5647
rect 966 5595 994 5614
rect 854 4186 938 4214
rect 126 3425 154 3430
rect 910 2618 938 4186
rect 1022 3290 1050 3295
rect 1022 3009 1050 3262
rect 1022 2983 1023 3009
rect 1049 2983 1050 3009
rect 1022 2977 1050 2983
rect 1022 2898 1050 2903
rect 966 2618 994 2623
rect 910 2617 994 2618
rect 910 2591 967 2617
rect 993 2591 994 2617
rect 910 2590 994 2591
rect 966 2585 994 2590
rect 910 2226 938 2231
rect 910 657 938 2198
rect 966 2226 994 2231
rect 1022 2226 1050 2870
rect 966 2225 1050 2226
rect 966 2199 967 2225
rect 993 2199 1050 2225
rect 966 2198 1050 2199
rect 966 2193 994 2198
rect 1078 1721 1106 6454
rect 1246 6425 1274 6566
rect 1246 6399 1247 6425
rect 1273 6399 1274 6425
rect 1246 6393 1274 6399
rect 1414 6146 1442 6151
rect 1134 5697 1162 5703
rect 1134 5671 1135 5697
rect 1161 5671 1162 5697
rect 1134 5306 1162 5671
rect 1134 5273 1162 5278
rect 1190 5586 1218 5591
rect 1190 4634 1218 5558
rect 1190 4601 1218 4606
rect 1414 4577 1442 6118
rect 1806 6145 1834 6734
rect 1862 6593 1890 6790
rect 1862 6567 1863 6593
rect 1889 6567 1890 6593
rect 1862 6561 1890 6567
rect 2086 6706 2114 6711
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 1806 6119 1807 6145
rect 1833 6119 1834 6145
rect 1806 6113 1834 6119
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 1414 4551 1415 4577
rect 1441 4551 1442 4577
rect 1414 4545 1442 4551
rect 1526 5250 1554 5255
rect 1526 3794 1554 5222
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 1638 4578 1666 4583
rect 1638 4521 1666 4550
rect 1638 4495 1639 4521
rect 1665 4495 1666 4521
rect 1638 4489 1666 4495
rect 2086 4242 2114 6678
rect 2142 6594 2170 7056
rect 2366 6762 2394 7056
rect 2366 6729 2394 6734
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 2142 6561 2170 6566
rect 2142 6482 2170 6487
rect 2142 6481 2450 6482
rect 2142 6455 2143 6481
rect 2169 6455 2450 6481
rect 2142 6454 2450 6455
rect 2142 6449 2170 6454
rect 2198 6034 2226 6039
rect 2198 5987 2226 6006
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 2310 5810 2338 5815
rect 2310 5763 2338 5782
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 2366 4242 2394 4247
rect 2086 4241 2394 4242
rect 2086 4215 2367 4241
rect 2393 4215 2394 4241
rect 2086 4214 2394 4215
rect 2366 4209 2394 4214
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 1526 3761 1554 3766
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 1302 3346 1330 3351
rect 1246 2842 1274 2847
rect 1246 2795 1274 2814
rect 1246 2674 1274 2679
rect 1302 2674 1330 3318
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 1246 2673 1330 2674
rect 1246 2647 1247 2673
rect 1273 2647 1330 2673
rect 1246 2646 1330 2647
rect 1246 2641 1274 2646
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 1190 2058 1218 2063
rect 1190 2011 1218 2030
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 1302 1778 1330 1783
rect 1302 1731 1330 1750
rect 1078 1695 1079 1721
rect 1105 1695 1106 1721
rect 1078 1689 1106 1695
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 966 1442 994 1447
rect 966 1049 994 1414
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 966 1023 967 1049
rect 993 1023 994 1049
rect 966 1017 994 1023
rect 1246 994 1274 999
rect 1246 947 1274 966
rect 910 631 911 657
rect 937 631 938 657
rect 910 625 938 631
rect 1470 826 1498 831
rect 1190 490 1218 495
rect 1190 443 1218 462
rect 1470 56 1498 798
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2422 770 2450 6454
rect 2590 5810 2618 7056
rect 2814 6818 2842 7056
rect 2814 6785 2842 6790
rect 2982 6594 3010 6599
rect 2982 6547 3010 6566
rect 2590 5777 2618 5782
rect 2926 6034 2954 6039
rect 2590 5697 2618 5703
rect 2590 5671 2591 5697
rect 2617 5671 2618 5697
rect 2590 5586 2618 5671
rect 2590 5553 2618 5558
rect 2590 5474 2618 5479
rect 2534 4634 2562 4639
rect 2534 4521 2562 4606
rect 2534 4495 2535 4521
rect 2561 4495 2562 4521
rect 2534 4489 2562 4495
rect 2590 2898 2618 5446
rect 2758 4802 2786 4807
rect 2758 4577 2786 4774
rect 2758 4551 2759 4577
rect 2785 4551 2786 4577
rect 2758 4545 2786 4551
rect 2646 4130 2674 4135
rect 2646 4083 2674 4102
rect 2926 3010 2954 6006
rect 3038 5641 3066 7056
rect 3262 6594 3290 7056
rect 3486 6594 3514 7056
rect 3262 6566 3402 6594
rect 3038 5615 3039 5641
rect 3065 5615 3066 5641
rect 3038 5609 3066 5615
rect 3262 6481 3290 6487
rect 3262 6455 3263 6481
rect 3289 6455 3290 6481
rect 2926 2977 2954 2982
rect 2590 2865 2618 2870
rect 3262 2618 3290 6455
rect 3318 5698 3346 5703
rect 3318 5651 3346 5670
rect 3374 5361 3402 6566
rect 3486 6561 3514 6566
rect 3486 6202 3514 6207
rect 3710 6202 3738 7056
rect 3766 6594 3794 6599
rect 3934 6594 3962 7056
rect 3934 6566 4130 6594
rect 3766 6547 3794 6566
rect 3486 6201 3738 6202
rect 3486 6175 3487 6201
rect 3513 6175 3738 6201
rect 3486 6174 3738 6175
rect 4046 6481 4074 6487
rect 4046 6455 4047 6481
rect 4073 6455 4074 6481
rect 3486 6169 3514 6174
rect 3766 6034 3794 6039
rect 3766 6033 3850 6034
rect 3766 6007 3767 6033
rect 3793 6007 3850 6033
rect 3766 6006 3850 6007
rect 3766 6001 3794 6006
rect 3374 5335 3375 5361
rect 3401 5335 3402 5361
rect 3374 5329 3402 5335
rect 3262 2585 3290 2590
rect 3766 5249 3794 5255
rect 3766 5223 3767 5249
rect 3793 5223 3794 5249
rect 3766 2450 3794 5223
rect 3766 2417 3794 2422
rect 2590 2114 2618 2119
rect 2590 1889 2618 2086
rect 2590 1863 2591 1889
rect 2617 1863 2618 1889
rect 2590 1857 2618 1863
rect 2870 1946 2898 1951
rect 2870 1833 2898 1918
rect 2870 1807 2871 1833
rect 2897 1807 2898 1833
rect 2870 1801 2898 1807
rect 3822 1050 3850 6006
rect 3878 5810 3906 5815
rect 3878 5763 3906 5782
rect 3878 5194 3906 5199
rect 3878 5025 3906 5166
rect 3878 4999 3879 5025
rect 3905 4999 3906 5025
rect 3878 4993 3906 4999
rect 4046 3682 4074 6455
rect 4102 5361 4130 6566
rect 4158 5810 4186 7056
rect 4382 6594 4410 7056
rect 4382 6561 4410 6566
rect 4270 6202 4298 6207
rect 4270 6155 4298 6174
rect 4550 6033 4578 6039
rect 4550 6007 4551 6033
rect 4577 6007 4578 6033
rect 4550 5978 4578 6007
rect 4550 5945 4578 5950
rect 4158 5777 4186 5782
rect 4158 5697 4186 5703
rect 4158 5671 4159 5697
rect 4185 5671 4186 5697
rect 4158 5530 4186 5671
rect 4158 5497 4186 5502
rect 4214 5586 4242 5591
rect 4102 5335 4103 5361
rect 4129 5335 4130 5361
rect 4102 5329 4130 5335
rect 4158 4858 4186 4863
rect 4158 4811 4186 4830
rect 4046 3649 4074 3654
rect 4046 3010 4074 3015
rect 4046 2963 4074 2982
rect 4214 1610 4242 5558
rect 4606 5418 4634 7056
rect 4830 6202 4858 7056
rect 4886 6650 4914 6655
rect 4886 6593 4914 6622
rect 4886 6567 4887 6593
rect 4913 6567 4914 6593
rect 4886 6561 4914 6567
rect 4998 6594 5026 6599
rect 4830 6169 4858 6174
rect 4998 6145 5026 6566
rect 5054 6314 5082 7056
rect 5278 6594 5306 7056
rect 5278 6561 5306 6566
rect 5166 6482 5194 6487
rect 5166 6481 5418 6482
rect 5166 6455 5167 6481
rect 5193 6455 5418 6481
rect 5166 6454 5418 6455
rect 5166 6449 5194 6454
rect 5054 6286 5138 6314
rect 4998 6119 4999 6145
rect 5025 6119 5026 6145
rect 4998 6113 5026 6119
rect 4830 5418 4858 5423
rect 4606 5417 4858 5418
rect 4606 5391 4831 5417
rect 4857 5391 4858 5417
rect 4606 5390 4858 5391
rect 4830 5385 4858 5390
rect 4550 5249 4578 5255
rect 4550 5223 4551 5249
rect 4577 5223 4578 5249
rect 4550 5082 4578 5223
rect 4550 5049 4578 5054
rect 5110 4858 5138 6286
rect 5334 6146 5362 6151
rect 5334 6089 5362 6118
rect 5334 6063 5335 6089
rect 5361 6063 5362 6089
rect 5334 6057 5362 6063
rect 5334 5249 5362 5255
rect 5334 5223 5335 5249
rect 5361 5223 5362 5249
rect 5334 5194 5362 5223
rect 5334 5161 5362 5166
rect 5390 4914 5418 6454
rect 5502 6146 5530 7056
rect 5670 6594 5698 6599
rect 5670 6547 5698 6566
rect 5502 6118 5642 6146
rect 5446 5810 5474 5815
rect 5446 5763 5474 5782
rect 5390 4881 5418 4886
rect 5446 5698 5474 5703
rect 5278 4858 5306 4863
rect 5110 4857 5306 4858
rect 5110 4831 5279 4857
rect 5305 4831 5306 4857
rect 5110 4830 5306 4831
rect 5278 4825 5306 4830
rect 4326 2954 4354 2959
rect 4326 2907 4354 2926
rect 5446 2338 5474 5670
rect 5614 5417 5642 6118
rect 5726 5810 5754 7056
rect 5950 6650 5978 7056
rect 5950 6617 5978 6622
rect 5950 6481 5978 6487
rect 5950 6455 5951 6481
rect 5977 6455 5978 6481
rect 5838 6202 5866 6207
rect 5838 6155 5866 6174
rect 5726 5777 5754 5782
rect 5614 5391 5615 5417
rect 5641 5391 5642 5417
rect 5614 5385 5642 5391
rect 5726 5697 5754 5703
rect 5726 5671 5727 5697
rect 5753 5671 5754 5697
rect 5726 3234 5754 5671
rect 5782 4913 5810 4919
rect 5782 4887 5783 4913
rect 5809 4887 5810 4913
rect 5782 3570 5810 4887
rect 5782 3537 5810 3542
rect 5726 3201 5754 3206
rect 5446 2305 5474 2310
rect 5894 2898 5922 2903
rect 4214 1577 4242 1582
rect 3822 1017 3850 1022
rect 4830 1498 4858 1503
rect 4830 1049 4858 1470
rect 4830 1023 4831 1049
rect 4857 1023 4858 1049
rect 4830 1017 4858 1023
rect 4550 993 4578 999
rect 4550 967 4551 993
rect 4577 967 4578 993
rect 4550 938 4578 967
rect 5054 994 5082 999
rect 5054 993 5138 994
rect 5054 967 5055 993
rect 5081 967 5138 993
rect 5054 966 5138 967
rect 5054 961 5082 966
rect 4550 905 4578 910
rect 2422 737 2450 742
rect 4382 658 4410 663
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2926 154 2954 159
rect 2926 56 2954 126
rect 4382 56 4410 630
rect 5054 601 5082 607
rect 5054 575 5055 601
rect 5081 575 5082 601
rect 5054 210 5082 575
rect 5110 266 5138 966
rect 5278 937 5306 943
rect 5278 911 5279 937
rect 5305 911 5306 937
rect 5278 882 5306 911
rect 5278 849 5306 854
rect 5894 826 5922 2870
rect 5950 1554 5978 6455
rect 6118 6033 6146 6039
rect 6118 6007 6119 6033
rect 6145 6007 6146 6033
rect 6118 5922 6146 6007
rect 6118 5889 6146 5894
rect 6062 5810 6090 5815
rect 5950 1521 5978 1526
rect 6006 2842 6034 2847
rect 6006 1442 6034 2814
rect 6006 1409 6034 1414
rect 5838 798 5922 826
rect 5950 1330 5978 1335
rect 5110 233 5138 238
rect 5278 545 5306 551
rect 5278 519 5279 545
rect 5305 519 5306 545
rect 5054 177 5082 182
rect 5278 154 5306 519
rect 5278 121 5306 126
rect 5838 56 5866 798
rect 5950 658 5978 1302
rect 5950 625 5978 630
rect 6062 210 6090 5782
rect 6174 5641 6202 7056
rect 6398 6202 6426 7056
rect 6622 6594 6650 7056
rect 6622 6561 6650 6566
rect 6454 6482 6482 6487
rect 6454 6435 6482 6454
rect 6398 6169 6426 6174
rect 6678 6202 6706 6207
rect 6174 5615 6175 5641
rect 6201 5615 6202 5641
rect 6174 5609 6202 5615
rect 6342 6034 6370 6039
rect 6286 5418 6314 5423
rect 6118 5250 6146 5255
rect 6118 5203 6146 5222
rect 6230 4129 6258 4135
rect 6230 4103 6231 4129
rect 6257 4103 6258 4129
rect 6174 4074 6202 4079
rect 6118 1386 6146 1391
rect 6118 434 6146 1358
rect 6174 1106 6202 4046
rect 6230 3010 6258 4103
rect 6286 3962 6314 5390
rect 6286 3929 6314 3934
rect 6230 2977 6258 2982
rect 6342 2226 6370 6006
rect 6510 5697 6538 5703
rect 6510 5671 6511 5697
rect 6537 5671 6538 5697
rect 6510 5362 6538 5671
rect 6510 5329 6538 5334
rect 6510 5193 6538 5199
rect 6510 5167 6511 5193
rect 6537 5167 6538 5193
rect 6454 5082 6482 5087
rect 6398 4298 6426 4303
rect 6398 2954 6426 4270
rect 6398 2921 6426 2926
rect 6342 2193 6370 2198
rect 6454 2002 6482 5054
rect 6510 4466 6538 5167
rect 6678 5026 6706 6174
rect 6734 5697 6762 5703
rect 6734 5671 6735 5697
rect 6761 5671 6762 5697
rect 6734 5474 6762 5671
rect 6734 5441 6762 5446
rect 6678 4993 6706 4998
rect 6790 5249 6818 5255
rect 6790 5223 6791 5249
rect 6817 5223 6818 5249
rect 6790 4858 6818 5223
rect 6846 4858 6874 7056
rect 6958 6426 6986 6431
rect 6958 6379 6986 6398
rect 7070 6146 7098 7056
rect 7070 6118 7154 6146
rect 7070 6034 7098 6039
rect 7070 5987 7098 6006
rect 7126 5418 7154 6118
rect 7182 5642 7210 5647
rect 7294 5642 7322 7056
rect 7406 6538 7434 6543
rect 7406 6425 7434 6510
rect 7406 6399 7407 6425
rect 7433 6399 7434 6425
rect 7406 6393 7434 6399
rect 7462 6482 7490 6487
rect 7462 6145 7490 6454
rect 7518 6426 7546 7056
rect 7518 6393 7546 6398
rect 7462 6119 7463 6145
rect 7489 6119 7490 6145
rect 7462 6113 7490 6119
rect 7350 5978 7378 5983
rect 7350 5698 7378 5950
rect 7518 5922 7546 5927
rect 7518 5754 7546 5894
rect 7518 5721 7546 5726
rect 7350 5665 7378 5670
rect 7462 5697 7490 5703
rect 7462 5671 7463 5697
rect 7489 5671 7490 5697
rect 7182 5641 7322 5642
rect 7182 5615 7183 5641
rect 7209 5615 7322 5641
rect 7182 5614 7322 5615
rect 7182 5609 7210 5614
rect 7350 5530 7378 5535
rect 7182 5418 7210 5423
rect 7126 5417 7210 5418
rect 7126 5391 7183 5417
rect 7209 5391 7210 5417
rect 7126 5390 7210 5391
rect 7182 5385 7210 5390
rect 7070 4858 7098 4863
rect 6846 4857 7098 4858
rect 6846 4831 7071 4857
rect 7097 4831 7098 4857
rect 6846 4830 7098 4831
rect 6790 4825 6818 4830
rect 7070 4825 7098 4830
rect 6734 4802 6762 4807
rect 6510 4433 6538 4438
rect 6622 4522 6650 4527
rect 6510 4074 6538 4079
rect 6510 4073 6594 4074
rect 6510 4047 6511 4073
rect 6537 4047 6594 4073
rect 6510 4046 6594 4047
rect 6510 4041 6538 4046
rect 6454 1969 6482 1974
rect 6510 2674 6538 2679
rect 6510 1890 6538 2646
rect 6510 1857 6538 1862
rect 6286 1554 6314 1559
rect 6230 1106 6258 1111
rect 6174 1105 6258 1106
rect 6174 1079 6231 1105
rect 6257 1079 6258 1105
rect 6174 1078 6258 1079
rect 6230 1073 6258 1078
rect 6286 1106 6314 1526
rect 6566 1554 6594 4046
rect 6622 4018 6650 4494
rect 6622 3985 6650 3990
rect 6678 4466 6706 4471
rect 6678 3738 6706 4438
rect 6734 3906 6762 4774
rect 6734 3873 6762 3878
rect 6846 4354 6874 4359
rect 6678 3705 6706 3710
rect 6846 1834 6874 4326
rect 7350 3458 7378 5502
rect 7406 3794 7434 3799
rect 7406 3747 7434 3766
rect 7350 3425 7378 3430
rect 7462 3290 7490 5671
rect 7742 5418 7770 7056
rect 7854 6482 7882 6487
rect 7966 6482 7994 7056
rect 8190 6706 8218 7056
rect 7854 6481 7938 6482
rect 7854 6455 7855 6481
rect 7881 6455 7938 6481
rect 7854 6454 7938 6455
rect 7854 6449 7882 6454
rect 7910 5530 7938 6454
rect 7966 6449 7994 6454
rect 8022 6678 8218 6706
rect 7966 5642 7994 5647
rect 8022 5642 8050 6678
rect 8190 6594 8218 6599
rect 8190 6201 8218 6566
rect 8414 6538 8442 7056
rect 8414 6505 8442 6510
rect 8582 6986 8610 6991
rect 8190 6175 8191 6201
rect 8217 6175 8218 6201
rect 8190 6169 8218 6175
rect 7966 5641 8050 5642
rect 7966 5615 7967 5641
rect 7993 5615 8050 5641
rect 7966 5614 8050 5615
rect 8470 6033 8498 6039
rect 8470 6007 8471 6033
rect 8497 6007 8498 6033
rect 7966 5609 7994 5614
rect 7910 5502 8330 5530
rect 8134 5418 8162 5423
rect 7742 5417 8162 5418
rect 7742 5391 8135 5417
rect 8161 5391 8162 5417
rect 7742 5390 8162 5391
rect 8134 5385 8162 5390
rect 7686 5249 7714 5255
rect 7686 5223 7687 5249
rect 7713 5223 7714 5249
rect 7462 3257 7490 3262
rect 7518 4913 7546 4919
rect 7518 4887 7519 4913
rect 7545 4887 7546 4913
rect 7406 3234 7434 3239
rect 7126 2730 7154 2735
rect 7126 2506 7154 2702
rect 7126 2473 7154 2478
rect 7406 2394 7434 3206
rect 7518 3234 7546 4887
rect 7574 4298 7602 4303
rect 7602 4270 7658 4298
rect 7574 4265 7602 4270
rect 7630 4186 7658 4270
rect 7630 4153 7658 4158
rect 7686 4074 7714 5223
rect 7854 5249 7882 5255
rect 7854 5223 7855 5249
rect 7881 5223 7882 5249
rect 7686 4041 7714 4046
rect 7742 4298 7770 4303
rect 7742 3962 7770 4270
rect 7630 3934 7770 3962
rect 7630 3737 7658 3934
rect 7630 3711 7631 3737
rect 7657 3711 7658 3737
rect 7630 3705 7658 3711
rect 7686 3738 7714 3743
rect 7518 3201 7546 3206
rect 7406 2361 7434 2366
rect 6846 1801 6874 1806
rect 7126 1722 7154 1727
rect 6566 1521 6594 1526
rect 6622 1666 6650 1671
rect 6286 1073 6314 1078
rect 6118 401 6146 406
rect 6510 937 6538 943
rect 6510 911 6511 937
rect 6537 911 6538 937
rect 6510 378 6538 911
rect 6622 714 6650 1638
rect 6678 938 6706 943
rect 6678 770 6706 910
rect 7126 826 7154 1694
rect 7686 1218 7714 3710
rect 7854 2842 7882 5223
rect 8246 4074 8274 4079
rect 7854 2809 7882 2814
rect 8078 2954 8106 2959
rect 7686 1185 7714 1190
rect 7798 1610 7826 1615
rect 7630 1106 7658 1111
rect 7630 1059 7658 1078
rect 7350 1050 7378 1055
rect 7350 1003 7378 1022
rect 7798 1049 7826 1582
rect 8078 1105 8106 2926
rect 8246 2225 8274 4046
rect 8302 3346 8330 5502
rect 8302 3313 8330 3318
rect 8358 3402 8386 3407
rect 8246 2199 8247 2225
rect 8273 2199 8274 2225
rect 8246 2193 8274 2199
rect 8358 2058 8386 3374
rect 8470 3066 8498 6007
rect 8470 3033 8498 3038
rect 8414 2505 8442 2511
rect 8414 2479 8415 2505
rect 8441 2479 8442 2505
rect 8414 2450 8442 2479
rect 8414 2417 8442 2422
rect 8358 2025 8386 2030
rect 8414 2338 8442 2343
rect 8414 1721 8442 2310
rect 8414 1695 8415 1721
rect 8441 1695 8442 1721
rect 8414 1689 8442 1695
rect 8526 2057 8554 2063
rect 8526 2031 8527 2057
rect 8553 2031 8554 2057
rect 8078 1079 8079 1105
rect 8105 1079 8106 1105
rect 8078 1073 8106 1079
rect 7798 1023 7799 1049
rect 7825 1023 7826 1049
rect 7798 1017 7826 1023
rect 7126 793 7154 798
rect 7574 994 7602 999
rect 6678 737 6706 742
rect 6622 681 6650 686
rect 7294 714 7322 719
rect 6510 345 6538 350
rect 6062 177 6090 182
rect 7294 56 7322 686
rect 7574 602 7602 966
rect 7686 882 7714 887
rect 7686 658 7714 854
rect 7686 625 7714 630
rect 7574 569 7602 574
rect 8526 322 8554 2031
rect 8582 1777 8610 6958
rect 8638 6594 8666 7056
rect 8638 6561 8666 6566
rect 8694 6650 8722 6655
rect 8694 6593 8722 6622
rect 8694 6567 8695 6593
rect 8721 6567 8722 6593
rect 8694 6561 8722 6567
rect 8638 5642 8666 5647
rect 8638 5305 8666 5614
rect 8862 5418 8890 7056
rect 8918 6481 8946 6487
rect 8918 6455 8919 6481
rect 8945 6455 8946 6481
rect 8918 5530 8946 6455
rect 8974 6370 9002 6375
rect 8974 6201 9002 6342
rect 8974 6175 8975 6201
rect 9001 6175 9002 6201
rect 8974 6169 9002 6175
rect 9086 5810 9114 7056
rect 9310 6202 9338 7056
rect 9478 6594 9506 6599
rect 9478 6547 9506 6566
rect 9534 6370 9562 7056
rect 9534 6337 9562 6342
rect 9702 6874 9730 6879
rect 9310 6174 9562 6202
rect 9198 6089 9226 6095
rect 9198 6063 9199 6089
rect 9225 6063 9226 6089
rect 9198 5922 9226 6063
rect 9422 6090 9450 6095
rect 9422 6043 9450 6062
rect 9198 5889 9226 5894
rect 9310 5810 9338 5815
rect 9086 5809 9338 5810
rect 9086 5783 9311 5809
rect 9337 5783 9338 5809
rect 9086 5782 9338 5783
rect 9310 5777 9338 5782
rect 9030 5697 9058 5703
rect 9030 5671 9031 5697
rect 9057 5671 9058 5697
rect 8918 5502 9002 5530
rect 8918 5418 8946 5423
rect 8862 5417 8946 5418
rect 8862 5391 8919 5417
rect 8945 5391 8946 5417
rect 8862 5390 8946 5391
rect 8918 5385 8946 5390
rect 8638 5279 8639 5305
rect 8665 5279 8666 5305
rect 8638 5273 8666 5279
rect 8974 4578 9002 5502
rect 8862 4550 9002 4578
rect 8638 4409 8666 4415
rect 8638 4383 8639 4409
rect 8665 4383 8666 4409
rect 8638 3178 8666 4383
rect 8638 3145 8666 3150
rect 8694 3458 8722 3463
rect 8638 2674 8666 2679
rect 8638 2627 8666 2646
rect 8582 1751 8583 1777
rect 8609 1751 8610 1777
rect 8582 1745 8610 1751
rect 8694 1442 8722 3430
rect 8750 3346 8778 3351
rect 8750 3299 8778 3318
rect 8862 3178 8890 4550
rect 8918 4465 8946 4471
rect 8918 4439 8919 4465
rect 8945 4439 8946 4465
rect 8918 4242 8946 4439
rect 8918 4209 8946 4214
rect 8974 4130 9002 4135
rect 8974 3345 9002 4102
rect 9030 3794 9058 5671
rect 9534 5417 9562 6174
rect 9534 5391 9535 5417
rect 9561 5391 9562 5417
rect 9534 5385 9562 5391
rect 9478 5250 9506 5255
rect 9478 5082 9506 5222
rect 9478 5049 9506 5054
rect 9198 4970 9226 4975
rect 9030 3761 9058 3766
rect 9086 3906 9114 3911
rect 8974 3319 8975 3345
rect 9001 3319 9002 3345
rect 8974 3313 9002 3319
rect 8862 3145 8890 3150
rect 8694 1409 8722 1414
rect 8750 2506 8778 2511
rect 8526 289 8554 294
rect 8750 56 8778 2478
rect 9030 1834 9058 1839
rect 9030 1498 9058 1806
rect 9030 1465 9058 1470
rect 9086 434 9114 3878
rect 9198 3402 9226 4942
rect 9198 3369 9226 3374
rect 9702 3122 9730 6846
rect 9758 6650 9786 7056
rect 9758 6617 9786 6622
rect 9814 6986 9842 6991
rect 9758 6482 9786 6487
rect 9758 6435 9786 6454
rect 9702 3089 9730 3094
rect 9366 2618 9394 2623
rect 9366 2571 9394 2590
rect 9646 2618 9674 2623
rect 9646 2571 9674 2590
rect 9142 2562 9170 2567
rect 9142 546 9170 2534
rect 9814 1694 9842 6958
rect 9870 6538 9898 6543
rect 9870 4130 9898 6510
rect 9926 6202 9954 6207
rect 9982 6202 10010 7056
rect 9926 6201 10010 6202
rect 9926 6175 9927 6201
rect 9953 6175 10010 6201
rect 9926 6174 10010 6175
rect 10038 6258 10066 6263
rect 9926 6169 9954 6174
rect 10038 5642 10066 6230
rect 10150 5810 10178 5815
rect 10206 5810 10234 7056
rect 10150 5809 10234 5810
rect 10150 5783 10151 5809
rect 10177 5783 10234 5809
rect 10150 5782 10234 5783
rect 10262 6818 10290 6823
rect 10150 5777 10178 5782
rect 10038 5609 10066 5614
rect 9982 5305 10010 5311
rect 9982 5279 9983 5305
rect 10009 5279 10010 5305
rect 9982 4634 10010 5279
rect 10094 5194 10122 5199
rect 9982 4601 10010 4606
rect 10038 4746 10066 4751
rect 9870 4097 9898 4102
rect 9982 4186 10010 4191
rect 9982 3738 10010 4158
rect 10038 4130 10066 4718
rect 10038 4097 10066 4102
rect 9982 3705 10010 3710
rect 10038 3570 10066 3575
rect 10038 2170 10066 3542
rect 10094 3290 10122 5166
rect 10262 4578 10290 6790
rect 10430 6594 10458 7056
rect 10430 6561 10458 6566
rect 10598 6594 10626 6599
rect 10598 6547 10626 6566
rect 10486 5978 10514 5983
rect 10262 4545 10290 4550
rect 10318 5697 10346 5703
rect 10318 5671 10319 5697
rect 10345 5671 10346 5697
rect 10094 3257 10122 3262
rect 10038 2137 10066 2142
rect 10262 1890 10290 1895
rect 10318 1890 10346 5671
rect 10486 5586 10514 5950
rect 10654 5642 10682 7056
rect 10878 6594 10906 7056
rect 11102 6594 11130 7056
rect 10878 6566 11074 6594
rect 10822 6481 10850 6487
rect 10822 6455 10823 6481
rect 10849 6455 10850 6481
rect 10710 5642 10738 5647
rect 10654 5641 10738 5642
rect 10654 5615 10711 5641
rect 10737 5615 10738 5641
rect 10654 5614 10738 5615
rect 10710 5609 10738 5614
rect 10486 5553 10514 5558
rect 10822 5418 10850 6455
rect 10822 5385 10850 5390
rect 10878 5866 10906 5871
rect 10766 5249 10794 5255
rect 10766 5223 10767 5249
rect 10793 5223 10794 5249
rect 10486 5193 10514 5199
rect 10486 5167 10487 5193
rect 10513 5167 10514 5193
rect 10430 5082 10458 5087
rect 10374 4522 10402 4527
rect 10374 3850 10402 4494
rect 10430 3906 10458 5054
rect 10430 3873 10458 3878
rect 10374 3817 10402 3822
rect 10486 3514 10514 5167
rect 10766 5194 10794 5223
rect 10766 5161 10794 5166
rect 10822 4466 10850 4471
rect 10822 4419 10850 4438
rect 10486 3481 10514 3486
rect 10766 4354 10794 4359
rect 10430 3458 10458 3463
rect 10430 2898 10458 3430
rect 10430 2865 10458 2870
rect 10654 3066 10682 3071
rect 10654 2617 10682 3038
rect 10766 3010 10794 4326
rect 10766 2977 10794 2982
rect 10822 3850 10850 3855
rect 10822 2674 10850 3822
rect 10878 3010 10906 5838
rect 11046 5418 11074 6566
rect 11102 6561 11130 6566
rect 11158 6762 11186 6767
rect 11158 5698 11186 6734
rect 11214 6202 11242 6207
rect 11326 6202 11354 7056
rect 11382 6594 11410 6599
rect 11382 6547 11410 6566
rect 11214 6201 11354 6202
rect 11214 6175 11215 6201
rect 11241 6175 11354 6201
rect 11214 6174 11354 6175
rect 11214 6169 11242 6174
rect 11494 6033 11522 6039
rect 11494 6007 11495 6033
rect 11521 6007 11522 6033
rect 11438 5866 11466 5871
rect 11158 5665 11186 5670
rect 11214 5697 11242 5703
rect 11214 5671 11215 5697
rect 11241 5671 11242 5697
rect 11102 5418 11130 5423
rect 11046 5417 11130 5418
rect 11046 5391 11103 5417
rect 11129 5391 11130 5417
rect 11046 5390 11130 5391
rect 11102 5385 11130 5390
rect 10990 4466 11018 4471
rect 10878 2977 10906 2982
rect 10934 3570 10962 3575
rect 10934 2954 10962 3542
rect 10934 2921 10962 2926
rect 10822 2641 10850 2646
rect 10934 2674 10962 2679
rect 10934 2627 10962 2646
rect 10654 2591 10655 2617
rect 10681 2591 10682 2617
rect 10654 2585 10682 2591
rect 10990 2506 11018 4438
rect 11102 4465 11130 4471
rect 11102 4439 11103 4465
rect 11129 4439 11130 4465
rect 11102 3402 11130 4439
rect 11102 3369 11130 3374
rect 10822 2478 11018 2506
rect 10374 1890 10402 1895
rect 10318 1862 10374 1890
rect 9814 1666 9898 1694
rect 9870 1106 9898 1666
rect 10262 1442 10290 1862
rect 10374 1857 10402 1862
rect 10262 1409 10290 1414
rect 9870 1073 9898 1078
rect 10654 1386 10682 1391
rect 10654 714 10682 1358
rect 10654 681 10682 686
rect 9254 546 9282 551
rect 9142 513 9170 518
rect 9198 518 9254 546
rect 9198 434 9226 518
rect 9254 513 9282 518
rect 10542 546 10570 551
rect 9086 406 9226 434
rect 10206 98 10234 103
rect 10206 56 10234 70
rect 10374 98 10402 103
rect 1456 0 1512 56
rect 2912 0 2968 56
rect 4368 0 4424 56
rect 5824 0 5880 56
rect 7280 0 7336 56
rect 8736 0 8792 56
rect 10192 0 10248 56
rect 10374 42 10402 70
rect 10542 42 10570 518
rect 10822 434 10850 2478
rect 11214 2282 11242 5671
rect 11214 2249 11242 2254
rect 11326 5138 11354 5143
rect 10878 1722 10906 1727
rect 10906 1694 10962 1722
rect 10878 1689 10906 1694
rect 10878 1274 10906 1279
rect 10878 770 10906 1246
rect 10878 737 10906 742
rect 10934 714 10962 1694
rect 11158 938 11186 943
rect 11158 891 11186 910
rect 10934 681 10962 686
rect 10822 401 10850 406
rect 11326 378 11354 5110
rect 11438 1105 11466 5838
rect 11494 2954 11522 6007
rect 11550 5641 11578 7056
rect 11662 6481 11690 6487
rect 11662 6455 11663 6481
rect 11689 6455 11690 6481
rect 11662 6370 11690 6455
rect 11662 6337 11690 6342
rect 11550 5615 11551 5641
rect 11577 5615 11578 5641
rect 11550 5609 11578 5615
rect 11774 5474 11802 7056
rect 11998 6594 12026 7056
rect 12222 6762 12250 7056
rect 11998 6561 12026 6566
rect 12166 6734 12250 6762
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11998 6202 12026 6207
rect 12166 6202 12194 6734
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 11998 6201 12194 6202
rect 11998 6175 11999 6201
rect 12025 6175 12194 6201
rect 11998 6174 12194 6175
rect 12446 6202 12474 7056
rect 12670 6706 12698 7056
rect 12502 6678 12698 6706
rect 12502 6593 12530 6678
rect 12502 6567 12503 6593
rect 12529 6567 12530 6593
rect 12502 6561 12530 6567
rect 12670 6482 12698 6487
rect 12558 6202 12586 6207
rect 12446 6201 12586 6202
rect 12446 6175 12559 6201
rect 12585 6175 12586 6201
rect 12446 6174 12586 6175
rect 11998 6169 12026 6174
rect 12558 6169 12586 6174
rect 12166 6089 12194 6095
rect 12166 6063 12167 6089
rect 12193 6063 12194 6089
rect 11998 5698 12026 5703
rect 11998 5651 12026 5670
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11774 5446 11858 5474
rect 11902 5469 12034 5474
rect 12110 5474 12138 5479
rect 11830 5418 11858 5446
rect 11998 5418 12026 5423
rect 11830 5417 12026 5418
rect 11830 5391 11999 5417
rect 12025 5391 12026 5417
rect 11830 5390 12026 5391
rect 11998 5385 12026 5390
rect 11774 5362 11802 5367
rect 11606 5306 11634 5311
rect 11606 5259 11634 5278
rect 11774 5026 11802 5334
rect 12110 5138 12138 5446
rect 12110 5105 12138 5110
rect 11774 4993 11802 4998
rect 12110 4746 12138 4751
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 12110 4354 12138 4718
rect 12166 4690 12194 6063
rect 12614 6090 12642 6095
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12446 5866 12474 5871
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12446 4746 12474 5838
rect 12614 5306 12642 6062
rect 12670 5418 12698 6454
rect 12782 6482 12810 6487
rect 12782 6481 12866 6482
rect 12782 6455 12783 6481
rect 12809 6455 12866 6481
rect 12782 6454 12866 6455
rect 12782 6449 12810 6454
rect 12782 5922 12810 5927
rect 12670 5385 12698 5390
rect 12726 5698 12754 5703
rect 12614 5273 12642 5278
rect 12502 5250 12530 5255
rect 12502 5249 12586 5250
rect 12502 5223 12503 5249
rect 12529 5223 12586 5249
rect 12502 5222 12586 5223
rect 12502 5217 12530 5222
rect 12558 5082 12586 5222
rect 12558 5054 12698 5082
rect 12446 4713 12474 4718
rect 12166 4657 12194 4662
rect 12614 4522 12642 4527
rect 12446 4354 12474 4359
rect 12110 4321 12138 4326
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 12446 4186 12474 4326
rect 12446 4153 12474 4158
rect 12558 4130 12586 4135
rect 12614 4130 12642 4494
rect 12586 4102 12642 4130
rect 12558 4097 12586 4102
rect 12614 4018 12642 4023
rect 12558 3990 12614 4018
rect 11902 3934 12034 3939
rect 11774 3906 11802 3911
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 11774 3066 11802 3878
rect 12222 3850 12250 3855
rect 12110 3822 12222 3850
rect 12110 3570 12138 3822
rect 12222 3817 12250 3822
rect 12558 3850 12586 3990
rect 12614 3985 12642 3990
rect 12558 3817 12586 3822
rect 12558 3738 12586 3743
rect 12446 3570 12474 3575
rect 12110 3537 12138 3542
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12446 3389 12474 3542
rect 12222 3361 12474 3389
rect 11830 3206 12138 3234
rect 11830 3178 11858 3206
rect 12110 3178 12138 3206
rect 11830 3145 11858 3150
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12110 3145 12138 3150
rect 11902 3117 12034 3122
rect 11774 3033 11802 3038
rect 11494 2921 11522 2926
rect 12222 2842 12250 3361
rect 12110 2814 12250 2842
rect 12446 3290 12474 3295
rect 12110 2730 12138 2814
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12110 2697 12138 2702
rect 12278 2618 12306 2623
rect 12446 2618 12474 3262
rect 12558 2673 12586 3710
rect 12670 2730 12698 5054
rect 12726 2786 12754 5670
rect 12782 3962 12810 5894
rect 12782 3929 12810 3934
rect 12726 2753 12754 2758
rect 12782 3794 12810 3799
rect 12670 2697 12698 2702
rect 12558 2647 12559 2673
rect 12585 2647 12586 2673
rect 12558 2641 12586 2647
rect 12278 2617 12474 2618
rect 12278 2591 12279 2617
rect 12305 2591 12474 2617
rect 12278 2590 12474 2591
rect 12278 2585 12306 2590
rect 12502 2562 12530 2567
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 11902 2333 12034 2338
rect 12110 2338 12138 2343
rect 11774 2002 11802 2007
rect 11774 1721 11802 1974
rect 11998 1890 12026 1895
rect 12110 1890 12138 2310
rect 12502 2002 12530 2534
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12502 1969 12530 1974
rect 12558 2114 12586 2119
rect 12232 1941 12364 1946
rect 11998 1889 12138 1890
rect 11998 1863 11999 1889
rect 12025 1863 12138 1889
rect 11998 1862 12138 1863
rect 11998 1857 12026 1862
rect 11774 1695 11775 1721
rect 11801 1695 11802 1721
rect 11774 1689 11802 1695
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 11438 1079 11439 1105
rect 11465 1079 11466 1105
rect 11438 1073 11466 1079
rect 12558 994 12586 2086
rect 12558 961 12586 966
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 12782 658 12810 3766
rect 12838 1050 12866 6454
rect 12894 5642 12922 7056
rect 13118 6146 13146 7056
rect 13286 6594 13314 6599
rect 13342 6594 13370 7056
rect 13566 6762 13594 7056
rect 13566 6729 13594 6734
rect 13286 6593 13370 6594
rect 13286 6567 13287 6593
rect 13313 6567 13370 6593
rect 13286 6566 13370 6567
rect 13286 6561 13314 6566
rect 13566 6481 13594 6487
rect 13566 6455 13567 6481
rect 13593 6455 13594 6481
rect 13118 6113 13146 6118
rect 13174 6258 13202 6263
rect 13062 6034 13090 6039
rect 13062 5987 13090 6006
rect 13118 5642 13146 5647
rect 12894 5641 13146 5642
rect 12894 5615 13119 5641
rect 13145 5615 13146 5641
rect 12894 5614 13146 5615
rect 13118 5609 13146 5614
rect 13174 2338 13202 6230
rect 13454 6146 13482 6151
rect 13454 6099 13482 6118
rect 13398 5642 13426 5647
rect 13398 4130 13426 5614
rect 13566 4746 13594 6455
rect 13734 6034 13762 6039
rect 13566 4713 13594 4718
rect 13622 5697 13650 5703
rect 13622 5671 13623 5697
rect 13649 5671 13650 5697
rect 13454 4578 13482 4583
rect 13454 4298 13482 4550
rect 13454 4265 13482 4270
rect 13398 4097 13426 4102
rect 13230 3934 13426 3962
rect 13230 2562 13258 3934
rect 13398 3850 13426 3934
rect 13566 3850 13594 3855
rect 13398 3822 13482 3850
rect 13454 3794 13482 3822
rect 13566 3794 13594 3822
rect 13454 3766 13594 3794
rect 13398 3654 13482 3682
rect 13286 3010 13314 3015
rect 13398 3010 13426 3654
rect 13454 3458 13482 3654
rect 13454 3425 13482 3430
rect 13566 3514 13594 3519
rect 13286 2963 13314 2982
rect 13342 2982 13426 3010
rect 13454 3346 13482 3351
rect 13454 3010 13482 3318
rect 13230 2529 13258 2534
rect 13342 2450 13370 2982
rect 13454 2977 13482 2982
rect 13566 2953 13594 3486
rect 13566 2927 13567 2953
rect 13593 2927 13594 2953
rect 13566 2921 13594 2927
rect 13398 2898 13426 2903
rect 13426 2870 13482 2898
rect 13398 2865 13426 2870
rect 13342 2417 13370 2422
rect 13398 2562 13426 2567
rect 13174 2305 13202 2310
rect 13398 1890 13426 2534
rect 13454 2450 13482 2870
rect 13454 2417 13482 2422
rect 13510 2506 13538 2511
rect 13398 1857 13426 1862
rect 13454 2058 13482 2063
rect 12838 1017 12866 1022
rect 13118 1834 13146 1839
rect 12782 625 12810 630
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 11326 345 11354 350
rect 11662 98 11690 103
rect 11662 56 11690 70
rect 13118 56 13146 1806
rect 13454 602 13482 2030
rect 13510 1386 13538 2478
rect 13510 1353 13538 1358
rect 13566 1554 13594 1559
rect 13454 569 13482 574
rect 13566 154 13594 1526
rect 13622 1106 13650 5671
rect 13678 5474 13706 5479
rect 13678 2674 13706 5446
rect 13734 4466 13762 6006
rect 13790 5978 13818 7056
rect 13958 6762 13986 6767
rect 13958 6425 13986 6734
rect 13958 6399 13959 6425
rect 13985 6399 13986 6425
rect 13958 6393 13986 6399
rect 13846 6034 13874 6039
rect 13846 5987 13874 6006
rect 13790 5945 13818 5950
rect 14014 5922 14042 7056
rect 13958 5894 14042 5922
rect 14126 6314 14154 6319
rect 13734 4433 13762 4438
rect 13790 5026 13818 5031
rect 13734 3346 13762 3351
rect 13734 2954 13762 3318
rect 13790 3178 13818 4998
rect 13790 3145 13818 3150
rect 13846 4970 13874 4975
rect 13734 2921 13762 2926
rect 13678 2641 13706 2646
rect 13846 2562 13874 4942
rect 13958 4018 13986 5894
rect 14014 5810 14042 5815
rect 14014 5763 14042 5782
rect 14070 5754 14098 5759
rect 14014 5698 14042 5703
rect 14014 4242 14042 5670
rect 14070 4970 14098 5726
rect 14070 4937 14098 4942
rect 14014 4209 14042 4214
rect 13958 3985 13986 3990
rect 14126 3906 14154 6286
rect 14238 5922 14266 7056
rect 14462 6874 14490 7056
rect 14462 6841 14490 6846
rect 14462 6481 14490 6487
rect 14462 6455 14463 6481
rect 14489 6455 14490 6481
rect 14238 5889 14266 5894
rect 14350 6370 14378 6375
rect 14294 5810 14322 5815
rect 14238 5642 14266 5647
rect 14238 5595 14266 5614
rect 14294 5474 14322 5782
rect 14294 5441 14322 5446
rect 14182 5418 14210 5423
rect 14182 4858 14210 5390
rect 14294 5362 14322 5367
rect 14182 4825 14210 4830
rect 14238 4914 14266 4919
rect 14126 3873 14154 3878
rect 14182 4746 14210 4751
rect 13846 2529 13874 2534
rect 14182 1162 14210 4718
rect 14238 4018 14266 4886
rect 14238 3985 14266 3990
rect 14294 2954 14322 5334
rect 14350 5082 14378 6342
rect 14462 6146 14490 6455
rect 14686 6202 14714 7056
rect 14910 6594 14938 7056
rect 14910 6566 14994 6594
rect 14462 6113 14490 6118
rect 14630 6174 14714 6202
rect 14910 6482 14938 6487
rect 14630 6034 14658 6174
rect 14910 6145 14938 6454
rect 14910 6119 14911 6145
rect 14937 6119 14938 6145
rect 14910 6113 14938 6119
rect 14350 5049 14378 5054
rect 14406 6006 14658 6034
rect 14686 6089 14714 6095
rect 14686 6063 14687 6089
rect 14713 6063 14714 6089
rect 14350 4354 14378 4359
rect 14350 4186 14378 4326
rect 14350 4153 14378 4158
rect 14406 3794 14434 6006
rect 14630 5362 14658 5367
rect 14518 4466 14546 4471
rect 14406 3761 14434 3766
rect 14462 4465 14546 4466
rect 14462 4439 14519 4465
rect 14545 4439 14546 4465
rect 14462 4438 14546 4439
rect 14294 2921 14322 2926
rect 14182 1129 14210 1134
rect 14238 2674 14266 2679
rect 13622 1073 13650 1078
rect 14238 266 14266 2646
rect 14462 1498 14490 4438
rect 14518 4433 14546 4438
rect 14518 3794 14546 3799
rect 14518 2617 14546 3766
rect 14518 2591 14519 2617
rect 14545 2591 14546 2617
rect 14518 2585 14546 2591
rect 14574 2786 14602 2791
rect 14462 1465 14490 1470
rect 14574 1498 14602 2758
rect 14630 2058 14658 5334
rect 14630 2025 14658 2030
rect 14686 1694 14714 6063
rect 14854 6090 14882 6095
rect 14798 4522 14826 4527
rect 14798 4475 14826 4494
rect 14854 3514 14882 6062
rect 14910 4746 14938 4751
rect 14910 3850 14938 4718
rect 14910 3817 14938 3822
rect 14966 3738 14994 6566
rect 15022 5194 15050 5199
rect 15022 3850 15050 5166
rect 15134 4522 15162 7056
rect 15358 6258 15386 7056
rect 15582 6986 15610 7056
rect 15582 6953 15610 6958
rect 15358 6225 15386 6230
rect 15470 6370 15498 6375
rect 15190 6146 15218 6151
rect 15190 6099 15218 6118
rect 15470 6089 15498 6342
rect 15470 6063 15471 6089
rect 15497 6063 15498 6089
rect 15470 6057 15498 6063
rect 15694 6034 15722 6039
rect 15358 5978 15386 5983
rect 15134 4489 15162 4494
rect 15190 4634 15218 4639
rect 15078 4130 15106 4135
rect 15078 3906 15106 4102
rect 15078 3873 15106 3878
rect 15022 3817 15050 3822
rect 14966 3705 14994 3710
rect 14854 3481 14882 3486
rect 15134 3290 15162 3295
rect 15190 3290 15218 4606
rect 15134 3289 15218 3290
rect 15134 3263 15135 3289
rect 15161 3263 15218 3289
rect 15134 3262 15218 3263
rect 15246 4354 15274 4359
rect 15134 3257 15162 3262
rect 14798 3234 14826 3239
rect 14798 3009 14826 3206
rect 14798 2983 14799 3009
rect 14825 2983 14826 3009
rect 14798 2977 14826 2983
rect 15078 2898 15106 2903
rect 15078 2851 15106 2870
rect 14798 2561 14826 2567
rect 14798 2535 14799 2561
rect 14825 2535 14826 2561
rect 14686 1666 14770 1694
rect 14574 1465 14602 1470
rect 14742 1330 14770 1666
rect 14742 1297 14770 1302
rect 14406 770 14434 775
rect 14406 546 14434 742
rect 14406 513 14434 518
rect 14238 233 14266 238
rect 14574 266 14602 271
rect 13566 121 13594 126
rect 14574 56 14602 238
rect 14798 98 14826 2535
rect 15246 2506 15274 4326
rect 15358 3457 15386 5950
rect 15414 5922 15442 5927
rect 15414 5586 15442 5894
rect 15414 5558 15554 5586
rect 15358 3431 15359 3457
rect 15385 3431 15386 3457
rect 15358 3425 15386 3431
rect 15470 5082 15498 5087
rect 15246 2473 15274 2478
rect 15414 2506 15442 2511
rect 15134 2226 15162 2231
rect 15134 546 15162 2198
rect 15414 1105 15442 2478
rect 15414 1079 15415 1105
rect 15441 1079 15442 1105
rect 15414 1073 15442 1079
rect 15246 993 15274 999
rect 15246 967 15247 993
rect 15273 967 15274 993
rect 15246 882 15274 967
rect 15246 849 15274 854
rect 15358 994 15386 999
rect 15358 882 15386 966
rect 15358 849 15386 854
rect 15470 826 15498 5054
rect 15526 1694 15554 5558
rect 15582 5362 15610 5367
rect 15582 3794 15610 5334
rect 15582 3761 15610 3766
rect 15526 1666 15610 1694
rect 15582 1554 15610 1666
rect 15582 1521 15610 1526
rect 15694 1218 15722 6006
rect 15806 2618 15834 7056
rect 16030 6314 16058 7056
rect 16254 7042 16282 7056
rect 16254 7009 16282 7014
rect 16030 6281 16058 6286
rect 15918 6034 15946 6039
rect 15918 5698 15946 6006
rect 15918 5665 15946 5670
rect 16198 5586 16226 5591
rect 15974 4410 16002 4415
rect 15974 4298 16002 4382
rect 16198 4354 16226 5558
rect 16198 4321 16226 4326
rect 16366 5530 16394 5535
rect 15974 4265 16002 4270
rect 15918 3458 15946 3463
rect 15918 3010 15946 3430
rect 15918 2977 15946 2982
rect 16310 3122 16338 3127
rect 15806 2585 15834 2590
rect 16310 1694 16338 3094
rect 16366 2786 16394 5502
rect 16366 2753 16394 2758
rect 16366 2618 16394 2623
rect 16366 2394 16394 2590
rect 16366 2361 16394 2366
rect 16478 2338 16506 7056
rect 16478 2305 16506 2310
rect 16534 6538 16562 6543
rect 16534 1694 16562 6510
rect 16310 1666 16394 1694
rect 16366 1610 16394 1666
rect 16366 1577 16394 1582
rect 16478 1666 16562 1694
rect 16590 6202 16618 6207
rect 15694 1185 15722 1190
rect 16478 1105 16506 1666
rect 16478 1079 16479 1105
rect 16505 1079 16506 1105
rect 16478 1073 16506 1079
rect 16198 938 16226 943
rect 16198 891 16226 910
rect 15470 793 15498 798
rect 16590 658 16618 6174
rect 16646 5530 16674 5535
rect 16646 5082 16674 5502
rect 16702 5138 16730 7056
rect 16814 6258 16842 6263
rect 16814 5250 16842 6230
rect 16814 5217 16842 5222
rect 16702 5110 16842 5138
rect 16646 5049 16674 5054
rect 16814 4858 16842 5110
rect 16814 4825 16842 4830
rect 16926 4858 16954 7056
rect 17150 5250 17178 7056
rect 17150 5217 17178 5222
rect 16926 4825 16954 4830
rect 16982 5138 17010 5143
rect 16702 4802 16730 4807
rect 16702 4746 16730 4774
rect 16982 4746 17010 5110
rect 16702 4718 16842 4746
rect 16814 3514 16842 4718
rect 16982 4713 17010 4718
rect 16870 4354 16898 4359
rect 16870 4186 16898 4326
rect 16870 4153 16898 4158
rect 16814 3481 16842 3486
rect 17374 3234 17402 7056
rect 17486 6706 17514 6711
rect 17486 4186 17514 6678
rect 17598 6594 17626 7056
rect 17598 6561 17626 6566
rect 17654 6089 17682 6095
rect 17654 6063 17655 6089
rect 17681 6063 17682 6089
rect 17654 5922 17682 6063
rect 17654 5889 17682 5894
rect 17822 5698 17850 7056
rect 17822 5665 17850 5670
rect 17878 6033 17906 6039
rect 17878 6007 17879 6033
rect 17905 6007 17906 6033
rect 17878 5306 17906 6007
rect 17878 5273 17906 5278
rect 17710 4970 17738 4975
rect 17598 4746 17626 4751
rect 17486 4153 17514 4158
rect 17542 4634 17570 4639
rect 17486 4074 17514 4079
rect 17430 3738 17458 3743
rect 17430 3691 17458 3710
rect 17374 3201 17402 3206
rect 16702 1946 16730 1951
rect 16702 1834 16730 1918
rect 16702 1801 16730 1806
rect 16814 1946 16842 1951
rect 16814 1722 16842 1918
rect 16814 1689 16842 1694
rect 16590 625 16618 630
rect 16758 938 16786 943
rect 15134 513 15162 518
rect 15974 434 16002 439
rect 15974 322 16002 406
rect 16086 322 16114 327
rect 15974 289 16002 294
rect 16030 294 16086 322
rect 14798 65 14826 70
rect 16030 56 16058 294
rect 16086 289 16114 294
rect 10374 14 10570 42
rect 11648 0 11704 56
rect 13104 0 13160 56
rect 14560 0 14616 56
rect 16016 0 16072 56
rect 16758 42 16786 910
rect 17486 490 17514 4046
rect 17542 3850 17570 4606
rect 17598 4018 17626 4718
rect 17598 3985 17626 3990
rect 17654 4634 17682 4639
rect 17654 3906 17682 4606
rect 17654 3873 17682 3878
rect 17542 3822 17626 3850
rect 17542 3738 17570 3743
rect 17542 2842 17570 3710
rect 17598 3570 17626 3822
rect 17710 3794 17738 4942
rect 18046 4970 18074 7056
rect 18270 6818 18298 7056
rect 18270 6785 18298 6790
rect 18046 4937 18074 4942
rect 18214 5250 18242 5255
rect 17766 4690 17794 4695
rect 17766 3906 17794 4662
rect 18214 4690 18242 5222
rect 18214 4657 18242 4662
rect 17766 3873 17794 3878
rect 18382 4410 18410 4415
rect 17710 3761 17738 3766
rect 17710 3682 17738 3687
rect 17710 3635 17738 3654
rect 17598 3542 17738 3570
rect 17542 2809 17570 2814
rect 17542 2002 17570 2007
rect 17542 602 17570 1974
rect 17654 1778 17682 1783
rect 17654 1274 17682 1750
rect 17598 1246 17682 1274
rect 17598 826 17626 1246
rect 17654 1162 17682 1167
rect 17654 1049 17682 1134
rect 17654 1023 17655 1049
rect 17681 1023 17682 1049
rect 17654 1017 17682 1023
rect 17598 793 17626 798
rect 17710 714 17738 3542
rect 18046 3458 18074 3463
rect 17990 2842 18018 2847
rect 17822 2282 17850 2287
rect 17822 770 17850 2254
rect 17934 1666 17962 1671
rect 17878 1610 17906 1615
rect 17878 1162 17906 1582
rect 17878 1129 17906 1134
rect 17934 1105 17962 1638
rect 17934 1079 17935 1105
rect 17961 1079 17962 1105
rect 17934 1073 17962 1079
rect 17990 938 18018 2814
rect 18046 1946 18074 3430
rect 18158 3290 18186 3295
rect 18158 3243 18186 3262
rect 18046 1913 18074 1918
rect 18214 2954 18242 2959
rect 18214 1610 18242 2926
rect 18382 2506 18410 4382
rect 18438 4298 18466 4303
rect 18438 3850 18466 4270
rect 18438 3817 18466 3822
rect 18438 3346 18466 3351
rect 18494 3346 18522 7056
rect 18662 6314 18690 6319
rect 18550 5474 18578 5479
rect 18550 4242 18578 5446
rect 18550 4209 18578 4214
rect 18606 4690 18634 4695
rect 18438 3345 18522 3346
rect 18438 3319 18439 3345
rect 18465 3319 18522 3345
rect 18438 3318 18522 3319
rect 18550 3682 18578 3687
rect 18438 3313 18466 3318
rect 18550 2954 18578 3654
rect 18606 3346 18634 4662
rect 18662 4410 18690 6286
rect 18718 6090 18746 7056
rect 18718 6057 18746 6062
rect 18942 5978 18970 7056
rect 18942 5945 18970 5950
rect 18998 6986 19026 6991
rect 18662 4377 18690 4382
rect 18606 3313 18634 3318
rect 18886 3402 18914 3407
rect 18382 2473 18410 2478
rect 18438 2926 18578 2954
rect 18214 1577 18242 1582
rect 18270 2450 18298 2455
rect 18158 1106 18186 1111
rect 18158 1049 18186 1078
rect 18158 1023 18159 1049
rect 18185 1023 18186 1049
rect 18158 1017 18186 1023
rect 17990 905 18018 910
rect 17822 737 17850 742
rect 17710 681 17738 686
rect 18270 658 18298 2422
rect 18438 2170 18466 2926
rect 18438 2137 18466 2142
rect 18438 1106 18466 1111
rect 18438 1059 18466 1078
rect 18774 1050 18802 1055
rect 18774 1003 18802 1022
rect 18886 1050 18914 3374
rect 18998 1694 19026 6958
rect 19110 6426 19138 6431
rect 19054 5978 19082 5983
rect 19054 5586 19082 5950
rect 19054 5553 19082 5558
rect 19110 3374 19138 6398
rect 19166 6034 19194 7056
rect 19390 6258 19418 7056
rect 19390 6225 19418 6230
rect 19166 6001 19194 6006
rect 19614 5810 19642 7056
rect 19838 6650 19866 7056
rect 19838 6617 19866 6622
rect 19614 5777 19642 5782
rect 19558 5698 19586 5703
rect 19446 5530 19474 5535
rect 19334 3570 19362 3575
rect 19110 3346 19250 3374
rect 18942 1666 19026 1694
rect 19222 1666 19250 3346
rect 19334 2226 19362 3542
rect 19334 2193 19362 2198
rect 19446 1890 19474 5502
rect 19502 4802 19530 4807
rect 19502 2674 19530 4774
rect 19558 3850 19586 5670
rect 20006 5194 20034 5199
rect 19558 3817 19586 3822
rect 19614 5138 19642 5143
rect 19502 2641 19530 2646
rect 19614 2282 19642 5110
rect 19782 4578 19810 4583
rect 19782 2954 19810 4550
rect 20006 3794 20034 5166
rect 20006 3761 20034 3766
rect 20062 3738 20090 7056
rect 20174 6202 20202 6207
rect 20174 5810 20202 6174
rect 20174 5777 20202 5782
rect 20062 3705 20090 3710
rect 20174 4690 20202 4695
rect 20118 3458 20146 3463
rect 20118 3290 20146 3430
rect 20118 3257 20146 3262
rect 19782 2921 19810 2926
rect 20174 2673 20202 4662
rect 20230 4466 20258 4471
rect 20230 4419 20258 4438
rect 20286 4074 20314 7056
rect 20510 6090 20538 7056
rect 20510 6057 20538 6062
rect 20678 6090 20706 6095
rect 20678 6043 20706 6062
rect 20398 5978 20426 5983
rect 20398 5931 20426 5950
rect 20566 4970 20594 4975
rect 20342 4634 20370 4639
rect 20342 4410 20370 4606
rect 20566 4634 20594 4942
rect 20566 4601 20594 4606
rect 20510 4522 20538 4527
rect 20510 4475 20538 4494
rect 20342 4377 20370 4382
rect 20286 4041 20314 4046
rect 20622 4298 20650 4303
rect 20622 3738 20650 4270
rect 20622 3705 20650 3710
rect 20678 4242 20706 4247
rect 20174 2647 20175 2673
rect 20201 2647 20202 2673
rect 20174 2641 20202 2647
rect 20454 3178 20482 3183
rect 20454 2617 20482 3150
rect 20454 2591 20455 2617
rect 20481 2591 20482 2617
rect 20454 2585 20482 2591
rect 19614 2249 19642 2254
rect 20230 2562 20258 2567
rect 19446 1857 19474 1862
rect 20174 1722 20202 1727
rect 20174 1675 20202 1694
rect 18942 1106 18970 1666
rect 19222 1633 19250 1638
rect 20230 1666 20258 2534
rect 20230 1633 20258 1638
rect 20342 2562 20370 2567
rect 19726 1386 19754 1391
rect 18942 1073 18970 1078
rect 19446 1218 19474 1223
rect 18886 1017 18914 1022
rect 19446 1049 19474 1190
rect 19726 1105 19754 1358
rect 20342 1274 20370 2534
rect 20398 2282 20426 2287
rect 20398 1889 20426 2254
rect 20398 1863 20399 1889
rect 20425 1863 20426 1889
rect 20398 1857 20426 1863
rect 20342 1246 20426 1274
rect 19726 1079 19727 1105
rect 19753 1079 19754 1105
rect 19726 1073 19754 1079
rect 19446 1023 19447 1049
rect 19473 1023 19474 1049
rect 19446 1017 19474 1023
rect 19054 994 19082 999
rect 19054 947 19082 966
rect 18270 625 18298 630
rect 18438 938 18466 943
rect 17542 569 17570 574
rect 18438 546 18466 910
rect 20286 938 20314 943
rect 20286 770 20314 910
rect 20286 737 20314 742
rect 18438 513 18466 518
rect 18942 658 18970 663
rect 17486 457 17514 462
rect 17486 154 17514 159
rect 17486 56 17514 126
rect 18942 56 18970 630
rect 20398 56 20426 1246
rect 20622 1050 20650 1055
rect 20622 1003 20650 1022
rect 20678 434 20706 4214
rect 20734 2002 20762 7056
rect 20958 6314 20986 7056
rect 20958 6281 20986 6286
rect 20958 6202 20986 6207
rect 20734 1969 20762 1974
rect 20790 5922 20818 5927
rect 20790 1218 20818 5894
rect 20958 4018 20986 6174
rect 20958 3985 20986 3990
rect 21126 5474 21154 5479
rect 20846 3906 20874 3911
rect 20846 3793 20874 3878
rect 20846 3767 20847 3793
rect 20873 3767 20874 3793
rect 20846 3761 20874 3767
rect 21126 3737 21154 5446
rect 21126 3711 21127 3737
rect 21153 3711 21154 3737
rect 21126 3705 21154 3711
rect 21182 2786 21210 7056
rect 21126 2758 21210 2786
rect 21238 5754 21266 5759
rect 20902 2730 20930 2735
rect 20902 2617 20930 2702
rect 20902 2591 20903 2617
rect 20929 2591 20930 2617
rect 20902 2585 20930 2591
rect 21014 2113 21042 2119
rect 21014 2087 21015 2113
rect 21041 2087 21042 2113
rect 21014 1778 21042 2087
rect 21014 1745 21042 1750
rect 20790 1185 20818 1190
rect 20902 1442 20930 1447
rect 20902 1105 20930 1414
rect 20902 1079 20903 1105
rect 20929 1079 20930 1105
rect 20902 1073 20930 1079
rect 21070 1330 21098 1335
rect 21070 1049 21098 1302
rect 21070 1023 21071 1049
rect 21097 1023 21098 1049
rect 21070 1017 21098 1023
rect 20678 401 20706 406
rect 21126 378 21154 2758
rect 21182 2674 21210 2679
rect 21182 2627 21210 2646
rect 21238 1778 21266 5726
rect 21406 2898 21434 7056
rect 21630 6538 21658 7056
rect 21630 6505 21658 6510
rect 21854 6370 21882 7056
rect 22078 6426 22106 7056
rect 22302 6762 22330 7056
rect 22526 6986 22554 7056
rect 22526 6953 22554 6958
rect 22302 6734 22442 6762
rect 22232 6678 22364 6683
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22232 6645 22364 6650
rect 22078 6393 22106 6398
rect 21854 6337 21882 6342
rect 21902 6286 22034 6291
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 21902 6253 22034 6258
rect 21798 6034 21826 6039
rect 21798 5987 21826 6006
rect 21518 5978 21546 5983
rect 21462 5977 21546 5978
rect 21462 5951 21519 5977
rect 21545 5951 21546 5977
rect 21462 5950 21546 5951
rect 22414 5978 22442 6734
rect 22638 6146 22666 6151
rect 22414 5950 22554 5978
rect 21462 5082 21490 5950
rect 21518 5945 21546 5950
rect 22232 5894 22364 5899
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22232 5861 22364 5866
rect 22470 5866 22498 5871
rect 21902 5502 22034 5507
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 21902 5469 22034 5474
rect 21798 5250 21826 5255
rect 21798 5203 21826 5222
rect 21518 5193 21546 5199
rect 21518 5167 21519 5193
rect 21545 5167 21546 5193
rect 21518 5138 21546 5167
rect 21518 5105 21546 5110
rect 22232 5110 22364 5115
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22232 5077 22364 5082
rect 21462 5049 21490 5054
rect 21902 4718 22034 4723
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 21902 4685 22034 4690
rect 22232 4326 22364 4331
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22232 4293 22364 4298
rect 21966 4129 21994 4135
rect 21966 4103 21967 4129
rect 21993 4103 21994 4129
rect 21742 4074 21770 4079
rect 21742 4027 21770 4046
rect 21966 4018 21994 4103
rect 21966 3985 21994 3990
rect 21902 3934 22034 3939
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 21902 3901 22034 3906
rect 22232 3542 22364 3547
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22232 3509 22364 3514
rect 21406 2865 21434 2870
rect 21742 3402 21770 3407
rect 21742 2617 21770 3374
rect 21902 3150 22034 3155
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 21902 3117 22034 3122
rect 22078 2898 22106 2903
rect 22078 2851 22106 2870
rect 22358 2898 22386 2903
rect 22358 2851 22386 2870
rect 22232 2758 22364 2763
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22232 2725 22364 2730
rect 22470 2674 22498 5838
rect 22470 2641 22498 2646
rect 21742 2591 21743 2617
rect 21769 2591 21770 2617
rect 21742 2585 21770 2591
rect 21462 2561 21490 2567
rect 21462 2535 21463 2561
rect 21489 2535 21490 2561
rect 21462 2338 21490 2535
rect 22470 2450 22498 2455
rect 21902 2366 22034 2371
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 21902 2333 22034 2338
rect 21462 2305 21490 2310
rect 21294 2170 21322 2175
rect 21294 2123 21322 2142
rect 22232 1974 22364 1979
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22232 1941 22364 1946
rect 22190 1834 22218 1839
rect 22190 1787 22218 1806
rect 22470 1833 22498 2422
rect 22470 1807 22471 1833
rect 22497 1807 22498 1833
rect 22470 1801 22498 1807
rect 21238 1745 21266 1750
rect 21518 1610 21546 1615
rect 21350 1330 21378 1335
rect 21350 1105 21378 1302
rect 21350 1079 21351 1105
rect 21377 1079 21378 1105
rect 21350 1073 21378 1079
rect 21518 1049 21546 1582
rect 21902 1582 22034 1587
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 21902 1549 22034 1554
rect 22078 1554 22106 1559
rect 21798 1106 21826 1111
rect 21798 1059 21826 1078
rect 22022 1106 22050 1111
rect 22078 1106 22106 1526
rect 22526 1386 22554 5950
rect 22582 5922 22610 5927
rect 22582 2170 22610 5894
rect 22638 5642 22666 6118
rect 22638 5609 22666 5614
rect 22638 4298 22666 4303
rect 22638 3290 22666 4270
rect 22638 3257 22666 3262
rect 22582 2137 22610 2142
rect 22526 1353 22554 1358
rect 22582 2002 22610 2007
rect 22232 1190 22364 1195
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22232 1157 22364 1162
rect 22050 1078 22106 1106
rect 22022 1073 22050 1078
rect 21518 1023 21519 1049
rect 21545 1023 21546 1049
rect 21518 1017 21546 1023
rect 21902 798 22034 803
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 21902 765 22034 770
rect 22582 658 22610 1974
rect 22638 1834 22666 1839
rect 22638 1442 22666 1806
rect 22638 1409 22666 1414
rect 22694 1498 22722 1503
rect 22582 625 22610 630
rect 22638 994 22666 999
rect 22232 406 22364 411
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22232 373 22364 378
rect 21126 345 21154 350
rect 22638 322 22666 966
rect 22694 937 22722 1470
rect 22750 1050 22778 7056
rect 22974 4522 23002 7056
rect 23142 5642 23170 5647
rect 23142 5595 23170 5614
rect 23198 5194 23226 7056
rect 23254 6594 23282 6599
rect 23254 5474 23282 6566
rect 23422 5922 23450 7056
rect 23422 5889 23450 5894
rect 23478 6202 23506 6207
rect 23254 5441 23282 5446
rect 23310 5866 23338 5871
rect 23198 5161 23226 5166
rect 23310 4858 23338 5838
rect 23366 5697 23394 5703
rect 23366 5671 23367 5697
rect 23393 5671 23394 5697
rect 23366 5082 23394 5671
rect 23478 5138 23506 6174
rect 23646 5978 23674 7056
rect 23646 5945 23674 5950
rect 23478 5105 23506 5110
rect 23646 5698 23674 5703
rect 23366 5049 23394 5054
rect 23310 4825 23338 4830
rect 22974 4489 23002 4494
rect 23422 4018 23450 4023
rect 23366 3402 23394 3407
rect 22750 1017 22778 1022
rect 22806 2842 22834 2847
rect 22694 911 22695 937
rect 22721 911 22722 937
rect 22694 905 22722 911
rect 22694 826 22722 831
rect 22694 658 22722 798
rect 22694 625 22722 630
rect 22638 289 22666 294
rect 22806 322 22834 2814
rect 23254 2058 23282 2063
rect 23254 1833 23282 2030
rect 23254 1807 23255 1833
rect 23281 1807 23282 1833
rect 23254 1801 23282 1807
rect 23366 1610 23394 3374
rect 23366 1577 23394 1582
rect 23422 1442 23450 3990
rect 23478 3794 23506 3799
rect 23478 3234 23506 3766
rect 23534 3346 23562 3351
rect 23534 3299 23562 3318
rect 23478 3206 23562 3234
rect 23478 2506 23506 2511
rect 23478 1777 23506 2478
rect 23478 1751 23479 1777
rect 23505 1751 23506 1777
rect 23478 1745 23506 1751
rect 23422 1409 23450 1414
rect 23534 1218 23562 3206
rect 23646 1834 23674 5670
rect 23814 4409 23842 4415
rect 23814 4383 23815 4409
rect 23841 4383 23842 4409
rect 23702 3289 23730 3295
rect 23702 3263 23703 3289
rect 23729 3263 23730 3289
rect 23702 3010 23730 3263
rect 23702 2977 23730 2982
rect 23814 2002 23842 4383
rect 23814 1969 23842 1974
rect 23646 1801 23674 1806
rect 23870 1330 23898 7056
rect 24094 5698 24122 7056
rect 24094 5665 24122 5670
rect 24318 5642 24346 7056
rect 24542 6650 24570 7056
rect 24206 5614 24346 5642
rect 24486 6622 24570 6650
rect 23982 5026 24010 5031
rect 23982 2338 24010 4998
rect 24094 5026 24122 5031
rect 24094 4577 24122 4998
rect 24094 4551 24095 4577
rect 24121 4551 24122 4577
rect 24094 4545 24122 4551
rect 24206 4214 24234 5614
rect 23982 2305 24010 2310
rect 24038 4186 24234 4214
rect 24262 4410 24290 4415
rect 24038 1554 24066 4186
rect 24262 2842 24290 4382
rect 24318 4298 24346 4303
rect 24318 3290 24346 4270
rect 24318 3257 24346 3262
rect 24262 2809 24290 2814
rect 24374 2898 24402 2903
rect 24038 1521 24066 1526
rect 24206 2674 24234 2679
rect 23870 1297 23898 1302
rect 23534 1185 23562 1190
rect 22918 1106 22946 1111
rect 22918 1059 22946 1078
rect 24038 993 24066 999
rect 24038 967 24039 993
rect 24065 967 24066 993
rect 23478 938 23506 943
rect 23478 490 23506 910
rect 23478 457 23506 462
rect 22806 289 22834 294
rect 24038 266 24066 967
rect 24206 826 24234 2646
rect 24318 2618 24346 2623
rect 24262 2114 24290 2119
rect 24262 2067 24290 2086
rect 24318 1834 24346 2590
rect 24374 2394 24402 2870
rect 24374 2361 24402 2366
rect 24318 1801 24346 1806
rect 24318 1498 24346 1503
rect 24318 1049 24346 1470
rect 24486 1106 24514 6622
rect 24766 4214 24794 7056
rect 24990 4214 25018 7056
rect 24542 4186 24794 4214
rect 24934 4186 25018 4214
rect 25158 4298 25186 4303
rect 24542 2169 24570 4186
rect 24934 2506 24962 4186
rect 25158 3402 25186 4270
rect 25214 4214 25242 7056
rect 25438 6593 25466 7056
rect 25438 6567 25439 6593
rect 25465 6567 25466 6593
rect 25438 6561 25466 6567
rect 25662 6594 25690 7056
rect 25662 6561 25690 6566
rect 25606 6481 25634 6487
rect 25606 6455 25607 6481
rect 25633 6455 25634 6481
rect 25550 5082 25578 5087
rect 25214 4186 25298 4214
rect 25158 3369 25186 3374
rect 25214 3345 25242 3351
rect 25214 3319 25215 3345
rect 25241 3319 25242 3345
rect 25214 2674 25242 3319
rect 24934 2473 24962 2478
rect 25158 2646 25242 2674
rect 25158 2450 25186 2646
rect 25214 2562 25242 2567
rect 25214 2515 25242 2534
rect 25158 2422 25242 2450
rect 24542 2143 24543 2169
rect 24569 2143 24570 2169
rect 24542 2137 24570 2143
rect 24766 2282 24794 2287
rect 24486 1073 24514 1078
rect 24318 1023 24319 1049
rect 24345 1023 24346 1049
rect 24318 1017 24346 1023
rect 24598 994 24626 999
rect 24598 947 24626 966
rect 24206 793 24234 798
rect 24038 233 24066 238
rect 23310 210 23338 215
rect 21854 98 21882 103
rect 21854 56 21882 70
rect 23310 56 23338 182
rect 24766 56 24794 2254
rect 24990 1890 25018 1895
rect 24990 1833 25018 1862
rect 24990 1807 24991 1833
rect 25017 1807 25018 1833
rect 24990 1801 25018 1807
rect 25214 1106 25242 2422
rect 25270 1889 25298 4186
rect 25494 3346 25522 3351
rect 25494 3299 25522 3318
rect 25438 3066 25466 3071
rect 25326 2786 25354 2791
rect 25326 2562 25354 2758
rect 25438 2617 25466 3038
rect 25438 2591 25439 2617
rect 25465 2591 25466 2617
rect 25438 2585 25466 2591
rect 25326 2529 25354 2534
rect 25270 1863 25271 1889
rect 25297 1863 25298 1889
rect 25270 1857 25298 1863
rect 25438 1610 25466 1615
rect 25214 1078 25298 1106
rect 24878 1050 24906 1055
rect 24878 1003 24906 1022
rect 25214 993 25242 999
rect 25214 967 25215 993
rect 25241 967 25242 993
rect 24878 434 24906 439
rect 24878 322 24906 406
rect 24878 289 24906 294
rect 25214 154 25242 967
rect 25214 121 25242 126
rect 25270 98 25298 1078
rect 25438 1049 25466 1582
rect 25438 1023 25439 1049
rect 25465 1023 25466 1049
rect 25438 1017 25466 1023
rect 25550 602 25578 5054
rect 25606 1666 25634 6455
rect 25774 6481 25802 6487
rect 25774 6455 25775 6481
rect 25801 6455 25802 6481
rect 25774 6146 25802 6455
rect 25886 6202 25914 7056
rect 26054 6594 26082 6599
rect 26054 6547 26082 6566
rect 25886 6169 25914 6174
rect 26054 6482 26082 6487
rect 25774 6113 25802 6118
rect 26054 6089 26082 6454
rect 26054 6063 26055 6089
rect 26081 6063 26082 6089
rect 26054 6057 26082 6063
rect 26110 5810 26138 7056
rect 26334 6538 26362 7056
rect 26558 6762 26586 7056
rect 26558 6729 26586 6734
rect 26334 6505 26362 6510
rect 26782 6370 26810 7056
rect 26782 6342 26866 6370
rect 26558 6258 26586 6263
rect 26278 6202 26306 6207
rect 26278 6155 26306 6174
rect 26502 5810 26530 5815
rect 26110 5809 26530 5810
rect 26110 5783 26503 5809
rect 26529 5783 26530 5809
rect 26110 5782 26530 5783
rect 26502 5777 26530 5782
rect 26222 5697 26250 5703
rect 26222 5671 26223 5697
rect 26249 5671 26250 5697
rect 26222 5306 26250 5671
rect 26222 5273 26250 5278
rect 26390 4634 26418 4639
rect 26390 4521 26418 4606
rect 26390 4495 26391 4521
rect 26417 4495 26418 4521
rect 26390 4489 26418 4495
rect 26558 4214 26586 6230
rect 26782 6090 26810 6095
rect 26782 6043 26810 6062
rect 26838 5866 26866 6342
rect 26838 5833 26866 5838
rect 26894 6202 26922 6207
rect 26614 5138 26642 5143
rect 26614 4577 26642 5110
rect 26614 4551 26615 4577
rect 26641 4551 26642 4577
rect 26614 4545 26642 4551
rect 26894 4410 26922 6174
rect 27006 6202 27034 7056
rect 27230 6594 27258 7056
rect 27454 6874 27482 7056
rect 27678 6930 27706 7056
rect 27678 6897 27706 6902
rect 27454 6841 27482 6846
rect 27230 6561 27258 6566
rect 27454 6762 27482 6767
rect 27454 6593 27482 6734
rect 27454 6567 27455 6593
rect 27481 6567 27482 6593
rect 27454 6561 27482 6567
rect 27006 6169 27034 6174
rect 27062 6538 27090 6543
rect 27062 6201 27090 6510
rect 27062 6175 27063 6201
rect 27089 6175 27090 6201
rect 27062 6169 27090 6175
rect 27174 6481 27202 6487
rect 27174 6455 27175 6481
rect 27201 6455 27202 6481
rect 27174 6034 27202 6455
rect 27902 6426 27930 7056
rect 27902 6393 27930 6398
rect 27958 6481 27986 6487
rect 27958 6455 27959 6481
rect 27985 6455 27986 6481
rect 27958 6258 27986 6455
rect 27958 6225 27986 6230
rect 27846 6202 27874 6207
rect 27846 6155 27874 6174
rect 28126 6146 28154 7056
rect 28126 6113 28154 6118
rect 28182 6930 28210 6935
rect 27174 6001 27202 6006
rect 27566 6033 27594 6039
rect 27566 6007 27567 6033
rect 27593 6007 27594 6033
rect 27286 5866 27314 5871
rect 27286 5809 27314 5838
rect 27286 5783 27287 5809
rect 27313 5783 27314 5809
rect 27286 5777 27314 5783
rect 27006 5697 27034 5703
rect 27006 5671 27007 5697
rect 27033 5671 27034 5697
rect 27006 5250 27034 5671
rect 27006 5217 27034 5222
rect 26894 4377 26922 4382
rect 26446 4186 26586 4214
rect 26446 2450 26474 4186
rect 26950 2730 26978 2735
rect 26446 2417 26474 2422
rect 26670 2506 26698 2511
rect 25606 1633 25634 1638
rect 26054 2226 26082 2231
rect 26054 1666 26082 2198
rect 26054 1633 26082 1638
rect 26054 1554 26082 1559
rect 26054 1441 26082 1526
rect 26670 1498 26698 2478
rect 26670 1465 26698 1470
rect 26054 1415 26055 1441
rect 26081 1415 26082 1441
rect 26054 1409 26082 1415
rect 26222 1442 26250 1447
rect 25550 569 25578 574
rect 26054 1162 26082 1167
rect 26054 490 26082 1134
rect 26054 457 26082 462
rect 25270 65 25298 70
rect 26222 56 26250 1414
rect 26278 1273 26306 1279
rect 26278 1247 26279 1273
rect 26305 1247 26306 1273
rect 26278 882 26306 1247
rect 26278 849 26306 854
rect 26894 994 26922 999
rect 26894 546 26922 966
rect 26950 826 26978 2702
rect 27174 2450 27202 2455
rect 27174 1610 27202 2422
rect 27566 2394 27594 6007
rect 28182 5810 28210 6902
rect 28238 6594 28266 6599
rect 28238 6547 28266 6566
rect 28350 6482 28378 7056
rect 28574 6538 28602 7056
rect 28574 6505 28602 6510
rect 28630 6874 28658 6879
rect 28350 6449 28378 6454
rect 28630 6201 28658 6846
rect 28630 6175 28631 6201
rect 28657 6175 28658 6201
rect 28630 6169 28658 6175
rect 28574 6146 28602 6151
rect 28350 6034 28378 6039
rect 28294 6033 28378 6034
rect 28294 6007 28351 6033
rect 28377 6007 28378 6033
rect 28294 6006 28378 6007
rect 28238 5810 28266 5815
rect 28182 5809 28266 5810
rect 28182 5783 28239 5809
rect 28265 5783 28266 5809
rect 28182 5782 28266 5783
rect 28238 5777 28266 5782
rect 28014 5697 28042 5703
rect 28014 5671 28015 5697
rect 28041 5671 28042 5697
rect 27734 5530 27762 5535
rect 27678 5306 27706 5311
rect 27678 5259 27706 5278
rect 27734 3122 27762 5502
rect 27958 4913 27986 4919
rect 27958 4887 27959 4913
rect 27985 4887 27986 4913
rect 27958 4298 27986 4887
rect 27958 4265 27986 4270
rect 27958 4130 27986 4135
rect 27958 4083 27986 4102
rect 27734 3089 27762 3094
rect 27566 2361 27594 2366
rect 27846 2226 27874 2231
rect 27846 2179 27874 2198
rect 27174 1577 27202 1582
rect 28014 1050 28042 5671
rect 28070 5250 28098 5255
rect 28070 5203 28098 5222
rect 28238 5249 28266 5255
rect 28238 5223 28239 5249
rect 28265 5223 28266 5249
rect 28238 5082 28266 5223
rect 28238 5049 28266 5054
rect 28126 4970 28154 4975
rect 28126 4521 28154 4942
rect 28238 4858 28266 4863
rect 28238 4811 28266 4830
rect 28126 4495 28127 4521
rect 28153 4495 28154 4521
rect 28126 4489 28154 4495
rect 28238 4466 28266 4471
rect 28238 4185 28266 4438
rect 28238 4159 28239 4185
rect 28265 4159 28266 4185
rect 28238 4153 28266 4159
rect 28294 2506 28322 6006
rect 28350 6001 28378 6006
rect 28462 5474 28490 5479
rect 28350 4578 28378 4583
rect 28350 4531 28378 4550
rect 28462 4241 28490 5446
rect 28574 5361 28602 6118
rect 28798 6146 28826 7056
rect 29022 6650 29050 7056
rect 29022 6617 29050 6622
rect 28798 6113 28826 6118
rect 29022 6482 29050 6487
rect 29022 5809 29050 6454
rect 29022 5783 29023 5809
rect 29049 5783 29050 5809
rect 29022 5777 29050 5783
rect 29078 6481 29106 6487
rect 29078 6455 29079 6481
rect 29105 6455 29106 6481
rect 28742 5698 28770 5703
rect 28574 5335 28575 5361
rect 28601 5335 28602 5361
rect 28574 5329 28602 5335
rect 28630 5697 28770 5698
rect 28630 5671 28743 5697
rect 28769 5671 28770 5697
rect 28630 5670 28770 5671
rect 28630 5026 28658 5670
rect 28742 5665 28770 5670
rect 28910 5698 28938 5703
rect 28574 4998 28658 5026
rect 28574 4634 28602 4998
rect 28686 4913 28714 4919
rect 28686 4887 28687 4913
rect 28713 4887 28714 4913
rect 28686 4746 28714 4887
rect 28686 4718 28826 4746
rect 28574 4606 28714 4634
rect 28574 4409 28602 4415
rect 28574 4383 28575 4409
rect 28601 4383 28602 4409
rect 28574 4354 28602 4383
rect 28574 4321 28602 4326
rect 28462 4215 28463 4241
rect 28489 4215 28490 4241
rect 28462 4209 28490 4215
rect 28630 4242 28658 4247
rect 28630 3514 28658 4214
rect 28630 3481 28658 3486
rect 28686 3066 28714 4606
rect 28798 4577 28826 4718
rect 28910 4690 28938 5670
rect 29022 5362 29050 5367
rect 29022 5305 29050 5334
rect 29022 5279 29023 5305
rect 29049 5279 29050 5305
rect 29022 5273 29050 5279
rect 28966 4970 28994 4975
rect 28966 4923 28994 4942
rect 28798 4551 28799 4577
rect 28825 4551 28826 4577
rect 28798 4545 28826 4551
rect 28854 4662 28938 4690
rect 28742 4410 28770 4415
rect 28742 4185 28770 4382
rect 28742 4159 28743 4185
rect 28769 4159 28770 4185
rect 28742 4153 28770 4159
rect 28854 4074 28882 4662
rect 28910 4186 28938 4191
rect 28910 4139 28938 4158
rect 28854 4041 28882 4046
rect 28910 3850 28938 3855
rect 28910 3737 28938 3822
rect 28910 3711 28911 3737
rect 28937 3711 28938 3737
rect 28910 3705 28938 3711
rect 28686 3033 28714 3038
rect 28966 3122 28994 3127
rect 28966 3009 28994 3094
rect 28966 2983 28967 3009
rect 28993 2983 28994 3009
rect 28966 2977 28994 2983
rect 28686 2842 28714 2847
rect 28686 2795 28714 2814
rect 28630 2730 28658 2735
rect 28630 2617 28658 2702
rect 28630 2591 28631 2617
rect 28657 2591 28658 2617
rect 28630 2585 28658 2591
rect 28294 2473 28322 2478
rect 28350 2561 28378 2567
rect 28350 2535 28351 2561
rect 28377 2535 28378 2561
rect 28070 2058 28098 2063
rect 28070 2011 28098 2030
rect 28014 1017 28042 1022
rect 26950 793 26978 798
rect 28350 658 28378 2535
rect 28910 2561 28938 2567
rect 28910 2535 28911 2561
rect 28937 2535 28938 2561
rect 28910 1666 28938 2535
rect 29078 2450 29106 6455
rect 29246 6370 29274 7056
rect 29470 6594 29498 7056
rect 29470 6561 29498 6566
rect 29414 6426 29442 6431
rect 29414 6379 29442 6398
rect 29246 6337 29274 6342
rect 29414 6146 29442 6151
rect 29302 5977 29330 5983
rect 29302 5951 29303 5977
rect 29329 5951 29330 5977
rect 29302 5922 29330 5951
rect 29302 5889 29330 5894
rect 29414 5361 29442 6118
rect 29694 6146 29722 7056
rect 29862 6481 29890 6487
rect 29862 6455 29863 6481
rect 29889 6455 29890 6481
rect 29694 6113 29722 6118
rect 29806 6370 29834 6375
rect 29582 6033 29610 6039
rect 29582 6007 29583 6033
rect 29609 6007 29610 6033
rect 29414 5335 29415 5361
rect 29441 5335 29442 5361
rect 29414 5329 29442 5335
rect 29470 5810 29498 5815
rect 29414 4914 29442 4919
rect 29414 4867 29442 4886
rect 29358 4690 29386 4695
rect 29358 4633 29386 4662
rect 29358 4607 29359 4633
rect 29385 4607 29386 4633
rect 29358 4601 29386 4607
rect 29190 4130 29218 4135
rect 29358 4130 29386 4135
rect 29190 4129 29386 4130
rect 29190 4103 29191 4129
rect 29217 4103 29359 4129
rect 29385 4103 29386 4129
rect 29190 4102 29386 4103
rect 29190 4097 29218 4102
rect 29358 4097 29386 4102
rect 29414 3737 29442 3743
rect 29414 3711 29415 3737
rect 29441 3711 29442 3737
rect 29190 3682 29218 3687
rect 29190 3635 29218 3654
rect 29414 3626 29442 3711
rect 29414 3593 29442 3598
rect 29246 3345 29274 3351
rect 29246 3319 29247 3345
rect 29273 3319 29274 3345
rect 29246 3234 29274 3319
rect 29470 3289 29498 5782
rect 29526 5698 29554 5703
rect 29526 5651 29554 5670
rect 29526 5250 29554 5255
rect 29526 4214 29554 5222
rect 29582 4521 29610 6007
rect 29806 5809 29834 6342
rect 29806 5783 29807 5809
rect 29833 5783 29834 5809
rect 29806 5777 29834 5783
rect 29750 4914 29778 4919
rect 29750 4867 29778 4886
rect 29582 4495 29583 4521
rect 29609 4495 29610 4521
rect 29582 4489 29610 4495
rect 29862 4214 29890 6455
rect 29918 6370 29946 7056
rect 30422 6986 30450 6991
rect 30310 6650 30338 6655
rect 30254 6538 30282 6543
rect 30254 6491 30282 6510
rect 29918 6337 29946 6342
rect 30310 6145 30338 6622
rect 30310 6119 30311 6145
rect 30337 6119 30338 6145
rect 30310 6113 30338 6119
rect 29526 4186 29610 4214
rect 29582 3793 29610 4186
rect 29582 3767 29583 3793
rect 29609 3767 29610 3793
rect 29582 3761 29610 3767
rect 29806 4186 29890 4214
rect 29918 6033 29946 6039
rect 29918 6007 29919 6033
rect 29945 6007 29946 6033
rect 29470 3263 29471 3289
rect 29497 3263 29498 3289
rect 29470 3257 29498 3263
rect 29526 3570 29554 3575
rect 29246 3201 29274 3206
rect 29414 2953 29442 2959
rect 29414 2927 29415 2953
rect 29441 2927 29442 2953
rect 29190 2618 29218 2623
rect 29190 2571 29218 2590
rect 29078 2417 29106 2422
rect 29414 2338 29442 2927
rect 29414 2305 29442 2310
rect 28910 1633 28938 1638
rect 29526 1554 29554 3542
rect 29806 3402 29834 4186
rect 29862 4130 29890 4135
rect 29862 4073 29890 4102
rect 29862 4047 29863 4073
rect 29889 4047 29890 4073
rect 29862 4041 29890 4047
rect 29806 3369 29834 3374
rect 29694 3345 29722 3351
rect 29694 3319 29695 3345
rect 29721 3319 29722 3345
rect 29694 3178 29722 3319
rect 29694 3145 29722 3150
rect 29638 3010 29666 3015
rect 29638 2963 29666 2982
rect 29694 2674 29722 2679
rect 29694 2627 29722 2646
rect 29694 1778 29722 1783
rect 29694 1731 29722 1750
rect 29918 1722 29946 6007
rect 30366 5697 30394 5703
rect 30366 5671 30367 5697
rect 30393 5671 30394 5697
rect 30310 5305 30338 5311
rect 30310 5279 30311 5305
rect 30337 5279 30338 5305
rect 30142 4913 30170 4919
rect 30142 4887 30143 4913
rect 30169 4887 30170 4913
rect 30142 4802 30170 4887
rect 30142 4769 30170 4774
rect 30198 4858 30226 4863
rect 30198 4129 30226 4830
rect 30254 4466 30282 4471
rect 30254 4419 30282 4438
rect 30198 4103 30199 4129
rect 30225 4103 30226 4129
rect 30198 4097 30226 4103
rect 30254 3738 30282 3743
rect 30254 3691 30282 3710
rect 30254 3458 30282 3463
rect 29974 3346 30002 3351
rect 29974 3299 30002 3318
rect 30142 3345 30170 3351
rect 30142 3319 30143 3345
rect 30169 3319 30170 3345
rect 30142 3290 30170 3319
rect 30142 3257 30170 3262
rect 30254 2953 30282 3430
rect 30310 3122 30338 5279
rect 30310 3089 30338 3094
rect 30254 2927 30255 2953
rect 30281 2927 30282 2953
rect 30254 2921 30282 2927
rect 30142 2730 30170 2735
rect 30142 2617 30170 2702
rect 30142 2591 30143 2617
rect 30169 2591 30170 2617
rect 30142 2585 30170 2591
rect 29974 2562 30002 2567
rect 29974 2515 30002 2534
rect 30366 2226 30394 5671
rect 30422 5306 30450 6958
rect 32102 6762 32130 6767
rect 31262 6594 31290 6599
rect 31262 6547 31290 6566
rect 31374 6538 31402 6543
rect 30982 6481 31010 6487
rect 30982 6455 30983 6481
rect 31009 6455 31010 6481
rect 30590 6370 30618 6375
rect 30590 5809 30618 6342
rect 30590 5783 30591 5809
rect 30617 5783 30618 5809
rect 30590 5777 30618 5783
rect 30702 6033 30730 6039
rect 30702 6007 30703 6033
rect 30729 6007 30730 6033
rect 30422 5273 30450 5278
rect 30646 4858 30674 4863
rect 30646 4811 30674 4830
rect 30702 4214 30730 6007
rect 30982 5642 31010 6455
rect 31094 6146 31122 6151
rect 31094 6099 31122 6118
rect 30982 5609 31010 5614
rect 31094 5697 31122 5703
rect 31094 5671 31095 5697
rect 31121 5671 31122 5697
rect 31094 5530 31122 5671
rect 31318 5642 31346 5647
rect 31094 5497 31122 5502
rect 31150 5641 31346 5642
rect 31150 5615 31319 5641
rect 31345 5615 31346 5641
rect 31150 5614 31346 5615
rect 31094 5418 31122 5423
rect 30758 5361 30786 5367
rect 30758 5335 30759 5361
rect 30785 5335 30786 5361
rect 30758 5082 30786 5335
rect 31094 5305 31122 5390
rect 31094 5279 31095 5305
rect 31121 5279 31122 5305
rect 31094 5273 31122 5279
rect 30758 5049 30786 5054
rect 31094 5194 31122 5199
rect 30982 4913 31010 4919
rect 30982 4887 30983 4913
rect 31009 4887 31010 4913
rect 30758 4634 30786 4639
rect 30758 4587 30786 4606
rect 30534 4186 30562 4191
rect 30534 4139 30562 4158
rect 30590 4186 30730 4214
rect 30590 3570 30618 4186
rect 30926 4130 30954 4135
rect 30870 4129 30954 4130
rect 30870 4103 30927 4129
rect 30953 4103 30954 4129
rect 30870 4102 30954 4103
rect 30590 3537 30618 3542
rect 30758 3793 30786 3799
rect 30758 3767 30759 3793
rect 30785 3767 30786 3793
rect 30758 3402 30786 3767
rect 30758 3369 30786 3374
rect 30646 3233 30674 3239
rect 30646 3207 30647 3233
rect 30673 3207 30674 3233
rect 30646 2954 30674 3207
rect 30758 3066 30786 3071
rect 30758 3019 30786 3038
rect 30870 3010 30898 4102
rect 30926 4097 30954 4102
rect 30982 3346 31010 4887
rect 31094 4858 31122 5166
rect 31094 4825 31122 4830
rect 31150 4521 31178 5614
rect 31318 5609 31346 5614
rect 31374 5530 31402 6510
rect 31822 6314 31850 6319
rect 31542 5866 31570 5871
rect 31262 5502 31402 5530
rect 31486 5642 31514 5647
rect 31262 4970 31290 5502
rect 31262 4937 31290 4942
rect 31318 5418 31346 5423
rect 31318 4634 31346 5390
rect 31430 5249 31458 5255
rect 31430 5223 31431 5249
rect 31457 5223 31458 5249
rect 31318 4601 31346 4606
rect 31374 4857 31402 4863
rect 31374 4831 31375 4857
rect 31401 4831 31402 4857
rect 31150 4495 31151 4521
rect 31177 4495 31178 4521
rect 31150 4489 31178 4495
rect 31374 4522 31402 4831
rect 31430 4746 31458 5223
rect 31486 4914 31514 5614
rect 31486 4881 31514 4886
rect 31430 4713 31458 4718
rect 31374 4489 31402 4494
rect 31430 4465 31458 4471
rect 31430 4439 31431 4465
rect 31457 4439 31458 4465
rect 31430 4298 31458 4439
rect 31430 4265 31458 4270
rect 31542 4186 31570 5838
rect 31542 4153 31570 4158
rect 31822 4130 31850 6286
rect 31878 6090 31906 6095
rect 31878 4690 31906 6062
rect 31878 4657 31906 4662
rect 31822 4097 31850 4102
rect 31542 4074 31570 4079
rect 31430 4017 31458 4023
rect 31430 3991 31431 4017
rect 31457 3991 31458 4017
rect 31430 3850 31458 3991
rect 31430 3817 31458 3822
rect 31542 3849 31570 4046
rect 31542 3823 31543 3849
rect 31569 3823 31570 3849
rect 31542 3817 31570 3823
rect 31150 3737 31178 3743
rect 31150 3711 31151 3737
rect 31177 3711 31178 3737
rect 31094 3514 31122 3519
rect 30982 3313 31010 3318
rect 31038 3345 31066 3351
rect 31038 3319 31039 3345
rect 31065 3319 31066 3345
rect 30870 2977 30898 2982
rect 30646 2921 30674 2926
rect 30534 2618 30562 2623
rect 30534 2571 30562 2590
rect 30926 2562 30954 2567
rect 30926 2515 30954 2534
rect 30366 2193 30394 2198
rect 30254 2113 30282 2119
rect 30254 2087 30255 2113
rect 30281 2087 30282 2113
rect 29974 1778 30002 1783
rect 30142 1778 30170 1783
rect 29974 1777 30170 1778
rect 29974 1751 29975 1777
rect 30001 1751 30143 1777
rect 30169 1751 30170 1777
rect 29974 1750 30170 1751
rect 29974 1745 30002 1750
rect 30142 1745 30170 1750
rect 29918 1689 29946 1694
rect 29526 1521 29554 1526
rect 29246 1442 29274 1447
rect 29190 1330 29218 1335
rect 29190 1283 29218 1302
rect 28910 1273 28938 1279
rect 28910 1247 28911 1273
rect 28937 1247 28938 1273
rect 28798 1050 28826 1055
rect 28798 1003 28826 1022
rect 28574 994 28602 999
rect 28574 947 28602 966
rect 28910 714 28938 1247
rect 29246 1049 29274 1414
rect 30254 1442 30282 2087
rect 30646 2113 30674 2119
rect 30646 2087 30647 2113
rect 30673 2087 30674 2113
rect 30254 1409 30282 1414
rect 30534 2058 30562 2063
rect 29414 1385 29442 1391
rect 29414 1359 29415 1385
rect 29441 1359 29442 1385
rect 29414 1274 29442 1359
rect 29638 1386 29666 1391
rect 29638 1339 29666 1358
rect 29414 1241 29442 1246
rect 30086 1330 30114 1335
rect 29694 1218 29722 1223
rect 29246 1023 29247 1049
rect 29273 1023 29274 1049
rect 29246 1017 29274 1023
rect 29414 1162 29442 1167
rect 28966 993 28994 999
rect 28966 967 28967 993
rect 28993 967 28994 993
rect 28966 938 28994 967
rect 28966 905 28994 910
rect 28910 681 28938 686
rect 29134 882 29162 887
rect 28350 625 28378 630
rect 26894 513 26922 518
rect 27678 602 27706 607
rect 27678 56 27706 574
rect 29134 56 29162 854
rect 29302 545 29330 551
rect 29302 519 29303 545
rect 29329 519 29330 545
rect 29302 378 29330 519
rect 29414 434 29442 1134
rect 29694 1105 29722 1190
rect 29694 1079 29695 1105
rect 29721 1079 29722 1105
rect 29694 1073 29722 1079
rect 29974 994 30002 999
rect 29974 947 30002 966
rect 29414 401 29442 406
rect 29806 657 29834 663
rect 29806 631 29807 657
rect 29833 631 29834 657
rect 29302 345 29330 350
rect 29806 266 29834 631
rect 30086 601 30114 1302
rect 30254 1329 30282 1335
rect 30254 1303 30255 1329
rect 30281 1303 30282 1329
rect 30142 1050 30170 1055
rect 30142 1003 30170 1022
rect 30254 770 30282 1303
rect 30254 737 30282 742
rect 30086 575 30087 601
rect 30113 575 30114 601
rect 30086 569 30114 575
rect 30534 378 30562 2030
rect 30646 1834 30674 2087
rect 30646 1801 30674 1806
rect 30926 1778 30954 1783
rect 30926 1731 30954 1750
rect 30646 1722 30674 1727
rect 30646 1675 30674 1694
rect 30646 1330 30674 1335
rect 30646 1283 30674 1302
rect 30926 994 30954 999
rect 30926 947 30954 966
rect 30646 882 30674 887
rect 30646 835 30674 854
rect 31038 826 31066 3319
rect 31094 2953 31122 3486
rect 31094 2927 31095 2953
rect 31121 2927 31122 2953
rect 31094 2921 31122 2927
rect 31094 2674 31122 2679
rect 31094 2169 31122 2646
rect 31094 2143 31095 2169
rect 31121 2143 31122 2169
rect 31094 2137 31122 2143
rect 31094 1386 31122 1391
rect 31094 1339 31122 1358
rect 31150 1162 31178 3711
rect 31430 3626 31458 3631
rect 31430 3289 31458 3598
rect 31430 3263 31431 3289
rect 31457 3263 31458 3289
rect 31430 3257 31458 3263
rect 31542 3178 31570 3183
rect 31542 3065 31570 3150
rect 31542 3039 31543 3065
rect 31569 3039 31570 3065
rect 31542 3033 31570 3039
rect 32102 3066 32130 6734
rect 32102 3033 32130 3038
rect 31318 2730 31346 2735
rect 31262 2618 31290 2623
rect 31262 2282 31290 2590
rect 31318 2617 31346 2702
rect 31318 2591 31319 2617
rect 31345 2591 31346 2617
rect 31318 2585 31346 2591
rect 31262 2249 31290 2254
rect 31542 2506 31570 2511
rect 31542 2281 31570 2478
rect 31542 2255 31543 2281
rect 31569 2255 31570 2281
rect 31542 2249 31570 2255
rect 31430 2058 31458 2063
rect 31318 1722 31346 1727
rect 31318 1386 31346 1694
rect 31430 1721 31458 2030
rect 31430 1695 31431 1721
rect 31457 1695 31458 1721
rect 31430 1689 31458 1695
rect 31542 1610 31570 1615
rect 31542 1497 31570 1582
rect 31542 1471 31543 1497
rect 31569 1471 31570 1497
rect 31542 1465 31570 1471
rect 31318 1353 31346 1358
rect 31150 1129 31178 1134
rect 31374 1330 31402 1335
rect 31038 793 31066 798
rect 30590 657 30618 663
rect 30590 631 30591 657
rect 30617 631 30618 657
rect 30590 490 30618 631
rect 31094 601 31122 607
rect 31094 575 31095 601
rect 31121 575 31122 601
rect 31094 546 31122 575
rect 31094 513 31122 518
rect 30590 457 30618 462
rect 30534 350 30618 378
rect 29806 233 29834 238
rect 30590 56 30618 350
rect 16758 9 16786 14
rect 17472 0 17528 56
rect 18928 0 18984 56
rect 20384 0 20440 56
rect 21840 0 21896 56
rect 23296 0 23352 56
rect 24752 0 24808 56
rect 26208 0 26264 56
rect 27664 0 27720 56
rect 29120 0 29176 56
rect 30576 0 30632 56
rect 31374 42 31402 1302
rect 31430 1162 31458 1167
rect 31430 937 31458 1134
rect 31430 911 31431 937
rect 31457 911 31458 937
rect 31430 905 31458 911
rect 31542 938 31570 943
rect 31542 713 31570 910
rect 31542 687 31543 713
rect 31569 687 31570 713
rect 31542 681 31570 687
rect 31374 9 31402 14
<< via2 >>
rect 126 6958 154 6986
rect 1862 6790 1890 6818
rect 1806 6734 1834 6762
rect 1246 6566 1274 6594
rect 798 6510 826 6538
rect 462 6286 490 6314
rect 462 5222 490 5250
rect 798 4998 826 5026
rect 1078 6454 1106 6482
rect 966 5641 994 5642
rect 966 5615 967 5641
rect 967 5615 993 5641
rect 993 5615 994 5641
rect 966 5614 994 5615
rect 126 3430 154 3458
rect 1022 3262 1050 3290
rect 1022 2870 1050 2898
rect 910 2198 938 2226
rect 1414 6118 1442 6146
rect 1134 5278 1162 5306
rect 1190 5558 1218 5586
rect 1190 4606 1218 4634
rect 2086 6678 2114 6706
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 1526 5222 1554 5250
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1638 4550 1666 4578
rect 2366 6734 2394 6762
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 2142 6566 2170 6594
rect 2198 6033 2226 6034
rect 2198 6007 2199 6033
rect 2199 6007 2225 6033
rect 2225 6007 2226 6033
rect 2198 6006 2226 6007
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 2310 5809 2338 5810
rect 2310 5783 2311 5809
rect 2311 5783 2337 5809
rect 2337 5783 2338 5809
rect 2310 5782 2338 5783
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 1526 3766 1554 3794
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1302 3318 1330 3346
rect 1246 2841 1274 2842
rect 1246 2815 1247 2841
rect 1247 2815 1273 2841
rect 1273 2815 1274 2841
rect 1246 2814 1274 2815
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 1190 2057 1218 2058
rect 1190 2031 1191 2057
rect 1191 2031 1217 2057
rect 1217 2031 1218 2057
rect 1190 2030 1218 2031
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 1302 1777 1330 1778
rect 1302 1751 1303 1777
rect 1303 1751 1329 1777
rect 1329 1751 1330 1777
rect 1302 1750 1330 1751
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 966 1414 994 1442
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 1246 993 1274 994
rect 1246 967 1247 993
rect 1247 967 1273 993
rect 1273 967 1274 993
rect 1246 966 1274 967
rect 1470 798 1498 826
rect 1190 489 1218 490
rect 1190 463 1191 489
rect 1191 463 1217 489
rect 1217 463 1218 489
rect 1190 462 1218 463
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2814 6790 2842 6818
rect 2982 6593 3010 6594
rect 2982 6567 2983 6593
rect 2983 6567 3009 6593
rect 3009 6567 3010 6593
rect 2982 6566 3010 6567
rect 2590 5782 2618 5810
rect 2926 6006 2954 6034
rect 2590 5558 2618 5586
rect 2590 5446 2618 5474
rect 2534 4606 2562 4634
rect 2758 4774 2786 4802
rect 2646 4129 2674 4130
rect 2646 4103 2647 4129
rect 2647 4103 2673 4129
rect 2673 4103 2674 4129
rect 2646 4102 2674 4103
rect 2926 2982 2954 3010
rect 2590 2870 2618 2898
rect 3318 5697 3346 5698
rect 3318 5671 3319 5697
rect 3319 5671 3345 5697
rect 3345 5671 3346 5697
rect 3318 5670 3346 5671
rect 3486 6566 3514 6594
rect 3766 6593 3794 6594
rect 3766 6567 3767 6593
rect 3767 6567 3793 6593
rect 3793 6567 3794 6593
rect 3766 6566 3794 6567
rect 3262 2590 3290 2618
rect 3766 2422 3794 2450
rect 2590 2086 2618 2114
rect 2870 1918 2898 1946
rect 3878 5809 3906 5810
rect 3878 5783 3879 5809
rect 3879 5783 3905 5809
rect 3905 5783 3906 5809
rect 3878 5782 3906 5783
rect 3878 5166 3906 5194
rect 4382 6566 4410 6594
rect 4270 6201 4298 6202
rect 4270 6175 4271 6201
rect 4271 6175 4297 6201
rect 4297 6175 4298 6201
rect 4270 6174 4298 6175
rect 4550 5950 4578 5978
rect 4158 5782 4186 5810
rect 4158 5502 4186 5530
rect 4214 5558 4242 5586
rect 4158 4857 4186 4858
rect 4158 4831 4159 4857
rect 4159 4831 4185 4857
rect 4185 4831 4186 4857
rect 4158 4830 4186 4831
rect 4046 3654 4074 3682
rect 4046 3009 4074 3010
rect 4046 2983 4047 3009
rect 4047 2983 4073 3009
rect 4073 2983 4074 3009
rect 4046 2982 4074 2983
rect 4886 6622 4914 6650
rect 4998 6566 5026 6594
rect 4830 6174 4858 6202
rect 5278 6566 5306 6594
rect 4550 5054 4578 5082
rect 5334 6118 5362 6146
rect 5334 5166 5362 5194
rect 5670 6593 5698 6594
rect 5670 6567 5671 6593
rect 5671 6567 5697 6593
rect 5697 6567 5698 6593
rect 5670 6566 5698 6567
rect 5446 5809 5474 5810
rect 5446 5783 5447 5809
rect 5447 5783 5473 5809
rect 5473 5783 5474 5809
rect 5446 5782 5474 5783
rect 5390 4886 5418 4914
rect 5446 5670 5474 5698
rect 4326 2953 4354 2954
rect 4326 2927 4327 2953
rect 4327 2927 4353 2953
rect 4353 2927 4354 2953
rect 4326 2926 4354 2927
rect 5950 6622 5978 6650
rect 5838 6201 5866 6202
rect 5838 6175 5839 6201
rect 5839 6175 5865 6201
rect 5865 6175 5866 6201
rect 5838 6174 5866 6175
rect 5726 5782 5754 5810
rect 5782 3542 5810 3570
rect 5726 3206 5754 3234
rect 5446 2310 5474 2338
rect 5894 2870 5922 2898
rect 4214 1582 4242 1610
rect 3822 1022 3850 1050
rect 4830 1470 4858 1498
rect 4550 910 4578 938
rect 2422 742 2450 770
rect 4382 630 4410 658
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 2926 126 2954 154
rect 5278 854 5306 882
rect 6118 5894 6146 5922
rect 6062 5782 6090 5810
rect 5950 1526 5978 1554
rect 6006 2814 6034 2842
rect 6006 1414 6034 1442
rect 5950 1302 5978 1330
rect 5110 238 5138 266
rect 5054 182 5082 210
rect 5278 126 5306 154
rect 5950 630 5978 658
rect 6622 6566 6650 6594
rect 6454 6481 6482 6482
rect 6454 6455 6455 6481
rect 6455 6455 6481 6481
rect 6481 6455 6482 6481
rect 6454 6454 6482 6455
rect 6398 6174 6426 6202
rect 6678 6174 6706 6202
rect 6342 6006 6370 6034
rect 6286 5390 6314 5418
rect 6118 5249 6146 5250
rect 6118 5223 6119 5249
rect 6119 5223 6145 5249
rect 6145 5223 6146 5249
rect 6118 5222 6146 5223
rect 6174 4046 6202 4074
rect 6118 1358 6146 1386
rect 6286 3934 6314 3962
rect 6230 2982 6258 3010
rect 6510 5334 6538 5362
rect 6454 5054 6482 5082
rect 6398 4270 6426 4298
rect 6398 2926 6426 2954
rect 6342 2198 6370 2226
rect 6734 5446 6762 5474
rect 6678 4998 6706 5026
rect 6790 4830 6818 4858
rect 6958 6425 6986 6426
rect 6958 6399 6959 6425
rect 6959 6399 6985 6425
rect 6985 6399 6986 6425
rect 6958 6398 6986 6399
rect 7070 6033 7098 6034
rect 7070 6007 7071 6033
rect 7071 6007 7097 6033
rect 7097 6007 7098 6033
rect 7070 6006 7098 6007
rect 7406 6510 7434 6538
rect 7462 6454 7490 6482
rect 7518 6398 7546 6426
rect 7350 5950 7378 5978
rect 7518 5894 7546 5922
rect 7518 5726 7546 5754
rect 7350 5670 7378 5698
rect 7350 5502 7378 5530
rect 6734 4774 6762 4802
rect 6510 4438 6538 4466
rect 6622 4494 6650 4522
rect 6454 1974 6482 2002
rect 6510 2646 6538 2674
rect 6510 1862 6538 1890
rect 6286 1526 6314 1554
rect 6622 3990 6650 4018
rect 6678 4438 6706 4466
rect 6734 3878 6762 3906
rect 6846 4326 6874 4354
rect 6678 3710 6706 3738
rect 7406 3793 7434 3794
rect 7406 3767 7407 3793
rect 7407 3767 7433 3793
rect 7433 3767 7434 3793
rect 7406 3766 7434 3767
rect 7350 3430 7378 3458
rect 7966 6454 7994 6482
rect 8190 6566 8218 6594
rect 8414 6510 8442 6538
rect 8582 6958 8610 6986
rect 7462 3262 7490 3290
rect 7406 3206 7434 3234
rect 7126 2702 7154 2730
rect 7126 2478 7154 2506
rect 7574 4270 7602 4298
rect 7630 4158 7658 4186
rect 7686 4046 7714 4074
rect 7742 4270 7770 4298
rect 7686 3710 7714 3738
rect 7518 3206 7546 3234
rect 7406 2366 7434 2394
rect 6846 1806 6874 1834
rect 7126 1694 7154 1722
rect 6566 1526 6594 1554
rect 6622 1638 6650 1666
rect 6286 1078 6314 1106
rect 6118 406 6146 434
rect 6678 910 6706 938
rect 8246 4046 8274 4074
rect 7854 2814 7882 2842
rect 8078 2926 8106 2954
rect 7686 1190 7714 1218
rect 7798 1582 7826 1610
rect 7630 1105 7658 1106
rect 7630 1079 7631 1105
rect 7631 1079 7657 1105
rect 7657 1079 7658 1105
rect 7630 1078 7658 1079
rect 7350 1049 7378 1050
rect 7350 1023 7351 1049
rect 7351 1023 7377 1049
rect 7377 1023 7378 1049
rect 7350 1022 7378 1023
rect 8302 3318 8330 3346
rect 8358 3374 8386 3402
rect 8470 3038 8498 3066
rect 8414 2422 8442 2450
rect 8358 2030 8386 2058
rect 8414 2310 8442 2338
rect 7126 798 7154 826
rect 7574 966 7602 994
rect 6678 742 6706 770
rect 6622 686 6650 714
rect 7294 686 7322 714
rect 6510 350 6538 378
rect 6062 182 6090 210
rect 7686 854 7714 882
rect 7686 630 7714 658
rect 7574 574 7602 602
rect 8638 6566 8666 6594
rect 8694 6622 8722 6650
rect 8638 5614 8666 5642
rect 8974 6342 9002 6370
rect 9478 6593 9506 6594
rect 9478 6567 9479 6593
rect 9479 6567 9505 6593
rect 9505 6567 9506 6593
rect 9478 6566 9506 6567
rect 9534 6342 9562 6370
rect 9702 6846 9730 6874
rect 9422 6089 9450 6090
rect 9422 6063 9423 6089
rect 9423 6063 9449 6089
rect 9449 6063 9450 6089
rect 9422 6062 9450 6063
rect 9198 5894 9226 5922
rect 8638 3150 8666 3178
rect 8694 3430 8722 3458
rect 8638 2673 8666 2674
rect 8638 2647 8639 2673
rect 8639 2647 8665 2673
rect 8665 2647 8666 2673
rect 8638 2646 8666 2647
rect 8750 3345 8778 3346
rect 8750 3319 8751 3345
rect 8751 3319 8777 3345
rect 8777 3319 8778 3345
rect 8750 3318 8778 3319
rect 8918 4214 8946 4242
rect 8974 4102 9002 4130
rect 9478 5222 9506 5250
rect 9478 5054 9506 5082
rect 9198 4942 9226 4970
rect 9030 3766 9058 3794
rect 9086 3878 9114 3906
rect 8862 3150 8890 3178
rect 8694 1414 8722 1442
rect 8750 2478 8778 2506
rect 8526 294 8554 322
rect 9030 1806 9058 1834
rect 9030 1470 9058 1498
rect 9198 3374 9226 3402
rect 9758 6622 9786 6650
rect 9814 6958 9842 6986
rect 9758 6481 9786 6482
rect 9758 6455 9759 6481
rect 9759 6455 9785 6481
rect 9785 6455 9786 6481
rect 9758 6454 9786 6455
rect 9702 3094 9730 3122
rect 9366 2617 9394 2618
rect 9366 2591 9367 2617
rect 9367 2591 9393 2617
rect 9393 2591 9394 2617
rect 9366 2590 9394 2591
rect 9646 2617 9674 2618
rect 9646 2591 9647 2617
rect 9647 2591 9673 2617
rect 9673 2591 9674 2617
rect 9646 2590 9674 2591
rect 9142 2534 9170 2562
rect 9870 6510 9898 6538
rect 10038 6230 10066 6258
rect 10262 6790 10290 6818
rect 10038 5614 10066 5642
rect 10094 5166 10122 5194
rect 9982 4606 10010 4634
rect 10038 4718 10066 4746
rect 9870 4102 9898 4130
rect 9982 4158 10010 4186
rect 10038 4102 10066 4130
rect 9982 3710 10010 3738
rect 10038 3542 10066 3570
rect 10430 6566 10458 6594
rect 10598 6593 10626 6594
rect 10598 6567 10599 6593
rect 10599 6567 10625 6593
rect 10625 6567 10626 6593
rect 10598 6566 10626 6567
rect 10486 5950 10514 5978
rect 10262 4550 10290 4578
rect 10094 3262 10122 3290
rect 10038 2142 10066 2170
rect 10262 1862 10290 1890
rect 10486 5558 10514 5586
rect 10822 5390 10850 5418
rect 10878 5838 10906 5866
rect 10430 5054 10458 5082
rect 10374 4494 10402 4522
rect 10430 3878 10458 3906
rect 10374 3822 10402 3850
rect 10766 5166 10794 5194
rect 10822 4465 10850 4466
rect 10822 4439 10823 4465
rect 10823 4439 10849 4465
rect 10849 4439 10850 4465
rect 10822 4438 10850 4439
rect 10486 3486 10514 3514
rect 10766 4326 10794 4354
rect 10430 3430 10458 3458
rect 10430 2870 10458 2898
rect 10654 3038 10682 3066
rect 10766 2982 10794 3010
rect 10822 3822 10850 3850
rect 11102 6566 11130 6594
rect 11158 6734 11186 6762
rect 11382 6593 11410 6594
rect 11382 6567 11383 6593
rect 11383 6567 11409 6593
rect 11409 6567 11410 6593
rect 11382 6566 11410 6567
rect 11438 5838 11466 5866
rect 11158 5670 11186 5698
rect 10990 4438 11018 4466
rect 10878 2982 10906 3010
rect 10934 3542 10962 3570
rect 10934 2926 10962 2954
rect 10822 2646 10850 2674
rect 10934 2673 10962 2674
rect 10934 2647 10935 2673
rect 10935 2647 10961 2673
rect 10961 2647 10962 2673
rect 10934 2646 10962 2647
rect 11102 3374 11130 3402
rect 10374 1862 10402 1890
rect 10262 1414 10290 1442
rect 9870 1078 9898 1106
rect 10654 1358 10682 1386
rect 10654 686 10682 714
rect 9142 518 9170 546
rect 9254 518 9282 546
rect 10542 518 10570 546
rect 10206 70 10234 98
rect 10374 70 10402 98
rect 11214 2254 11242 2282
rect 11326 5110 11354 5138
rect 10878 1694 10906 1722
rect 10878 1246 10906 1274
rect 10878 742 10906 770
rect 11158 937 11186 938
rect 11158 911 11159 937
rect 11159 911 11185 937
rect 11185 911 11186 937
rect 11158 910 11186 911
rect 10934 686 10962 714
rect 10822 406 10850 434
rect 11662 6342 11690 6370
rect 11998 6566 12026 6594
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 12670 6454 12698 6482
rect 11998 5697 12026 5698
rect 11998 5671 11999 5697
rect 11999 5671 12025 5697
rect 12025 5671 12026 5697
rect 11998 5670 12026 5671
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 12110 5446 12138 5474
rect 11774 5334 11802 5362
rect 11606 5305 11634 5306
rect 11606 5279 11607 5305
rect 11607 5279 11633 5305
rect 11633 5279 11634 5305
rect 11606 5278 11634 5279
rect 12110 5110 12138 5138
rect 11774 4998 11802 5026
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 12110 4718 12138 4746
rect 12614 6062 12642 6090
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12446 5838 12474 5866
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12782 5894 12810 5922
rect 12670 5390 12698 5418
rect 12726 5670 12754 5698
rect 12614 5278 12642 5306
rect 12446 4718 12474 4746
rect 12166 4662 12194 4690
rect 12614 4494 12642 4522
rect 12110 4326 12138 4354
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12446 4326 12474 4354
rect 12446 4158 12474 4186
rect 12558 4102 12586 4130
rect 12614 3990 12642 4018
rect 11902 3933 11930 3934
rect 11774 3878 11802 3906
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12222 3822 12250 3850
rect 12558 3822 12586 3850
rect 12558 3710 12586 3738
rect 12110 3542 12138 3570
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12446 3542 12474 3570
rect 11830 3150 11858 3178
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12110 3150 12138 3178
rect 12006 3122 12034 3123
rect 11774 3038 11802 3066
rect 11494 2926 11522 2954
rect 12446 3262 12474 3290
rect 12110 2702 12138 2730
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 12782 3934 12810 3962
rect 12726 2758 12754 2786
rect 12782 3766 12810 3794
rect 12670 2702 12698 2730
rect 12502 2534 12530 2562
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12006 2338 12034 2339
rect 12110 2310 12138 2338
rect 11774 1974 11802 2002
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12502 1974 12530 2002
rect 12558 2086 12586 2114
rect 12336 1946 12364 1947
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12558 966 12586 994
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 13566 6734 13594 6762
rect 13118 6118 13146 6146
rect 13174 6230 13202 6258
rect 13062 6033 13090 6034
rect 13062 6007 13063 6033
rect 13063 6007 13089 6033
rect 13089 6007 13090 6033
rect 13062 6006 13090 6007
rect 13454 6145 13482 6146
rect 13454 6119 13455 6145
rect 13455 6119 13481 6145
rect 13481 6119 13482 6145
rect 13454 6118 13482 6119
rect 13398 5614 13426 5642
rect 13734 6006 13762 6034
rect 13566 4718 13594 4746
rect 13454 4550 13482 4578
rect 13454 4270 13482 4298
rect 13398 4102 13426 4130
rect 13566 3822 13594 3850
rect 13454 3430 13482 3458
rect 13566 3486 13594 3514
rect 13286 3009 13314 3010
rect 13286 2983 13287 3009
rect 13287 2983 13313 3009
rect 13313 2983 13314 3009
rect 13286 2982 13314 2983
rect 13454 3318 13482 3346
rect 13454 2982 13482 3010
rect 13230 2534 13258 2562
rect 13398 2870 13426 2898
rect 13342 2422 13370 2450
rect 13398 2534 13426 2562
rect 13174 2310 13202 2338
rect 13454 2422 13482 2450
rect 13510 2478 13538 2506
rect 13398 1862 13426 1890
rect 13454 2030 13482 2058
rect 12838 1022 12866 1050
rect 13118 1806 13146 1834
rect 12782 630 12810 658
rect 11326 350 11354 378
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 11662 70 11690 98
rect 13510 1358 13538 1386
rect 13566 1526 13594 1554
rect 13454 574 13482 602
rect 13678 5446 13706 5474
rect 13958 6734 13986 6762
rect 13846 6033 13874 6034
rect 13846 6007 13847 6033
rect 13847 6007 13873 6033
rect 13873 6007 13874 6033
rect 13846 6006 13874 6007
rect 13790 5950 13818 5978
rect 14126 6286 14154 6314
rect 13734 4438 13762 4466
rect 13790 4998 13818 5026
rect 13734 3318 13762 3346
rect 13790 3150 13818 3178
rect 13846 4942 13874 4970
rect 13734 2926 13762 2954
rect 13678 2646 13706 2674
rect 14014 5809 14042 5810
rect 14014 5783 14015 5809
rect 14015 5783 14041 5809
rect 14041 5783 14042 5809
rect 14014 5782 14042 5783
rect 14070 5726 14098 5754
rect 14014 5670 14042 5698
rect 14070 4942 14098 4970
rect 14014 4214 14042 4242
rect 13958 3990 13986 4018
rect 14462 6846 14490 6874
rect 14238 5894 14266 5922
rect 14350 6342 14378 6370
rect 14294 5782 14322 5810
rect 14238 5641 14266 5642
rect 14238 5615 14239 5641
rect 14239 5615 14265 5641
rect 14265 5615 14266 5641
rect 14238 5614 14266 5615
rect 14294 5446 14322 5474
rect 14182 5390 14210 5418
rect 14294 5334 14322 5362
rect 14182 4830 14210 4858
rect 14238 4886 14266 4914
rect 14126 3878 14154 3906
rect 14182 4718 14210 4746
rect 13846 2534 13874 2562
rect 14238 3990 14266 4018
rect 14462 6118 14490 6146
rect 14910 6454 14938 6482
rect 14350 5054 14378 5082
rect 14350 4326 14378 4354
rect 14350 4158 14378 4186
rect 14630 5334 14658 5362
rect 14406 3766 14434 3794
rect 14294 2926 14322 2954
rect 14182 1134 14210 1162
rect 14238 2646 14266 2674
rect 13622 1078 13650 1106
rect 14518 3766 14546 3794
rect 14574 2758 14602 2786
rect 14462 1470 14490 1498
rect 14630 2030 14658 2058
rect 14854 6062 14882 6090
rect 14798 4521 14826 4522
rect 14798 4495 14799 4521
rect 14799 4495 14825 4521
rect 14825 4495 14826 4521
rect 14798 4494 14826 4495
rect 14910 4718 14938 4746
rect 14910 3822 14938 3850
rect 15022 5166 15050 5194
rect 15582 6958 15610 6986
rect 15358 6230 15386 6258
rect 15470 6342 15498 6370
rect 15190 6145 15218 6146
rect 15190 6119 15191 6145
rect 15191 6119 15217 6145
rect 15217 6119 15218 6145
rect 15190 6118 15218 6119
rect 15694 6006 15722 6034
rect 15358 5950 15386 5978
rect 15134 4494 15162 4522
rect 15190 4606 15218 4634
rect 15078 4102 15106 4130
rect 15078 3878 15106 3906
rect 15022 3822 15050 3850
rect 14966 3710 14994 3738
rect 14854 3486 14882 3514
rect 15246 4326 15274 4354
rect 14798 3206 14826 3234
rect 15078 2897 15106 2898
rect 15078 2871 15079 2897
rect 15079 2871 15105 2897
rect 15105 2871 15106 2897
rect 15078 2870 15106 2871
rect 14574 1470 14602 1498
rect 14742 1302 14770 1330
rect 14406 742 14434 770
rect 14406 518 14434 546
rect 14238 238 14266 266
rect 14574 238 14602 266
rect 13566 126 13594 154
rect 15414 5894 15442 5922
rect 15470 5054 15498 5082
rect 15246 2478 15274 2506
rect 15414 2478 15442 2506
rect 15134 2198 15162 2226
rect 15246 854 15274 882
rect 15358 966 15386 994
rect 15358 854 15386 882
rect 15582 5334 15610 5362
rect 15582 3766 15610 3794
rect 15582 1526 15610 1554
rect 16254 7014 16282 7042
rect 16030 6286 16058 6314
rect 15918 6006 15946 6034
rect 15918 5670 15946 5698
rect 16198 5558 16226 5586
rect 15974 4382 16002 4410
rect 16198 4326 16226 4354
rect 16366 5502 16394 5530
rect 15974 4270 16002 4298
rect 15918 3430 15946 3458
rect 15918 2982 15946 3010
rect 16310 3094 16338 3122
rect 15806 2590 15834 2618
rect 16366 2758 16394 2786
rect 16366 2590 16394 2618
rect 16366 2366 16394 2394
rect 16478 2310 16506 2338
rect 16534 6510 16562 6538
rect 16366 1582 16394 1610
rect 16590 6174 16618 6202
rect 15694 1190 15722 1218
rect 16198 937 16226 938
rect 16198 911 16199 937
rect 16199 911 16225 937
rect 16225 911 16226 937
rect 16198 910 16226 911
rect 15470 798 15498 826
rect 16646 5502 16674 5530
rect 16814 6230 16842 6258
rect 16814 5222 16842 5250
rect 16646 5054 16674 5082
rect 16814 4830 16842 4858
rect 17150 5222 17178 5250
rect 16926 4830 16954 4858
rect 16982 5110 17010 5138
rect 16702 4774 16730 4802
rect 16982 4718 17010 4746
rect 16870 4326 16898 4354
rect 16870 4158 16898 4186
rect 16814 3486 16842 3514
rect 17486 6678 17514 6706
rect 17598 6566 17626 6594
rect 17654 5894 17682 5922
rect 17822 5670 17850 5698
rect 17878 5278 17906 5306
rect 17710 4942 17738 4970
rect 17598 4718 17626 4746
rect 17486 4158 17514 4186
rect 17542 4606 17570 4634
rect 17486 4046 17514 4074
rect 17430 3737 17458 3738
rect 17430 3711 17431 3737
rect 17431 3711 17457 3737
rect 17457 3711 17458 3737
rect 17430 3710 17458 3711
rect 17374 3206 17402 3234
rect 16702 1918 16730 1946
rect 16702 1806 16730 1834
rect 16814 1918 16842 1946
rect 16814 1694 16842 1722
rect 16590 630 16618 658
rect 16758 910 16786 938
rect 15134 518 15162 546
rect 15974 406 16002 434
rect 15974 294 16002 322
rect 16086 294 16114 322
rect 14798 70 14826 98
rect 17598 3990 17626 4018
rect 17654 4606 17682 4634
rect 17654 3878 17682 3906
rect 17542 3710 17570 3738
rect 18270 6790 18298 6818
rect 18046 4942 18074 4970
rect 18214 5222 18242 5250
rect 17766 4662 17794 4690
rect 18214 4662 18242 4690
rect 17766 3878 17794 3906
rect 18382 4382 18410 4410
rect 17710 3766 17738 3794
rect 17710 3681 17738 3682
rect 17710 3655 17711 3681
rect 17711 3655 17737 3681
rect 17737 3655 17738 3681
rect 17710 3654 17738 3655
rect 17542 2814 17570 2842
rect 17542 1974 17570 2002
rect 17654 1750 17682 1778
rect 17654 1134 17682 1162
rect 17598 798 17626 826
rect 18046 3430 18074 3458
rect 17990 2814 18018 2842
rect 17822 2254 17850 2282
rect 17934 1638 17962 1666
rect 17878 1582 17906 1610
rect 17878 1134 17906 1162
rect 18158 3289 18186 3290
rect 18158 3263 18159 3289
rect 18159 3263 18185 3289
rect 18185 3263 18186 3289
rect 18158 3262 18186 3263
rect 18046 1918 18074 1946
rect 18214 2926 18242 2954
rect 18438 4270 18466 4298
rect 18438 3822 18466 3850
rect 18662 6286 18690 6314
rect 18550 5446 18578 5474
rect 18550 4214 18578 4242
rect 18606 4662 18634 4690
rect 18550 3654 18578 3682
rect 18718 6062 18746 6090
rect 18942 5950 18970 5978
rect 18998 6958 19026 6986
rect 18662 4382 18690 4410
rect 18606 3318 18634 3346
rect 18886 3374 18914 3402
rect 18382 2478 18410 2506
rect 18214 1582 18242 1610
rect 18270 2422 18298 2450
rect 18158 1078 18186 1106
rect 17990 910 18018 938
rect 17822 742 17850 770
rect 17710 686 17738 714
rect 18438 2142 18466 2170
rect 18438 1105 18466 1106
rect 18438 1079 18439 1105
rect 18439 1079 18465 1105
rect 18465 1079 18466 1105
rect 18438 1078 18466 1079
rect 18774 1049 18802 1050
rect 18774 1023 18775 1049
rect 18775 1023 18801 1049
rect 18801 1023 18802 1049
rect 18774 1022 18802 1023
rect 19110 6398 19138 6426
rect 19054 5950 19082 5978
rect 19054 5558 19082 5586
rect 19390 6230 19418 6258
rect 19166 6006 19194 6034
rect 19838 6622 19866 6650
rect 19614 5782 19642 5810
rect 19558 5670 19586 5698
rect 19446 5502 19474 5530
rect 19334 3542 19362 3570
rect 19334 2198 19362 2226
rect 19502 4774 19530 4802
rect 20006 5166 20034 5194
rect 19558 3822 19586 3850
rect 19614 5110 19642 5138
rect 19502 2646 19530 2674
rect 19782 4550 19810 4578
rect 20006 3766 20034 3794
rect 20174 6174 20202 6202
rect 20174 5782 20202 5810
rect 20062 3710 20090 3738
rect 20174 4662 20202 4690
rect 20118 3430 20146 3458
rect 20118 3262 20146 3290
rect 19782 2926 19810 2954
rect 20230 4465 20258 4466
rect 20230 4439 20231 4465
rect 20231 4439 20257 4465
rect 20257 4439 20258 4465
rect 20230 4438 20258 4439
rect 20510 6062 20538 6090
rect 20678 6089 20706 6090
rect 20678 6063 20679 6089
rect 20679 6063 20705 6089
rect 20705 6063 20706 6089
rect 20678 6062 20706 6063
rect 20398 5977 20426 5978
rect 20398 5951 20399 5977
rect 20399 5951 20425 5977
rect 20425 5951 20426 5977
rect 20398 5950 20426 5951
rect 20566 4942 20594 4970
rect 20342 4606 20370 4634
rect 20566 4606 20594 4634
rect 20510 4521 20538 4522
rect 20510 4495 20511 4521
rect 20511 4495 20537 4521
rect 20537 4495 20538 4521
rect 20510 4494 20538 4495
rect 20342 4382 20370 4410
rect 20286 4046 20314 4074
rect 20622 4270 20650 4298
rect 20622 3710 20650 3738
rect 20678 4214 20706 4242
rect 20454 3150 20482 3178
rect 19614 2254 19642 2282
rect 20230 2534 20258 2562
rect 19446 1862 19474 1890
rect 20174 1721 20202 1722
rect 20174 1695 20175 1721
rect 20175 1695 20201 1721
rect 20201 1695 20202 1721
rect 20174 1694 20202 1695
rect 19222 1638 19250 1666
rect 20230 1638 20258 1666
rect 20342 2534 20370 2562
rect 19726 1358 19754 1386
rect 18942 1078 18970 1106
rect 19446 1190 19474 1218
rect 18886 1022 18914 1050
rect 20398 2254 20426 2282
rect 19054 993 19082 994
rect 19054 967 19055 993
rect 19055 967 19081 993
rect 19081 967 19082 993
rect 19054 966 19082 967
rect 18270 630 18298 658
rect 18438 910 18466 938
rect 17542 574 17570 602
rect 20286 910 20314 938
rect 20286 742 20314 770
rect 18438 518 18466 546
rect 18942 630 18970 658
rect 17486 462 17514 490
rect 17486 126 17514 154
rect 20622 1049 20650 1050
rect 20622 1023 20623 1049
rect 20623 1023 20649 1049
rect 20649 1023 20650 1049
rect 20622 1022 20650 1023
rect 20958 6286 20986 6314
rect 20958 6174 20986 6202
rect 20734 1974 20762 2002
rect 20790 5894 20818 5922
rect 20958 3990 20986 4018
rect 21126 5446 21154 5474
rect 20846 3878 20874 3906
rect 21238 5726 21266 5754
rect 20902 2702 20930 2730
rect 21014 1750 21042 1778
rect 20790 1190 20818 1218
rect 20902 1414 20930 1442
rect 21070 1302 21098 1330
rect 20678 406 20706 434
rect 21182 2673 21210 2674
rect 21182 2647 21183 2673
rect 21183 2647 21209 2673
rect 21209 2647 21210 2673
rect 21182 2646 21210 2647
rect 21630 6510 21658 6538
rect 22526 6958 22554 6986
rect 22232 6677 22260 6678
rect 22232 6651 22233 6677
rect 22233 6651 22259 6677
rect 22259 6651 22260 6677
rect 22232 6650 22260 6651
rect 22284 6677 22312 6678
rect 22284 6651 22285 6677
rect 22285 6651 22311 6677
rect 22311 6651 22312 6677
rect 22284 6650 22312 6651
rect 22336 6677 22364 6678
rect 22336 6651 22337 6677
rect 22337 6651 22363 6677
rect 22363 6651 22364 6677
rect 22336 6650 22364 6651
rect 22078 6398 22106 6426
rect 21854 6342 21882 6370
rect 21902 6285 21930 6286
rect 21902 6259 21903 6285
rect 21903 6259 21929 6285
rect 21929 6259 21930 6285
rect 21902 6258 21930 6259
rect 21954 6285 21982 6286
rect 21954 6259 21955 6285
rect 21955 6259 21981 6285
rect 21981 6259 21982 6285
rect 21954 6258 21982 6259
rect 22006 6285 22034 6286
rect 22006 6259 22007 6285
rect 22007 6259 22033 6285
rect 22033 6259 22034 6285
rect 22006 6258 22034 6259
rect 21798 6033 21826 6034
rect 21798 6007 21799 6033
rect 21799 6007 21825 6033
rect 21825 6007 21826 6033
rect 21798 6006 21826 6007
rect 22638 6118 22666 6146
rect 22232 5893 22260 5894
rect 22232 5867 22233 5893
rect 22233 5867 22259 5893
rect 22259 5867 22260 5893
rect 22232 5866 22260 5867
rect 22284 5893 22312 5894
rect 22284 5867 22285 5893
rect 22285 5867 22311 5893
rect 22311 5867 22312 5893
rect 22284 5866 22312 5867
rect 22336 5893 22364 5894
rect 22336 5867 22337 5893
rect 22337 5867 22363 5893
rect 22363 5867 22364 5893
rect 22336 5866 22364 5867
rect 22470 5838 22498 5866
rect 21902 5501 21930 5502
rect 21902 5475 21903 5501
rect 21903 5475 21929 5501
rect 21929 5475 21930 5501
rect 21902 5474 21930 5475
rect 21954 5501 21982 5502
rect 21954 5475 21955 5501
rect 21955 5475 21981 5501
rect 21981 5475 21982 5501
rect 21954 5474 21982 5475
rect 22006 5501 22034 5502
rect 22006 5475 22007 5501
rect 22007 5475 22033 5501
rect 22033 5475 22034 5501
rect 22006 5474 22034 5475
rect 21798 5249 21826 5250
rect 21798 5223 21799 5249
rect 21799 5223 21825 5249
rect 21825 5223 21826 5249
rect 21798 5222 21826 5223
rect 21518 5110 21546 5138
rect 22232 5109 22260 5110
rect 21462 5054 21490 5082
rect 22232 5083 22233 5109
rect 22233 5083 22259 5109
rect 22259 5083 22260 5109
rect 22232 5082 22260 5083
rect 22284 5109 22312 5110
rect 22284 5083 22285 5109
rect 22285 5083 22311 5109
rect 22311 5083 22312 5109
rect 22284 5082 22312 5083
rect 22336 5109 22364 5110
rect 22336 5083 22337 5109
rect 22337 5083 22363 5109
rect 22363 5083 22364 5109
rect 22336 5082 22364 5083
rect 21902 4717 21930 4718
rect 21902 4691 21903 4717
rect 21903 4691 21929 4717
rect 21929 4691 21930 4717
rect 21902 4690 21930 4691
rect 21954 4717 21982 4718
rect 21954 4691 21955 4717
rect 21955 4691 21981 4717
rect 21981 4691 21982 4717
rect 21954 4690 21982 4691
rect 22006 4717 22034 4718
rect 22006 4691 22007 4717
rect 22007 4691 22033 4717
rect 22033 4691 22034 4717
rect 22006 4690 22034 4691
rect 22232 4325 22260 4326
rect 22232 4299 22233 4325
rect 22233 4299 22259 4325
rect 22259 4299 22260 4325
rect 22232 4298 22260 4299
rect 22284 4325 22312 4326
rect 22284 4299 22285 4325
rect 22285 4299 22311 4325
rect 22311 4299 22312 4325
rect 22284 4298 22312 4299
rect 22336 4325 22364 4326
rect 22336 4299 22337 4325
rect 22337 4299 22363 4325
rect 22363 4299 22364 4325
rect 22336 4298 22364 4299
rect 21742 4073 21770 4074
rect 21742 4047 21743 4073
rect 21743 4047 21769 4073
rect 21769 4047 21770 4073
rect 21742 4046 21770 4047
rect 21966 3990 21994 4018
rect 21902 3933 21930 3934
rect 21902 3907 21903 3933
rect 21903 3907 21929 3933
rect 21929 3907 21930 3933
rect 21902 3906 21930 3907
rect 21954 3933 21982 3934
rect 21954 3907 21955 3933
rect 21955 3907 21981 3933
rect 21981 3907 21982 3933
rect 21954 3906 21982 3907
rect 22006 3933 22034 3934
rect 22006 3907 22007 3933
rect 22007 3907 22033 3933
rect 22033 3907 22034 3933
rect 22006 3906 22034 3907
rect 22232 3541 22260 3542
rect 22232 3515 22233 3541
rect 22233 3515 22259 3541
rect 22259 3515 22260 3541
rect 22232 3514 22260 3515
rect 22284 3541 22312 3542
rect 22284 3515 22285 3541
rect 22285 3515 22311 3541
rect 22311 3515 22312 3541
rect 22284 3514 22312 3515
rect 22336 3541 22364 3542
rect 22336 3515 22337 3541
rect 22337 3515 22363 3541
rect 22363 3515 22364 3541
rect 22336 3514 22364 3515
rect 21406 2870 21434 2898
rect 21742 3374 21770 3402
rect 21902 3149 21930 3150
rect 21902 3123 21903 3149
rect 21903 3123 21929 3149
rect 21929 3123 21930 3149
rect 21902 3122 21930 3123
rect 21954 3149 21982 3150
rect 21954 3123 21955 3149
rect 21955 3123 21981 3149
rect 21981 3123 21982 3149
rect 21954 3122 21982 3123
rect 22006 3149 22034 3150
rect 22006 3123 22007 3149
rect 22007 3123 22033 3149
rect 22033 3123 22034 3149
rect 22006 3122 22034 3123
rect 22078 2897 22106 2898
rect 22078 2871 22079 2897
rect 22079 2871 22105 2897
rect 22105 2871 22106 2897
rect 22078 2870 22106 2871
rect 22358 2897 22386 2898
rect 22358 2871 22359 2897
rect 22359 2871 22385 2897
rect 22385 2871 22386 2897
rect 22358 2870 22386 2871
rect 22232 2757 22260 2758
rect 22232 2731 22233 2757
rect 22233 2731 22259 2757
rect 22259 2731 22260 2757
rect 22232 2730 22260 2731
rect 22284 2757 22312 2758
rect 22284 2731 22285 2757
rect 22285 2731 22311 2757
rect 22311 2731 22312 2757
rect 22284 2730 22312 2731
rect 22336 2757 22364 2758
rect 22336 2731 22337 2757
rect 22337 2731 22363 2757
rect 22363 2731 22364 2757
rect 22336 2730 22364 2731
rect 22470 2646 22498 2674
rect 22470 2422 22498 2450
rect 21462 2310 21490 2338
rect 21902 2365 21930 2366
rect 21902 2339 21903 2365
rect 21903 2339 21929 2365
rect 21929 2339 21930 2365
rect 21902 2338 21930 2339
rect 21954 2365 21982 2366
rect 21954 2339 21955 2365
rect 21955 2339 21981 2365
rect 21981 2339 21982 2365
rect 21954 2338 21982 2339
rect 22006 2365 22034 2366
rect 22006 2339 22007 2365
rect 22007 2339 22033 2365
rect 22033 2339 22034 2365
rect 22006 2338 22034 2339
rect 21294 2169 21322 2170
rect 21294 2143 21295 2169
rect 21295 2143 21321 2169
rect 21321 2143 21322 2169
rect 21294 2142 21322 2143
rect 22232 1973 22260 1974
rect 22232 1947 22233 1973
rect 22233 1947 22259 1973
rect 22259 1947 22260 1973
rect 22232 1946 22260 1947
rect 22284 1973 22312 1974
rect 22284 1947 22285 1973
rect 22285 1947 22311 1973
rect 22311 1947 22312 1973
rect 22284 1946 22312 1947
rect 22336 1973 22364 1974
rect 22336 1947 22337 1973
rect 22337 1947 22363 1973
rect 22363 1947 22364 1973
rect 22336 1946 22364 1947
rect 22190 1833 22218 1834
rect 22190 1807 22191 1833
rect 22191 1807 22217 1833
rect 22217 1807 22218 1833
rect 22190 1806 22218 1807
rect 21238 1750 21266 1778
rect 21518 1582 21546 1610
rect 21350 1302 21378 1330
rect 21902 1581 21930 1582
rect 21902 1555 21903 1581
rect 21903 1555 21929 1581
rect 21929 1555 21930 1581
rect 21902 1554 21930 1555
rect 21954 1581 21982 1582
rect 21954 1555 21955 1581
rect 21955 1555 21981 1581
rect 21981 1555 21982 1581
rect 21954 1554 21982 1555
rect 22006 1581 22034 1582
rect 22006 1555 22007 1581
rect 22007 1555 22033 1581
rect 22033 1555 22034 1581
rect 22006 1554 22034 1555
rect 22078 1526 22106 1554
rect 21798 1105 21826 1106
rect 21798 1079 21799 1105
rect 21799 1079 21825 1105
rect 21825 1079 21826 1105
rect 21798 1078 21826 1079
rect 22582 5894 22610 5922
rect 22638 5614 22666 5642
rect 22638 4270 22666 4298
rect 22638 3262 22666 3290
rect 22582 2142 22610 2170
rect 22526 1358 22554 1386
rect 22582 1974 22610 2002
rect 22232 1189 22260 1190
rect 22232 1163 22233 1189
rect 22233 1163 22259 1189
rect 22259 1163 22260 1189
rect 22232 1162 22260 1163
rect 22284 1189 22312 1190
rect 22284 1163 22285 1189
rect 22285 1163 22311 1189
rect 22311 1163 22312 1189
rect 22284 1162 22312 1163
rect 22336 1189 22364 1190
rect 22336 1163 22337 1189
rect 22337 1163 22363 1189
rect 22363 1163 22364 1189
rect 22336 1162 22364 1163
rect 22022 1078 22050 1106
rect 21902 797 21930 798
rect 21902 771 21903 797
rect 21903 771 21929 797
rect 21929 771 21930 797
rect 21902 770 21930 771
rect 21954 797 21982 798
rect 21954 771 21955 797
rect 21955 771 21981 797
rect 21981 771 21982 797
rect 21954 770 21982 771
rect 22006 797 22034 798
rect 22006 771 22007 797
rect 22007 771 22033 797
rect 22033 771 22034 797
rect 22006 770 22034 771
rect 22638 1806 22666 1834
rect 22638 1414 22666 1442
rect 22694 1470 22722 1498
rect 22582 630 22610 658
rect 22638 966 22666 994
rect 21126 350 21154 378
rect 22232 405 22260 406
rect 22232 379 22233 405
rect 22233 379 22259 405
rect 22259 379 22260 405
rect 22232 378 22260 379
rect 22284 405 22312 406
rect 22284 379 22285 405
rect 22285 379 22311 405
rect 22311 379 22312 405
rect 22284 378 22312 379
rect 22336 405 22364 406
rect 22336 379 22337 405
rect 22337 379 22363 405
rect 22363 379 22364 405
rect 22336 378 22364 379
rect 23142 5641 23170 5642
rect 23142 5615 23143 5641
rect 23143 5615 23169 5641
rect 23169 5615 23170 5641
rect 23142 5614 23170 5615
rect 23254 6566 23282 6594
rect 23422 5894 23450 5922
rect 23478 6174 23506 6202
rect 23254 5446 23282 5474
rect 23310 5838 23338 5866
rect 23198 5166 23226 5194
rect 23646 5950 23674 5978
rect 23478 5110 23506 5138
rect 23646 5670 23674 5698
rect 23366 5054 23394 5082
rect 23310 4830 23338 4858
rect 22974 4494 23002 4522
rect 23422 3990 23450 4018
rect 23366 3374 23394 3402
rect 22750 1022 22778 1050
rect 22806 2814 22834 2842
rect 22694 798 22722 826
rect 22694 630 22722 658
rect 22638 294 22666 322
rect 23254 2030 23282 2058
rect 23366 1582 23394 1610
rect 23478 3766 23506 3794
rect 23534 3345 23562 3346
rect 23534 3319 23535 3345
rect 23535 3319 23561 3345
rect 23561 3319 23562 3345
rect 23534 3318 23562 3319
rect 23478 2478 23506 2506
rect 23422 1414 23450 1442
rect 23702 2982 23730 3010
rect 23814 1974 23842 2002
rect 23646 1806 23674 1834
rect 24094 5670 24122 5698
rect 23982 4998 24010 5026
rect 24094 4998 24122 5026
rect 23982 2310 24010 2338
rect 24262 4382 24290 4410
rect 24318 4270 24346 4298
rect 24318 3262 24346 3290
rect 24262 2814 24290 2842
rect 24374 2870 24402 2898
rect 24038 1526 24066 1554
rect 24206 2646 24234 2674
rect 23870 1302 23898 1330
rect 23534 1190 23562 1218
rect 22918 1105 22946 1106
rect 22918 1079 22919 1105
rect 22919 1079 22945 1105
rect 22945 1079 22946 1105
rect 22918 1078 22946 1079
rect 23478 910 23506 938
rect 23478 462 23506 490
rect 22806 294 22834 322
rect 24318 2590 24346 2618
rect 24262 2113 24290 2114
rect 24262 2087 24263 2113
rect 24263 2087 24289 2113
rect 24289 2087 24290 2113
rect 24262 2086 24290 2087
rect 24374 2366 24402 2394
rect 24318 1806 24346 1834
rect 24318 1470 24346 1498
rect 25158 4270 25186 4298
rect 25662 6566 25690 6594
rect 25550 5054 25578 5082
rect 25158 3374 25186 3402
rect 24934 2478 24962 2506
rect 25214 2561 25242 2562
rect 25214 2535 25215 2561
rect 25215 2535 25241 2561
rect 25241 2535 25242 2561
rect 25214 2534 25242 2535
rect 24766 2254 24794 2282
rect 24486 1078 24514 1106
rect 24598 993 24626 994
rect 24598 967 24599 993
rect 24599 967 24625 993
rect 24625 967 24626 993
rect 24598 966 24626 967
rect 24206 798 24234 826
rect 24038 238 24066 266
rect 23310 182 23338 210
rect 21854 70 21882 98
rect 24990 1862 25018 1890
rect 25494 3345 25522 3346
rect 25494 3319 25495 3345
rect 25495 3319 25521 3345
rect 25521 3319 25522 3345
rect 25494 3318 25522 3319
rect 25438 3038 25466 3066
rect 25326 2758 25354 2786
rect 25326 2534 25354 2562
rect 25438 1582 25466 1610
rect 24878 1049 24906 1050
rect 24878 1023 24879 1049
rect 24879 1023 24905 1049
rect 24905 1023 24906 1049
rect 24878 1022 24906 1023
rect 24878 406 24906 434
rect 24878 294 24906 322
rect 25214 126 25242 154
rect 26054 6593 26082 6594
rect 26054 6567 26055 6593
rect 26055 6567 26081 6593
rect 26081 6567 26082 6593
rect 26054 6566 26082 6567
rect 25886 6174 25914 6202
rect 26054 6454 26082 6482
rect 25774 6118 25802 6146
rect 26558 6734 26586 6762
rect 26334 6510 26362 6538
rect 26558 6230 26586 6258
rect 26278 6201 26306 6202
rect 26278 6175 26279 6201
rect 26279 6175 26305 6201
rect 26305 6175 26306 6201
rect 26278 6174 26306 6175
rect 26222 5278 26250 5306
rect 26390 4606 26418 4634
rect 26782 6089 26810 6090
rect 26782 6063 26783 6089
rect 26783 6063 26809 6089
rect 26809 6063 26810 6089
rect 26782 6062 26810 6063
rect 26838 5838 26866 5866
rect 26894 6174 26922 6202
rect 26614 5110 26642 5138
rect 27678 6902 27706 6930
rect 27454 6846 27482 6874
rect 27230 6566 27258 6594
rect 27454 6734 27482 6762
rect 27006 6174 27034 6202
rect 27062 6510 27090 6538
rect 27902 6398 27930 6426
rect 27958 6230 27986 6258
rect 27846 6201 27874 6202
rect 27846 6175 27847 6201
rect 27847 6175 27873 6201
rect 27873 6175 27874 6201
rect 27846 6174 27874 6175
rect 28126 6118 28154 6146
rect 28182 6902 28210 6930
rect 27174 6006 27202 6034
rect 27286 5838 27314 5866
rect 27006 5222 27034 5250
rect 26894 4382 26922 4410
rect 26950 2702 26978 2730
rect 26446 2422 26474 2450
rect 26670 2478 26698 2506
rect 25606 1638 25634 1666
rect 26054 2198 26082 2226
rect 26054 1638 26082 1666
rect 26054 1526 26082 1554
rect 26670 1470 26698 1498
rect 26222 1414 26250 1442
rect 25550 574 25578 602
rect 26054 1134 26082 1162
rect 26054 462 26082 490
rect 25270 70 25298 98
rect 26278 854 26306 882
rect 26894 966 26922 994
rect 27174 2422 27202 2450
rect 28238 6593 28266 6594
rect 28238 6567 28239 6593
rect 28239 6567 28265 6593
rect 28265 6567 28266 6593
rect 28238 6566 28266 6567
rect 28574 6510 28602 6538
rect 28630 6846 28658 6874
rect 28350 6454 28378 6482
rect 28574 6118 28602 6146
rect 27734 5502 27762 5530
rect 27678 5305 27706 5306
rect 27678 5279 27679 5305
rect 27679 5279 27705 5305
rect 27705 5279 27706 5305
rect 27678 5278 27706 5279
rect 27958 4270 27986 4298
rect 27958 4129 27986 4130
rect 27958 4103 27959 4129
rect 27959 4103 27985 4129
rect 27985 4103 27986 4129
rect 27958 4102 27986 4103
rect 27734 3094 27762 3122
rect 27566 2366 27594 2394
rect 27846 2225 27874 2226
rect 27846 2199 27847 2225
rect 27847 2199 27873 2225
rect 27873 2199 27874 2225
rect 27846 2198 27874 2199
rect 27174 1582 27202 1610
rect 28070 5249 28098 5250
rect 28070 5223 28071 5249
rect 28071 5223 28097 5249
rect 28097 5223 28098 5249
rect 28070 5222 28098 5223
rect 28238 5054 28266 5082
rect 28126 4942 28154 4970
rect 28238 4857 28266 4858
rect 28238 4831 28239 4857
rect 28239 4831 28265 4857
rect 28265 4831 28266 4857
rect 28238 4830 28266 4831
rect 28238 4438 28266 4466
rect 28462 5446 28490 5474
rect 28350 4577 28378 4578
rect 28350 4551 28351 4577
rect 28351 4551 28377 4577
rect 28377 4551 28378 4577
rect 28350 4550 28378 4551
rect 29022 6622 29050 6650
rect 28798 6118 28826 6146
rect 29022 6454 29050 6482
rect 28910 5670 28938 5698
rect 28574 4326 28602 4354
rect 28630 4214 28658 4242
rect 28630 3486 28658 3514
rect 29022 5334 29050 5362
rect 28966 4969 28994 4970
rect 28966 4943 28967 4969
rect 28967 4943 28993 4969
rect 28993 4943 28994 4969
rect 28966 4942 28994 4943
rect 28742 4382 28770 4410
rect 28910 4185 28938 4186
rect 28910 4159 28911 4185
rect 28911 4159 28937 4185
rect 28937 4159 28938 4185
rect 28910 4158 28938 4159
rect 28854 4046 28882 4074
rect 28910 3822 28938 3850
rect 28686 3038 28714 3066
rect 28966 3094 28994 3122
rect 28686 2841 28714 2842
rect 28686 2815 28687 2841
rect 28687 2815 28713 2841
rect 28713 2815 28714 2841
rect 28686 2814 28714 2815
rect 28630 2702 28658 2730
rect 28294 2478 28322 2506
rect 28070 2057 28098 2058
rect 28070 2031 28071 2057
rect 28071 2031 28097 2057
rect 28097 2031 28098 2057
rect 28070 2030 28098 2031
rect 28014 1022 28042 1050
rect 26950 798 26978 826
rect 29470 6566 29498 6594
rect 29414 6425 29442 6426
rect 29414 6399 29415 6425
rect 29415 6399 29441 6425
rect 29441 6399 29442 6425
rect 29414 6398 29442 6399
rect 29246 6342 29274 6370
rect 29414 6118 29442 6146
rect 29302 5894 29330 5922
rect 29694 6118 29722 6146
rect 29806 6342 29834 6370
rect 29470 5782 29498 5810
rect 29414 4913 29442 4914
rect 29414 4887 29415 4913
rect 29415 4887 29441 4913
rect 29441 4887 29442 4913
rect 29414 4886 29442 4887
rect 29358 4662 29386 4690
rect 29190 3681 29218 3682
rect 29190 3655 29191 3681
rect 29191 3655 29217 3681
rect 29217 3655 29218 3681
rect 29190 3654 29218 3655
rect 29414 3598 29442 3626
rect 29526 5697 29554 5698
rect 29526 5671 29527 5697
rect 29527 5671 29553 5697
rect 29553 5671 29554 5697
rect 29526 5670 29554 5671
rect 29526 5222 29554 5250
rect 29750 4913 29778 4914
rect 29750 4887 29751 4913
rect 29751 4887 29777 4913
rect 29777 4887 29778 4913
rect 29750 4886 29778 4887
rect 30422 6958 30450 6986
rect 30310 6622 30338 6650
rect 30254 6537 30282 6538
rect 30254 6511 30255 6537
rect 30255 6511 30281 6537
rect 30281 6511 30282 6537
rect 30254 6510 30282 6511
rect 29918 6342 29946 6370
rect 29526 3542 29554 3570
rect 29246 3206 29274 3234
rect 29190 2617 29218 2618
rect 29190 2591 29191 2617
rect 29191 2591 29217 2617
rect 29217 2591 29218 2617
rect 29190 2590 29218 2591
rect 29078 2422 29106 2450
rect 29414 2310 29442 2338
rect 28910 1638 28938 1666
rect 29862 4102 29890 4130
rect 29806 3374 29834 3402
rect 29694 3150 29722 3178
rect 29638 3009 29666 3010
rect 29638 2983 29639 3009
rect 29639 2983 29665 3009
rect 29665 2983 29666 3009
rect 29638 2982 29666 2983
rect 29694 2673 29722 2674
rect 29694 2647 29695 2673
rect 29695 2647 29721 2673
rect 29721 2647 29722 2673
rect 29694 2646 29722 2647
rect 29694 1777 29722 1778
rect 29694 1751 29695 1777
rect 29695 1751 29721 1777
rect 29721 1751 29722 1777
rect 29694 1750 29722 1751
rect 30142 4774 30170 4802
rect 30198 4830 30226 4858
rect 30254 4465 30282 4466
rect 30254 4439 30255 4465
rect 30255 4439 30281 4465
rect 30281 4439 30282 4465
rect 30254 4438 30282 4439
rect 30254 3737 30282 3738
rect 30254 3711 30255 3737
rect 30255 3711 30281 3737
rect 30281 3711 30282 3737
rect 30254 3710 30282 3711
rect 30254 3430 30282 3458
rect 29974 3345 30002 3346
rect 29974 3319 29975 3345
rect 29975 3319 30001 3345
rect 30001 3319 30002 3345
rect 29974 3318 30002 3319
rect 30142 3262 30170 3290
rect 30310 3094 30338 3122
rect 30142 2702 30170 2730
rect 29974 2561 30002 2562
rect 29974 2535 29975 2561
rect 29975 2535 30001 2561
rect 30001 2535 30002 2561
rect 29974 2534 30002 2535
rect 32102 6734 32130 6762
rect 31262 6593 31290 6594
rect 31262 6567 31263 6593
rect 31263 6567 31289 6593
rect 31289 6567 31290 6593
rect 31262 6566 31290 6567
rect 31374 6510 31402 6538
rect 30590 6342 30618 6370
rect 30422 5278 30450 5306
rect 30646 4857 30674 4858
rect 30646 4831 30647 4857
rect 30647 4831 30673 4857
rect 30673 4831 30674 4857
rect 30646 4830 30674 4831
rect 31094 6145 31122 6146
rect 31094 6119 31095 6145
rect 31095 6119 31121 6145
rect 31121 6119 31122 6145
rect 31094 6118 31122 6119
rect 30982 5614 31010 5642
rect 31094 5502 31122 5530
rect 31094 5390 31122 5418
rect 30758 5054 30786 5082
rect 31094 5166 31122 5194
rect 30758 4633 30786 4634
rect 30758 4607 30759 4633
rect 30759 4607 30785 4633
rect 30785 4607 30786 4633
rect 30758 4606 30786 4607
rect 30534 4185 30562 4186
rect 30534 4159 30535 4185
rect 30535 4159 30561 4185
rect 30561 4159 30562 4185
rect 30534 4158 30562 4159
rect 30590 3542 30618 3570
rect 30758 3374 30786 3402
rect 30758 3065 30786 3066
rect 30758 3039 30759 3065
rect 30759 3039 30785 3065
rect 30785 3039 30786 3065
rect 30758 3038 30786 3039
rect 31094 4830 31122 4858
rect 31822 6286 31850 6314
rect 31542 5838 31570 5866
rect 31486 5614 31514 5642
rect 31262 4942 31290 4970
rect 31318 5390 31346 5418
rect 31318 4606 31346 4634
rect 31486 4886 31514 4914
rect 31430 4718 31458 4746
rect 31374 4494 31402 4522
rect 31430 4270 31458 4298
rect 31542 4158 31570 4186
rect 31878 6062 31906 6090
rect 31878 4662 31906 4690
rect 31822 4102 31850 4130
rect 31542 4046 31570 4074
rect 31430 3822 31458 3850
rect 31094 3486 31122 3514
rect 30982 3318 31010 3346
rect 30870 2982 30898 3010
rect 30646 2926 30674 2954
rect 30534 2617 30562 2618
rect 30534 2591 30535 2617
rect 30535 2591 30561 2617
rect 30561 2591 30562 2617
rect 30534 2590 30562 2591
rect 30926 2561 30954 2562
rect 30926 2535 30927 2561
rect 30927 2535 30953 2561
rect 30953 2535 30954 2561
rect 30926 2534 30954 2535
rect 30366 2198 30394 2226
rect 29918 1694 29946 1722
rect 29526 1526 29554 1554
rect 29246 1414 29274 1442
rect 29190 1329 29218 1330
rect 29190 1303 29191 1329
rect 29191 1303 29217 1329
rect 29217 1303 29218 1329
rect 29190 1302 29218 1303
rect 28798 1049 28826 1050
rect 28798 1023 28799 1049
rect 28799 1023 28825 1049
rect 28825 1023 28826 1049
rect 28798 1022 28826 1023
rect 28574 993 28602 994
rect 28574 967 28575 993
rect 28575 967 28601 993
rect 28601 967 28602 993
rect 28574 966 28602 967
rect 30254 1414 30282 1442
rect 30534 2030 30562 2058
rect 29638 1385 29666 1386
rect 29638 1359 29639 1385
rect 29639 1359 29665 1385
rect 29665 1359 29666 1385
rect 29638 1358 29666 1359
rect 29414 1246 29442 1274
rect 30086 1302 30114 1330
rect 29694 1190 29722 1218
rect 29414 1134 29442 1162
rect 28966 910 28994 938
rect 28910 686 28938 714
rect 29134 854 29162 882
rect 28350 630 28378 658
rect 26894 518 26922 546
rect 27678 574 27706 602
rect 29974 993 30002 994
rect 29974 967 29975 993
rect 29975 967 30001 993
rect 30001 967 30002 993
rect 29974 966 30002 967
rect 29414 406 29442 434
rect 29302 350 29330 378
rect 30142 1049 30170 1050
rect 30142 1023 30143 1049
rect 30143 1023 30169 1049
rect 30169 1023 30170 1049
rect 30142 1022 30170 1023
rect 30254 742 30282 770
rect 30646 1806 30674 1834
rect 30926 1777 30954 1778
rect 30926 1751 30927 1777
rect 30927 1751 30953 1777
rect 30953 1751 30954 1777
rect 30926 1750 30954 1751
rect 30646 1721 30674 1722
rect 30646 1695 30647 1721
rect 30647 1695 30673 1721
rect 30673 1695 30674 1721
rect 30646 1694 30674 1695
rect 30646 1329 30674 1330
rect 30646 1303 30647 1329
rect 30647 1303 30673 1329
rect 30673 1303 30674 1329
rect 30646 1302 30674 1303
rect 30926 993 30954 994
rect 30926 967 30927 993
rect 30927 967 30953 993
rect 30953 967 30954 993
rect 30926 966 30954 967
rect 30646 881 30674 882
rect 30646 855 30647 881
rect 30647 855 30673 881
rect 30673 855 30674 881
rect 30646 854 30674 855
rect 31094 2646 31122 2674
rect 31094 1385 31122 1386
rect 31094 1359 31095 1385
rect 31095 1359 31121 1385
rect 31121 1359 31122 1385
rect 31094 1358 31122 1359
rect 31430 3598 31458 3626
rect 31542 3150 31570 3178
rect 32102 3038 32130 3066
rect 31318 2702 31346 2730
rect 31262 2590 31290 2618
rect 31262 2254 31290 2282
rect 31542 2478 31570 2506
rect 31430 2030 31458 2058
rect 31318 1694 31346 1722
rect 31542 1582 31570 1610
rect 31318 1358 31346 1386
rect 31150 1134 31178 1162
rect 31374 1302 31402 1330
rect 31038 798 31066 826
rect 31094 518 31122 546
rect 30590 462 30618 490
rect 29806 238 29834 266
rect 16758 14 16786 42
rect 31430 1134 31458 1162
rect 31542 910 31570 938
rect 31374 14 31402 42
<< metal3 >>
rect 8582 7014 16254 7042
rect 16282 7014 16287 7042
rect 0 6986 56 7000
rect 8582 6986 8610 7014
rect 32144 6986 32200 7000
rect 0 6958 126 6986
rect 154 6958 159 6986
rect 8577 6958 8582 6986
rect 8610 6958 8615 6986
rect 9809 6958 9814 6986
rect 9842 6958 15582 6986
rect 15610 6958 15615 6986
rect 18993 6958 18998 6986
rect 19026 6958 22526 6986
rect 22554 6958 22559 6986
rect 30417 6958 30422 6986
rect 30450 6958 32200 6986
rect 0 6944 56 6958
rect 32144 6944 32200 6958
rect 27673 6902 27678 6930
rect 27706 6902 28182 6930
rect 28210 6902 28215 6930
rect 9697 6846 9702 6874
rect 9730 6846 14462 6874
rect 14490 6846 14495 6874
rect 27449 6846 27454 6874
rect 27482 6846 28630 6874
rect 28658 6846 28663 6874
rect 1857 6790 1862 6818
rect 1890 6790 2814 6818
rect 2842 6790 2847 6818
rect 10257 6790 10262 6818
rect 10290 6790 18270 6818
rect 18298 6790 18303 6818
rect 0 6762 56 6776
rect 32144 6762 32200 6776
rect 0 6734 1218 6762
rect 1801 6734 1806 6762
rect 1834 6734 2366 6762
rect 2394 6734 2399 6762
rect 11153 6734 11158 6762
rect 11186 6734 13454 6762
rect 13561 6734 13566 6762
rect 13594 6734 13958 6762
rect 13986 6734 13991 6762
rect 26553 6734 26558 6762
rect 26586 6734 27454 6762
rect 27482 6734 27487 6762
rect 32097 6734 32102 6762
rect 32130 6734 32200 6762
rect 0 6720 56 6734
rect 1190 6706 1218 6734
rect 13426 6706 13454 6734
rect 32144 6720 32200 6734
rect 1190 6678 2086 6706
rect 2114 6678 2119 6706
rect 13426 6678 17486 6706
rect 17514 6678 17519 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 22227 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22369 6678
rect 4881 6622 4886 6650
rect 4914 6622 5950 6650
rect 5978 6622 5983 6650
rect 8689 6622 8694 6650
rect 8722 6622 9758 6650
rect 9786 6622 9791 6650
rect 13426 6622 19838 6650
rect 19866 6622 19871 6650
rect 29017 6622 29022 6650
rect 29050 6622 30310 6650
rect 30338 6622 30343 6650
rect 1241 6566 1246 6594
rect 1274 6566 2142 6594
rect 2170 6566 2175 6594
rect 2977 6566 2982 6594
rect 3010 6566 3486 6594
rect 3514 6566 3519 6594
rect 3761 6566 3766 6594
rect 3794 6566 4382 6594
rect 4410 6566 4415 6594
rect 4993 6566 4998 6594
rect 5026 6566 5278 6594
rect 5306 6566 5311 6594
rect 5665 6566 5670 6594
rect 5698 6566 6622 6594
rect 6650 6566 6655 6594
rect 8185 6566 8190 6594
rect 8218 6566 8638 6594
rect 8666 6566 8671 6594
rect 9473 6566 9478 6594
rect 9506 6566 10430 6594
rect 10458 6566 10463 6594
rect 10593 6566 10598 6594
rect 10626 6566 11102 6594
rect 11130 6566 11135 6594
rect 11377 6566 11382 6594
rect 11410 6566 11998 6594
rect 12026 6566 12031 6594
rect 0 6538 56 6552
rect 13426 6538 13454 6622
rect 17593 6566 17598 6594
rect 17626 6566 23254 6594
rect 23282 6566 23287 6594
rect 25657 6566 25662 6594
rect 25690 6566 26054 6594
rect 26082 6566 26087 6594
rect 27225 6566 27230 6594
rect 27258 6566 28238 6594
rect 28266 6566 28271 6594
rect 29465 6566 29470 6594
rect 29498 6566 31262 6594
rect 31290 6566 31295 6594
rect 32144 6538 32200 6552
rect 0 6510 798 6538
rect 826 6510 831 6538
rect 7401 6510 7406 6538
rect 7434 6510 8414 6538
rect 8442 6510 8447 6538
rect 9865 6510 9870 6538
rect 9898 6510 13454 6538
rect 16529 6510 16534 6538
rect 16562 6510 21630 6538
rect 21658 6510 21663 6538
rect 26329 6510 26334 6538
rect 26362 6510 27062 6538
rect 27090 6510 27095 6538
rect 28569 6510 28574 6538
rect 28602 6510 30254 6538
rect 30282 6510 30287 6538
rect 31369 6510 31374 6538
rect 31402 6510 32200 6538
rect 0 6496 56 6510
rect 32144 6496 32200 6510
rect 1073 6454 1078 6482
rect 1106 6454 6454 6482
rect 6482 6454 6487 6482
rect 7457 6454 7462 6482
rect 7490 6454 7966 6482
rect 7994 6454 7999 6482
rect 9753 6454 9758 6482
rect 9786 6454 12670 6482
rect 12698 6454 12703 6482
rect 14905 6454 14910 6482
rect 14938 6454 26054 6482
rect 26082 6454 26087 6482
rect 28345 6454 28350 6482
rect 28378 6454 29022 6482
rect 29050 6454 29055 6482
rect 6953 6398 6958 6426
rect 6986 6398 7518 6426
rect 7546 6398 7551 6426
rect 14009 6398 14014 6426
rect 14042 6398 18942 6426
rect 18970 6398 18975 6426
rect 19105 6398 19110 6426
rect 19138 6398 22078 6426
rect 22106 6398 22111 6426
rect 27897 6398 27902 6426
rect 27930 6398 29414 6426
rect 29442 6398 29447 6426
rect 8969 6342 8974 6370
rect 9002 6342 9534 6370
rect 9562 6342 9567 6370
rect 11657 6342 11662 6370
rect 11690 6342 14350 6370
rect 14378 6342 14383 6370
rect 15465 6342 15470 6370
rect 15498 6342 21854 6370
rect 21882 6342 21887 6370
rect 29241 6342 29246 6370
rect 29274 6342 29806 6370
rect 29834 6342 29839 6370
rect 29913 6342 29918 6370
rect 29946 6342 30590 6370
rect 30618 6342 30623 6370
rect 0 6314 56 6328
rect 32144 6314 32200 6328
rect 0 6286 462 6314
rect 490 6286 495 6314
rect 14121 6286 14126 6314
rect 14154 6286 16030 6314
rect 16058 6286 16063 6314
rect 18657 6286 18662 6314
rect 18690 6286 20958 6314
rect 20986 6286 20991 6314
rect 31817 6286 31822 6314
rect 31850 6286 32200 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 21897 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22039 6286
rect 32144 6272 32200 6286
rect 6225 6230 6230 6258
rect 6258 6230 10038 6258
rect 10066 6230 10071 6258
rect 13169 6230 13174 6258
rect 13202 6230 15358 6258
rect 15386 6230 15391 6258
rect 16809 6230 16814 6258
rect 16842 6230 19390 6258
rect 19418 6230 19423 6258
rect 22521 6230 22526 6258
rect 22554 6230 26418 6258
rect 26553 6230 26558 6258
rect 26586 6230 27958 6258
rect 27986 6230 27991 6258
rect 26390 6202 26418 6230
rect 4265 6174 4270 6202
rect 4298 6174 4830 6202
rect 4858 6174 4863 6202
rect 5833 6174 5838 6202
rect 5866 6174 6398 6202
rect 6426 6174 6431 6202
rect 6673 6174 6678 6202
rect 6706 6174 7462 6202
rect 7490 6174 7495 6202
rect 7546 6174 15890 6202
rect 16585 6174 16590 6202
rect 16618 6174 18830 6202
rect 18858 6174 18863 6202
rect 18937 6174 18942 6202
rect 18970 6174 20174 6202
rect 20202 6174 20207 6202
rect 20953 6174 20958 6202
rect 20986 6174 23478 6202
rect 23506 6174 23511 6202
rect 25881 6174 25886 6202
rect 25914 6174 26278 6202
rect 26306 6174 26311 6202
rect 26390 6174 26894 6202
rect 26922 6174 26927 6202
rect 27001 6174 27006 6202
rect 27034 6174 27846 6202
rect 27874 6174 27879 6202
rect 7546 6146 7574 6174
rect 15862 6146 15890 6174
rect 1409 6118 1414 6146
rect 1442 6118 4298 6146
rect 5329 6118 5334 6146
rect 5362 6118 7574 6146
rect 13113 6118 13118 6146
rect 13146 6118 13454 6146
rect 13482 6118 13487 6146
rect 14457 6118 14462 6146
rect 14490 6118 15190 6146
rect 15218 6118 15223 6146
rect 15862 6118 22526 6146
rect 22554 6118 22559 6146
rect 22633 6118 22638 6146
rect 22666 6118 25774 6146
rect 25802 6118 25807 6146
rect 28121 6118 28126 6146
rect 28154 6118 28574 6146
rect 28602 6118 28607 6146
rect 28793 6118 28798 6146
rect 28826 6118 29414 6146
rect 29442 6118 29447 6146
rect 29689 6118 29694 6146
rect 29722 6118 31094 6146
rect 31122 6118 31127 6146
rect 0 6090 56 6104
rect 4270 6090 4298 6118
rect 32144 6090 32200 6104
rect 0 6062 4214 6090
rect 4270 6062 9422 6090
rect 9450 6062 9455 6090
rect 12609 6062 12614 6090
rect 12642 6062 14518 6090
rect 14546 6062 14551 6090
rect 14849 6062 14854 6090
rect 14882 6062 18718 6090
rect 18746 6062 18751 6090
rect 18825 6062 18830 6090
rect 18858 6062 20510 6090
rect 20538 6062 20543 6090
rect 20673 6062 20678 6090
rect 20706 6062 26782 6090
rect 26810 6062 26815 6090
rect 31873 6062 31878 6090
rect 31906 6062 32200 6090
rect 0 6048 56 6062
rect 4186 6034 4214 6062
rect 32144 6048 32200 6062
rect 2193 6006 2198 6034
rect 2226 6006 2926 6034
rect 2954 6006 2959 6034
rect 4186 6006 6230 6034
rect 6258 6006 6263 6034
rect 6337 6006 6342 6034
rect 6370 6006 7070 6034
rect 7098 6006 7103 6034
rect 13057 6006 13062 6034
rect 13090 6006 13734 6034
rect 13762 6006 13767 6034
rect 13841 6006 13846 6034
rect 13874 6006 15694 6034
rect 15722 6006 15727 6034
rect 15913 6006 15918 6034
rect 15946 6006 19166 6034
rect 19194 6006 19199 6034
rect 21793 6006 21798 6034
rect 21826 6006 27174 6034
rect 27202 6006 27207 6034
rect 4545 5950 4550 5978
rect 4578 5950 7350 5978
rect 7378 5950 7383 5978
rect 7457 5950 7462 5978
rect 7490 5950 10486 5978
rect 10514 5950 10519 5978
rect 12166 5950 13790 5978
rect 13818 5950 13823 5978
rect 15353 5950 15358 5978
rect 15386 5950 18942 5978
rect 18970 5950 18975 5978
rect 19049 5950 19054 5978
rect 19082 5950 20398 5978
rect 20426 5950 20431 5978
rect 22470 5950 23646 5978
rect 23674 5950 23679 5978
rect 6113 5894 6118 5922
rect 6146 5894 7518 5922
rect 7546 5894 7551 5922
rect 9193 5894 9198 5922
rect 9226 5894 9231 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 9198 5866 9226 5894
rect 12166 5866 12194 5950
rect 12777 5894 12782 5922
rect 12810 5894 14238 5922
rect 14266 5894 14271 5922
rect 14513 5894 14518 5922
rect 14546 5894 15414 5922
rect 15442 5894 15447 5922
rect 15526 5894 17654 5922
rect 17682 5894 17687 5922
rect 18041 5894 18046 5922
rect 18074 5894 20790 5922
rect 20818 5894 20823 5922
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 15526 5866 15554 5894
rect 22227 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22369 5894
rect 22470 5866 22498 5950
rect 22577 5894 22582 5922
rect 22610 5894 23422 5922
rect 23450 5894 23455 5922
rect 23534 5894 29302 5922
rect 29330 5894 29335 5922
rect 23534 5866 23562 5894
rect 32144 5866 32200 5880
rect 0 5838 2086 5866
rect 2114 5838 2119 5866
rect 9198 5838 10878 5866
rect 10906 5838 10911 5866
rect 11433 5838 11438 5866
rect 11466 5838 12194 5866
rect 12441 5838 12446 5866
rect 12474 5838 15554 5866
rect 22465 5838 22470 5866
rect 22498 5838 22503 5866
rect 23305 5838 23310 5866
rect 23338 5838 23562 5866
rect 26833 5838 26838 5866
rect 26866 5838 27286 5866
rect 27314 5838 27319 5866
rect 31537 5838 31542 5866
rect 31570 5838 32200 5866
rect 0 5824 56 5838
rect 32144 5824 32200 5838
rect 2305 5782 2310 5810
rect 2338 5782 2590 5810
rect 2618 5782 2623 5810
rect 3873 5782 3878 5810
rect 3906 5782 4158 5810
rect 4186 5782 4191 5810
rect 5441 5782 5446 5810
rect 5474 5782 5726 5810
rect 5754 5782 5759 5810
rect 6057 5782 6062 5810
rect 6090 5782 14014 5810
rect 14042 5782 14047 5810
rect 14289 5782 14294 5810
rect 14322 5782 19614 5810
rect 19642 5782 19647 5810
rect 20169 5782 20174 5810
rect 20202 5782 29470 5810
rect 29498 5782 29503 5810
rect 7513 5726 7518 5754
rect 7546 5726 14070 5754
rect 14098 5726 14103 5754
rect 14849 5726 14854 5754
rect 14882 5726 21238 5754
rect 21266 5726 21271 5754
rect 3313 5670 3318 5698
rect 3346 5670 5446 5698
rect 5474 5670 5479 5698
rect 7345 5670 7350 5698
rect 7378 5670 11158 5698
rect 11186 5670 11191 5698
rect 11993 5670 11998 5698
rect 12026 5670 12726 5698
rect 12754 5670 12759 5698
rect 14009 5670 14014 5698
rect 14042 5670 15918 5698
rect 15946 5670 15951 5698
rect 17817 5670 17822 5698
rect 17850 5670 19558 5698
rect 19586 5670 19591 5698
rect 23641 5670 23646 5698
rect 23674 5670 24094 5698
rect 24122 5670 24127 5698
rect 28905 5670 28910 5698
rect 28938 5670 29526 5698
rect 29554 5670 29559 5698
rect 0 5642 56 5656
rect 32144 5642 32200 5656
rect 0 5614 882 5642
rect 961 5614 966 5642
rect 994 5614 8638 5642
rect 8666 5614 8671 5642
rect 10033 5614 10038 5642
rect 10066 5614 13398 5642
rect 13426 5614 13431 5642
rect 14233 5614 14238 5642
rect 14266 5614 22638 5642
rect 22666 5614 22671 5642
rect 23137 5614 23142 5642
rect 23170 5614 30982 5642
rect 31010 5614 31015 5642
rect 31481 5614 31486 5642
rect 31514 5614 32200 5642
rect 0 5600 56 5614
rect 854 5586 882 5614
rect 32144 5600 32200 5614
rect 854 5558 1190 5586
rect 1218 5558 1223 5586
rect 2585 5558 2590 5586
rect 2618 5558 4214 5586
rect 4242 5558 4247 5586
rect 10481 5558 10486 5586
rect 10514 5558 15918 5586
rect 15946 5558 15951 5586
rect 16193 5558 16198 5586
rect 16226 5558 19054 5586
rect 19082 5558 19087 5586
rect 4153 5502 4158 5530
rect 4186 5502 7350 5530
rect 7378 5502 7383 5530
rect 13426 5502 16366 5530
rect 16394 5502 16399 5530
rect 16641 5502 16646 5530
rect 16674 5502 19446 5530
rect 19474 5502 19479 5530
rect 27729 5502 27734 5530
rect 27762 5502 31094 5530
rect 31122 5502 31127 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 13426 5474 13454 5502
rect 21897 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22039 5502
rect 2585 5446 2590 5474
rect 2618 5446 6734 5474
rect 6762 5446 6767 5474
rect 12105 5446 12110 5474
rect 12138 5446 13454 5474
rect 13673 5446 13678 5474
rect 13706 5446 14294 5474
rect 14322 5446 14327 5474
rect 15185 5446 15190 5474
rect 15218 5446 18550 5474
rect 18578 5446 18583 5474
rect 21121 5446 21126 5474
rect 21154 5446 21798 5474
rect 21826 5446 21831 5474
rect 23249 5446 23254 5474
rect 23282 5446 28462 5474
rect 28490 5446 28495 5474
rect 0 5418 56 5432
rect 32144 5418 32200 5432
rect 0 5390 6286 5418
rect 6314 5390 6319 5418
rect 10817 5390 10822 5418
rect 10850 5390 12194 5418
rect 12665 5390 12670 5418
rect 12698 5390 14070 5418
rect 14098 5390 14103 5418
rect 14177 5390 14182 5418
rect 14210 5390 31094 5418
rect 31122 5390 31127 5418
rect 31313 5390 31318 5418
rect 31346 5390 32200 5418
rect 0 5376 56 5390
rect 12166 5362 12194 5390
rect 32144 5376 32200 5390
rect 6505 5334 6510 5362
rect 6538 5334 11774 5362
rect 11802 5334 11807 5362
rect 12166 5334 14294 5362
rect 14322 5334 14327 5362
rect 14401 5334 14406 5362
rect 14434 5334 14630 5362
rect 14658 5334 14663 5362
rect 15577 5334 15582 5362
rect 15610 5334 29022 5362
rect 29050 5334 29055 5362
rect 1129 5278 1134 5306
rect 1162 5278 10066 5306
rect 11601 5278 11606 5306
rect 11634 5278 12614 5306
rect 12642 5278 12647 5306
rect 13393 5278 13398 5306
rect 13426 5278 14854 5306
rect 14882 5278 14887 5306
rect 17873 5278 17878 5306
rect 17906 5278 26222 5306
rect 26250 5278 26255 5306
rect 27673 5278 27678 5306
rect 27706 5278 30422 5306
rect 30450 5278 30455 5306
rect 10038 5250 10066 5278
rect 457 5222 462 5250
rect 490 5222 1526 5250
rect 1554 5222 1559 5250
rect 2081 5222 2086 5250
rect 2114 5222 4214 5250
rect 6113 5222 6118 5250
rect 6146 5222 9478 5250
rect 9506 5222 9511 5250
rect 10038 5222 16814 5250
rect 16842 5222 16847 5250
rect 17145 5222 17150 5250
rect 17178 5222 18214 5250
rect 18242 5222 18247 5250
rect 18489 5222 18494 5250
rect 18522 5222 21658 5250
rect 21793 5222 21798 5250
rect 21826 5222 27006 5250
rect 27034 5222 27039 5250
rect 28065 5222 28070 5250
rect 28098 5222 29526 5250
rect 29554 5222 29559 5250
rect 0 5194 56 5208
rect 0 5166 3878 5194
rect 3906 5166 3911 5194
rect 0 5152 56 5166
rect 4186 5138 4214 5222
rect 5329 5166 5334 5194
rect 5362 5166 10094 5194
rect 10122 5166 10127 5194
rect 10761 5166 10766 5194
rect 10794 5166 15022 5194
rect 15050 5166 15055 5194
rect 16809 5166 16814 5194
rect 16842 5166 20006 5194
rect 20034 5166 20039 5194
rect 21630 5138 21658 5222
rect 32144 5194 32200 5208
rect 21793 5166 21798 5194
rect 21826 5166 23198 5194
rect 23226 5166 23231 5194
rect 31089 5166 31094 5194
rect 31122 5166 32200 5194
rect 32144 5152 32200 5166
rect 4186 5110 11018 5138
rect 11321 5110 11326 5138
rect 11354 5110 12110 5138
rect 12138 5110 12143 5138
rect 12609 5110 12614 5138
rect 12642 5110 16842 5138
rect 16977 5110 16982 5138
rect 17010 5110 19334 5138
rect 19609 5110 19614 5138
rect 19642 5110 21518 5138
rect 21546 5110 21551 5138
rect 21630 5110 21854 5138
rect 23473 5110 23478 5138
rect 23506 5110 26614 5138
rect 26642 5110 26647 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 4545 5054 4550 5082
rect 4578 5054 6454 5082
rect 6482 5054 6487 5082
rect 9473 5054 9478 5082
rect 9506 5054 10430 5082
rect 10458 5054 10463 5082
rect 793 4998 798 5026
rect 826 4998 6678 5026
rect 6706 4998 6711 5026
rect 0 4970 56 4984
rect 10990 4970 11018 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 14345 5054 14350 5082
rect 14378 5054 15470 5082
rect 15498 5054 15503 5082
rect 15582 5054 16646 5082
rect 16674 5054 16679 5082
rect 15582 5026 15610 5054
rect 11769 4998 11774 5026
rect 11802 4998 13790 5026
rect 13818 4998 13823 5026
rect 13902 4998 15610 5026
rect 16814 5026 16842 5110
rect 19306 5082 19334 5110
rect 18438 5054 18494 5082
rect 18522 5054 18527 5082
rect 19306 5054 21462 5082
rect 21490 5054 21495 5082
rect 18438 5026 18466 5054
rect 21826 5026 21854 5110
rect 22227 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22369 5110
rect 23361 5054 23366 5082
rect 23394 5054 25550 5082
rect 25578 5054 25583 5082
rect 27706 5054 28238 5082
rect 28266 5054 28271 5082
rect 30753 5054 30758 5082
rect 30786 5054 31402 5082
rect 27706 5026 27734 5054
rect 16814 4998 18466 5026
rect 18545 4998 18550 5026
rect 18578 4998 20706 5026
rect 21826 4998 23982 5026
rect 24010 4998 24015 5026
rect 24089 4998 24094 5026
rect 24122 4998 27734 5026
rect 13902 4970 13930 4998
rect 20678 4970 20706 4998
rect 31374 4970 31402 5054
rect 32144 4970 32200 4984
rect 0 4942 9198 4970
rect 9226 4942 9231 4970
rect 10990 4942 13734 4970
rect 13762 4942 13767 4970
rect 13841 4942 13846 4970
rect 13874 4942 13930 4970
rect 14065 4942 14070 4970
rect 14098 4942 17710 4970
rect 17738 4942 17743 4970
rect 18041 4942 18046 4970
rect 18074 4942 20566 4970
rect 20594 4942 20599 4970
rect 20678 4942 28126 4970
rect 28154 4942 28159 4970
rect 28961 4942 28966 4970
rect 28994 4942 31262 4970
rect 31290 4942 31295 4970
rect 31374 4942 32200 4970
rect 0 4928 56 4942
rect 32144 4928 32200 4942
rect 5385 4886 5390 4914
rect 5418 4886 14238 4914
rect 14266 4886 14271 4914
rect 14681 4886 14686 4914
rect 14714 4886 29414 4914
rect 29442 4886 29447 4914
rect 29745 4886 29750 4914
rect 29778 4886 31486 4914
rect 31514 4886 31519 4914
rect 4153 4830 4158 4858
rect 4186 4830 5474 4858
rect 6785 4830 6790 4858
rect 6818 4830 14182 4858
rect 14210 4830 14215 4858
rect 16809 4830 16814 4858
rect 16842 4830 16847 4858
rect 16921 4830 16926 4858
rect 16954 4830 18550 4858
rect 18578 4830 18583 4858
rect 18657 4830 18662 4858
rect 18690 4830 19334 4858
rect 20169 4830 20174 4858
rect 20202 4830 23310 4858
rect 23338 4830 23343 4858
rect 28233 4830 28238 4858
rect 28266 4830 30198 4858
rect 30226 4830 30231 4858
rect 30641 4830 30646 4858
rect 30674 4830 31094 4858
rect 31122 4830 31127 4858
rect 5446 4802 5474 4830
rect 16814 4802 16842 4830
rect 2753 4774 2758 4802
rect 2786 4774 4214 4802
rect 5446 4774 6734 4802
rect 6762 4774 6767 4802
rect 7569 4774 7574 4802
rect 7602 4774 12698 4802
rect 0 4746 56 4760
rect 4186 4746 4214 4774
rect 12670 4746 12698 4774
rect 13426 4774 16702 4802
rect 16730 4774 16735 4802
rect 16814 4774 18802 4802
rect 13426 4746 13454 4774
rect 0 4718 1806 4746
rect 1834 4718 1839 4746
rect 4186 4718 10038 4746
rect 10066 4718 10071 4746
rect 12105 4718 12110 4746
rect 12138 4718 12446 4746
rect 12474 4718 12479 4746
rect 12670 4718 13454 4746
rect 13561 4718 13566 4746
rect 13594 4718 14182 4746
rect 14210 4718 14215 4746
rect 14905 4718 14910 4746
rect 14938 4718 16982 4746
rect 17010 4718 17015 4746
rect 17593 4718 17598 4746
rect 17626 4718 18606 4746
rect 18634 4718 18639 4746
rect 0 4704 56 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 18774 4690 18802 4774
rect 19306 4746 19334 4830
rect 19497 4774 19502 4802
rect 19530 4774 30142 4802
rect 30170 4774 30175 4802
rect 32144 4746 32200 4760
rect 19306 4718 20482 4746
rect 31425 4718 31430 4746
rect 31458 4718 32200 4746
rect 12161 4662 12166 4690
rect 12194 4662 17766 4690
rect 17794 4662 17799 4690
rect 18209 4662 18214 4690
rect 18242 4662 18606 4690
rect 18634 4662 18639 4690
rect 18774 4662 20174 4690
rect 20202 4662 20207 4690
rect 1185 4606 1190 4634
rect 1218 4606 2534 4634
rect 2562 4606 2567 4634
rect 9977 4606 9982 4634
rect 10010 4606 15190 4634
rect 15218 4606 15223 4634
rect 15302 4606 17542 4634
rect 17570 4606 17575 4634
rect 17649 4606 17654 4634
rect 17682 4606 20342 4634
rect 20370 4606 20375 4634
rect 15302 4578 15330 4606
rect 20454 4578 20482 4718
rect 21897 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22039 4718
rect 32144 4704 32200 4718
rect 29353 4662 29358 4690
rect 29386 4662 31878 4690
rect 31906 4662 31911 4690
rect 20561 4606 20566 4634
rect 20594 4606 26390 4634
rect 26418 4606 26423 4634
rect 30753 4606 30758 4634
rect 30786 4606 31318 4634
rect 31346 4606 31351 4634
rect 1633 4550 1638 4578
rect 1666 4550 10262 4578
rect 10290 4550 10295 4578
rect 10481 4550 10486 4578
rect 10514 4550 13454 4578
rect 13482 4550 13487 4578
rect 13617 4550 13622 4578
rect 13650 4550 15330 4578
rect 15857 4550 15862 4578
rect 15890 4550 19782 4578
rect 19810 4550 19815 4578
rect 20454 4550 28350 4578
rect 28378 4550 28383 4578
rect 0 4522 56 4536
rect 32144 4522 32200 4536
rect 0 4494 6622 4522
rect 6650 4494 6655 4522
rect 10369 4494 10374 4522
rect 10402 4494 12502 4522
rect 12530 4494 12535 4522
rect 12609 4494 12614 4522
rect 12642 4494 14686 4522
rect 14714 4494 14719 4522
rect 14793 4494 14798 4522
rect 14826 4494 15134 4522
rect 15162 4494 15167 4522
rect 15969 4494 15974 4522
rect 16002 4494 20370 4522
rect 20505 4494 20510 4522
rect 20538 4494 22974 4522
rect 23002 4494 23007 4522
rect 31369 4494 31374 4522
rect 31402 4494 32200 4522
rect 0 4480 56 4494
rect 20342 4466 20370 4494
rect 32144 4480 32200 4494
rect 1801 4438 1806 4466
rect 1834 4438 6510 4466
rect 6538 4438 6543 4466
rect 6673 4438 6678 4466
rect 6706 4438 10822 4466
rect 10850 4438 10855 4466
rect 10985 4438 10990 4466
rect 11018 4438 13398 4466
rect 13426 4438 13431 4466
rect 13729 4438 13734 4466
rect 13762 4438 20230 4466
rect 20258 4438 20263 4466
rect 20342 4438 24794 4466
rect 28233 4438 28238 4466
rect 28266 4438 30254 4466
rect 30282 4438 30287 4466
rect 4186 4382 15862 4410
rect 15890 4382 15895 4410
rect 15969 4382 15974 4410
rect 16002 4382 18158 4410
rect 18186 4382 18191 4410
rect 18377 4382 18382 4410
rect 18410 4382 18662 4410
rect 18690 4382 18695 4410
rect 20337 4382 20342 4410
rect 20370 4382 24262 4410
rect 24290 4382 24295 4410
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 0 4270 2114 4298
rect 0 4256 56 4270
rect 2086 4242 2114 4270
rect 4186 4242 4214 4382
rect 24766 4354 24794 4438
rect 26889 4382 26894 4410
rect 26922 4382 28742 4410
rect 28770 4382 28775 4410
rect 6841 4326 6846 4354
rect 6874 4326 10486 4354
rect 10514 4326 10519 4354
rect 10761 4326 10766 4354
rect 10794 4326 12110 4354
rect 12138 4326 12143 4354
rect 12441 4326 12446 4354
rect 12474 4326 14350 4354
rect 14378 4326 14383 4354
rect 15241 4326 15246 4354
rect 15274 4326 16198 4354
rect 16226 4326 16231 4354
rect 16865 4326 16870 4354
rect 16898 4326 21854 4354
rect 24766 4326 28574 4354
rect 28602 4326 28607 4354
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 6393 4270 6398 4298
rect 6426 4270 7574 4298
rect 7602 4270 7607 4298
rect 7737 4270 7742 4298
rect 7770 4270 10962 4298
rect 13449 4270 13454 4298
rect 13482 4270 15974 4298
rect 16002 4270 16007 4298
rect 18433 4270 18438 4298
rect 18466 4270 20622 4298
rect 20650 4270 20655 4298
rect 10934 4242 10962 4270
rect 21826 4242 21854 4326
rect 22227 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22369 4326
rect 32144 4298 32200 4312
rect 22633 4270 22638 4298
rect 22666 4270 24318 4298
rect 24346 4270 24351 4298
rect 25153 4270 25158 4298
rect 25186 4270 27958 4298
rect 27986 4270 27991 4298
rect 31425 4270 31430 4298
rect 31458 4270 32200 4298
rect 32144 4256 32200 4270
rect 2086 4214 4214 4242
rect 7518 4214 7574 4242
rect 7602 4214 7607 4242
rect 8913 4214 8918 4242
rect 8946 4214 10906 4242
rect 10934 4214 14014 4242
rect 14042 4214 14047 4242
rect 15073 4214 15078 4242
rect 15106 4214 18466 4242
rect 18545 4214 18550 4242
rect 18578 4214 20678 4242
rect 20706 4214 20711 4242
rect 21826 4214 28630 4242
rect 28658 4214 28663 4242
rect 7518 4130 7546 4214
rect 10878 4186 10906 4214
rect 18438 4186 18466 4214
rect 7625 4158 7630 4186
rect 7658 4158 9982 4186
rect 10010 4158 10015 4186
rect 10878 4158 12446 4186
rect 12474 4158 12479 4186
rect 12553 4158 12558 4186
rect 12586 4158 13538 4186
rect 14345 4158 14350 4186
rect 14378 4158 16870 4186
rect 16898 4158 16903 4186
rect 17481 4158 17486 4186
rect 17514 4158 17822 4186
rect 17850 4158 17855 4186
rect 18438 4158 28910 4186
rect 28938 4158 28943 4186
rect 30529 4158 30534 4186
rect 30562 4158 31542 4186
rect 31570 4158 31575 4186
rect 13510 4130 13538 4158
rect 2641 4102 2646 4130
rect 2674 4102 7546 4130
rect 8969 4102 8974 4130
rect 9002 4102 9870 4130
rect 9898 4102 9903 4130
rect 10033 4102 10038 4130
rect 10066 4102 12558 4130
rect 12586 4102 12591 4130
rect 13379 4102 13398 4130
rect 13426 4102 13431 4130
rect 13510 4102 15078 4130
rect 15106 4102 15111 4130
rect 16366 4102 27958 4130
rect 27986 4102 27991 4130
rect 29857 4102 29862 4130
rect 29890 4102 31822 4130
rect 31850 4102 31855 4130
rect 0 4074 56 4088
rect 16366 4074 16394 4102
rect 32144 4074 32200 4088
rect 0 4046 6174 4074
rect 6202 4046 6207 4074
rect 7681 4046 7686 4074
rect 7714 4046 8246 4074
rect 8274 4046 8279 4074
rect 10481 4046 10486 4074
rect 10514 4046 16394 4074
rect 17481 4046 17486 4074
rect 17514 4046 20286 4074
rect 20314 4046 20319 4074
rect 21737 4046 21742 4074
rect 21770 4046 28854 4074
rect 28882 4046 28887 4074
rect 31537 4046 31542 4074
rect 31570 4046 32200 4074
rect 0 4032 56 4046
rect 32144 4032 32200 4046
rect 6617 3990 6622 4018
rect 6650 3990 12502 4018
rect 12530 3990 12535 4018
rect 12609 3990 12614 4018
rect 12642 3990 13958 4018
rect 13986 3990 13991 4018
rect 14233 3990 14238 4018
rect 14266 3990 17598 4018
rect 17626 3990 17631 4018
rect 17817 3990 17822 4018
rect 17850 3990 20958 4018
rect 20986 3990 20991 4018
rect 21961 3990 21966 4018
rect 21994 3990 23422 4018
rect 23450 3990 23455 4018
rect 6281 3934 6286 3962
rect 6314 3934 10486 3962
rect 10514 3934 10519 3962
rect 12105 3934 12110 3962
rect 12138 3934 12782 3962
rect 12810 3934 12815 3962
rect 13449 3934 13454 3962
rect 13482 3934 20174 3962
rect 20202 3934 20207 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 21897 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22039 3934
rect 6729 3878 6734 3906
rect 6762 3878 9086 3906
rect 9114 3878 9119 3906
rect 10425 3878 10430 3906
rect 10458 3878 11774 3906
rect 11802 3878 11807 3906
rect 12110 3878 14126 3906
rect 14154 3878 14159 3906
rect 15073 3878 15078 3906
rect 15106 3878 17654 3906
rect 17682 3878 17687 3906
rect 17761 3878 17766 3906
rect 17794 3878 20846 3906
rect 20874 3878 20879 3906
rect 0 3850 56 3864
rect 12110 3850 12138 3878
rect 32144 3850 32200 3864
rect 0 3822 10374 3850
rect 10402 3822 10407 3850
rect 10817 3822 10822 3850
rect 10850 3822 12138 3850
rect 12217 3822 12222 3850
rect 12250 3822 12558 3850
rect 12586 3822 12591 3850
rect 13449 3822 13454 3850
rect 13482 3822 13487 3850
rect 13561 3822 13566 3850
rect 13594 3822 14910 3850
rect 14938 3822 14943 3850
rect 15017 3822 15022 3850
rect 15050 3822 18438 3850
rect 18466 3822 18471 3850
rect 19553 3822 19558 3850
rect 19586 3822 28910 3850
rect 28938 3822 28943 3850
rect 31425 3822 31430 3850
rect 31458 3822 32200 3850
rect 0 3808 56 3822
rect 13454 3794 13482 3822
rect 32144 3808 32200 3822
rect 1521 3766 1526 3794
rect 1554 3766 7154 3794
rect 7401 3766 7406 3794
rect 7434 3766 9030 3794
rect 9058 3766 9063 3794
rect 12777 3766 12782 3794
rect 12810 3766 13482 3794
rect 13510 3766 14406 3794
rect 14434 3766 14439 3794
rect 14513 3766 14518 3794
rect 14546 3766 15582 3794
rect 15610 3766 15615 3794
rect 17705 3766 17710 3794
rect 17738 3766 18998 3794
rect 19026 3766 19031 3794
rect 20001 3766 20006 3794
rect 20034 3766 23478 3794
rect 23506 3766 23511 3794
rect 7126 3738 7154 3766
rect 13510 3738 13538 3766
rect 1862 3710 6678 3738
rect 6706 3710 6711 3738
rect 7126 3710 7686 3738
rect 7714 3710 7719 3738
rect 9977 3710 9982 3738
rect 10010 3710 12110 3738
rect 12138 3710 12143 3738
rect 12553 3710 12558 3738
rect 12586 3710 13538 3738
rect 13617 3710 13622 3738
rect 13650 3710 14854 3738
rect 14882 3710 14887 3738
rect 14961 3710 14966 3738
rect 14994 3710 17430 3738
rect 17458 3710 17463 3738
rect 17537 3710 17542 3738
rect 17570 3710 20062 3738
rect 20090 3710 20095 3738
rect 20617 3710 20622 3738
rect 20650 3710 30254 3738
rect 30282 3710 30287 3738
rect 0 3626 56 3640
rect 1862 3626 1890 3710
rect 4041 3654 4046 3682
rect 4074 3654 17710 3682
rect 17738 3654 17743 3682
rect 18545 3654 18550 3682
rect 18578 3654 29190 3682
rect 29218 3654 29223 3682
rect 32144 3626 32200 3640
rect 0 3598 1890 3626
rect 4186 3598 29414 3626
rect 29442 3598 29447 3626
rect 31425 3598 31430 3626
rect 31458 3598 32200 3626
rect 0 3584 56 3598
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 4186 3458 4214 3598
rect 32144 3584 32200 3598
rect 5777 3542 5782 3570
rect 5810 3542 10038 3570
rect 10066 3542 10071 3570
rect 10929 3542 10934 3570
rect 10962 3542 12110 3570
rect 12138 3542 12143 3570
rect 12441 3542 12446 3570
rect 12474 3542 19334 3570
rect 19362 3542 19367 3570
rect 29521 3542 29526 3570
rect 29554 3542 30590 3570
rect 30618 3542 30623 3570
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 22227 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22369 3542
rect 121 3430 126 3458
rect 154 3430 4214 3458
rect 7126 3486 10486 3514
rect 10514 3486 10519 3514
rect 13561 3486 13566 3514
rect 13594 3486 14854 3514
rect 14882 3486 14887 3514
rect 14961 3486 14966 3514
rect 14994 3486 16058 3514
rect 16809 3486 16814 3514
rect 16842 3486 21854 3514
rect 28625 3486 28630 3514
rect 28658 3486 31094 3514
rect 31122 3486 31127 3514
rect 0 3402 56 3416
rect 7126 3402 7154 3486
rect 16030 3458 16058 3486
rect 21826 3458 21854 3486
rect 7345 3430 7350 3458
rect 7378 3430 8694 3458
rect 8722 3430 8727 3458
rect 8806 3430 10430 3458
rect 10458 3430 10463 3458
rect 13449 3430 13454 3458
rect 13482 3430 15918 3458
rect 15946 3430 15951 3458
rect 16030 3430 16814 3458
rect 16842 3430 16847 3458
rect 18041 3430 18046 3458
rect 18074 3430 20118 3458
rect 20146 3430 20151 3458
rect 21826 3430 30254 3458
rect 30282 3430 30287 3458
rect 8806 3402 8834 3430
rect 32144 3402 32200 3416
rect 0 3374 7154 3402
rect 8353 3374 8358 3402
rect 8386 3374 8834 3402
rect 9193 3374 9198 3402
rect 9226 3374 10094 3402
rect 11097 3374 11102 3402
rect 11130 3374 13454 3402
rect 13482 3374 13487 3402
rect 13673 3374 13678 3402
rect 13706 3374 15134 3402
rect 15162 3374 15167 3402
rect 15246 3374 18886 3402
rect 18914 3374 18919 3402
rect 18993 3374 18998 3402
rect 19026 3374 21742 3402
rect 21770 3374 21775 3402
rect 23361 3374 23366 3402
rect 23394 3374 25158 3402
rect 25186 3374 25191 3402
rect 28742 3374 29806 3402
rect 29834 3374 29839 3402
rect 30753 3374 30758 3402
rect 30786 3374 32200 3402
rect 0 3360 56 3374
rect 10066 3346 10094 3374
rect 15246 3346 15274 3374
rect 28742 3346 28770 3374
rect 32144 3360 32200 3374
rect 1297 3318 1302 3346
rect 1330 3318 7070 3346
rect 7098 3318 7103 3346
rect 8297 3318 8302 3346
rect 8330 3318 8750 3346
rect 8778 3318 8783 3346
rect 10066 3318 12558 3346
rect 12586 3318 12591 3346
rect 12833 3318 12838 3346
rect 12866 3318 13454 3346
rect 13482 3318 13487 3346
rect 13729 3318 13734 3346
rect 13762 3318 15274 3346
rect 18601 3318 18606 3346
rect 18634 3318 23534 3346
rect 23562 3318 23567 3346
rect 25489 3318 25494 3346
rect 25522 3318 28770 3346
rect 29969 3318 29974 3346
rect 30002 3318 30982 3346
rect 31010 3318 31015 3346
rect 1017 3262 1022 3290
rect 1050 3262 7462 3290
rect 7490 3262 7495 3290
rect 10089 3262 10094 3290
rect 10122 3262 12446 3290
rect 12474 3262 12479 3290
rect 12670 3262 18158 3290
rect 18186 3262 18191 3290
rect 20113 3262 20118 3290
rect 20146 3262 22638 3290
rect 22666 3262 22671 3290
rect 24313 3262 24318 3290
rect 24346 3262 30142 3290
rect 30170 3262 30175 3290
rect 1806 3206 4214 3234
rect 5721 3206 5726 3234
rect 5754 3206 7406 3234
rect 7434 3206 7439 3234
rect 7513 3206 7518 3234
rect 7546 3206 12558 3234
rect 12586 3206 12591 3234
rect 0 3178 56 3192
rect 1806 3178 1834 3206
rect 0 3150 1834 3178
rect 4186 3178 4214 3206
rect 12670 3178 12698 3262
rect 12777 3206 12782 3234
rect 12810 3206 14798 3234
rect 14826 3206 14831 3234
rect 17369 3206 17374 3234
rect 17402 3206 29246 3234
rect 29274 3206 29279 3234
rect 32144 3178 32200 3192
rect 4186 3150 8638 3178
rect 8666 3150 8671 3178
rect 8857 3150 8862 3178
rect 8890 3150 11830 3178
rect 11858 3150 11863 3178
rect 12105 3150 12110 3178
rect 12138 3150 12698 3178
rect 13785 3150 13790 3178
rect 13818 3150 20454 3178
rect 20482 3150 20487 3178
rect 24766 3150 29694 3178
rect 29722 3150 29727 3178
rect 31537 3150 31542 3178
rect 31570 3150 32200 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 21897 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22039 3150
rect 7065 3094 7070 3122
rect 7098 3094 9702 3122
rect 9730 3094 9735 3122
rect 12110 3094 12838 3122
rect 12866 3094 12871 3122
rect 13729 3094 13734 3122
rect 13762 3094 16310 3122
rect 16338 3094 16343 3122
rect 12110 3066 12138 3094
rect 24766 3066 24794 3150
rect 32144 3136 32200 3150
rect 8465 3038 8470 3066
rect 8498 3038 10654 3066
rect 10682 3038 10687 3066
rect 11769 3038 11774 3066
rect 11802 3038 12138 3066
rect 12497 3038 12502 3066
rect 12530 3038 24794 3066
rect 24822 3094 27734 3122
rect 27762 3094 27767 3122
rect 28961 3094 28966 3122
rect 28994 3094 30310 3122
rect 30338 3094 30343 3122
rect 2921 2982 2926 3010
rect 2954 2982 4046 3010
rect 4074 2982 4079 3010
rect 4186 2982 6230 3010
rect 6258 2982 6263 3010
rect 7546 2982 10766 3010
rect 10794 2982 10799 3010
rect 10873 2982 10878 3010
rect 10906 2982 13286 3010
rect 13314 2982 13319 3010
rect 13449 2982 13454 3010
rect 13482 2982 14014 3010
rect 14042 2982 14047 3010
rect 15913 2982 15918 3010
rect 15946 2982 23702 3010
rect 23730 2982 23735 3010
rect 0 2954 56 2968
rect 4186 2954 4214 2982
rect 0 2926 4214 2954
rect 4321 2926 4326 2954
rect 4354 2926 6398 2954
rect 6426 2926 6431 2954
rect 0 2912 56 2926
rect 7546 2898 7574 2982
rect 24822 2954 24850 3094
rect 25433 3038 25438 3066
rect 25466 3038 28686 3066
rect 28714 3038 28719 3066
rect 30753 3038 30758 3066
rect 30786 3038 32102 3066
rect 32130 3038 32135 3066
rect 29633 2982 29638 3010
rect 29666 2982 30870 3010
rect 30898 2982 30903 3010
rect 32144 2954 32200 2968
rect 8073 2926 8078 2954
rect 8106 2926 10934 2954
rect 10962 2926 10967 2954
rect 11489 2926 11494 2954
rect 11522 2926 13734 2954
rect 13762 2926 13767 2954
rect 14289 2926 14294 2954
rect 14322 2926 18214 2954
rect 18242 2926 18247 2954
rect 19777 2926 19782 2954
rect 19810 2926 24850 2954
rect 30641 2926 30646 2954
rect 30674 2926 32200 2954
rect 32144 2912 32200 2926
rect 1017 2870 1022 2898
rect 1050 2870 2590 2898
rect 2618 2870 2623 2898
rect 5889 2870 5894 2898
rect 5922 2870 7574 2898
rect 10425 2870 10430 2898
rect 10458 2870 13398 2898
rect 13426 2870 13431 2898
rect 15073 2870 15078 2898
rect 15106 2870 21406 2898
rect 21434 2870 21439 2898
rect 21826 2870 22078 2898
rect 22106 2870 22111 2898
rect 22353 2870 22358 2898
rect 22386 2870 24374 2898
rect 24402 2870 24407 2898
rect 21826 2842 21854 2870
rect 1241 2814 1246 2842
rect 1274 2814 4214 2842
rect 6001 2814 6006 2842
rect 6034 2814 7854 2842
rect 7882 2814 7887 2842
rect 10486 2814 17542 2842
rect 17570 2814 17575 2842
rect 17985 2814 17990 2842
rect 18018 2814 21854 2842
rect 21966 2814 22806 2842
rect 22834 2814 22839 2842
rect 24257 2814 24262 2842
rect 24290 2814 28686 2842
rect 28714 2814 28719 2842
rect 4186 2786 4214 2814
rect 10486 2786 10514 2814
rect 21966 2786 21994 2814
rect 4186 2758 10514 2786
rect 12721 2758 12726 2786
rect 12754 2758 14574 2786
rect 14602 2758 14607 2786
rect 16361 2758 16366 2786
rect 16394 2758 21994 2786
rect 22409 2758 22414 2786
rect 22442 2758 25326 2786
rect 25354 2758 25359 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 22227 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22369 2758
rect 32144 2730 32200 2744
rect 0 2702 2114 2730
rect 7121 2702 7126 2730
rect 7154 2702 12110 2730
rect 12138 2702 12143 2730
rect 12665 2702 12670 2730
rect 12698 2702 20902 2730
rect 20930 2702 20935 2730
rect 22582 2702 26950 2730
rect 26978 2702 26983 2730
rect 28625 2702 28630 2730
rect 28658 2702 30142 2730
rect 30170 2702 30175 2730
rect 31313 2702 31318 2730
rect 31346 2702 32200 2730
rect 0 2688 56 2702
rect 2086 2674 2114 2702
rect 2086 2646 6510 2674
rect 6538 2646 6543 2674
rect 8633 2646 8638 2674
rect 8666 2646 10822 2674
rect 10850 2646 10855 2674
rect 10929 2646 10934 2674
rect 10962 2646 13678 2674
rect 13706 2646 13711 2674
rect 14233 2646 14238 2674
rect 14266 2646 19502 2674
rect 19530 2646 19535 2674
rect 21177 2646 21182 2674
rect 21210 2646 22470 2674
rect 22498 2646 22503 2674
rect 22582 2618 22610 2702
rect 32144 2688 32200 2702
rect 24201 2646 24206 2674
rect 24234 2646 29694 2674
rect 29722 2646 29727 2674
rect 30422 2646 31094 2674
rect 31122 2646 31127 2674
rect 30422 2618 30450 2646
rect 3257 2590 3262 2618
rect 3290 2590 9366 2618
rect 9394 2590 9399 2618
rect 9641 2590 9646 2618
rect 9674 2590 15806 2618
rect 15834 2590 15839 2618
rect 16361 2590 16366 2618
rect 16394 2590 22610 2618
rect 22750 2590 24318 2618
rect 24346 2590 24351 2618
rect 29185 2590 29190 2618
rect 29218 2590 30450 2618
rect 30529 2590 30534 2618
rect 30562 2590 31262 2618
rect 31290 2590 31295 2618
rect 9137 2534 9142 2562
rect 9170 2534 12502 2562
rect 12530 2534 12535 2562
rect 12614 2534 13230 2562
rect 13258 2534 13263 2562
rect 13393 2534 13398 2562
rect 13426 2534 13846 2562
rect 13874 2534 13879 2562
rect 17654 2534 20230 2562
rect 20258 2534 20263 2562
rect 20337 2534 20342 2562
rect 20370 2534 22414 2562
rect 22442 2534 22447 2562
rect 0 2506 56 2520
rect 12614 2506 12642 2534
rect 17654 2506 17682 2534
rect 22750 2506 22778 2590
rect 25209 2534 25214 2562
rect 25242 2534 25326 2562
rect 25354 2534 25359 2562
rect 29969 2534 29974 2562
rect 30002 2534 30926 2562
rect 30954 2534 30959 2562
rect 32144 2506 32200 2520
rect 0 2478 7126 2506
rect 7154 2478 7159 2506
rect 8745 2478 8750 2506
rect 8778 2478 12642 2506
rect 13505 2478 13510 2506
rect 13538 2478 15246 2506
rect 15274 2478 15279 2506
rect 15409 2478 15414 2506
rect 15442 2478 17682 2506
rect 17710 2478 18382 2506
rect 18410 2478 18415 2506
rect 21826 2478 22778 2506
rect 23473 2478 23478 2506
rect 23506 2478 24934 2506
rect 24962 2478 24967 2506
rect 26665 2478 26670 2506
rect 26698 2478 28294 2506
rect 28322 2478 28327 2506
rect 31537 2478 31542 2506
rect 31570 2478 32200 2506
rect 0 2464 56 2478
rect 17710 2450 17738 2478
rect 21826 2450 21854 2478
rect 32144 2464 32200 2478
rect 3761 2422 3766 2450
rect 3794 2422 8414 2450
rect 8442 2422 8447 2450
rect 10486 2422 13342 2450
rect 13370 2422 13375 2450
rect 13449 2422 13454 2450
rect 13482 2422 17738 2450
rect 18265 2422 18270 2450
rect 18298 2422 21854 2450
rect 22465 2422 22470 2450
rect 22498 2422 26446 2450
rect 26474 2422 26479 2450
rect 27169 2422 27174 2450
rect 27202 2422 29078 2450
rect 29106 2422 29111 2450
rect 10486 2394 10514 2422
rect 7401 2366 7406 2394
rect 7434 2366 10514 2394
rect 13449 2366 13454 2394
rect 13482 2366 16366 2394
rect 16394 2366 16399 2394
rect 24369 2366 24374 2394
rect 24402 2366 27566 2394
rect 27594 2366 27599 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 21897 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22039 2366
rect 5441 2310 5446 2338
rect 5474 2310 8414 2338
rect 8442 2310 8447 2338
rect 12105 2310 12110 2338
rect 12138 2310 13174 2338
rect 13202 2310 13207 2338
rect 16473 2310 16478 2338
rect 16506 2310 21462 2338
rect 21490 2310 21495 2338
rect 23977 2310 23982 2338
rect 24010 2310 29414 2338
rect 29442 2310 29447 2338
rect 0 2282 56 2296
rect 32144 2282 32200 2296
rect 0 2254 6706 2282
rect 11209 2254 11214 2282
rect 11242 2254 12670 2282
rect 12698 2254 12703 2282
rect 17817 2254 17822 2282
rect 17850 2254 19614 2282
rect 19642 2254 19647 2282
rect 20393 2254 20398 2282
rect 20426 2254 24766 2282
rect 24794 2254 24799 2282
rect 31257 2254 31262 2282
rect 31290 2254 32200 2282
rect 0 2240 56 2254
rect 6678 2226 6706 2254
rect 32144 2240 32200 2254
rect 905 2198 910 2226
rect 938 2198 6342 2226
rect 6370 2198 6375 2226
rect 6678 2198 15134 2226
rect 15162 2198 15167 2226
rect 19329 2198 19334 2226
rect 19362 2198 26054 2226
rect 26082 2198 26087 2226
rect 27841 2198 27846 2226
rect 27874 2198 30366 2226
rect 30394 2198 30399 2226
rect 10033 2142 10038 2170
rect 10066 2142 18438 2170
rect 18466 2142 18471 2170
rect 21289 2142 21294 2170
rect 21322 2142 22582 2170
rect 22610 2142 22615 2170
rect 1078 2086 2590 2114
rect 2618 2086 2623 2114
rect 6673 2086 6678 2114
rect 6706 2086 12558 2114
rect 12586 2086 12591 2114
rect 12665 2086 12670 2114
rect 12698 2086 24262 2114
rect 24290 2086 24295 2114
rect 0 2058 56 2072
rect 1078 2058 1106 2086
rect 32144 2058 32200 2072
rect 0 2030 1106 2058
rect 1185 2030 1190 2058
rect 1218 2030 8358 2058
rect 8386 2030 8391 2058
rect 11886 2030 13454 2058
rect 13482 2030 13487 2058
rect 14625 2030 14630 2058
rect 14658 2030 23254 2058
rect 23282 2030 23287 2058
rect 28065 2030 28070 2058
rect 28098 2030 30534 2058
rect 30562 2030 30567 2058
rect 31425 2030 31430 2058
rect 31458 2030 32200 2058
rect 0 2016 56 2030
rect 6449 1974 6454 2002
rect 6482 1974 11774 2002
rect 11802 1974 11807 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 11886 1946 11914 2030
rect 32144 2016 32200 2030
rect 12497 1974 12502 2002
rect 12530 1974 17542 2002
rect 17570 1974 17575 2002
rect 19306 1974 20734 2002
rect 20762 1974 20767 2002
rect 22577 1974 22582 2002
rect 22610 1974 23814 2002
rect 23842 1974 23847 2002
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 2865 1918 2870 1946
rect 2898 1918 11914 1946
rect 12441 1918 12446 1946
rect 12474 1918 13678 1946
rect 13706 1918 13711 1946
rect 15946 1918 16702 1946
rect 16730 1918 16735 1946
rect 16809 1918 16814 1946
rect 16842 1918 18046 1946
rect 18074 1918 18079 1946
rect 6505 1862 6510 1890
rect 6538 1862 10262 1890
rect 10290 1862 10295 1890
rect 10369 1862 10374 1890
rect 10402 1862 13398 1890
rect 13426 1862 13431 1890
rect 0 1834 56 1848
rect 15946 1834 15974 1918
rect 19306 1890 19334 1974
rect 22227 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22369 1974
rect 0 1806 6846 1834
rect 6874 1806 6879 1834
rect 9025 1806 9030 1834
rect 9058 1806 12446 1834
rect 12474 1806 12479 1834
rect 13113 1806 13118 1834
rect 13146 1806 15974 1834
rect 16366 1862 19334 1890
rect 19441 1862 19446 1890
rect 19474 1862 24990 1890
rect 25018 1862 25023 1890
rect 0 1792 56 1806
rect 16366 1778 16394 1862
rect 32144 1834 32200 1848
rect 16697 1806 16702 1834
rect 16730 1806 22190 1834
rect 22218 1806 22223 1834
rect 22633 1806 22638 1834
rect 22666 1806 23646 1834
rect 23674 1806 23679 1834
rect 24313 1806 24318 1834
rect 24346 1806 29834 1834
rect 30641 1806 30646 1834
rect 30674 1806 32200 1834
rect 29806 1778 29834 1806
rect 32144 1792 32200 1806
rect 1297 1750 1302 1778
rect 1330 1750 16394 1778
rect 17649 1750 17654 1778
rect 17682 1750 21014 1778
rect 21042 1750 21047 1778
rect 21233 1750 21238 1778
rect 21266 1750 29694 1778
rect 29722 1750 29727 1778
rect 29806 1750 30926 1778
rect 30954 1750 30959 1778
rect 7121 1694 7126 1722
rect 7154 1694 10878 1722
rect 10906 1694 10911 1722
rect 11718 1694 14322 1722
rect 16809 1694 16814 1722
rect 16842 1694 16847 1722
rect 17313 1694 17318 1722
rect 17346 1694 18494 1722
rect 18522 1694 18527 1722
rect 20169 1694 20174 1722
rect 20202 1694 29918 1722
rect 29946 1694 29951 1722
rect 30641 1694 30646 1722
rect 30674 1694 31318 1722
rect 31346 1694 31351 1722
rect 1806 1638 6622 1666
rect 6650 1638 6655 1666
rect 0 1610 56 1624
rect 1806 1610 1834 1638
rect 11718 1610 11746 1694
rect 14294 1666 14322 1694
rect 16814 1666 16842 1694
rect 11825 1638 11830 1666
rect 11858 1638 13622 1666
rect 13650 1638 13655 1666
rect 14294 1638 16842 1666
rect 17929 1638 17934 1666
rect 17962 1638 19222 1666
rect 19250 1638 19255 1666
rect 20225 1638 20230 1666
rect 20258 1638 25606 1666
rect 25634 1638 25639 1666
rect 26049 1638 26054 1666
rect 26082 1638 28910 1666
rect 28938 1638 28943 1666
rect 32144 1610 32200 1624
rect 0 1582 1834 1610
rect 4209 1582 4214 1610
rect 4242 1582 7798 1610
rect 7826 1582 7831 1610
rect 10066 1582 11746 1610
rect 16361 1582 16366 1610
rect 16394 1582 17878 1610
rect 17906 1582 17911 1610
rect 18209 1582 18214 1610
rect 18242 1582 21518 1610
rect 21546 1582 21551 1610
rect 22129 1582 22134 1610
rect 22162 1582 23366 1610
rect 23394 1582 23399 1610
rect 25433 1582 25438 1610
rect 25466 1582 27174 1610
rect 27202 1582 27207 1610
rect 31537 1582 31542 1610
rect 31570 1582 32200 1610
rect 0 1568 56 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 10066 1554 10094 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 21897 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22039 1582
rect 32144 1568 32200 1582
rect 5945 1526 5950 1554
rect 5978 1526 6286 1554
rect 6314 1526 6319 1554
rect 6561 1526 6566 1554
rect 6594 1526 10094 1554
rect 13561 1526 13566 1554
rect 13594 1526 15190 1554
rect 15218 1526 15223 1554
rect 15577 1526 15582 1554
rect 15610 1526 18914 1554
rect 22073 1526 22078 1554
rect 22106 1526 24038 1554
rect 24066 1526 24071 1554
rect 26049 1526 26054 1554
rect 26082 1526 29526 1554
rect 29554 1526 29559 1554
rect 18886 1498 18914 1526
rect 4825 1470 4830 1498
rect 4858 1470 9030 1498
rect 9058 1470 9063 1498
rect 10066 1470 14462 1498
rect 14490 1470 14495 1498
rect 14569 1470 14574 1498
rect 14602 1470 18578 1498
rect 18886 1470 22694 1498
rect 22722 1470 22727 1498
rect 24313 1470 24318 1498
rect 24346 1470 26670 1498
rect 26698 1470 26703 1498
rect 10066 1442 10094 1470
rect 961 1414 966 1442
rect 994 1414 6006 1442
rect 6034 1414 6039 1442
rect 8689 1414 8694 1442
rect 8722 1414 10094 1442
rect 10257 1414 10262 1442
rect 10290 1414 17318 1442
rect 17346 1414 17351 1442
rect 0 1386 56 1400
rect 0 1358 6118 1386
rect 6146 1358 6151 1386
rect 10649 1358 10654 1386
rect 10682 1358 13510 1386
rect 13538 1358 13543 1386
rect 0 1344 56 1358
rect 18550 1330 18578 1470
rect 20897 1414 20902 1442
rect 20930 1414 22638 1442
rect 22666 1414 22671 1442
rect 23417 1414 23422 1442
rect 23450 1414 26222 1442
rect 26250 1414 26255 1442
rect 29241 1414 29246 1442
rect 29274 1414 30254 1442
rect 30282 1414 30287 1442
rect 32144 1386 32200 1400
rect 19721 1358 19726 1386
rect 19754 1358 22526 1386
rect 22554 1358 22559 1386
rect 29633 1358 29638 1386
rect 29666 1358 31094 1386
rect 31122 1358 31127 1386
rect 31313 1358 31318 1386
rect 31346 1358 32200 1386
rect 32144 1344 32200 1358
rect 5945 1302 5950 1330
rect 5978 1302 14742 1330
rect 14770 1302 14775 1330
rect 18550 1302 21070 1330
rect 21098 1302 21103 1330
rect 21345 1302 21350 1330
rect 21378 1302 23870 1330
rect 23898 1302 23903 1330
rect 29185 1302 29190 1330
rect 29218 1302 30086 1330
rect 30114 1302 30119 1330
rect 30641 1302 30646 1330
rect 30674 1302 31374 1330
rect 31402 1302 31407 1330
rect 10873 1246 10878 1274
rect 10906 1246 29414 1274
rect 29442 1246 29447 1274
rect 7681 1190 7686 1218
rect 7714 1190 12194 1218
rect 12446 1190 15078 1218
rect 15106 1190 15111 1218
rect 15689 1190 15694 1218
rect 15722 1190 19446 1218
rect 19474 1190 19479 1218
rect 20785 1190 20790 1218
rect 20818 1190 22162 1218
rect 23529 1190 23534 1218
rect 23562 1190 29694 1218
rect 29722 1190 29727 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 0 1134 2114 1162
rect 0 1120 56 1134
rect 2086 1106 2114 1134
rect 2422 1134 11830 1162
rect 11858 1134 11863 1162
rect 2422 1106 2450 1134
rect 12166 1106 12194 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 12446 1106 12474 1190
rect 14177 1134 14182 1162
rect 14210 1134 17654 1162
rect 17682 1134 17687 1162
rect 17873 1134 17878 1162
rect 17906 1134 20762 1162
rect 2086 1078 2450 1106
rect 6281 1078 6286 1106
rect 6314 1078 7490 1106
rect 7625 1078 7630 1106
rect 7658 1078 9870 1106
rect 9898 1078 9903 1106
rect 12166 1078 12474 1106
rect 13617 1078 13622 1106
rect 13650 1078 18158 1106
rect 18186 1078 18191 1106
rect 18433 1078 18438 1106
rect 18466 1078 18942 1106
rect 18970 1078 18975 1106
rect 7462 1050 7490 1078
rect 20734 1050 20762 1134
rect 22134 1106 22162 1190
rect 22227 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22369 1190
rect 32144 1162 32200 1176
rect 22414 1134 26054 1162
rect 26082 1134 26087 1162
rect 29409 1134 29414 1162
rect 29442 1134 31150 1162
rect 31178 1134 31183 1162
rect 31425 1134 31430 1162
rect 31458 1134 32200 1162
rect 22414 1106 22442 1134
rect 32144 1120 32200 1134
rect 21793 1078 21798 1106
rect 21826 1078 22022 1106
rect 22050 1078 22055 1106
rect 22134 1078 22442 1106
rect 22913 1078 22918 1106
rect 22946 1078 24486 1106
rect 24514 1078 24519 1106
rect 3817 1022 3822 1050
rect 3850 1022 7350 1050
rect 7378 1022 7383 1050
rect 7462 1022 8190 1050
rect 8218 1022 8223 1050
rect 12833 1022 12838 1050
rect 12866 1022 18774 1050
rect 18802 1022 18807 1050
rect 18881 1022 18886 1050
rect 18914 1022 20622 1050
rect 20650 1022 20655 1050
rect 20734 1022 22134 1050
rect 22162 1022 22167 1050
rect 22302 1022 22750 1050
rect 22778 1022 22783 1050
rect 24873 1022 24878 1050
rect 24906 1022 28014 1050
rect 28042 1022 28047 1050
rect 28793 1022 28798 1050
rect 28826 1022 30142 1050
rect 30170 1022 30175 1050
rect 22302 994 22330 1022
rect 1241 966 1246 994
rect 1274 966 7574 994
rect 7602 966 7607 994
rect 12553 966 12558 994
rect 12586 966 15358 994
rect 15386 966 15391 994
rect 19049 966 19054 994
rect 19082 966 22330 994
rect 22633 966 22638 994
rect 22666 966 24598 994
rect 24626 966 24631 994
rect 26889 966 26894 994
rect 26922 966 28574 994
rect 28602 966 28607 994
rect 29969 966 29974 994
rect 30002 966 30926 994
rect 30954 966 30959 994
rect 0 938 56 952
rect 32144 938 32200 952
rect 0 910 4550 938
rect 4578 910 4583 938
rect 6673 910 6678 938
rect 6706 910 11158 938
rect 11186 910 11191 938
rect 11998 910 16198 938
rect 16226 910 16231 938
rect 16753 910 16758 938
rect 16786 910 17990 938
rect 18018 910 18023 938
rect 18433 910 18438 938
rect 18466 910 20202 938
rect 20281 910 20286 938
rect 20314 910 22834 938
rect 23473 910 23478 938
rect 23506 910 28966 938
rect 28994 910 28999 938
rect 31537 910 31542 938
rect 31570 910 32200 938
rect 0 896 56 910
rect 11998 882 12026 910
rect 20174 882 20202 910
rect 1694 854 4214 882
rect 5273 854 5278 882
rect 5306 854 7686 882
rect 7714 854 7719 882
rect 8185 854 8190 882
rect 8218 854 12026 882
rect 14294 854 15246 882
rect 15274 854 15279 882
rect 15353 854 15358 882
rect 15386 854 20146 882
rect 20174 854 22722 882
rect 1694 826 1722 854
rect 1465 798 1470 826
rect 1498 798 1722 826
rect 4186 826 4214 854
rect 14294 826 14322 854
rect 20118 826 20146 854
rect 22694 826 22722 854
rect 22806 826 22834 910
rect 32144 896 32200 910
rect 26273 854 26278 882
rect 26306 854 29134 882
rect 29162 854 29167 882
rect 30641 854 30646 882
rect 30674 854 31290 882
rect 4186 798 7126 826
rect 7154 798 7159 826
rect 12110 798 14322 826
rect 15465 798 15470 826
rect 15498 798 17598 826
rect 17626 798 17631 826
rect 20118 798 21854 826
rect 22689 798 22694 826
rect 22722 798 22727 826
rect 22806 798 24206 826
rect 24234 798 24239 826
rect 26945 798 26950 826
rect 26978 798 31038 826
rect 31066 798 31071 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 2417 742 2422 770
rect 2450 742 6678 770
rect 6706 742 6711 770
rect 7126 742 10878 770
rect 10906 742 10911 770
rect 0 714 56 728
rect 7126 714 7154 742
rect 12110 714 12138 798
rect 14401 742 14406 770
rect 14434 742 17822 770
rect 17850 742 17855 770
rect 18489 742 18494 770
rect 18522 742 20286 770
rect 20314 742 20319 770
rect 21826 714 21854 798
rect 21897 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22039 798
rect 22129 742 22134 770
rect 22162 742 30254 770
rect 30282 742 30287 770
rect 31262 714 31290 854
rect 32144 714 32200 728
rect 0 686 4214 714
rect 6617 686 6622 714
rect 6650 686 7154 714
rect 7289 686 7294 714
rect 7322 686 10654 714
rect 10682 686 10687 714
rect 10929 686 10934 714
rect 10962 686 12138 714
rect 17705 686 17710 714
rect 17738 686 18858 714
rect 21826 686 28910 714
rect 28938 686 28943 714
rect 31262 686 32200 714
rect 0 672 56 686
rect 4186 546 4214 686
rect 4377 630 4382 658
rect 4410 630 5950 658
rect 5978 630 5983 658
rect 7681 630 7686 658
rect 7714 630 12782 658
rect 12810 630 12815 658
rect 13006 630 16590 658
rect 16618 630 16623 658
rect 17206 630 18270 658
rect 18298 630 18303 658
rect 13006 602 13034 630
rect 17206 602 17234 630
rect 7569 574 7574 602
rect 7602 574 13034 602
rect 13449 574 13454 602
rect 13482 574 17234 602
rect 17537 574 17542 602
rect 17570 574 18746 602
rect 18718 546 18746 574
rect 18830 546 18858 686
rect 32144 672 32200 686
rect 18937 630 18942 658
rect 18970 630 22582 658
rect 22610 630 22615 658
rect 22689 630 22694 658
rect 22722 630 28350 658
rect 28378 630 28383 658
rect 18937 574 18942 602
rect 18970 574 24850 602
rect 25545 574 25550 602
rect 25578 574 27678 602
rect 27706 574 27711 602
rect 24822 546 24850 574
rect 4186 518 9142 546
rect 9170 518 9175 546
rect 9249 518 9254 546
rect 9282 518 10430 546
rect 10458 518 10463 546
rect 10537 518 10542 546
rect 10570 518 14406 546
rect 14434 518 14439 546
rect 15129 518 15134 546
rect 15162 518 18438 546
rect 18466 518 18471 546
rect 18713 518 18718 546
rect 18746 518 18751 546
rect 18830 518 24682 546
rect 24822 518 26894 546
rect 26922 518 26927 546
rect 27706 518 31094 546
rect 31122 518 31127 546
rect 0 490 56 504
rect 0 462 602 490
rect 1185 462 1190 490
rect 1218 462 17486 490
rect 17514 462 17519 490
rect 18153 462 18158 490
rect 18186 462 23478 490
rect 23506 462 23511 490
rect 0 448 56 462
rect 574 322 602 462
rect 6113 406 6118 434
rect 6146 406 10822 434
rect 10850 406 10855 434
rect 15969 406 15974 434
rect 16002 406 18634 434
rect 20673 406 20678 434
rect 20706 406 22134 434
rect 22162 406 22167 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 18606 378 18634 406
rect 22227 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22369 406
rect 24654 378 24682 518
rect 27706 490 27734 518
rect 32144 490 32200 504
rect 26049 462 26054 490
rect 26082 462 27734 490
rect 30585 462 30590 490
rect 30618 462 32200 490
rect 32144 448 32200 462
rect 24873 406 24878 434
rect 24906 406 29414 434
rect 29442 406 29447 434
rect 6505 350 6510 378
rect 6538 350 11326 378
rect 11354 350 11359 378
rect 15129 350 15134 378
rect 15162 350 18046 378
rect 18074 350 18079 378
rect 18606 350 21126 378
rect 21154 350 21159 378
rect 24654 350 29302 378
rect 29330 350 29335 378
rect 574 294 6678 322
rect 6706 294 6711 322
rect 8521 294 8526 322
rect 8554 294 15974 322
rect 16002 294 16007 322
rect 16081 294 16086 322
rect 16114 294 22638 322
rect 22666 294 22671 322
rect 22801 294 22806 322
rect 22834 294 24878 322
rect 24906 294 24911 322
rect 0 266 56 280
rect 32144 266 32200 280
rect 0 238 5110 266
rect 5138 238 5143 266
rect 10425 238 10430 266
rect 10458 238 14238 266
rect 14266 238 14271 266
rect 14569 238 14574 266
rect 14602 238 24038 266
rect 24066 238 24071 266
rect 29801 238 29806 266
rect 29834 238 32200 266
rect 0 224 56 238
rect 32144 224 32200 238
rect 2142 182 5054 210
rect 5082 182 5087 210
rect 5166 182 6062 210
rect 6090 182 6095 210
rect 15946 182 23310 210
rect 23338 182 23343 210
rect 0 42 56 56
rect 2142 42 2170 182
rect 5166 154 5194 182
rect 2921 126 2926 154
rect 2954 126 5194 154
rect 5273 126 5278 154
rect 5306 126 13566 154
rect 13594 126 13599 154
rect 15946 98 15974 182
rect 17481 126 17486 154
rect 17514 126 25214 154
rect 25242 126 25247 154
rect 10201 70 10206 98
rect 10234 70 10374 98
rect 10402 70 10407 98
rect 11657 70 11662 98
rect 11690 70 11695 98
rect 14793 70 14798 98
rect 14826 70 15974 98
rect 21849 70 21854 98
rect 21882 70 25270 98
rect 25298 70 25303 98
rect 0 14 2170 42
rect 11662 42 11690 70
rect 32144 42 32200 56
rect 11662 14 16758 42
rect 16786 14 16791 42
rect 31369 14 31374 42
rect 31402 14 32200 42
rect 0 0 56 14
rect 32144 0 32200 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 22232 6650 22260 6678
rect 22284 6650 22312 6678
rect 22336 6650 22364 6678
rect 14014 6398 14042 6426
rect 18942 6398 18970 6426
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 21902 6258 21930 6286
rect 21954 6258 21982 6286
rect 22006 6258 22034 6286
rect 6230 6230 6258 6258
rect 22526 6230 22554 6258
rect 7462 6174 7490 6202
rect 18830 6174 18858 6202
rect 18942 6174 18970 6202
rect 22526 6118 22554 6146
rect 14518 6062 14546 6090
rect 18830 6062 18858 6090
rect 6230 6006 6258 6034
rect 7462 5950 7490 5978
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 14518 5894 14546 5922
rect 18046 5894 18074 5922
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 22232 5866 22260 5894
rect 22284 5866 22312 5894
rect 22336 5866 22364 5894
rect 2086 5838 2114 5866
rect 14854 5726 14882 5754
rect 15918 5558 15946 5586
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 21902 5474 21930 5502
rect 21954 5474 21982 5502
rect 22006 5474 22034 5502
rect 15190 5446 15218 5474
rect 21798 5446 21826 5474
rect 14070 5390 14098 5418
rect 14406 5334 14434 5362
rect 13398 5278 13426 5306
rect 14854 5278 14882 5306
rect 2086 5222 2114 5250
rect 18494 5222 18522 5250
rect 16814 5166 16842 5194
rect 21798 5166 21826 5194
rect 12614 5110 12642 5138
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 18494 5054 18522 5082
rect 22232 5082 22260 5110
rect 22284 5082 22312 5110
rect 22336 5082 22364 5110
rect 18550 4998 18578 5026
rect 13734 4942 13762 4970
rect 14686 4886 14714 4914
rect 18550 4830 18578 4858
rect 18662 4830 18690 4858
rect 20174 4830 20202 4858
rect 7574 4774 7602 4802
rect 1806 4718 1834 4746
rect 18606 4718 18634 4746
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 21902 4690 21930 4718
rect 21954 4690 21982 4718
rect 22006 4690 22034 4718
rect 10486 4550 10514 4578
rect 13622 4550 13650 4578
rect 15862 4550 15890 4578
rect 12502 4494 12530 4522
rect 14686 4494 14714 4522
rect 15974 4494 16002 4522
rect 1806 4438 1834 4466
rect 13398 4438 13426 4466
rect 15862 4382 15890 4410
rect 18158 4382 18186 4410
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 10486 4326 10514 4354
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 22232 4298 22260 4326
rect 22284 4298 22312 4326
rect 22336 4298 22364 4326
rect 7574 4214 7602 4242
rect 15078 4214 15106 4242
rect 12558 4158 12586 4186
rect 17822 4158 17850 4186
rect 13398 4102 13426 4130
rect 10486 4046 10514 4074
rect 12502 3990 12530 4018
rect 17822 3990 17850 4018
rect 10486 3934 10514 3962
rect 12110 3934 12138 3962
rect 13454 3934 13482 3962
rect 20174 3934 20202 3962
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 21902 3906 21930 3934
rect 21954 3906 21982 3934
rect 22006 3906 22034 3934
rect 13454 3822 13482 3850
rect 18998 3766 19026 3794
rect 12110 3710 12138 3738
rect 13622 3710 13650 3738
rect 14854 3710 14882 3738
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 22232 3514 22260 3542
rect 22284 3514 22312 3542
rect 22336 3514 22364 3542
rect 14966 3486 14994 3514
rect 16814 3430 16842 3458
rect 13454 3374 13482 3402
rect 13678 3374 13706 3402
rect 15134 3374 15162 3402
rect 18998 3374 19026 3402
rect 7070 3318 7098 3346
rect 12558 3318 12586 3346
rect 12838 3318 12866 3346
rect 12558 3206 12586 3234
rect 12782 3206 12810 3234
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 21902 3122 21930 3150
rect 21954 3122 21982 3150
rect 22006 3122 22034 3150
rect 7070 3094 7098 3122
rect 12838 3094 12866 3122
rect 13734 3094 13762 3122
rect 12502 3038 12530 3066
rect 14014 2982 14042 3010
rect 22414 2758 22442 2786
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 22232 2730 22260 2758
rect 22284 2730 22312 2758
rect 22336 2730 22364 2758
rect 22414 2534 22442 2562
rect 13454 2366 13482 2394
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 21902 2338 21930 2366
rect 21954 2338 21982 2366
rect 22006 2338 22034 2366
rect 12670 2254 12698 2282
rect 6678 2086 6706 2114
rect 12670 2086 12698 2114
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 12446 1918 12474 1946
rect 13678 1918 13706 1946
rect 22232 1946 22260 1974
rect 22284 1946 22312 1974
rect 22336 1946 22364 1974
rect 12446 1806 12474 1834
rect 17318 1694 17346 1722
rect 18494 1694 18522 1722
rect 11830 1638 11858 1666
rect 13622 1638 13650 1666
rect 22134 1582 22162 1610
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 21902 1554 21930 1582
rect 21954 1554 21982 1582
rect 22006 1554 22034 1582
rect 15190 1526 15218 1554
rect 17318 1414 17346 1442
rect 15078 1190 15106 1218
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 11830 1134 11858 1162
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 22232 1162 22260 1190
rect 22284 1162 22312 1190
rect 22336 1162 22364 1190
rect 8190 1022 8218 1050
rect 22134 1022 22162 1050
rect 8190 854 8218 882
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 18494 742 18522 770
rect 21902 770 21930 798
rect 21954 770 21982 798
rect 22006 770 22034 798
rect 22134 742 22162 770
rect 18942 574 18970 602
rect 10430 518 10458 546
rect 18718 518 18746 546
rect 18158 462 18186 490
rect 22134 406 22162 434
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 22232 378 22260 406
rect 22284 378 22312 406
rect 22336 378 22364 406
rect 15134 350 15162 378
rect 18046 350 18074 378
rect 6678 294 6706 322
rect 10430 238 10458 266
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 11888 6286 12048 7112
rect 6230 6258 6258 6263
rect 6230 6034 6258 6230
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 6230 6001 6258 6006
rect 7462 6202 7490 6207
rect 7462 5978 7490 6174
rect 7462 5945 7490 5950
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1806 4746 1834 4751
rect 1806 4466 1834 4718
rect 1806 4433 1834 4438
rect 1888 4718 2048 5474
rect 2086 5866 2114 5871
rect 2086 5250 2114 5838
rect 2086 5217 2114 5222
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 5110 2378 5866
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 7574 4802 7602 4807
rect 7574 4242 7602 4774
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 10486 4578 10514 4583
rect 10486 4354 10514 4550
rect 10486 4321 10514 4326
rect 7574 4209 7602 4214
rect 10486 4074 10514 4079
rect 10486 3962 10514 4046
rect 10486 3929 10514 3934
rect 11888 3934 12048 4690
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 14014 6426 14042 6431
rect 13398 5306 13426 5311
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 12614 5138 12642 5143
rect 12614 4559 12642 5110
rect 12502 4531 12642 4559
rect 12502 4522 12530 4531
rect 12502 4489 12530 4494
rect 13398 4466 13426 5278
rect 13734 4970 13762 4975
rect 13398 4433 13426 4438
rect 13622 4578 13650 4583
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 7070 3346 7098 3351
rect 7070 3122 7098 3318
rect 7070 3089 7098 3094
rect 11888 3150 12048 3906
rect 12110 3962 12138 3967
rect 12110 3738 12138 3934
rect 12110 3705 12138 3710
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 6678 2114 6706 2119
rect 6678 322 6706 2086
rect 11830 1666 11858 1671
rect 11830 1162 11858 1638
rect 11830 1129 11858 1134
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 8190 1050 8218 1055
rect 8190 882 8218 1022
rect 8190 849 8218 854
rect 11888 798 12048 1554
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 6678 289 6706 294
rect 10430 546 10458 551
rect 10430 266 10458 518
rect 10430 233 10458 238
rect 11888 0 12048 770
rect 12218 3542 12378 4298
rect 12558 4186 12586 4191
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12502 4018 12530 4023
rect 12502 3066 12530 3990
rect 12558 3346 12586 4158
rect 13398 4130 13426 4135
rect 13426 4102 13482 4109
rect 13398 4081 13482 4102
rect 13454 3962 13482 4081
rect 13454 3929 13482 3934
rect 13454 3850 13482 3855
rect 13622 3839 13650 4550
rect 13482 3822 13650 3839
rect 13454 3811 13650 3822
rect 13622 3738 13650 3743
rect 13454 3402 13482 3407
rect 12558 3313 12586 3318
rect 12838 3346 12866 3351
rect 12558 3234 12586 3239
rect 12782 3234 12810 3239
rect 12586 3206 12782 3209
rect 12558 3181 12810 3206
rect 12838 3122 12866 3318
rect 12838 3089 12866 3094
rect 12502 3033 12530 3038
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 13454 2394 13482 3374
rect 13454 2361 13482 2366
rect 12670 2282 12698 2287
rect 12670 2114 12698 2254
rect 12670 2081 12698 2086
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12446 1946 12474 1951
rect 12446 1834 12474 1918
rect 12446 1801 12474 1806
rect 13622 1666 13650 3710
rect 13678 3402 13706 3407
rect 13678 1946 13706 3374
rect 13734 3122 13762 4942
rect 13734 3089 13762 3094
rect 14014 3010 14042 6398
rect 18942 6426 18970 6431
rect 18830 6202 18858 6207
rect 14518 6090 14546 6095
rect 14518 5922 14546 6062
rect 18830 6090 18858 6174
rect 18942 6202 18970 6398
rect 18942 6169 18970 6174
rect 21888 6286 22048 7112
rect 21888 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22048 6286
rect 18830 6057 18858 6062
rect 14518 5889 14546 5894
rect 18046 5922 18074 5927
rect 14854 5754 14882 5759
rect 14070 5418 14098 5423
rect 14070 5369 14098 5390
rect 14070 5362 14434 5369
rect 14070 5341 14406 5362
rect 14406 5329 14434 5334
rect 14854 5306 14882 5726
rect 15918 5586 15946 5591
rect 14854 5273 14882 5278
rect 15190 5474 15218 5479
rect 14686 4914 14714 4919
rect 14686 4522 14714 4886
rect 14686 4489 14714 4494
rect 15078 4242 15106 4247
rect 14854 3738 14882 3743
rect 14854 3659 14882 3710
rect 14854 3631 14994 3659
rect 14966 3514 14994 3631
rect 14966 3481 14994 3486
rect 14014 2977 14042 2982
rect 13678 1913 13706 1918
rect 13622 1633 13650 1638
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 15078 1218 15106 4214
rect 15078 1185 15106 1190
rect 15134 3402 15162 3407
rect 12218 406 12378 1162
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 15134 378 15162 3374
rect 15190 1554 15218 5446
rect 15862 4578 15890 4583
rect 15862 4410 15890 4550
rect 15918 4559 15946 5558
rect 16814 5194 16842 5199
rect 15918 4531 16002 4559
rect 15974 4522 16002 4531
rect 15974 4489 16002 4494
rect 15862 4377 15890 4382
rect 16814 3458 16842 5166
rect 17822 4186 17850 4191
rect 17822 4018 17850 4158
rect 17822 3985 17850 3990
rect 16814 3425 16842 3430
rect 15190 1521 15218 1526
rect 17318 1722 17346 1727
rect 17318 1442 17346 1694
rect 17318 1409 17346 1414
rect 15134 345 15162 350
rect 18046 378 18074 5894
rect 21888 5502 22048 6258
rect 21798 5474 21826 5479
rect 18494 5250 18522 5255
rect 18494 5082 18522 5222
rect 21798 5194 21826 5446
rect 21798 5161 21826 5166
rect 21888 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22048 5502
rect 18494 5049 18522 5054
rect 18550 5026 18578 5031
rect 18550 4858 18578 4998
rect 18550 4825 18578 4830
rect 18662 4858 18690 4863
rect 18662 4829 18690 4830
rect 18606 4801 18690 4829
rect 20174 4858 20202 4863
rect 18606 4746 18634 4801
rect 18606 4713 18634 4718
rect 18158 4410 18186 4415
rect 18158 490 18186 4382
rect 20174 3962 20202 4830
rect 20174 3929 20202 3934
rect 21888 4718 22048 5474
rect 21888 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22048 4718
rect 21888 3934 22048 4690
rect 21888 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22048 3934
rect 18998 3794 19026 3799
rect 18998 3402 19026 3766
rect 18998 3369 19026 3374
rect 21888 3150 22048 3906
rect 21888 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22048 3150
rect 21888 2366 22048 3122
rect 21888 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22048 2366
rect 18494 1722 18522 1727
rect 18494 770 18522 1694
rect 18494 737 18522 742
rect 21888 1582 22048 2338
rect 22218 6678 22378 7112
rect 22218 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22378 6678
rect 22218 5894 22378 6650
rect 22526 6258 22554 6263
rect 22526 6146 22554 6230
rect 22526 6113 22554 6118
rect 22218 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22378 5894
rect 22218 5110 22378 5866
rect 22218 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22378 5110
rect 22218 4326 22378 5082
rect 22218 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22378 4326
rect 22218 3542 22378 4298
rect 22218 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22378 3542
rect 22218 2758 22378 3514
rect 22218 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22378 2758
rect 22218 1974 22378 2730
rect 22414 2786 22442 2791
rect 22414 2562 22442 2758
rect 22414 2529 22442 2534
rect 22218 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22378 1974
rect 21888 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22048 1582
rect 21888 798 22048 1554
rect 22134 1610 22162 1615
rect 22134 1050 22162 1582
rect 22134 1017 22162 1022
rect 22218 1190 22378 1946
rect 22218 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22378 1190
rect 21888 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22048 798
rect 18942 602 18970 607
rect 18718 574 18942 599
rect 18718 571 18970 574
rect 18718 546 18746 571
rect 18942 569 18970 571
rect 18718 513 18746 518
rect 18158 457 18186 462
rect 18046 345 18074 350
rect 21888 0 22048 770
rect 22134 770 22162 775
rect 22134 434 22162 742
rect 22134 401 22162 406
rect 22218 406 22378 1162
rect 22218 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22378 406
rect 22218 0 22378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 4928 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 4928 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 28840 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 28448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 4480 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 29624 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 29624 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 29288 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 28896 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 2520 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 28280 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 28840 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 29624 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 6160 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 8568 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 10416 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 10752 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 29288 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 6160 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 31024 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 29624 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 6440 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 28616 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 3808 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 27888 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 27888 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 29232 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 28840 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 28504 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 2296 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 29288 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 13944 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 14560 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform 1 0 17528 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 20328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 21448 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 21448 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform 1 0 22008 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform 1 0 22120 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform 1 0 23968 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform 1 0 24528 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform 1 0 25088 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform 1 0 23744 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform 1 0 25088 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform 1 0 25144 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 14896 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 20496 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 22064 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 23464 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 26376 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 28168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 1344 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform -1 0 4424 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform -1 0 8176 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform -1 0 11536 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform -1 0 8736 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform -1 0 8736 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform -1 0 9744 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform -1 0 7728 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform -1 0 12096 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform -1 0 14896 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 17360 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform -1 0 12656 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 26320 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 28840 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 28392 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 29176 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 23408 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 28056 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 20104 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 21392 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 16576 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform -1 0 15176 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform -1 0 8624 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform -1 0 1288 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 1400 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform -1 0 1344 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 1288 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform -1 0 1344 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 9128 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform -1 0 11032 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 1288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform -1 0 7728 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 15456 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 13664 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 18536 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 1736 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform -1 0 25368 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform -1 0 23632 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 24640 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 23016 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 21896 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 21000 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 21448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 21280 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 21392 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 21224 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 20608 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 19152 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 18536 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 19824 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 18032 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 15568 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform 1 0 15176 0 -1 1176
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6
timestamp 1486834041
transform 1 0 672 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8
timestamp 1486834041
transform 1 0 784 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17
timestamp 1486834041
transform 1 0 1288 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33
timestamp 1486834041
transform 1 0 2184 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78
timestamp 1486834041
transform 1 0 4704 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90
timestamp 1486834041
transform 1 0 5376 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98
timestamp 1486834041
transform 1 0 5824 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 15680 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 17584 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 19488 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 21392 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_410
timestamp 1486834041
transform 1 0 23296 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_444
timestamp 1486834041
transform 1 0 25200 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_478
timestamp 1486834041
transform 1 0 27104 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_512
timestamp 1486834041
transform 1 0 29008 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_546
timestamp 1486834041
transform 1 0 30912 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_18
timestamp 1486834041
transform 1 0 1344 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_50
timestamp 1486834041
transform 1 0 3136 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 4032 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_90
timestamp 1486834041
transform 1 0 5376 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_98
timestamp 1486834041
transform 1 0 5824 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_102
timestamp 1486834041
transform 1 0 6048 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_112
timestamp 1486834041
transform 1 0 6608 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_120
timestamp 1486834041
transform 1 0 7056 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_174
timestamp 1486834041
transform 1 0 10080 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_190
timestamp 1486834041
transform 1 0 10976 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_200
timestamp 1486834041
transform 1 0 11536 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_208
timestamp 1486834041
transform 1 0 11984 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_244
timestamp 1486834041
transform 1 0 14000 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_260
timestamp 1486834041
transform 1 0 14896 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_264
timestamp 1486834041
transform 1 0 15120 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_271
timestamp 1486834041
transform 1 0 15512 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_279
timestamp 1486834041
transform 1 0 15960 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_290
timestamp 1486834041
transform 1 0 16576 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_306
timestamp 1486834041
transform 1 0 17472 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_316
timestamp 1486834041
transform 1 0 18032 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_325
timestamp 1486834041
transform 1 0 18536 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_327
timestamp 1486834041
transform 1 0 18648 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_336
timestamp 1486834041
transform 1 0 19152 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_348
timestamp 1486834041
transform 1 0 19824 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_352
timestamp 1486834041
transform 1 0 20048 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_360
timestamp 1486834041
transform 1 0 20496 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_385
timestamp 1486834041
transform 1 0 21896 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_393
timestamp 1486834041
transform 1 0 22344 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_405
timestamp 1486834041
transform 1 0 23016 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_413
timestamp 1486834041
transform 1 0 23464 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1486834041
transform 1 0 23688 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1486834041
transform 1 0 23800 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_430
timestamp 1486834041
transform 1 0 24416 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_440
timestamp 1486834041
transform 1 0 24976 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_450
timestamp 1486834041
transform 1 0 25536 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_482
timestamp 1486834041
transform 1 0 27328 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_492
timestamp 1486834041
transform 1 0 27888 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_500
timestamp 1486834041
transform 1 0 28336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_518
timestamp 1486834041
transform 1 0 29344 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_522
timestamp 1486834041
transform 1 0 29568 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 13832 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_247
timestamp 1486834041
transform 1 0 14168 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1486834041
transform 1 0 17752 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_317
timestamp 1486834041
transform 1 0 18088 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_381
timestamp 1486834041
transform 1 0 21672 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_387
timestamp 1486834041
transform 1 0 22008 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 25592 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_465
timestamp 1486834041
transform 1 0 26376 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_497
timestamp 1486834041
transform 1 0 28168 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_505
timestamp 1486834041
transform 1 0 28616 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1486834041
transform 1 0 29848 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_531
timestamp 1486834041
transform 1 0 30072 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_10
timestamp 1486834041
transform 1 0 896 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_19
timestamp 1486834041
transform 1 0 1400 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_35
timestamp 1486834041
transform 1 0 2296 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_47
timestamp 1486834041
transform 1 0 2968 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_63
timestamp 1486834041
transform 1 0 3864 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_67
timestamp 1486834041
transform 1 0 4088 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_69
timestamp 1486834041
transform 1 0 4200 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 7952 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_150
timestamp 1486834041
transform 1 0 8736 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_182
timestamp 1486834041
transform 1 0 10528 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_198
timestamp 1486834041
transform 1 0 11424 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_212
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_276
timestamp 1486834041
transform 1 0 15792 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_282
timestamp 1486834041
transform 1 0 16128 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_346
timestamp 1486834041
transform 1 0 19712 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_360
timestamp 1486834041
transform 1 0 20496 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_376
timestamp 1486834041
transform 1 0 21392 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_384
timestamp 1486834041
transform 1 0 21840 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_388
timestamp 1486834041
transform 1 0 22064 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_397
timestamp 1486834041
transform 1 0 22568 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_405
timestamp 1486834041
transform 1 0 23016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_407
timestamp 1486834041
transform 1 0 23128 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 23632 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_422
timestamp 1486834041
transform 1 0 23968 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_438
timestamp 1486834041
transform 1 0 24864 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_447
timestamp 1486834041
transform 1 0 25368 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_479
timestamp 1486834041
transform 1 0 27160 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_487
timestamp 1486834041
transform 1 0 27608 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_489
timestamp 1486834041
transform 1 0 27720 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_492
timestamp 1486834041
transform 1 0 27888 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_508
timestamp 1486834041
transform 1 0 28784 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_516
timestamp 1486834041
transform 1 0 29232 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_520
timestamp 1486834041
transform 1 0 29456 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_522
timestamp 1486834041
transform 1 0 29568 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1486834041
transform 1 0 672 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_8
timestamp 1486834041
transform 1 0 784 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_17
timestamp 1486834041
transform 1 0 1288 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_33
timestamp 1486834041
transform 1 0 2184 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_139
timestamp 1486834041
transform 1 0 8120 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_148
timestamp 1486834041
transform 1 0 8624 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_164
timestamp 1486834041
transform 1 0 9520 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_172
timestamp 1486834041
transform 1 0 9968 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_174
timestamp 1486834041
transform 1 0 10080 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 13832 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 17752 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_317
timestamp 1486834041
transform 1 0 18088 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_349
timestamp 1486834041
transform 1 0 19880 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_365
timestamp 1486834041
transform 1 0 20776 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_367
timestamp 1486834041
transform 1 0 20888 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_376
timestamp 1486834041
transform 1 0 21392 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_384
timestamp 1486834041
transform 1 0 21840 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_387
timestamp 1486834041
transform 1 0 22008 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_419
timestamp 1486834041
transform 1 0 23800 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_423
timestamp 1486834041
transform 1 0 24024 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_425
timestamp 1486834041
transform 1 0 24136 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_434
timestamp 1486834041
transform 1 0 24640 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_450
timestamp 1486834041
transform 1 0 25536 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_454
timestamp 1486834041
transform 1 0 25760 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_457
timestamp 1486834041
transform 1 0 25928 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_497
timestamp 1486834041
transform 1 0 28168 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_513
timestamp 1486834041
transform 1 0 29064 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_521
timestamp 1486834041
transform 1 0 29512 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1486834041
transform 1 0 29848 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_531
timestamp 1486834041
transform 1 0 30072 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_18
timestamp 1486834041
transform 1 0 1344 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_50
timestamp 1486834041
transform 1 0 3136 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 4032 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 7952 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_150
timestamp 1486834041
transform 1 0 8736 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_158
timestamp 1486834041
transform 1 0 9184 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_168
timestamp 1486834041
transform 1 0 9744 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_176
timestamp 1486834041
transform 1 0 10192 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_180
timestamp 1486834041
transform 1 0 10416 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_182
timestamp 1486834041
transform 1 0 10528 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_191
timestamp 1486834041
transform 1 0 11032 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_207
timestamp 1486834041
transform 1 0 11928 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_220
timestamp 1486834041
transform 1 0 12656 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_260
timestamp 1486834041
transform 1 0 14896 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_276
timestamp 1486834041
transform 1 0 15792 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_282
timestamp 1486834041
transform 1 0 16128 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_346
timestamp 1486834041
transform 1 0 19712 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_352
timestamp 1486834041
transform 1 0 20048 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_361
timestamp 1486834041
transform 1 0 20552 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_365
timestamp 1486834041
transform 1 0 20776 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_374
timestamp 1486834041
transform 1 0 21280 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_384
timestamp 1486834041
transform 1 0 21840 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 23632 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_422
timestamp 1486834041
transform 1 0 23968 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_438
timestamp 1486834041
transform 1 0 24864 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_450
timestamp 1486834041
transform 1 0 25536 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_482
timestamp 1486834041
transform 1 0 27328 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 27888 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 28112 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 28224 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_507
timestamp 1486834041
transform 1 0 28728 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_517
timestamp 1486834041
transform 1 0 29288 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_521
timestamp 1486834041
transform 1 0 29512 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_18
timestamp 1486834041
transform 1 0 1344 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1486834041
transform 1 0 3304 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_61
timestamp 1486834041
transform 1 0 3752 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_73
timestamp 1486834041
transform 1 0 4424 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 9912 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_209
timestamp 1486834041
transform 1 0 12040 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_225
timestamp 1486834041
transform 1 0 12936 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_229
timestamp 1486834041
transform 1 0 13160 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_238
timestamp 1486834041
transform 1 0 13664 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1486834041
transform 1 0 13888 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1486834041
transform 1 0 14000 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_255
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_265
timestamp 1486834041
transform 1 0 15176 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_297
timestamp 1486834041
transform 1 0 16968 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_313
timestamp 1486834041
transform 1 0 17864 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_317
timestamp 1486834041
transform 1 0 18088 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_381
timestamp 1486834041
transform 1 0 21672 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_395
timestamp 1486834041
transform 1 0 22456 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_427
timestamp 1486834041
transform 1 0 24248 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_443
timestamp 1486834041
transform 1 0 25144 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_451
timestamp 1486834041
transform 1 0 25592 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_457
timestamp 1486834041
transform 1 0 25928 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_489
timestamp 1486834041
transform 1 0 27720 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_513
timestamp 1486834041
transform 1 0 29064 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1486834041
transform 1 0 29848 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_531
timestamp 1486834041
transform 1 0 30072 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 4032 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1486834041
transform 1 0 7952 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_142
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_146
timestamp 1486834041
transform 1 0 8512 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_148
timestamp 1486834041
transform 1 0 8624 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_157
timestamp 1486834041
transform 1 0 9128 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_189
timestamp 1486834041
transform 1 0 10920 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_205
timestamp 1486834041
transform 1 0 11816 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_209
timestamp 1486834041
transform 1 0 12040 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_244
timestamp 1486834041
transform 1 0 14000 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_260
timestamp 1486834041
transform 1 0 14896 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_270
timestamp 1486834041
transform 1 0 15456 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_278
timestamp 1486834041
transform 1 0 15904 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_282
timestamp 1486834041
transform 1 0 16128 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1486834041
transform 1 0 17920 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_316
timestamp 1486834041
transform 1 0 18032 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_325
timestamp 1486834041
transform 1 0 18536 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_341
timestamp 1486834041
transform 1 0 19432 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_349
timestamp 1486834041
transform 1 0 19880 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_352
timestamp 1486834041
transform 1 0 20048 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_384
timestamp 1486834041
transform 1 0 21840 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_400
timestamp 1486834041
transform 1 0 22736 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_408
timestamp 1486834041
transform 1 0 23184 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_422
timestamp 1486834041
transform 1 0 23968 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_438
timestamp 1486834041
transform 1 0 24864 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_442
timestamp 1486834041
transform 1 0 25088 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_451
timestamp 1486834041
transform 1 0 25592 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_483
timestamp 1486834041
transform 1 0 27384 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_487
timestamp 1486834041
transform 1 0 27608 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_489
timestamp 1486834041
transform 1 0 27720 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_492
timestamp 1486834041
transform 1 0 27888 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_508
timestamp 1486834041
transform 1 0 28784 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_512
timestamp 1486834041
transform 1 0 29008 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_514
timestamp 1486834041
transform 1 0 29120 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 5992 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_123
timestamp 1486834041
transform 1 0 7224 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_132
timestamp 1486834041
transform 1 0 7728 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_164
timestamp 1486834041
transform 1 0 9520 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_172
timestamp 1486834041
transform 1 0 9968 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 10080 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 13832 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_279
timestamp 1486834041
transform 1 0 15960 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_295
timestamp 1486834041
transform 1 0 16856 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_303
timestamp 1486834041
transform 1 0 17304 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_312
timestamp 1486834041
transform 1 0 17808 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 17920 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_317
timestamp 1486834041
transform 1 0 18088 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_349
timestamp 1486834041
transform 1 0 19880 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_373
timestamp 1486834041
transform 1 0 21224 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 21672 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_387
timestamp 1486834041
transform 1 0 22008 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_451
timestamp 1486834041
transform 1 0 25592 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_457
timestamp 1486834041
transform 1 0 25928 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_489
timestamp 1486834041
transform 1 0 27720 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_505
timestamp 1486834041
transform 1 0 28616 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1486834041
transform 1 0 29848 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_531
timestamp 1486834041
transform 1 0 30072 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_34
timestamp 1486834041
transform 1 0 2240 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_43
timestamp 1486834041
transform 1 0 2744 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_59
timestamp 1486834041
transform 1 0 3640 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_67
timestamp 1486834041
transform 1 0 4088 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_69
timestamp 1486834041
transform 1 0 4200 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_112
timestamp 1486834041
transform 1 0 6608 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_128
timestamp 1486834041
transform 1 0 7504 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 7952 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 11872 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_276
timestamp 1486834041
transform 1 0 15792 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_282
timestamp 1486834041
transform 1 0 16128 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 19712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_352
timestamp 1486834041
transform 1 0 20048 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_368
timestamp 1486834041
transform 1 0 20944 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_376
timestamp 1486834041
transform 1 0 21392 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_388
timestamp 1486834041
transform 1 0 22064 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_422
timestamp 1486834041
transform 1 0 23968 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_486
timestamp 1486834041
transform 1 0 27552 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_500
timestamp 1486834041
transform 1 0 28336 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_10
timestamp 1486834041
transform 1 0 896 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_14
timestamp 1486834041
transform 1 0 1120 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_16
timestamp 1486834041
transform 1 0 1232 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_25
timestamp 1486834041
transform 1 0 1736 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1486834041
transform 1 0 2184 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_45
timestamp 1486834041
transform 1 0 2856 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_77
timestamp 1486834041
transform 1 0 4648 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_93
timestamp 1486834041
transform 1 0 5544 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 5992 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_139
timestamp 1486834041
transform 1 0 8120 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_155
timestamp 1486834041
transform 1 0 9016 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_185
timestamp 1486834041
transform 1 0 10696 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_194
timestamp 1486834041
transform 1 0 11200 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_226
timestamp 1486834041
transform 1 0 12992 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_242
timestamp 1486834041
transform 1 0 13888 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_244
timestamp 1486834041
transform 1 0 14000 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_247
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_251
timestamp 1486834041
transform 1 0 14392 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_260
timestamp 1486834041
transform 1 0 14896 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_292
timestamp 1486834041
transform 1 0 16688 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_308
timestamp 1486834041
transform 1 0 17584 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_312
timestamp 1486834041
transform 1 0 17808 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_314
timestamp 1486834041
transform 1 0 17920 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_317
timestamp 1486834041
transform 1 0 18088 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_349
timestamp 1486834041
transform 1 0 19880 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_353
timestamp 1486834041
transform 1 0 20104 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_362
timestamp 1486834041
transform 1 0 20608 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_378
timestamp 1486834041
transform 1 0 21504 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_382
timestamp 1486834041
transform 1 0 21728 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_384
timestamp 1486834041
transform 1 0 21840 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_387
timestamp 1486834041
transform 1 0 22008 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_403
timestamp 1486834041
transform 1 0 22904 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_411
timestamp 1486834041
transform 1 0 23352 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_415
timestamp 1486834041
transform 1 0 23576 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_417
timestamp 1486834041
transform 1 0 23688 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_426
timestamp 1486834041
transform 1 0 24192 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_442
timestamp 1486834041
transform 1 0 25088 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_450
timestamp 1486834041
transform 1 0 25536 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_454
timestamp 1486834041
transform 1 0 25760 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_457
timestamp 1486834041
transform 1 0 25928 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_461
timestamp 1486834041
transform 1 0 26152 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1486834041
transform 1 0 26264 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_472
timestamp 1486834041
transform 1 0 26768 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_488
timestamp 1486834041
transform 1 0 27664 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_492
timestamp 1486834041
transform 1 0 27888 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_494
timestamp 1486834041
transform 1 0 28000 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1486834041
transform 1 0 29848 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_531
timestamp 1486834041
transform 1 0 30072 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_34
timestamp 1486834041
transform 1 0 2240 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_50
timestamp 1486834041
transform 1 0 3136 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_58
timestamp 1486834041
transform 1 0 3584 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_80
timestamp 1486834041
transform 1 0 4816 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_84
timestamp 1486834041
transform 1 0 5040 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_99
timestamp 1486834041
transform 1 0 5880 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_115
timestamp 1486834041
transform 1 0 6776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 7672 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 8120 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 11872 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 15792 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_282
timestamp 1486834041
transform 1 0 16128 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 19712 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_352
timestamp 1486834041
transform 1 0 20048 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1486834041
transform 1 0 23632 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_422
timestamp 1486834041
transform 1 0 23968 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_486
timestamp 1486834041
transform 1 0 27552 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_500
timestamp 1486834041
transform 1 0 28336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_502
timestamp 1486834041
transform 1 0 28448 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_45
timestamp 1486834041
transform 1 0 2856 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_107
timestamp 1486834041
transform 1 0 6328 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_117
timestamp 1486834041
transform 1 0 6888 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1486834041
transform 1 0 10360 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_188
timestamp 1486834041
transform 1 0 10864 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_203
timestamp 1486834041
transform 1 0 11704 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_219
timestamp 1486834041
transform 1 0 12600 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_235
timestamp 1486834041
transform 1 0 13496 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1486834041
transform 1 0 13944 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 17752 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_317
timestamp 1486834041
transform 1 0 18088 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_349
timestamp 1486834041
transform 1 0 19880 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_365
timestamp 1486834041
transform 1 0 20776 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_373
timestamp 1486834041
transform 1 0 21224 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_387
timestamp 1486834041
transform 1 0 22008 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_451
timestamp 1486834041
transform 1 0 25592 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_457
timestamp 1486834041
transform 1 0 25928 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_473
timestamp 1486834041
transform 1 0 26824 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_481
timestamp 1486834041
transform 1 0 27272 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1486834041
transform 1 0 29848 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_531
timestamp 1486834041
transform 1 0 30072 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_6
timestamp 1486834041
transform 1 0 672 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_8
timestamp 1486834041
transform 1 0 784 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_17
timestamp 1486834041
transform 1 0 1288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_25
timestamp 1486834041
transform 1 0 1736 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_27
timestamp 1486834041
transform 1 0 1848 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 4816 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_150
timestamp 1486834041
transform 1 0 8736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_212
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_220
timestamp 1486834041
transform 1 0 12656 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_224
timestamp 1486834041
transform 1 0 12880 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_239
timestamp 1486834041
transform 1 0 13720 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_251
timestamp 1486834041
transform 1 0 14392 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_267
timestamp 1486834041
transform 1 0 15288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_275
timestamp 1486834041
transform 1 0 15736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 15960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_282
timestamp 1486834041
transform 1 0 16128 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_346
timestamp 1486834041
transform 1 0 19712 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 20048 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_384
timestamp 1486834041
transform 1 0 21840 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_400
timestamp 1486834041
transform 1 0 22736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_404
timestamp 1486834041
transform 1 0 22960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1486834041
transform 1 0 23464 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1486834041
transform 1 0 23688 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1486834041
transform 1 0 23800 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_422
timestamp 1486834041
transform 1 0 23968 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_454
timestamp 1486834041
transform 1 0 25760 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_458
timestamp 1486834041
transform 1 0 25984 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_460
timestamp 1486834041
transform 1 0 26096 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 27720 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_556
timestamp 1486834041
transform 1 0 31472 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_558
timestamp 1486834041
transform 1 0 31584 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_18
timestamp 1486834041
transform 1 0 1344 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_20
timestamp 1486834041
transform 1 0 1456 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_45
timestamp 1486834041
transform 1 0 2856 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_115
timestamp 1486834041
transform 1 0 6776 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_177
timestamp 1486834041
transform 1 0 10248 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_185
timestamp 1486834041
transform 1 0 10696 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_243
timestamp 1486834041
transform 1 0 13944 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_247
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_251
timestamp 1486834041
transform 1 0 14392 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_253
timestamp 1486834041
transform 1 0 14504 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_262
timestamp 1486834041
transform 1 0 15008 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_272
timestamp 1486834041
transform 1 0 15568 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_304
timestamp 1486834041
transform 1 0 17360 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_306
timestamp 1486834041
transform 1 0 17472 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_317
timestamp 1486834041
transform 1 0 18088 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_349
timestamp 1486834041
transform 1 0 19880 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_365
timestamp 1486834041
transform 1 0 20776 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_373
timestamp 1486834041
transform 1 0 21224 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_387
timestamp 1486834041
transform 1 0 22008 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 25592 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_513
timestamp 1486834041
transform 1 0 29064 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_515
timestamp 1486834041
transform 1 0 29176 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_524
timestamp 1486834041
transform 1 0 29680 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_555
timestamp 1486834041
transform 1 0 31416 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_559
timestamp 1486834041
transform 1 0 31640 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_206
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_254
timestamp 1486834041
transform 1 0 14560 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_270
timestamp 1486834041
transform 1 0 15456 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 15680 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_308
timestamp 1486834041
transform 1 0 17584 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_342
timestamp 1486834041
transform 1 0 19488 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_376
timestamp 1486834041
transform 1 0 21392 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_410
timestamp 1486834041
transform 1 0 23296 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_444
timestamp 1486834041
transform 1 0 25200 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_446
timestamp 1486834041
transform 1 0 25312 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_467
timestamp 1486834041
transform 1 0 26488 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_475
timestamp 1486834041
transform 1 0 26936 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_506
timestamp 1486834041
transform 1 0 28672 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_540
timestamp 1486834041
transform 1 0 30576 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_560
timestamp 1486834041
transform 1 0 31696 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 30184 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 30072 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 30968 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 30856 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 30072 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 30968 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 30184 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 30856 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 30856 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 30968 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 30968 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 29232 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 30856 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 30968 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 30184 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 30072 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 30184 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 29288 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 30072 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform -1 0 29736 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 29288 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 28504 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 30016 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 30184 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform -1 0 28168 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 30072 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 30968 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 30856 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 30072 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 30968 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 30184 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 30856 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 25704 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 29008 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 28168 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 28672 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 29792 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 28952 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 29848 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 29456 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 30912 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 30632 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 30240 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 25928 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 26152 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 26712 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 27104 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 26936 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 27496 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 27888 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 28280 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 27888 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 672 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 2296 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 2688 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 2240 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 3472 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 3864 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 3360 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 3864 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 4648 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 4144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 5432 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 4648 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 5880 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 6216 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 5824 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 6608 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 6216 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 6048 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 8568 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 8960 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 10136 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 9352 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 9072 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 9352 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 7672 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 7784 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 6608 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 6384 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 7784 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 7000 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform 1 0 7392 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 7952 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 8568 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 10528 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 13160 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 12880 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 13720 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform -1 0 13944 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform -1 0 13664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 14560 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 9856 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform -1 0 11312 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 11704 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform -1 0 10976 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform -1 0 11592 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 12096 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 12600 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform -1 0 11760 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 12376 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 25704 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 31864 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 31864 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 31864 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 31864 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 31864 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 31864 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 31864 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 31864 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 31864 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 31864 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 31864 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 31864 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 31864 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 31864 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 31864 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 31864 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 15568 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 17472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 19376 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 21280 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 23184 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 25088 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 26992 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_46
timestamp 1486834041
transform 1 0 28896 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_47
timestamp 1486834041
transform 1 0 30800 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 16016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_53
timestamp 1486834041
transform 1 0 23856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_54
timestamp 1486834041
transform 1 0 27776 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_55
timestamp 1486834041
transform 1 0 31640 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_60
timestamp 1486834041
transform 1 0 17976 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_61
timestamp 1486834041
transform 1 0 21896 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_62
timestamp 1486834041
transform 1 0 25816 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_63
timestamp 1486834041
transform 1 0 29736 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_67
timestamp 1486834041
transform 1 0 16016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_68
timestamp 1486834041
transform 1 0 19936 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_69
timestamp 1486834041
transform 1 0 23856 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_70
timestamp 1486834041
transform 1 0 27776 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_71
timestamp 1486834041
transform 1 0 31640 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_74
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_75
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1486834041
transform 1 0 17976 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1486834041
transform 1 0 21896 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1486834041
transform 1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_79
timestamp 1486834041
transform 1 0 29736 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_82
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_83
timestamp 1486834041
transform 1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_84
timestamp 1486834041
transform 1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_85
timestamp 1486834041
transform 1 0 23856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_86
timestamp 1486834041
transform 1 0 27776 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_87
timestamp 1486834041
transform 1 0 31640 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_88
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_89
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_90
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_91
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_92
timestamp 1486834041
transform 1 0 17976 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_93
timestamp 1486834041
transform 1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_94
timestamp 1486834041
transform 1 0 25816 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_95
timestamp 1486834041
transform 1 0 29736 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_96
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_97
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_98
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_99
timestamp 1486834041
transform 1 0 16016 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_100
timestamp 1486834041
transform 1 0 19936 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_101
timestamp 1486834041
transform 1 0 23856 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_102
timestamp 1486834041
transform 1 0 27776 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_103
timestamp 1486834041
transform 1 0 31640 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_104
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_105
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_106
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_107
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_108
timestamp 1486834041
transform 1 0 17976 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_109
timestamp 1486834041
transform 1 0 21896 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1486834041
transform 1 0 25816 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1486834041
transform 1 0 29736 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_112
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_113
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1486834041
transform 1 0 16016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_116
timestamp 1486834041
transform 1 0 19936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_117
timestamp 1486834041
transform 1 0 23856 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_118
timestamp 1486834041
transform 1 0 27776 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_119
timestamp 1486834041
transform 1 0 31640 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_120
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_121
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_122
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_123
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_124
timestamp 1486834041
transform 1 0 17976 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_125
timestamp 1486834041
transform 1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_126
timestamp 1486834041
transform 1 0 25816 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_127
timestamp 1486834041
transform 1 0 29736 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_128
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_129
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_130
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_131
timestamp 1486834041
transform 1 0 16016 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_132
timestamp 1486834041
transform 1 0 19936 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_133
timestamp 1486834041
transform 1 0 23856 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_134
timestamp 1486834041
transform 1 0 27776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_135
timestamp 1486834041
transform 1 0 31640 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_136
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_137
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_138
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_139
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_140
timestamp 1486834041
transform 1 0 17976 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_141
timestamp 1486834041
transform 1 0 21896 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_142
timestamp 1486834041
transform 1 0 25816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_143
timestamp 1486834041
transform 1 0 29736 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_144
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_145
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_146
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_147
timestamp 1486834041
transform 1 0 16016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_148
timestamp 1486834041
transform 1 0 19936 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1486834041
transform 1 0 23856 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1486834041
transform 1 0 27776 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1486834041
transform 1 0 31640 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_152
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1486834041
transform 1 0 17976 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1486834041
transform 1 0 21896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1486834041
transform 1 0 25816 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1486834041
transform 1 0 29736 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_162
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_167
timestamp 1486834041
transform 1 0 15568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_168
timestamp 1486834041
transform 1 0 17472 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_169
timestamp 1486834041
transform 1 0 19376 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_170
timestamp 1486834041
transform 1 0 21280 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_171
timestamp 1486834041
transform 1 0 23184 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_172
timestamp 1486834041
transform 1 0 25088 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1486834041
transform 1 0 26992 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1486834041
transform 1 0 28896 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_175
timestamp 1486834041
transform 1 0 30800 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 32144 0 32200 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 32144 2240 32200 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 32144 2464 32200 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 32144 2688 32200 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 32144 2912 32200 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 32144 3136 32200 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 32144 3360 32200 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 32144 3584 32200 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 32144 3808 32200 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 32144 4032 32200 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 32144 4256 32200 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 32144 224 32200 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 32144 4480 32200 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 32144 4704 32200 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 32144 4928 32200 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 32144 5152 32200 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 32144 5376 32200 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 32144 5600 32200 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 32144 5824 32200 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 32144 6048 32200 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 32144 6272 32200 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 32144 6496 32200 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 32144 448 32200 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 32144 6720 32200 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 32144 6944 32200 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 32144 672 32200 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 32144 896 32200 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 32144 1120 32200 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 32144 1344 32200 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 32144 1568 32200 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 32144 1792 32200 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 32144 2016 32200 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 2912 0 2968 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 17472 0 17528 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 18928 0 18984 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 20384 0 20440 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 21840 0 21896 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 23296 0 23352 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 24752 0 24808 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 26208 0 26264 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 27664 0 27720 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 29120 0 29176 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 30576 0 30632 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 4368 0 4424 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 5824 0 5880 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 8736 0 8792 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 11648 0 11704 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 13104 0 13160 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 14560 0 14616 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 16016 0 16072 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 25648 7056 25704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 27888 7056 27944 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 28112 7056 28168 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 28336 7056 28392 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 28560 7056 28616 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 28784 7056 28840 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 29008 7056 29064 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 29232 7056 29288 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 29456 7056 29512 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 29680 7056 29736 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 29904 7056 29960 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 25872 7056 25928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 26096 7056 26152 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 26320 7056 26376 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 26544 7056 26600 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 26768 7056 26824 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 26992 7056 27048 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 27216 7056 27272 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 27440 7056 27496 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 27664 7056 27720 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2128 7056 2184 7112 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 2352 7056 2408 7112 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2576 7056 2632 7112 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 2800 7056 2856 7112 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3024 7056 3080 7112 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 3248 7056 3304 7112 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 3472 7056 3528 7112 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 3696 7056 3752 7112 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3920 7056 3976 7112 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 4144 7056 4200 7112 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 4368 7056 4424 7112 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 4592 7056 4648 7112 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4816 7056 4872 7112 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 5040 7056 5096 7112 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 5264 7056 5320 7112 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 5488 7056 5544 7112 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 5712 7056 5768 7112 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 5936 7056 5992 7112 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 6160 7056 6216 7112 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 6384 7056 6440 7112 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 6608 7056 6664 7112 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 8848 7056 8904 7112 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 9072 7056 9128 7112 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 9296 7056 9352 7112 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 9520 7056 9576 7112 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 9744 7056 9800 7112 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 9968 7056 10024 7112 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 6832 7056 6888 7112 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 7056 7056 7112 7112 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 7280 7056 7336 7112 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 7504 7056 7560 7112 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 7728 7056 7784 7112 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 7952 7056 8008 7112 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 8176 7056 8232 7112 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 8400 7056 8456 7112 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 8624 7056 8680 7112 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 10192 7056 10248 7112 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 12432 7056 12488 7112 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 12656 7056 12712 7112 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 12880 7056 12936 7112 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 13104 7056 13160 7112 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 13328 7056 13384 7112 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 13552 7056 13608 7112 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 10416 7056 10472 7112 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 10640 7056 10696 7112 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 10864 7056 10920 7112 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 11088 7056 11144 7112 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 11312 7056 11368 7112 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 11536 7056 11592 7112 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 11760 7056 11816 7112 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 11984 7056 12040 7112 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 12208 7056 12264 7112 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 13776 7056 13832 7112 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 14000 7056 14056 7112 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 14224 7056 14280 7112 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 14448 7056 14504 7112 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 16464 7056 16520 7112 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 16688 7056 16744 7112 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 16912 7056 16968 7112 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 17136 7056 17192 7112 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 17360 7056 17416 7112 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 17584 7056 17640 7112 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 17808 7056 17864 7112 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 18032 7056 18088 7112 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 14672 7056 14728 7112 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 14896 7056 14952 7112 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 15120 7056 15176 7112 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 15344 7056 15400 7112 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 15568 7056 15624 7112 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 15792 7056 15848 7112 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 16016 7056 16072 7112 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 16240 7056 16296 7112 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 18256 7056 18312 7112 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 20496 7056 20552 7112 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 20720 7056 20776 7112 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 20944 7056 21000 7112 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 21168 7056 21224 7112 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 21392 7056 21448 7112 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 21616 7056 21672 7112 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 18480 7056 18536 7112 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 18704 7056 18760 7112 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 18928 7056 18984 7112 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 19152 7056 19208 7112 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 19376 7056 19432 7112 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 19600 7056 19656 7112 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 19824 7056 19880 7112 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 20048 7056 20104 7112 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 20272 7056 20328 7112 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 21840 7056 21896 7112 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 24080 7056 24136 7112 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 24304 7056 24360 7112 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 24528 7056 24584 7112 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 24752 7056 24808 7112 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 24976 7056 25032 7112 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 25200 7056 25256 7112 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 22064 7056 22120 7112 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 22288 7056 22344 7112 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 22512 7056 22568 7112 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 22736 7056 22792 7112 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 22960 7056 23016 7112 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 23184 7056 23240 7112 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 23408 7056 23464 7112 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 23632 7056 23688 7112 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 23856 7056 23912 7112 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1456 0 1512 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 25424 7056 25480 7112 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 7084 22048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 7084 22378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 16100 6272 16100 6272 0 VDD
rlabel metal1 16100 6664 16100 6664 0 VSS
rlabel metal3 1099 28 1099 28 0 FrameData[0]
rlabel metal3 22708 840 22708 840 0 FrameData[10]
rlabel metal2 26068 1932 26068 1932 0 FrameData[11]
rlabel metal3 1071 2716 1071 2716 0 FrameData[12]
rlabel metal3 2121 2940 2121 2940 0 FrameData[13]
rlabel metal3 931 3164 931 3164 0 FrameData[14]
rlabel metal3 7140 3444 7140 3444 0 FrameData[15]
rlabel metal3 959 3612 959 3612 0 FrameData[16]
rlabel metal2 23996 3668 23996 3668 0 FrameData[17]
rlabel metal2 6188 2576 6188 2576 0 FrameData[18]
rlabel metal3 24836 3024 24836 3024 0 FrameData[19]
rlabel metal2 5124 616 5124 616 0 FrameData[1]
rlabel metal3 24780 3108 24780 3108 0 FrameData[20]
rlabel metal3 931 4732 931 4732 0 FrameData[21]
rlabel metal2 24276 3612 24276 3612 0 FrameData[22]
rlabel metal3 1967 5180 1967 5180 0 FrameData[23]
rlabel metal3 3171 5404 3171 5404 0 FrameData[24]
rlabel metal2 2548 4564 2548 4564 0 FrameData[25]
rlabel metal4 22148 1316 22148 1316 0 FrameData[26]
rlabel metal2 23324 5348 23324 5348 0 FrameData[27]
rlabel metal3 12180 1148 12180 1148 0 FrameData[28]
rlabel metal3 427 6524 427 6524 0 FrameData[29]
rlabel metal3 315 476 315 476 0 FrameData[2]
rlabel metal2 2240 4228 2240 4228 0 FrameData[30]
rlabel metal3 91 6972 91 6972 0 FrameData[31]
rlabel metal3 24836 560 24836 560 0 FrameData[3]
rlabel metal2 4564 952 4564 952 0 FrameData[4]
rlabel metal3 1071 1148 1071 1148 0 FrameData[5]
rlabel metal2 6132 896 6132 896 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal2 23492 700 23492 700 0 FrameData[8]
rlabel metal3 567 2044 567 2044 0 FrameData[9]
rlabel metal3 31773 28 31773 28 0 FrameData_O[0]
rlabel metal3 31717 2268 31717 2268 0 FrameData_O[10]
rlabel metal2 31556 2380 31556 2380 0 FrameData_O[11]
rlabel metal2 31332 2660 31332 2660 0 FrameData_O[12]
rlabel metal3 31409 2940 31409 2940 0 FrameData_O[13]
rlabel metal2 31556 3108 31556 3108 0 FrameData_O[14]
rlabel metal3 31465 3388 31465 3388 0 FrameData_O[15]
rlabel metal2 31444 3444 31444 3444 0 FrameData_O[16]
rlabel metal3 31801 3836 31801 3836 0 FrameData_O[17]
rlabel metal2 31556 3948 31556 3948 0 FrameData_O[18]
rlabel metal3 31801 4284 31801 4284 0 FrameData_O[19]
rlabel metal3 30989 252 30989 252 0 FrameData_O[1]
rlabel metal3 31773 4508 31773 4508 0 FrameData_O[20]
rlabel metal3 31801 4732 31801 4732 0 FrameData_O[21]
rlabel metal3 31773 4956 31773 4956 0 FrameData_O[22]
rlabel metal3 30884 4844 30884 4844 0 FrameData_O[23]
rlabel metal3 31052 4620 31052 4620 0 FrameData_O[24]
rlabel metal3 30632 4900 30632 4900 0 FrameData_O[25]
rlabel metal3 31052 4172 31052 4172 0 FrameData_O[26]
rlabel metal3 32025 6076 32025 6076 0 FrameData_O[27]
rlabel metal2 29876 4088 29876 4088 0 FrameData_O[28]
rlabel metal3 30128 4956 30128 4956 0 FrameData_O[29]
rlabel metal3 31381 476 31381 476 0 FrameData_O[2]
rlabel metal3 31444 3052 31444 3052 0 FrameData_O[30]
rlabel metal3 31297 6972 31297 6972 0 FrameData_O[31]
rlabel metal3 31717 700 31717 700 0 FrameData_O[3]
rlabel metal2 31556 812 31556 812 0 FrameData_O[4]
rlabel metal2 31444 1036 31444 1036 0 FrameData_O[5]
rlabel metal3 31745 1372 31745 1372 0 FrameData_O[6]
rlabel metal2 31556 1540 31556 1540 0 FrameData_O[7]
rlabel metal3 31409 1820 31409 1820 0 FrameData_O[8]
rlabel metal2 31444 1876 31444 1876 0 FrameData_O[9]
rlabel metal2 2940 91 2940 91 0 FrameStrobe[0]
rlabel metal2 25228 560 25228 560 0 FrameStrobe[10]
rlabel metal2 22596 1316 22596 1316 0 FrameStrobe[11]
rlabel metal4 22428 2660 22428 2660 0 FrameStrobe[12]
rlabel metal2 21868 63 21868 63 0 FrameStrobe[13]
rlabel metal2 23324 119 23324 119 0 FrameStrobe[14]
rlabel metal2 24780 1155 24780 1155 0 FrameStrobe[15]
rlabel metal2 26236 735 26236 735 0 FrameStrobe[16]
rlabel metal2 27692 315 27692 315 0 FrameStrobe[17]
rlabel metal2 26292 1064 26292 1064 0 FrameStrobe[18]
rlabel metal2 30604 203 30604 203 0 FrameStrobe[19]
rlabel metal2 4396 343 4396 343 0 FrameStrobe[1]
rlabel metal2 5852 427 5852 427 0 FrameStrobe[2]
rlabel metal2 10668 1036 10668 1036 0 FrameStrobe[3]
rlabel metal2 21476 5516 21476 5516 0 FrameStrobe[4]
rlabel metal2 10220 63 10220 63 0 FrameStrobe[5]
rlabel metal2 11676 63 11676 63 0 FrameStrobe[6]
rlabel metal2 13132 931 13132 931 0 FrameStrobe[7]
rlabel metal2 14588 147 14588 147 0 FrameStrobe[8]
rlabel metal2 22652 644 22652 644 0 FrameStrobe[9]
rlabel metal2 25676 6825 25676 6825 0 FrameStrobe_O[0]
rlabel metal2 27916 6741 27916 6741 0 FrameStrobe_O[10]
rlabel metal2 28140 6601 28140 6601 0 FrameStrobe_O[11]
rlabel metal2 28364 6769 28364 6769 0 FrameStrobe_O[12]
rlabel metal2 28588 6797 28588 6797 0 FrameStrobe_O[13]
rlabel metal2 28812 6601 28812 6601 0 FrameStrobe_O[14]
rlabel metal2 29036 6853 29036 6853 0 FrameStrobe_O[15]
rlabel metal2 29260 6713 29260 6713 0 FrameStrobe_O[16]
rlabel metal2 29484 6825 29484 6825 0 FrameStrobe_O[17]
rlabel metal2 29708 6601 29708 6601 0 FrameStrobe_O[18]
rlabel metal2 29932 6713 29932 6713 0 FrameStrobe_O[19]
rlabel metal2 25900 6629 25900 6629 0 FrameStrobe_O[1]
rlabel metal2 26124 6433 26124 6433 0 FrameStrobe_O[2]
rlabel metal2 26348 6797 26348 6797 0 FrameStrobe_O[3]
rlabel metal2 26572 6909 26572 6909 0 FrameStrobe_O[4]
rlabel metal2 26796 6713 26796 6713 0 FrameStrobe_O[5]
rlabel metal2 27020 6629 27020 6629 0 FrameStrobe_O[6]
rlabel metal2 27244 6825 27244 6825 0 FrameStrobe_O[7]
rlabel metal2 27468 6965 27468 6965 0 FrameStrobe_O[8]
rlabel metal2 27692 6993 27692 6993 0 FrameStrobe_O[9]
rlabel metal2 1260 6496 1260 6496 0 N1BEG[0]
rlabel metal2 2380 6909 2380 6909 0 N1BEG[1]
rlabel metal3 2464 5796 2464 5796 0 N1BEG[2]
rlabel metal2 1876 6692 1876 6692 0 N1BEG[3]
rlabel metal2 3052 6349 3052 6349 0 N2BEG[0]
rlabel metal2 3388 5964 3388 5964 0 N2BEG[1]
rlabel metal3 3248 6580 3248 6580 0 N2BEG[2]
rlabel metal2 3724 6629 3724 6629 0 N2BEG[3]
rlabel metal2 4116 5964 4116 5964 0 N2BEG[4]
rlabel metal3 4032 5796 4032 5796 0 N2BEG[5]
rlabel metal2 4396 6825 4396 6825 0 N2BEG[6]
rlabel metal2 4732 5404 4732 5404 0 N2BEG[7]
rlabel metal3 4564 6188 4564 6188 0 N2BEGb[0]
rlabel metal2 5068 6685 5068 6685 0 N2BEGb[1]
rlabel metal2 5292 6825 5292 6825 0 N2BEGb[2]
rlabel metal2 5628 5768 5628 5768 0 N2BEGb[3]
rlabel metal3 5600 5796 5600 5796 0 N2BEGb[4]
rlabel metal2 4900 6608 4900 6608 0 N2BEGb[5]
rlabel metal2 6188 6349 6188 6349 0 N2BEGb[6]
rlabel metal2 6412 6629 6412 6629 0 N2BEGb[7]
rlabel metal3 6160 6580 6160 6580 0 N4BEG[0]
rlabel metal2 8876 6237 8876 6237 0 N4BEG[10]
rlabel metal2 9100 6433 9100 6433 0 N4BEG[11]
rlabel metal2 9548 5796 9548 5796 0 N4BEG[12]
rlabel metal2 9548 6713 9548 6713 0 N4BEG[13]
rlabel metal2 8708 6608 8708 6608 0 N4BEG[14]
rlabel metal2 9968 6188 9968 6188 0 N4BEG[15]
rlabel metal2 6860 5957 6860 5957 0 N4BEG[1]
rlabel metal2 7168 5404 7168 5404 0 N4BEG[2]
rlabel metal2 7252 5628 7252 5628 0 N4BEG[3]
rlabel metal3 7252 6412 7252 6412 0 N4BEG[4]
rlabel metal2 7756 6237 7756 6237 0 N4BEG[5]
rlabel metal2 7476 6300 7476 6300 0 N4BEG[6]
rlabel metal2 8008 5628 8008 5628 0 N4BEG[7]
rlabel metal2 7420 6468 7420 6468 0 N4BEG[8]
rlabel metal2 8652 6825 8652 6825 0 N4BEG[9]
rlabel metal2 10192 5796 10192 5796 0 NN4BEG[0]
rlabel metal2 12516 6188 12516 6188 0 NN4BEG[10]
rlabel metal2 12516 6636 12516 6636 0 NN4BEG[11]
rlabel metal2 12908 6349 12908 6349 0 NN4BEG[12]
rlabel metal2 13132 6601 13132 6601 0 NN4BEG[13]
rlabel metal2 13328 6580 13328 6580 0 NN4BEG[14]
rlabel metal2 13580 6909 13580 6909 0 NN4BEG[15]
rlabel metal3 9968 6580 9968 6580 0 NN4BEG[1]
rlabel metal2 10668 6349 10668 6349 0 NN4BEG[2]
rlabel metal2 11088 5404 11088 5404 0 NN4BEG[3]
rlabel metal3 10864 6580 10864 6580 0 NN4BEG[4]
rlabel metal2 11340 6629 11340 6629 0 NN4BEG[5]
rlabel metal2 11564 6349 11564 6349 0 NN4BEG[6]
rlabel metal2 11928 5404 11928 5404 0 NN4BEG[7]
rlabel metal3 11704 6580 11704 6580 0 NN4BEG[8]
rlabel metal2 12236 6909 12236 6909 0 NN4BEG[9]
rlabel metal3 11816 5852 11816 5852 0 S1END[0]
rlabel metal3 9520 2940 9520 2940 0 S1END[1]
rlabel metal3 5376 2940 5376 2940 0 S1END[2]
rlabel metal2 1316 2996 1316 2996 0 S1END[3]
rlabel metal2 21476 2436 21476 2436 0 S2END[0]
rlabel metal2 20188 3668 20188 3668 0 S2END[1]
rlabel metal3 20692 4984 20692 4984 0 S2END[2]
rlabel metal2 17164 6153 17164 6153 0 S2END[3]
rlabel metal2 29260 3276 29260 3276 0 S2END[4]
rlabel metal2 23268 6020 23268 6020 0 S2END[5]
rlabel metal2 28924 3780 28924 3780 0 S2END[6]
rlabel metal2 26404 4564 26404 4564 0 S2END[7]
rlabel metal2 12572 3192 12572 3192 0 S2MID[0]
rlabel metal3 16212 3724 16212 3724 0 S2MID[1]
rlabel metal3 14980 4508 14980 4508 0 S2MID[2]
rlabel metal2 13188 4284 13188 4284 0 S2MID[3]
rlabel metal3 8764 1092 8764 1092 0 S2MID[4]
rlabel metal2 15820 4837 15820 4837 0 S2MID[5]
rlabel metal3 12124 3864 12124 3864 0 S2MID[6]
rlabel metal3 8596 7000 8596 7000 0 S2MID[7]
rlabel metal2 1652 4536 1652 4536 0 S4END[0]
rlabel metal3 13020 616 13020 616 0 S4END[10]
rlabel metal2 20748 4529 20748 4529 0 S4END[11]
rlabel metal2 20972 6685 20972 6685 0 S4END[12]
rlabel metal2 15988 364 15988 364 0 S4END[13]
rlabel metal2 21420 4977 21420 4977 0 S4END[14]
rlabel metal2 21644 6797 21644 6797 0 S4END[15]
rlabel metal2 18508 5201 18508 5201 0 S4END[1]
rlabel metal2 13580 3220 13580 3220 0 S4END[2]
rlabel metal2 18956 6517 18956 6517 0 S4END[3]
rlabel metal2 7644 3836 7644 3836 0 S4END[4]
rlabel metal2 1148 5488 1148 5488 0 S4END[5]
rlabel metal2 19628 6433 19628 6433 0 S4END[6]
rlabel metal2 19852 6853 19852 6853 0 S4END[7]
rlabel metal3 2730 2828 2730 2828 0 S4END[8]
rlabel metal3 9352 476 9352 476 0 S4END[9]
rlabel metal2 21868 6713 21868 6713 0 SS4END[0]
rlabel metal2 22652 1624 22652 1624 0 SS4END[10]
rlabel metal2 22064 1092 22064 1092 0 SS4END[11]
rlabel metal3 23716 1092 23716 1092 0 SS4END[12]
rlabel metal2 24556 3178 24556 3178 0 SS4END[13]
rlabel metal3 24220 2492 24220 2492 0 SS4END[14]
rlabel metal2 25284 3038 25284 3038 0 SS4END[15]
rlabel metal2 22092 6741 22092 6741 0 SS4END[1]
rlabel metal2 22316 6909 22316 6909 0 SS4END[2]
rlabel metal2 22540 7021 22540 7021 0 SS4END[3]
rlabel metal3 22316 1008 22316 1008 0 SS4END[4]
rlabel metal2 22988 5789 22988 5789 0 SS4END[5]
rlabel metal2 23212 6125 23212 6125 0 SS4END[6]
rlabel metal2 23436 6489 23436 6489 0 SS4END[7]
rlabel metal2 23660 6517 23660 6517 0 SS4END[8]
rlabel metal2 23884 4193 23884 4193 0 SS4END[9]
rlabel metal2 1484 427 1484 427 0 UserCLK
rlabel metal2 25452 6825 25452 6825 0 UserCLKo
rlabel metal2 13580 840 13580 840 0 net1
rlabel metal3 21980 2800 21980 2800 0 net10
rlabel metal3 19768 1036 19768 1036 0 net100
rlabel metal3 18564 1400 18564 1400 0 net101
rlabel metal2 20916 2660 20916 2660 0 net102
rlabel metal2 17612 1036 17612 1036 0 net103
rlabel metal2 20860 3836 20860 3836 0 net104
rlabel metal2 25620 4060 25620 4060 0 net105
rlabel metal2 31164 5068 31164 5068 0 net11
rlabel metal3 24668 448 24668 448 0 net12
rlabel metal3 30492 3332 30492 3332 0 net13
rlabel metal2 6804 5040 6804 5040 0 net14
rlabel metal2 28980 3052 28980 3052 0 net15
rlabel metal4 10444 392 10444 392 0 net16
rlabel metal3 29260 4452 29260 4452 0 net17
rlabel metal2 2772 4676 2772 4676 0 net18
rlabel metal3 29232 4844 29232 4844 0 net19
rlabel metal2 28644 2660 28644 2660 0 net2
rlabel metal2 29596 5264 29596 5264 0 net20
rlabel metal2 29288 4116 29288 4116 0 net21
rlabel metal2 28812 4648 28812 4648 0 net22
rlabel metal2 30100 952 30100 952 0 net23
rlabel metal3 5096 4116 5096 4116 0 net24
rlabel metal2 29596 3990 29596 3990 0 net25
rlabel metal3 29484 1036 29484 1036 0 net26
rlabel metal3 22148 1148 22148 1148 0 net27
rlabel metal3 30464 980 30464 980 0 net28
rlabel metal2 30072 1764 30072 1764 0 net29
rlabel metal2 31108 2408 31108 2408 0 net3
rlabel metal3 30380 1372 30380 1372 0 net30
rlabel metal2 29260 1232 29260 1232 0 net31
rlabel metal2 2884 1876 2884 1876 0 net32
rlabel metal2 22652 5880 22652 5880 0 net33
rlabel metal2 27188 2016 27188 2016 0 net34
rlabel metal2 24108 4788 24108 4788 0 net35
rlabel metal2 25452 2828 25452 2828 0 net36
rlabel metal3 28756 3360 28756 3360 0 net37
rlabel metal2 29036 5320 29036 5320 0 net38
rlabel metal3 25060 1708 25060 1708 0 net39
rlabel metal3 30464 2548 30464 2548 0 net4
rlabel metal3 25312 4060 25312 4060 0 net40
rlabel metal2 30996 6048 30996 6048 0 net41
rlabel metal2 26068 1484 26068 1484 0 net42
rlabel metal3 29120 2212 29120 2212 0 net43
rlabel metal2 26068 6272 26068 6272 0 net44
rlabel metal2 26236 5488 26236 5488 0 net45
rlabel metal3 23744 6076 23744 6076 0 net46
rlabel metal2 27188 6244 27188 6244 0 net47
rlabel metal2 27020 5460 27020 5460 0 net48
rlabel metal3 23380 2884 23380 2884 0 net49
rlabel metal3 23492 4284 23492 4284 0 net5
rlabel metal3 24472 2436 24472 2436 0 net50
rlabel metal2 26684 1988 26684 1988 0 net51
rlabel metal3 26460 1036 26460 1036 0 net52
rlabel metal2 952 2604 952 2604 0 net53
rlabel metal3 3500 2996 3500 2996 0 net54
rlabel metal2 2604 5628 2604 5628 0 net55
rlabel metal2 2296 6468 2296 6468 0 net56
rlabel metal3 4396 5684 4396 5684 0 net57
rlabel metal2 3780 3836 3780 3836 0 net58
rlabel metal2 3276 4536 3276 4536 0 net59
rlabel metal3 29876 3500 29876 3500 0 net6
rlabel metal2 3808 6020 3808 6020 0 net60
rlabel metal3 5516 5068 5516 5068 0 net61
rlabel metal2 4172 5600 4172 5600 0 net62
rlabel metal2 4060 5068 4060 5068 0 net63
rlabel metal2 5348 5208 5348 5208 0 net64
rlabel metal2 26628 4844 26628 4844 0 net65
rlabel metal2 5796 4228 5796 4228 0 net66
rlabel metal4 22540 6188 22540 6188 0 net67
rlabel metal2 20188 5992 20188 5992 0 net68
rlabel metal2 23716 3136 23716 3136 0 net69
rlabel metal3 25452 3724 25452 3724 0 net7
rlabel metal2 5404 5684 5404 5684 0 net70
rlabel metal2 20468 2884 20468 2884 0 net71
rlabel metal2 21756 2996 21756 2996 0 net72
rlabel metal3 12012 896 12012 896 0 net73
rlabel metal2 8652 5460 8652 5460 0 net74
rlabel metal2 9044 4732 9044 4732 0 net75
rlabel metal2 9996 4956 9996 4956 0 net76
rlabel metal3 12096 2996 12096 2996 0 net77
rlabel metal3 12684 3220 12684 3220 0 net78
rlabel metal2 1428 5348 1428 5348 0 net79
rlabel metal3 22596 2660 22596 2660 0 net8
rlabel metal2 7532 4060 7532 4060 0 net80
rlabel metal2 8260 3136 8260 3136 0 net81
rlabel metal2 1008 2212 1008 2212 0 net82
rlabel metal2 1092 4088 1092 4088 0 net83
rlabel metal2 980 1232 980 1232 0 net84
rlabel metal2 924 1428 924 1428 0 net85
rlabel metal2 1036 3136 1036 3136 0 net86
rlabel metal3 8540 3332 8540 3332 0 net87
rlabel metal2 10668 2828 10668 2828 0 net88
rlabel metal2 25004 1848 25004 1848 0 net89
rlabel metal3 30268 2996 30268 2996 0 net9
rlabel metal2 13748 5236 13748 5236 0 net90
rlabel metal3 15820 1036 15820 1036 0 net91
rlabel metal2 18172 1064 18172 1064 0 net92
rlabel metal2 19460 1120 19460 1120 0 net93
rlabel metal2 17668 1092 17668 1092 0 net94
rlabel metal3 14840 6132 14840 6132 0 net95
rlabel metal2 23268 1932 23268 1932 0 net96
rlabel metal4 12684 2184 12684 2184 0 net97
rlabel metal2 22708 1204 22708 1204 0 net98
rlabel metal3 19880 1596 19880 1596 0 net99
<< properties >>
string FIXED_BBOX 0 0 32200 7112
<< end >>
