* NGSPICE file created from S_WARMBOOT.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

.subckt S_WARMBOOT BOOT_top CONFIGURED_top Co FrameData[0] FrameData[10] FrameData[11]
+ FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17]
+ FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22]
+ FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28]
+ FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4]
+ FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13]
+ N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7]
+ N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14]
+ NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7]
+ NN4BEG[8] NN4BEG[9] RESET_top S1END[0] S1END[1] S1END[2] S1END[3] S2END[0] S2END[1]
+ S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2]
+ S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11] S4END[12]
+ S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6]
+ S4END[7] S4END[8] S4END[9] SLOT_top0 SLOT_top1 SLOT_top2 SLOT_top3 SS4END[0] SS4END[10]
+ SS4END[11] SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3]
+ SS4END[4] SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VDD
+ VSS
XTAP_TAPCELL_ROW_9_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_062_ _021_ _023_ _026_ _027_ _011_ net56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_7_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_131_ net7 net64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_200_ net42 net133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_045_ net1 _011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput64 net66 FrameData_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput75 net77 FrameData_O[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput97 net99 FrameStrobe_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput86 net88 FrameData_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_9_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_130_ net4 net63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_061_ _009_ _024_ _010_ _027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_044_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q _010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_113_ net22 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_5_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput87 net89 FrameStrobe_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput98 net100 FrameStrobe_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput76 net78 FrameData_O[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput65 net67 FrameData_O[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput54 net56 BOOT_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_060_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q _025_ _026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ S4END[13] net137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_112_ net21 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_11_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_043_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q _009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput99 net101 FrameStrobe_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput88 net90 FrameStrobe_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput77 net79 FrameData_O[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput55 net57 FrameData_O[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput66 net68 FrameData_O[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_12_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_188_ S4END[14] net136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_12_Left_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_111_ net20 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput89 net91 FrameStrobe_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput67 net69 FrameData_O[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput78 net80 FrameData_O[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput56 net58 FrameData_O[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_15_Left_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_187_ S4END[15] net129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_110_ net19 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_6_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput57 net59 FrameData_O[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput68 net70 FrameData_O[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput79 net81 FrameData_O[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_3_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_186_ net28 net128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_169_ Inst_S_WARMBOOT_switch_matrix.N1BEG2 net111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput69 net71 FrameData_O[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_12_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput58 net60 FrameData_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XS_WARMBOOT_164 Co VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_185_ net29 net127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_099_ net8 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_168_ Inst_S_WARMBOOT_switch_matrix.N1BEG1 net110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput59 net61 FrameData_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_184_ net30 net126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_0_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_167_ Inst_S_WARMBOOT_switch_matrix.N1BEG0 net109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_098_ net7 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_1_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_219_ UserCLK net165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_183_ net31 net125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_0_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_166_ FrameStrobe[19] net99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_097_ net4 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_6_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_218_ net48 net151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_149_ FrameStrobe[2] net101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_182_ net32 net124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_096_ net3 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
X_165_ FrameStrobe[18] net98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_217_ net49 net150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_148_ FrameStrobe[1] net100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_079_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q _041_ _042_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_181_ net33 net123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_164_ FrameStrobe[17] net97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_095_ net2 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_10_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_147_ net6 net89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_216_ net50 net149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_078_ net49 net53 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q _041_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_180_ net34 net122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_163_ FrameStrobe[16] net96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_094_ net27 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q Inst_S_WARMBOOT_switch_matrix.N1BEG0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_215_ net51 net148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_11_Left_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_146_ net22 net81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_077_ net41 net45 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q _040_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_129_ net3 net62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Left_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_093_ net26 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q Inst_S_WARMBOOT_switch_matrix.N1BEG1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_162_ FrameStrobe[15] net95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 CONFIGURED_top net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_145_ net21 net80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_076_ _036_ _037_ _039_ net163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_214_ net52 net147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_059_ net51 net55 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q _025_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_128_ net2 net61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_161_ FrameStrobe[14] net94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_092_ net25 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q Inst_S_WARMBOOT_switch_matrix.N1BEG2
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput2 FrameData[13] net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_213_ net53 net146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_075_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q _038_ _039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_144_ net20 net78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_127_ FrameData[12] net60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_058_ net43 net47 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q _024_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_160_ FrameStrobe[13] net93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_091_ net24 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q Inst_S_WARMBOOT_switch_matrix.N1BEG3
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput3 FrameData[14] net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_212_ net54 net160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_074_ net26 net38 net30 net34 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
+ _038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_143_ net19 net77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_126_ FrameData[11] net59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_057_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q _022_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
+ _023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput50 SS4END[4] net52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_109_ net18 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_10_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_090_ _005_ _006_ _008_ net161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput4 FrameData[15] net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_211_ net55 net159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_142_ net18 net76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_073_ _014_ _034_ _015_ _037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_056_ net31 net35 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q _022_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_125_ FrameData[10] net58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput160 net162 SLOT_top1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_6_Left_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput51 SS4END[5] net53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput40 S4END[2] net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_108_ net17 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTAP_TAPCELL_ROW_13_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_465 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 FrameData[16] net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_141_ net17 net75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_072_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q _035_ _036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_210_ SS4END[8] net158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_124_ FrameData[9] net88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput150 net152 NN4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_055_ _009_ _020_ _021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput161 net163 SLOT_top2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput41 S4END[3] net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput30 S2END[4] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput52 SS4END[6] net54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_107_ net16 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_7_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 FrameData[17] net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_071_ net50 net54 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q _035_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_140_ net16 net74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput140 net142 N4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput151 net153 NN4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput162 net164 SLOT_top3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput31 S2END[5] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_123_ FrameData[8] net87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_054_ net27 net39 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q _020_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput20 FrameData[31] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput42 S4END[4] net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput53 SS4END[7] net55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_106_ net15 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_8_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput7 FrameData[18] net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_070_ net42 net46 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q _034_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_199_ net43 net132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput141 net143 N4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput130 net132 N4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput152 net154 NN4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput163 net165 UserCLKo VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_122_ FrameData[7] net86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_053_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q _019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput43 S4END[5] net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput32 S2END[6] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput10 FrameData[21] net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput21 RESET_top net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_13_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ net14 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_8_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 FrameData[19] net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_1_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_198_ net44 net131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput153 net155 NN4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput131 net133 N4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput142 net144 N4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput120 net122 N2BEGb[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_121_ FrameData[6] net85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_052_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q _018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput33 S2END[7] net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput44 S4END[6] net46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput22 S1END[0] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput11 FrameData[22] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_10_Left_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_104_ net13 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_3_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 FrameData[20] net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_197_ net45 net130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput143 net145 NN4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput132 net134 N4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput121 net123 N2BEGb[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput110 net112 N1BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_120_ FrameData[5] net84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput154 net156 NN4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_051_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q _017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput34 S2MID[0] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput45 S4END[7] net47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput23 S1END[1] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput12 FrameData[23] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_103_ net12 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_8_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net46 net144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput122 net124 N2BEGb[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput155 net157 NN4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput100 net102 FrameStrobe_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput144 net146 NN4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput111 net113 N2BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput133 net135 N4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_050_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q _016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput46 SS4END[0] net48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput35 S2MID[1] net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput24 S1END[2] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_179_ net35 net121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput13 FrameData[24] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_102_ net11 net6 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_15_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_195_ net47 net143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput101 net103 FrameStrobe_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput156 net158 NN4BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput145 net147 NN4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput134 net136 N4BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput123 net125 N2BEGb[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput112 net114 N2BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput36 S2MID[2] net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput25 S1END[3] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput14 FrameData[25] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput47 SS4END[1] net49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_178_ net36 net120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_101_ net10 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_6_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_2_Left_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_194_ S4END[8] net142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput102 net104 FrameStrobe_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput146 net148 NN4BEG[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput124 net126 N2BEGb[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput113 net115 N2BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput157 net159 NN4BEG[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput135 net137 N4BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput48 SS4END[2] net50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput26 S2END[0] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput37 S2MID[3] net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 FrameData[26] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_177_ net37 net119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_100_ net9 net5 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_193_ S4END[9] net141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput147 net149 NN4BEG[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput136 net138 N4BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput103 net105 FrameStrobe_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput125 net127 N2BEGb[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput158 net160 NN4BEG[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput114 net116 N2BEG[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput49 SS4END[3] net51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput38 S4END[0] net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput27 S2END[1] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_176_ net38 net118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput16 FrameData[27] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_159_ FrameStrobe[12] net92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_460 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_192_ S4END[10] net140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput115 net117 N2BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput148 net150 NN4BEG[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput137 net139 N4BEG[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput104 net106 FrameStrobe_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput126 net128 N2BEGb[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput159 net161 SLOT_top0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_11_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput39 S4END[1] net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput28 S2END[2] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_175_ net39 net117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput17 FrameData[28] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_15_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_158_ FrameStrobe[11] net91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_089_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q _007_ _008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_191_ S4END[11] net139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput149 net151 NN4BEG[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput138 net140 N4BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput127 net129 N4BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput105 net107 FrameStrobe_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput116 net118 N2BEG[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput29 S2END[3] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_174_ S2MID[4] net116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 FrameData[29] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_15_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_157_ FrameStrobe[10] net90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_088_ net24 net36 net28 net32 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
+ _007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Left_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_209_ SS4END[9] net157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ S4END[12] net138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput106 net108 FrameStrobe_O[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput139 net141 N4BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput128 net130 N4BEG[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput117 net119 N2BEG[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_173_ S2MID[5] net115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 FrameData[30] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_15_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_087_ _018_ _003_ _019_ _006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_156_ FrameStrobe[9] net108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_208_ SS4END[10] net156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_139_ net15 net73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput118 net120 N2BEG[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput129 net131 N4BEG[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput107 net109 N1BEG[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_15_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_172_ S2MID[6] net114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_086_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q _004_ _005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_155_ FrameStrobe[8] net107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_207_ SS4END[11] net155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_138_ net14 net72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_069_ _030_ _031_ _033_ net164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput90 net92 FrameStrobe_O[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput119 net121 N2BEGb[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput108 net110 N1BEG[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_171_ S2MID[7] net113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_15_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_154_ FrameStrobe[7] net106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_085_ net48 net52 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q _004_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_137_ net13 net71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_206_ SS4END[12] net154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_068_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q _032_ _033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput109 net111 N1BEG[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput91 net93 FrameStrobe_O[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput80 net82 FrameData_O[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_170_ Inst_S_WARMBOOT_switch_matrix.N1BEG3 net112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_153_ FrameStrobe[6] net105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_084_ net40 net44 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q _003_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_205_ SS4END[13] net153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_136_ net12 net70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_13_Left_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_067_ net27 net39 net31 net35 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
+ _032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_119_ FrameData[4] net83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput92 net94 FrameStrobe_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput70 net72 FrameData_O[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput81 net83 FrameData_O[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_152_ FrameStrobe[5] net104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_083_ _042_ _000_ _002_ net162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_8_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Left_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_204_ SS4END[14] net152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_135_ net11 net69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_066_ _012_ _028_ _013_ _031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_049_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q _015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_7_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_118_ FrameData[3] net82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_484 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput93 net95 FrameStrobe_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput71 net73 FrameData_O[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput60 net62 FrameData_O[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput82 net84 FrameData_O[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_151_ FrameStrobe[4] net103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_082_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q _001_ _002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_203_ SS4END[15] net145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_134_ net10 net67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_065_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q _029_ _030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_117_ FrameData[2] net79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_048_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q _014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_1_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput94 net96 FrameStrobe_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_13_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput72 net74 FrameData_O[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput61 net63 FrameData_O[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput83 net85 FrameData_O[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_150_ FrameStrobe[3] net102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_081_ net25 net37 net29 net33 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
+ _001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_064_ net51 net55 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q _029_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_202_ net40 net135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_133_ net9 net66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_116_ FrameData[1] net68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_047_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q _013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xfanout5 FrameStrobe[0] net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput73 net75 FrameData_O[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_9_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput62 net64 FrameData_O[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput95 net97 FrameStrobe_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput84 net86 FrameData_O[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_9_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_080_ _016_ _040_ _017_ _000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_132_ net8 net65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_063_ net43 net47 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q _028_ VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_201_ net41 net134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_115_ FrameData[0] net57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_046_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q _012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_5_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout6 FrameStrobe[0] net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net98 FrameStrobe_O[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput63 net65 FrameData_O[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput74 net76 FrameData_O[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput85 net87 FrameData_O[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
.ends

