module W_IO (A_I_top,
    A_O_top,
    A_T_top,
    B_I_top,
    B_O_top,
    B_T_top,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_IO_switch_matrix.E1BEG0 ;
 wire \Inst_W_IO_switch_matrix.E1BEG1 ;
 wire \Inst_W_IO_switch_matrix.E1BEG2 ;
 wire \Inst_W_IO_switch_matrix.E1BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG0 ;
 wire \Inst_W_IO_switch_matrix.E2BEG1 ;
 wire \Inst_W_IO_switch_matrix.E2BEG2 ;
 wire \Inst_W_IO_switch_matrix.E2BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG4 ;
 wire \Inst_W_IO_switch_matrix.E2BEG5 ;
 wire \Inst_W_IO_switch_matrix.E2BEG6 ;
 wire \Inst_W_IO_switch_matrix.E2BEG7 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb0 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb1 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb2 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb3 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb4 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb5 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb6 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG0 ;
 wire \Inst_W_IO_switch_matrix.E6BEG1 ;
 wire \Inst_W_IO_switch_matrix.E6BEG10 ;
 wire \Inst_W_IO_switch_matrix.E6BEG11 ;
 wire \Inst_W_IO_switch_matrix.E6BEG2 ;
 wire \Inst_W_IO_switch_matrix.E6BEG3 ;
 wire \Inst_W_IO_switch_matrix.E6BEG4 ;
 wire \Inst_W_IO_switch_matrix.E6BEG5 ;
 wire \Inst_W_IO_switch_matrix.E6BEG6 ;
 wire \Inst_W_IO_switch_matrix.E6BEG7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG8 ;
 wire \Inst_W_IO_switch_matrix.E6BEG9 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG0 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG1 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG10 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG11 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG12 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG13 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG14 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG15 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG2 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG3 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG4 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG5 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG6 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG7 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG8 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG9 ;
 wire net204;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net205;
 wire net206;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _042_ (.I(net69),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _043_ (.I(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _044_ (.I(net56),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _045_ (.I(net57),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _046_ (.I(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _047_ (.I(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _048_ (.I(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _049_ (.I0(net56),
    .I1(net57),
    .I2(net58),
    .I3(net59),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _050_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_007_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _051_ (.I0(net60),
    .I1(net61),
    .I2(net62),
    .I3(net63),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _052_ (.A1(_001_),
    .A2(_009_),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _053_ (.I0(net64),
    .I1(net65),
    .I2(net66),
    .I3(net67),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _054_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_011_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _055_ (.I0(net70),
    .I1(net71),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _056_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(net68),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _057_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_000_),
    .B(_014_),
    .C(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _058_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_013_),
    .B(_015_),
    .C(_001_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _059_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_012_),
    .A3(_016_),
    .B1(_008_),
    .B2(_010_),
    .ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _060_ (.I0(net56),
    .I1(net57),
    .I2(net58),
    .I3(net59),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _061_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(_017_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _062_ (.I0(net60),
    .I1(net61),
    .I2(net62),
    .I3(net63),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _063_ (.A1(_004_),
    .A2(_019_),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _064_ (.I0(net64),
    .I1(net65),
    .I2(net66),
    .I3(net67),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _065_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(_021_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _066_ (.I0(net70),
    .I1(net71),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _067_ (.A1(net68),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _068_ (.A1(_000_),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .C(_024_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _069_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_023_),
    .B(_025_),
    .C(_004_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _070_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .A2(_022_),
    .A3(_026_),
    .B1(_018_),
    .B2(_020_),
    .ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _071_ (.I0(net52),
    .I1(net84),
    .I2(net72),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG11 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _072_ (.I0(net53),
    .I1(net91),
    .I2(net75),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG10 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _073_ (.I0(net94),
    .I1(net87),
    .I2(net78),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG9 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _074_ (.I0(net95),
    .I1(net88),
    .I2(net79),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG8 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _075_ (.I0(net52),
    .I1(net98),
    .I2(net82),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _076_ (.I0(net53),
    .I1(net99),
    .I2(net83),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _077_ (.I0(net55),
    .I1(net92),
    .I2(net76),
    .I3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _078_ (.I0(net54),
    .I1(net93),
    .I2(net77),
    .I3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _079_ (.I0(net96),
    .I1(net89),
    .I2(net80),
    .I3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _080_ (.I0(net97),
    .I1(net90),
    .I2(net81),
    .I3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _081_ (.I0(net55),
    .I1(net85),
    .I2(net73),
    .I3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _082_ (.I0(net54),
    .I1(net86),
    .I2(net74),
    .I3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .Z(\Inst_W_IO_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _083_ (.I0(net65),
    .I1(net69),
    .I2(net67),
    .I3(net71),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG15 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _084_ (.I0(net64),
    .I1(net68),
    .I2(net66),
    .I3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG14 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _085_ (.I0(net81),
    .I1(net74),
    .I2(net83),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG13 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _086_ (.I0(net75),
    .I1(net79),
    .I2(net77),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG12 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _087_ (.I0(net80),
    .I1(net73),
    .I2(net82),
    .I3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG11 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _088_ (.I0(net72),
    .I1(net78),
    .I2(net76),
    .I3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG10 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _089_ (.I0(net75),
    .I1(net79),
    .I2(net77),
    .I3(net81),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG9 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _090_ (.I0(net78),
    .I1(net82),
    .I2(net80),
    .I3(net73),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG8 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _091_ (.I0(net65),
    .I1(net69),
    .I2(net67),
    .I3(net71),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _092_ (.I0(net64),
    .I1(net68),
    .I2(net66),
    .I3(net70),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _093_ (.I0(net57),
    .I1(net59),
    .I2(net61),
    .I3(net63),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _094_ (.I0(net56),
    .I1(net58),
    .I2(net60),
    .I3(net62),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _095_ (.I0(net81),
    .I1(net74),
    .I2(net83),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _096_ (.I0(net75),
    .I1(net79),
    .I2(net77),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _097_ (.I0(net80),
    .I1(net73),
    .I2(net82),
    .I3(net2),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _098_ (.I0(net72),
    .I1(net78),
    .I2(net76),
    .I3(net1),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(\Inst_W_IO_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _099_ (.I0(net56),
    .I1(net84),
    .I2(net98),
    .I3(net72),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _100_ (.I0(net57),
    .I1(net91),
    .I2(net99),
    .I3(net75),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _101_ (.I0(net58),
    .I1(net92),
    .I2(net85),
    .I3(net76),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _102_ (.I0(net59),
    .I1(net93),
    .I2(net86),
    .I3(net77),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _103_ (.I0(net60),
    .I1(net94),
    .I2(net87),
    .I3(net78),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _104_ (.I0(net61),
    .I1(net95),
    .I2(net88),
    .I3(net79),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _105_ (.I0(net62),
    .I1(net96),
    .I2(net89),
    .I3(net80),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _106_ (.I0(net63),
    .I1(net97),
    .I2(net90),
    .I3(net81),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEGb0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _107_ (.I0(net64),
    .I1(net84),
    .I2(net98),
    .I3(net72),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _108_ (.I0(net65),
    .I1(net91),
    .I2(net99),
    .I3(net75),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _109_ (.I0(net66),
    .I1(net92),
    .I2(net85),
    .I3(net76),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _110_ (.I0(net67),
    .I1(net93),
    .I2(net86),
    .I3(net77),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _111_ (.I0(net68),
    .I1(net94),
    .I2(net87),
    .I3(net78),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _112_ (.I0(net69),
    .I1(net95),
    .I2(net88),
    .I3(net79),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _113_ (.I0(net70),
    .I1(net96),
    .I2(net89),
    .I3(net80),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _114_ (.I0(net71),
    .I1(net97),
    .I2(net90),
    .I3(net81),
    .S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(\Inst_W_IO_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _115_ (.I0(net52),
    .I1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(\Inst_W_IO_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _116_ (.I0(net53),
    .I1(net2),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .Z(\Inst_W_IO_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _117_ (.I0(net54),
    .I1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(\Inst_W_IO_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _118_ (.I0(net55),
    .I1(net1),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .Z(\Inst_W_IO_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _119_ (.A1(net71),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _120_ (.A1(_003_),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .C(_027_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _121_ (.A1(net59),
    .A2(_005_),
    .A3(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _122_ (.A1(_002_),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A3(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _123_ (.A1(net60),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _124_ (.A1(net58),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _125_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_031_),
    .A3(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _126_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_028_),
    .A3(_029_),
    .B1(_030_),
    .B2(_033_),
    .ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _127_ (.A1(net70),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _128_ (.A1(_002_),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .C(_034_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _129_ (.A1(net61),
    .A2(_006_),
    .A3(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _130_ (.A1(net71),
    .A2(_006_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _131_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _132_ (.A1(net62),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _133_ (.A1(net60),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _134_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_039_),
    .A3(_040_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _135_ (.A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_035_),
    .A3(_036_),
    .B1(_038_),
    .B2(_041_),
    .ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _136_ (.D(net17),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _137_ (.D(net18),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _138_ (.D(net19),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _139_ (.D(net20),
    .E(net51),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _140_ (.D(net21),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _141_ (.D(net22),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _142_ (.D(net23),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _143_ (.D(net24),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _144_ (.D(net26),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _145_ (.D(net42),
    .E(net27),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _146_ (.D(net3),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _147_ (.D(net14),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _148_ (.D(net25),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _149_ (.D(net43),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _150_ (.D(net44),
    .E(net29),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _151_ (.D(net45),
    .E(net29),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _152_ (.D(net46),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _153_ (.D(net47),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _154_ (.D(net48),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _155_ (.D(net49),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _156_ (.D(net4),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _157_ (.D(net5),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _158_ (.D(net6),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _159_ (.D(net7),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _160_ (.D(net8),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _161_ (.D(net9),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _162_ (.D(net10),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _163_ (.D(net11),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _164_ (.D(net12),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _165_ (.D(net13),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _166_ (.D(net15),
    .E(net29),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _167_ (.D(net16),
    .E(net29),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _168_ (.D(net17),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _169_ (.D(net18),
    .E(net30),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _170_ (.D(net19),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _171_ (.D(net20),
    .E(net28),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _172_ (.D(net21),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _173_ (.D(net22),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _174_ (.D(net23),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _175_ (.D(net24),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _176_ (.D(net26),
    .E(net31),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _177_ (.D(net42),
    .E(net50),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _178_ (.D(net3),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _179_ (.D(net14),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _180_ (.D(net25),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _181_ (.D(net43),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _182_ (.D(net44),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _183_ (.D(net45),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _184_ (.D(net46),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _185_ (.D(net47),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _186_ (.D(net48),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _187_ (.D(net49),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _188_ (.D(net4),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _189_ (.D(net5),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _190_ (.D(net6),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _191_ (.D(net7),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _192_ (.D(net8),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _193_ (.D(net9),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _194_ (.D(net10),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _195_ (.D(net11),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _196_ (.D(net12),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _197_ (.D(net13),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _198_ (.D(net15),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _199_ (.D(net16),
    .E(net35),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _200_ (.D(net17),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _201_ (.D(net18),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _202_ (.D(net19),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _203_ (.D(net20),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _204_ (.D(net21),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _205_ (.D(net22),
    .E(net34),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _206_ (.D(net23),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _207_ (.D(net24),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _208_ (.D(net26),
    .E(net33),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _209_ (.D(net42),
    .E(net32),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _210_ (.D(net3),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _211_ (.D(net14),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _212_ (.D(net25),
    .E(net39),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _213_ (.D(net43),
    .E(net39),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _214_ (.D(net44),
    .E(net39),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _215_ (.D(net45),
    .E(net39),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _216_ (.D(net46),
    .E(net41),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _217_ (.D(net47),
    .E(net41),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _218_ (.D(net48),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _219_ (.D(net49),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _220_ (.D(net4),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _221_ (.D(net5),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _222_ (.D(net6),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _223_ (.D(net7),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _224_ (.D(net8),
    .E(net41),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _225_ (.D(net9),
    .E(net41),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _226_ (.D(net10),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _227_ (.D(net11),
    .E(net40),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _228_ (.D(net12),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _229_ (.D(net13),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _230_ (.D(net15),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _231_ (.D(net16),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _232_ (.D(net17),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _233_ (.D(net18),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _234_ (.D(net19),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _235_ (.D(net20),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _236_ (.D(net21),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _237_ (.D(net22),
    .E(net37),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _238_ (.D(net23),
    .E(net38),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _239_ (.D(net24),
    .E(net38),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _240_ (.D(net26),
    .E(net38),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _241_ (.D(net42),
    .E(net38),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _242_ (.D(net1),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _243_ (.D(net2),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _244_ (.I(\Inst_W_IO_switch_matrix.EE4BEG2 ),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _245_ (.I(\Inst_W_IO_switch_matrix.EE4BEG3 ),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _246_ (.I(\Inst_W_IO_switch_matrix.EE4BEG4 ),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _247_ (.I(\Inst_W_IO_switch_matrix.EE4BEG5 ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _248_ (.I(\Inst_W_IO_switch_matrix.EE4BEG6 ),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _249_ (.I(\Inst_W_IO_switch_matrix.EE4BEG7 ),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _250_ (.I(\Inst_W_IO_switch_matrix.EE4BEG8 ),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _251_ (.I(\Inst_W_IO_switch_matrix.EE4BEG9 ),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _252_ (.I(\Inst_W_IO_switch_matrix.EE4BEG10 ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _253_ (.I(\Inst_W_IO_switch_matrix.EE4BEG11 ),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _254_ (.I(\Inst_W_IO_switch_matrix.EE4BEG12 ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _255_ (.I(\Inst_W_IO_switch_matrix.EE4BEG13 ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _256_ (.I(\Inst_W_IO_switch_matrix.EE4BEG14 ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _257_ (.I(\Inst_W_IO_switch_matrix.EE4BEG15 ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _258_ (.I(net3),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _259_ (.I(net14),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _260_ (.I(net25),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _261_ (.I(net43),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _262_ (.I(net44),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _263_ (.I(net45),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _264_ (.I(net46),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _265_ (.I(net47),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _266_ (.I(net48),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _267_ (.I(net49),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _268_ (.I(net4),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _269_ (.I(net5),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _270_ (.I(net6),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _271_ (.I(net7),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _272_ (.I(net8),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _273_ (.I(net9),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _274_ (.I(net10),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _275_ (.I(net11),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _276_ (.I(net12),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _277_ (.I(net13),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _278_ (.I(net15),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _279_ (.I(net16),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _280_ (.I(net17),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _281_ (.I(net18),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _282_ (.I(net19),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _283_ (.I(net20),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _284_ (.I(net21),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _285_ (.I(net22),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _286_ (.I(net23),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _287_ (.I(net24),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _288_ (.I(net26),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _289_ (.I(net42),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _290_ (.I(net41),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _291_ (.I(net36),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _292_ (.I(net50),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _293_ (.I(net27),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _294_ (.I(FrameStrobe[4]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _295_ (.I(FrameStrobe[5]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _296_ (.I(FrameStrobe[6]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _297_ (.I(FrameStrobe[7]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _298_ (.I(FrameStrobe[8]),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _299_ (.I(FrameStrobe[9]),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _300_ (.I(FrameStrobe[10]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _301_ (.I(FrameStrobe[11]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _302_ (.I(FrameStrobe[12]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _303_ (.I(FrameStrobe[13]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _304_ (.I(FrameStrobe[14]),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _305_ (.I(FrameStrobe[15]),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _306_ (.I(FrameStrobe[16]),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _307_ (.I(FrameStrobe[17]),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _308_ (.I(FrameStrobe[18]),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _309_ (.I(FrameStrobe[19]),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _310_ (.I(clknet_1_0__leaf_UserCLK),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _311_ (.I(\Inst_W_IO_switch_matrix.E1BEG0 ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _312_ (.I(\Inst_W_IO_switch_matrix.E1BEG1 ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _313_ (.I(\Inst_W_IO_switch_matrix.E1BEG2 ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _314_ (.I(\Inst_W_IO_switch_matrix.E1BEG3 ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _315_ (.I(\Inst_W_IO_switch_matrix.E2BEG0 ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _316_ (.I(\Inst_W_IO_switch_matrix.E2BEG1 ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _317_ (.I(\Inst_W_IO_switch_matrix.E2BEG2 ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _318_ (.I(\Inst_W_IO_switch_matrix.E2BEG3 ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _319_ (.I(\Inst_W_IO_switch_matrix.E2BEG4 ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _320_ (.I(\Inst_W_IO_switch_matrix.E2BEG5 ),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _321_ (.I(\Inst_W_IO_switch_matrix.E2BEG6 ),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _322_ (.I(\Inst_W_IO_switch_matrix.E2BEG7 ),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _323_ (.I(\Inst_W_IO_switch_matrix.E2BEGb0 ),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _324_ (.I(\Inst_W_IO_switch_matrix.E2BEGb1 ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _325_ (.I(\Inst_W_IO_switch_matrix.E2BEGb2 ),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _326_ (.I(\Inst_W_IO_switch_matrix.E2BEGb3 ),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _327_ (.I(\Inst_W_IO_switch_matrix.E2BEGb4 ),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _328_ (.I(\Inst_W_IO_switch_matrix.E2BEGb5 ),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _329_ (.I(\Inst_W_IO_switch_matrix.E2BEGb6 ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _330_ (.I(\Inst_W_IO_switch_matrix.E2BEGb7 ),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _331_ (.I(\Inst_W_IO_switch_matrix.E6BEG0 ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _332_ (.I(\Inst_W_IO_switch_matrix.E6BEG1 ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _333_ (.I(\Inst_W_IO_switch_matrix.E6BEG2 ),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _334_ (.I(\Inst_W_IO_switch_matrix.E6BEG3 ),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _335_ (.I(\Inst_W_IO_switch_matrix.E6BEG4 ),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _336_ (.I(\Inst_W_IO_switch_matrix.E6BEG5 ),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _337_ (.I(\Inst_W_IO_switch_matrix.E6BEG6 ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _338_ (.I(\Inst_W_IO_switch_matrix.E6BEG7 ),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _339_ (.I(\Inst_W_IO_switch_matrix.E6BEG8 ),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _340_ (.I(\Inst_W_IO_switch_matrix.E6BEG9 ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _341_ (.I(\Inst_W_IO_switch_matrix.E6BEG10 ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _342_ (.I(\Inst_W_IO_switch_matrix.E6BEG11 ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _343_ (.I(\Inst_W_IO_switch_matrix.EE4BEG0 ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _344_ (.I(\Inst_W_IO_switch_matrix.EE4BEG1 ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_362 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout27 (.I(net51),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout28 (.I(net29),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout29 (.I(net30),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout30 (.I(net50),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout31 (.I(net50),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout32 (.I(net36),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout33 (.I(net36),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout34 (.I(net36),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout36 (.I(FrameStrobe[1]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout39 (.I(FrameStrobe[0]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout40 (.I(FrameStrobe[0]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout41 (.I(FrameStrobe[0]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(A_O_top),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(B_O_top),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(FrameData[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(FrameData[10]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(FrameData[11]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(FrameData[12]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(FrameData[13]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(FrameData[14]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(FrameData[15]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(FrameData[16]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(FrameData[17]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(FrameData[18]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(FrameData[19]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(FrameData[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(FrameData[20]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(FrameData[21]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(FrameData[22]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(FrameData[23]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(FrameData[24]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(FrameData[25]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(FrameData[26]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input22 (.I(FrameData[27]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(FrameData[28]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(FrameData[29]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(FrameData[2]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(FrameData[30]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(FrameData[31]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(FrameData[3]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(FrameData[4]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(FrameData[5]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(FrameData[6]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(FrameData[7]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(FrameData[8]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(FrameData[9]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input35 (.I(FrameStrobe[2]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input36 (.I(FrameStrobe[3]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input37 (.I(W1END[0]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input38 (.I(W1END[1]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input39 (.I(W1END[2]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(W1END[3]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input41 (.I(W2END[0]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(W2END[1]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(W2END[2]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input44 (.I(W2END[3]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(W2END[4]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(W2END[5]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(W2END[6]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(W2END[7]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(W2MID[0]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input50 (.I(W2MID[1]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input51 (.I(W2MID[2]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input52 (.I(W2MID[3]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input53 (.I(W2MID[4]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input54 (.I(W2MID[5]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input55 (.I(W2MID[6]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input56 (.I(W2MID[7]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input57 (.I(W6END[0]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input58 (.I(W6END[10]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input59 (.I(W6END[11]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input60 (.I(W6END[1]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input61 (.I(W6END[2]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(W6END[3]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input63 (.I(W6END[4]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input64 (.I(W6END[5]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input65 (.I(W6END[6]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input66 (.I(W6END[7]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input67 (.I(W6END[8]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input68 (.I(W6END[9]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input69 (.I(WW4END[0]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input70 (.I(WW4END[10]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input71 (.I(WW4END[11]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input72 (.I(WW4END[12]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input73 (.I(WW4END[13]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input74 (.I(WW4END[14]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input75 (.I(WW4END[15]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input76 (.I(WW4END[1]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input77 (.I(WW4END[2]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input78 (.I(WW4END[3]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input79 (.I(WW4END[4]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input80 (.I(WW4END[5]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input81 (.I(WW4END[6]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input82 (.I(WW4END[7]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input83 (.I(WW4END[8]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input84 (.I(WW4END[9]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output85 (.I(net100),
    .Z(A_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output86 (.I(net206),
    .Z(A_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output87 (.I(net205),
    .Z(B_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output88 (.I(net103),
    .Z(B_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output89 (.I(net104),
    .Z(E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output90 (.I(net105),
    .Z(E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output91 (.I(net106),
    .Z(E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output92 (.I(net107),
    .Z(E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output93 (.I(net108),
    .Z(E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output94 (.I(net109),
    .Z(E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output95 (.I(net110),
    .Z(E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output96 (.I(net111),
    .Z(E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output97 (.I(net112),
    .Z(E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output98 (.I(net113),
    .Z(E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output99 (.I(net114),
    .Z(E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output100 (.I(net115),
    .Z(E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output101 (.I(net116),
    .Z(E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output102 (.I(net117),
    .Z(E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output103 (.I(net118),
    .Z(E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output104 (.I(net119),
    .Z(E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output105 (.I(net120),
    .Z(E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output106 (.I(net121),
    .Z(E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output107 (.I(net122),
    .Z(E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output108 (.I(net123),
    .Z(E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output109 (.I(net124),
    .Z(E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output110 (.I(net125),
    .Z(E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output111 (.I(net126),
    .Z(E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output112 (.I(net127),
    .Z(E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output113 (.I(net128),
    .Z(E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output114 (.I(net129),
    .Z(E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output115 (.I(net130),
    .Z(E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output116 (.I(net131),
    .Z(E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output117 (.I(net132),
    .Z(E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output118 (.I(net133),
    .Z(E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output119 (.I(net134),
    .Z(E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output120 (.I(net135),
    .Z(E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output121 (.I(net136),
    .Z(EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output122 (.I(net137),
    .Z(EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output123 (.I(net138),
    .Z(EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output124 (.I(net139),
    .Z(EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output125 (.I(net140),
    .Z(EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output126 (.I(net141),
    .Z(EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output127 (.I(net142),
    .Z(EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output128 (.I(net143),
    .Z(EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output129 (.I(net144),
    .Z(EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output130 (.I(net145),
    .Z(EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output131 (.I(net146),
    .Z(EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output132 (.I(net147),
    .Z(EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output133 (.I(net148),
    .Z(EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output134 (.I(net149),
    .Z(EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output135 (.I(net150),
    .Z(EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output136 (.I(net151),
    .Z(EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output137 (.I(net152),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output138 (.I(net153),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output139 (.I(net154),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output140 (.I(net155),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output141 (.I(net156),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output142 (.I(net157),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output143 (.I(net158),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output144 (.I(net159),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output145 (.I(net160),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output146 (.I(net161),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output147 (.I(net162),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output148 (.I(net163),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output149 (.I(net164),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output150 (.I(net165),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output151 (.I(net166),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output152 (.I(net167),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output153 (.I(net168),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output154 (.I(net169),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output155 (.I(net170),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output156 (.I(net171),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output157 (.I(net172),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output158 (.I(net173),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output159 (.I(net174),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output160 (.I(net175),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output161 (.I(net176),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output162 (.I(net177),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output163 (.I(net178),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output164 (.I(net179),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output165 (.I(net180),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output166 (.I(net181),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output167 (.I(net182),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output168 (.I(net183),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output169 (.I(net184),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output170 (.I(net185),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output171 (.I(net186),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output172 (.I(net187),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output173 (.I(net188),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output174 (.I(net189),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output175 (.I(net190),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output176 (.I(net191),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output177 (.I(net192),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output178 (.I(net193),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output179 (.I(net194),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output180 (.I(net195),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output181 (.I(net196),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output182 (.I(net197),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output183 (.I(net198),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output184 (.I(net199),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output185 (.I(net200),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output186 (.I(net201),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output187 (.I(net202),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output188 (.I(net203),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net204),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire190 (.I(net102),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire191 (.I(net101),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_UserCLK (.I(UserCLK),
    .Z(UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK (.I(UserCLK),
    .Z(clknet_0_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK (.I(clknet_0_UserCLK),
    .Z(clknet_1_0__leaf_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK_regs (.I(UserCLK_regs),
    .Z(clknet_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_0__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_1__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_240 ();
endmodule
