VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_single
  CLASS BLOCK ;
  FOREIGN S_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 287.280 BY 71.120 ;
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 70.560 120.400 71.120 ;
    END
  END Co
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 0.560 0.560 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 0.560 22.960 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 0.560 25.200 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 0.560 27.440 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 0.560 29.680 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 0.560 31.920 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 0.560 34.160 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.840 0.560 36.400 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.080 0.560 38.640 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 0.560 40.880 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 0.560 43.120 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2.240 0.560 2.800 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 0.560 45.360 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 0.560 47.600 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.280 0.560 49.840 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 0.560 52.080 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 0.560 54.320 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 0.560 56.560 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 0.560 58.800 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 0.560 61.040 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.720 0.560 63.280 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 0.560 65.520 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 4.480 0.560 5.040 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 0.560 67.760 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 0.560 70.000 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 0.560 7.280 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.960 0.560 9.520 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 0.560 11.760 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 0.560 14.000 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 0.560 16.240 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.920 0.560 18.480 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 0.560 20.720 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 0.000 287.280 0.560 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 22.400 287.280 22.960 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 24.640 287.280 25.200 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 26.880 287.280 27.440 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 29.120 287.280 29.680 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 31.360 287.280 31.920 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 33.600 287.280 34.160 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 35.840 287.280 36.400 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 38.080 287.280 38.640 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 40.320 287.280 40.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 42.560 287.280 43.120 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 2.240 287.280 2.800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 44.800 287.280 45.360 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 47.040 287.280 47.600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 49.280 287.280 49.840 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 51.520 287.280 52.080 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 53.760 287.280 54.320 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 56.000 287.280 56.560 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 58.240 287.280 58.800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 60.480 287.280 61.040 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 62.720 287.280 63.280 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 64.960 287.280 65.520 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 4.480 287.280 5.040 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 67.200 287.280 67.760 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 69.440 287.280 70.000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 6.720 287.280 7.280 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 8.960 287.280 9.520 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 11.200 287.280 11.760 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 13.440 287.280 14.000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 15.680 287.280 16.240 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 17.920 287.280 18.480 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 286.720 20.160 287.280 20.720 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 0.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 0.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 0.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 0.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 0.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 0.560 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 0.000 224.560 0.560 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 0.560 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 0.000 251.440 0.560 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 0.000 264.880 0.560 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 0.560 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 0.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 0.560 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 0.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 0.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 0.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 0.560 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 0.560 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 0.000 130.480 0.560 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 0.560 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 70.560 241.360 71.120 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 70.560 263.760 71.120 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 70.560 266.000 71.120 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 70.560 268.240 71.120 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 70.560 270.480 71.120 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 70.560 272.720 71.120 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 70.560 274.960 71.120 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 70.560 277.200 71.120 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 70.560 279.440 71.120 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 70.560 281.680 71.120 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 70.560 283.920 71.120 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 70.560 243.600 71.120 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 70.560 245.840 71.120 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 70.560 248.080 71.120 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 70.560 250.320 71.120 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 70.560 252.560 71.120 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 70.560 254.800 71.120 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 70.560 257.040 71.120 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 70.560 259.280 71.120 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 70.560 261.520 71.120 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 70.560 3.920 71.120 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 70.560 6.160 71.120 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 70.560 8.400 71.120 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 70.560 10.640 71.120 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 70.560 12.880 71.120 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 70.560 15.120 71.120 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 70.560 17.360 71.120 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 70.560 19.600 71.120 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 70.560 21.840 71.120 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 70.560 24.080 71.120 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 70.560 26.320 71.120 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 70.560 28.560 71.120 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 70.560 30.800 71.120 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 70.560 33.040 71.120 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 70.560 35.280 71.120 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 70.560 37.520 71.120 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 70.560 39.760 71.120 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 70.560 42.000 71.120 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 70.560 44.240 71.120 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 70.560 46.480 71.120 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 70.560 48.720 71.120 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 70.560 71.120 71.120 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 70.560 73.360 71.120 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 70.560 75.600 71.120 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 70.560 77.840 71.120 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 70.560 80.080 71.120 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 70.560 82.320 71.120 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 70.560 50.960 71.120 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 70.560 53.200 71.120 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 70.560 55.440 71.120 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 70.560 57.680 71.120 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 70.560 59.920 71.120 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 70.560 62.160 71.120 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 70.560 64.400 71.120 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 70.560 66.640 71.120 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 70.560 68.880 71.120 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 70.560 84.560 71.120 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 70.560 106.960 71.120 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 70.560 109.200 71.120 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 70.560 111.440 71.120 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 70.560 113.680 71.120 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 70.560 115.920 71.120 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 70.560 118.160 71.120 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 70.560 86.800 71.120 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 70.560 89.040 71.120 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 70.560 91.280 71.120 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 70.560 93.520 71.120 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 70.560 95.760 71.120 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 70.560 98.000 71.120 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 70.560 100.240 71.120 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 70.560 102.480 71.120 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 70.560 104.720 71.120 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 70.560 122.640 71.120 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 70.560 124.880 71.120 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 70.560 127.120 71.120 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 70.560 129.360 71.120 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 70.560 149.520 71.120 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 70.560 151.760 71.120 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 70.560 154.000 71.120 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 70.560 156.240 71.120 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 70.560 158.480 71.120 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 70.560 160.720 71.120 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 70.560 162.960 71.120 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 70.560 165.200 71.120 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 70.560 131.600 71.120 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 70.560 133.840 71.120 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 70.560 136.080 71.120 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 70.560 138.320 71.120 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 70.560 140.560 71.120 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 70.560 142.800 71.120 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 70.560 145.040 71.120 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 70.560 147.280 71.120 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 70.560 167.440 71.120 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 70.560 189.840 71.120 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 70.560 192.080 71.120 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 70.560 194.320 71.120 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 70.560 196.560 71.120 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 70.560 198.800 71.120 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 70.560 201.040 71.120 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 70.560 169.680 71.120 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 70.560 171.920 71.120 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 70.560 174.160 71.120 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 70.560 176.400 71.120 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 70.560 178.640 71.120 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 70.560 180.880 71.120 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 70.560 183.120 71.120 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 70.560 185.360 71.120 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 70.560 187.600 71.120 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 70.560 203.280 71.120 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 70.560 225.680 71.120 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 70.560 227.920 71.120 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 70.560 230.160 71.120 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 70.560 232.400 71.120 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 70.560 234.640 71.120 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 70.560 236.880 71.120 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 70.560 205.520 71.120 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 70.560 207.760 71.120 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 70.560 210.000 71.120 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 70.560 212.240 71.120 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 70.560 214.480 71.120 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 70.560 216.720 71.120 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 70.560 218.960 71.120 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 70.560 221.200 71.120 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 70.560 223.440 71.120 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 0.000 9.520 0.560 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 70.560 239.120 71.120 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 0.000 20.480 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.880 0.000 120.480 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.880 0.000 220.480 71.120 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 0.000 23.780 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.180 0.000 123.780 71.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 222.180 0.000 223.780 71.120 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 284.350 67.070 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 283.920 66.940 ;
      LAYER Metal2 ;
        RECT 0.700 70.260 3.060 70.560 ;
        RECT 4.220 70.260 5.300 70.560 ;
        RECT 6.460 70.260 7.540 70.560 ;
        RECT 8.700 70.260 9.780 70.560 ;
        RECT 10.940 70.260 12.020 70.560 ;
        RECT 13.180 70.260 14.260 70.560 ;
        RECT 15.420 70.260 16.500 70.560 ;
        RECT 17.660 70.260 18.740 70.560 ;
        RECT 19.900 70.260 20.980 70.560 ;
        RECT 22.140 70.260 23.220 70.560 ;
        RECT 24.380 70.260 25.460 70.560 ;
        RECT 26.620 70.260 27.700 70.560 ;
        RECT 28.860 70.260 29.940 70.560 ;
        RECT 31.100 70.260 32.180 70.560 ;
        RECT 33.340 70.260 34.420 70.560 ;
        RECT 35.580 70.260 36.660 70.560 ;
        RECT 37.820 70.260 38.900 70.560 ;
        RECT 40.060 70.260 41.140 70.560 ;
        RECT 42.300 70.260 43.380 70.560 ;
        RECT 44.540 70.260 45.620 70.560 ;
        RECT 46.780 70.260 47.860 70.560 ;
        RECT 49.020 70.260 50.100 70.560 ;
        RECT 51.260 70.260 52.340 70.560 ;
        RECT 53.500 70.260 54.580 70.560 ;
        RECT 55.740 70.260 56.820 70.560 ;
        RECT 57.980 70.260 59.060 70.560 ;
        RECT 60.220 70.260 61.300 70.560 ;
        RECT 62.460 70.260 63.540 70.560 ;
        RECT 64.700 70.260 65.780 70.560 ;
        RECT 66.940 70.260 68.020 70.560 ;
        RECT 69.180 70.260 70.260 70.560 ;
        RECT 71.420 70.260 72.500 70.560 ;
        RECT 73.660 70.260 74.740 70.560 ;
        RECT 75.900 70.260 76.980 70.560 ;
        RECT 78.140 70.260 79.220 70.560 ;
        RECT 80.380 70.260 81.460 70.560 ;
        RECT 82.620 70.260 83.700 70.560 ;
        RECT 84.860 70.260 85.940 70.560 ;
        RECT 87.100 70.260 88.180 70.560 ;
        RECT 89.340 70.260 90.420 70.560 ;
        RECT 91.580 70.260 92.660 70.560 ;
        RECT 93.820 70.260 94.900 70.560 ;
        RECT 96.060 70.260 97.140 70.560 ;
        RECT 98.300 70.260 99.380 70.560 ;
        RECT 100.540 70.260 101.620 70.560 ;
        RECT 102.780 70.260 103.860 70.560 ;
        RECT 105.020 70.260 106.100 70.560 ;
        RECT 107.260 70.260 108.340 70.560 ;
        RECT 109.500 70.260 110.580 70.560 ;
        RECT 111.740 70.260 112.820 70.560 ;
        RECT 113.980 70.260 115.060 70.560 ;
        RECT 116.220 70.260 117.300 70.560 ;
        RECT 118.460 70.260 119.540 70.560 ;
        RECT 120.700 70.260 121.780 70.560 ;
        RECT 122.940 70.260 124.020 70.560 ;
        RECT 125.180 70.260 126.260 70.560 ;
        RECT 127.420 70.260 128.500 70.560 ;
        RECT 129.660 70.260 130.740 70.560 ;
        RECT 131.900 70.260 132.980 70.560 ;
        RECT 134.140 70.260 135.220 70.560 ;
        RECT 136.380 70.260 137.460 70.560 ;
        RECT 138.620 70.260 139.700 70.560 ;
        RECT 140.860 70.260 141.940 70.560 ;
        RECT 143.100 70.260 144.180 70.560 ;
        RECT 145.340 70.260 146.420 70.560 ;
        RECT 147.580 70.260 148.660 70.560 ;
        RECT 149.820 70.260 150.900 70.560 ;
        RECT 152.060 70.260 153.140 70.560 ;
        RECT 154.300 70.260 155.380 70.560 ;
        RECT 156.540 70.260 157.620 70.560 ;
        RECT 158.780 70.260 159.860 70.560 ;
        RECT 161.020 70.260 162.100 70.560 ;
        RECT 163.260 70.260 164.340 70.560 ;
        RECT 165.500 70.260 166.580 70.560 ;
        RECT 167.740 70.260 168.820 70.560 ;
        RECT 169.980 70.260 171.060 70.560 ;
        RECT 172.220 70.260 173.300 70.560 ;
        RECT 174.460 70.260 175.540 70.560 ;
        RECT 176.700 70.260 177.780 70.560 ;
        RECT 178.940 70.260 180.020 70.560 ;
        RECT 181.180 70.260 182.260 70.560 ;
        RECT 183.420 70.260 184.500 70.560 ;
        RECT 185.660 70.260 186.740 70.560 ;
        RECT 187.900 70.260 188.980 70.560 ;
        RECT 190.140 70.260 191.220 70.560 ;
        RECT 192.380 70.260 193.460 70.560 ;
        RECT 194.620 70.260 195.700 70.560 ;
        RECT 196.860 70.260 197.940 70.560 ;
        RECT 199.100 70.260 200.180 70.560 ;
        RECT 201.340 70.260 202.420 70.560 ;
        RECT 203.580 70.260 204.660 70.560 ;
        RECT 205.820 70.260 206.900 70.560 ;
        RECT 208.060 70.260 209.140 70.560 ;
        RECT 210.300 70.260 211.380 70.560 ;
        RECT 212.540 70.260 213.620 70.560 ;
        RECT 214.780 70.260 215.860 70.560 ;
        RECT 217.020 70.260 218.100 70.560 ;
        RECT 219.260 70.260 220.340 70.560 ;
        RECT 221.500 70.260 222.580 70.560 ;
        RECT 223.740 70.260 224.820 70.560 ;
        RECT 225.980 70.260 227.060 70.560 ;
        RECT 228.220 70.260 229.300 70.560 ;
        RECT 230.460 70.260 231.540 70.560 ;
        RECT 232.700 70.260 233.780 70.560 ;
        RECT 234.940 70.260 236.020 70.560 ;
        RECT 237.180 70.260 238.260 70.560 ;
        RECT 239.420 70.260 240.500 70.560 ;
        RECT 241.660 70.260 242.740 70.560 ;
        RECT 243.900 70.260 244.980 70.560 ;
        RECT 246.140 70.260 247.220 70.560 ;
        RECT 248.380 70.260 249.460 70.560 ;
        RECT 250.620 70.260 251.700 70.560 ;
        RECT 252.860 70.260 253.940 70.560 ;
        RECT 255.100 70.260 256.180 70.560 ;
        RECT 257.340 70.260 258.420 70.560 ;
        RECT 259.580 70.260 260.660 70.560 ;
        RECT 261.820 70.260 262.900 70.560 ;
        RECT 264.060 70.260 265.140 70.560 ;
        RECT 266.300 70.260 267.380 70.560 ;
        RECT 268.540 70.260 269.620 70.560 ;
        RECT 270.780 70.260 271.860 70.560 ;
        RECT 273.020 70.260 274.100 70.560 ;
        RECT 275.260 70.260 276.340 70.560 ;
        RECT 277.500 70.260 278.580 70.560 ;
        RECT 279.740 70.260 280.820 70.560 ;
        RECT 281.980 70.260 283.060 70.560 ;
        RECT 284.220 70.260 286.580 70.560 ;
        RECT 0.700 0.860 286.580 70.260 ;
        RECT 0.700 0.090 8.660 0.860 ;
        RECT 9.820 0.090 22.100 0.860 ;
        RECT 23.260 0.090 35.540 0.860 ;
        RECT 36.700 0.090 48.980 0.860 ;
        RECT 50.140 0.090 62.420 0.860 ;
        RECT 63.580 0.090 75.860 0.860 ;
        RECT 77.020 0.090 89.300 0.860 ;
        RECT 90.460 0.090 102.740 0.860 ;
        RECT 103.900 0.090 116.180 0.860 ;
        RECT 117.340 0.090 129.620 0.860 ;
        RECT 130.780 0.090 143.060 0.860 ;
        RECT 144.220 0.090 156.500 0.860 ;
        RECT 157.660 0.090 169.940 0.860 ;
        RECT 171.100 0.090 183.380 0.860 ;
        RECT 184.540 0.090 196.820 0.860 ;
        RECT 197.980 0.090 210.260 0.860 ;
        RECT 211.420 0.090 223.700 0.860 ;
        RECT 224.860 0.090 237.140 0.860 ;
        RECT 238.300 0.090 250.580 0.860 ;
        RECT 251.740 0.090 264.020 0.860 ;
        RECT 265.180 0.090 277.460 0.860 ;
        RECT 278.620 0.090 286.580 0.860 ;
      LAYER Metal3 ;
        RECT 0.560 70.300 286.720 70.980 ;
        RECT 0.860 69.140 286.420 70.300 ;
        RECT 0.560 68.060 286.720 69.140 ;
        RECT 0.860 66.900 286.420 68.060 ;
        RECT 0.560 65.820 286.720 66.900 ;
        RECT 0.860 64.660 286.420 65.820 ;
        RECT 0.560 63.580 286.720 64.660 ;
        RECT 0.860 62.420 286.420 63.580 ;
        RECT 0.560 61.340 286.720 62.420 ;
        RECT 0.860 60.180 286.420 61.340 ;
        RECT 0.560 59.100 286.720 60.180 ;
        RECT 0.860 57.940 286.420 59.100 ;
        RECT 0.560 56.860 286.720 57.940 ;
        RECT 0.860 55.700 286.420 56.860 ;
        RECT 0.560 54.620 286.720 55.700 ;
        RECT 0.860 53.460 286.420 54.620 ;
        RECT 0.560 52.380 286.720 53.460 ;
        RECT 0.860 51.220 286.420 52.380 ;
        RECT 0.560 50.140 286.720 51.220 ;
        RECT 0.860 48.980 286.420 50.140 ;
        RECT 0.560 47.900 286.720 48.980 ;
        RECT 0.860 46.740 286.420 47.900 ;
        RECT 0.560 45.660 286.720 46.740 ;
        RECT 0.860 44.500 286.420 45.660 ;
        RECT 0.560 43.420 286.720 44.500 ;
        RECT 0.860 42.260 286.420 43.420 ;
        RECT 0.560 41.180 286.720 42.260 ;
        RECT 0.860 40.020 286.420 41.180 ;
        RECT 0.560 38.940 286.720 40.020 ;
        RECT 0.860 37.780 286.420 38.940 ;
        RECT 0.560 36.700 286.720 37.780 ;
        RECT 0.860 35.540 286.420 36.700 ;
        RECT 0.560 34.460 286.720 35.540 ;
        RECT 0.860 33.300 286.420 34.460 ;
        RECT 0.560 32.220 286.720 33.300 ;
        RECT 0.860 31.060 286.420 32.220 ;
        RECT 0.560 29.980 286.720 31.060 ;
        RECT 0.860 28.820 286.420 29.980 ;
        RECT 0.560 27.740 286.720 28.820 ;
        RECT 0.860 26.580 286.420 27.740 ;
        RECT 0.560 25.500 286.720 26.580 ;
        RECT 0.860 24.340 286.420 25.500 ;
        RECT 0.560 23.260 286.720 24.340 ;
        RECT 0.860 22.100 286.420 23.260 ;
        RECT 0.560 21.020 286.720 22.100 ;
        RECT 0.860 19.860 286.420 21.020 ;
        RECT 0.560 18.780 286.720 19.860 ;
        RECT 0.860 17.620 286.420 18.780 ;
        RECT 0.560 16.540 286.720 17.620 ;
        RECT 0.860 15.380 286.420 16.540 ;
        RECT 0.560 14.300 286.720 15.380 ;
        RECT 0.860 13.140 286.420 14.300 ;
        RECT 0.560 12.060 286.720 13.140 ;
        RECT 0.860 10.900 286.420 12.060 ;
        RECT 0.560 9.820 286.720 10.900 ;
        RECT 0.860 8.660 286.420 9.820 ;
        RECT 0.560 7.580 286.720 8.660 ;
        RECT 0.860 6.420 286.420 7.580 ;
        RECT 0.560 5.340 286.720 6.420 ;
        RECT 0.860 4.180 286.420 5.340 ;
        RECT 0.560 3.100 286.720 4.180 ;
        RECT 0.860 1.940 286.420 3.100 ;
        RECT 0.560 0.860 286.720 1.940 ;
        RECT 0.860 0.140 286.420 0.860 ;
      LAYER Metal4 ;
        RECT 11.340 0.090 18.580 71.030 ;
        RECT 20.780 0.090 21.880 71.030 ;
        RECT 24.080 0.090 118.580 71.030 ;
        RECT 120.780 0.090 121.880 71.030 ;
        RECT 124.080 0.090 218.580 71.030 ;
        RECT 220.780 0.090 221.880 71.030 ;
        RECT 224.080 0.090 244.580 71.030 ;
  END
END S_term_single
END LIBRARY

