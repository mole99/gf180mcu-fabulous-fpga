magic
tech gf180mcuD
magscale 1 10
timestamp 1764323307
<< metal1 >>
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 2158 13186 2210 13198
rect 2158 13122 2210 13134
rect 3726 13186 3778 13198
rect 3726 13122 3778 13134
rect 5966 13186 6018 13198
rect 5966 13122 6018 13134
rect 7534 13186 7586 13198
rect 7534 13122 7586 13134
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 21198 13186 21250 13198
rect 21198 13122 21250 13134
rect 22654 13186 22706 13198
rect 22654 13122 22706 13134
rect 25454 13186 25506 13198
rect 25454 13122 25506 13134
rect 48974 13186 49026 13198
rect 48974 13122 49026 13134
rect 51102 13186 51154 13198
rect 51102 13122 51154 13134
rect 54910 13186 54962 13198
rect 54910 13122 54962 13134
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 17490 13022 17502 13074
rect 17554 13022 17566 13074
rect 52882 13022 52894 13074
rect 52946 13022 52958 13074
rect 2594 12910 2606 12962
rect 2658 12910 2670 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 6514 12910 6526 12962
rect 6578 12910 6590 12962
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 12898 12910 12910 12962
rect 12962 12910 12974 12962
rect 15586 12910 15598 12962
rect 15650 12910 15662 12962
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 18274 12910 18286 12962
rect 18338 12910 18350 12962
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 25106 12910 25118 12962
rect 25170 12910 25182 12962
rect 44930 12910 44942 12962
rect 44994 12910 45006 12962
rect 46834 12910 46846 12962
rect 46898 12910 46910 12962
rect 48402 12910 48414 12962
rect 48466 12910 48478 12962
rect 50530 12910 50542 12962
rect 50594 12910 50606 12962
rect 52322 12910 52334 12962
rect 52386 12910 52398 12962
rect 54338 12910 54350 12962
rect 54402 12910 54414 12962
rect 13918 12850 13970 12862
rect 13918 12786 13970 12798
rect 19294 12850 19346 12862
rect 19294 12786 19346 12798
rect 24110 12850 24162 12862
rect 24110 12786 24162 12798
rect 45950 12850 46002 12862
rect 45950 12786 46002 12798
rect 47854 12850 47906 12862
rect 47854 12786 47906 12798
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 2270 12402 2322 12414
rect 2270 12338 2322 12350
rect 6974 12402 7026 12414
rect 6974 12338 7026 12350
rect 8542 12402 8594 12414
rect 8542 12338 8594 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 22318 12402 22370 12414
rect 22318 12338 22370 12350
rect 23886 12402 23938 12414
rect 23886 12338 23938 12350
rect 49422 12402 49474 12414
rect 49422 12338 49474 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 54126 12402 54178 12414
rect 54126 12338 54178 12350
rect 55694 12402 55746 12414
rect 55694 12338 55746 12350
rect 5406 12290 5458 12302
rect 27918 12290 27970 12302
rect 3602 12238 3614 12290
rect 3666 12238 3678 12290
rect 18162 12238 18174 12290
rect 18226 12238 18238 12290
rect 19506 12238 19518 12290
rect 19570 12238 19582 12290
rect 21074 12238 21086 12290
rect 21138 12238 21150 12290
rect 28578 12238 28590 12290
rect 28642 12238 28654 12290
rect 38098 12238 38110 12290
rect 38162 12238 38174 12290
rect 5406 12226 5458 12238
rect 27918 12226 27970 12238
rect 20638 12178 20690 12190
rect 36878 12178 36930 12190
rect 2706 12126 2718 12178
rect 2770 12126 2782 12178
rect 5842 12126 5854 12178
rect 5906 12126 5918 12178
rect 18834 12126 18846 12178
rect 18898 12126 18910 12178
rect 21970 12126 21982 12178
rect 22034 12126 22046 12178
rect 23314 12126 23326 12178
rect 23378 12126 23390 12178
rect 20638 12114 20690 12126
rect 36878 12114 36930 12126
rect 44718 12178 44770 12190
rect 44718 12114 44770 12126
rect 46398 12178 46450 12190
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 46398 12114 46450 12126
rect 12798 12066 12850 12078
rect 29038 12066 29090 12078
rect 4386 12014 4398 12066
rect 4450 12014 4462 12066
rect 7522 12014 7534 12066
rect 7586 12014 7598 12066
rect 9090 12014 9102 12066
rect 9154 12014 9166 12066
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 12226 12014 12238 12066
rect 12290 12014 12302 12066
rect 15362 12014 15374 12066
rect 15426 12014 15438 12066
rect 15698 12014 15710 12066
rect 15762 12014 15774 12066
rect 17266 12014 17278 12066
rect 17330 12014 17342 12066
rect 12798 12002 12850 12014
rect 29038 12002 29090 12014
rect 36318 12066 36370 12078
rect 36318 12002 36370 12014
rect 45278 12066 45330 12078
rect 45278 12002 45330 12014
rect 46958 12066 47010 12078
rect 50990 12066 51042 12078
rect 48514 12014 48526 12066
rect 48578 12014 48590 12066
rect 48850 12014 48862 12066
rect 48914 12014 48926 12066
rect 53554 12014 53566 12066
rect 53618 12014 53630 12066
rect 55122 12014 55134 12066
rect 55186 12014 55198 12066
rect 46958 12002 47010 12014
rect 50990 12002 51042 12014
rect 13358 11954 13410 11966
rect 13358 11890 13410 11902
rect 27358 11954 27410 11966
rect 27358 11890 27410 11902
rect 37662 11954 37714 11966
rect 37662 11890 37714 11902
rect 47966 11954 48018 11966
rect 47966 11890 48018 11902
rect 50430 11954 50482 11966
rect 50430 11890 50482 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 4622 11618 4674 11630
rect 4622 11554 4674 11566
rect 6190 11618 6242 11630
rect 6190 11554 6242 11566
rect 7758 11618 7810 11630
rect 7758 11554 7810 11566
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 13918 11618 13970 11630
rect 13918 11554 13970 11566
rect 15486 11618 15538 11630
rect 15486 11554 15538 11566
rect 17390 11618 17442 11630
rect 17390 11554 17442 11566
rect 20526 11618 20578 11630
rect 20526 11554 20578 11566
rect 30942 11618 30994 11630
rect 30942 11554 30994 11566
rect 47182 11618 47234 11630
rect 50318 11618 50370 11630
rect 47506 11566 47518 11618
rect 47570 11566 47582 11618
rect 47182 11554 47234 11566
rect 50318 11554 50370 11566
rect 51886 11618 51938 11630
rect 51886 11554 51938 11566
rect 53454 11618 53506 11630
rect 53454 11554 53506 11566
rect 25118 11506 25170 11518
rect 2818 11454 2830 11506
rect 2882 11454 2894 11506
rect 8306 11454 8318 11506
rect 8370 11454 8382 11506
rect 25118 11442 25170 11454
rect 24558 11394 24610 11406
rect 1922 11342 1934 11394
rect 1986 11342 1998 11394
rect 3602 11342 3614 11394
rect 3666 11342 3678 11394
rect 5170 11342 5182 11394
rect 5234 11342 5246 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 13010 11342 13022 11394
rect 13074 11342 13086 11394
rect 13570 11342 13582 11394
rect 13634 11342 13646 11394
rect 14914 11342 14926 11394
rect 14978 11342 14990 11394
rect 16818 11342 16830 11394
rect 16882 11342 16894 11394
rect 18610 11342 18622 11394
rect 18674 11342 18686 11394
rect 19954 11342 19966 11394
rect 20018 11342 20030 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 24558 11330 24610 11342
rect 34414 11394 34466 11406
rect 54462 11394 54514 11406
rect 48290 11342 48302 11394
rect 48354 11342 48366 11394
rect 49746 11342 49758 11394
rect 49810 11342 49822 11394
rect 51314 11342 51326 11394
rect 51378 11342 51390 11394
rect 52882 11342 52894 11394
rect 52946 11342 52958 11394
rect 34414 11330 34466 11342
rect 54462 11330 54514 11342
rect 21758 11282 21810 11294
rect 34974 11282 35026 11294
rect 1586 11230 1598 11282
rect 1650 11230 1662 11282
rect 12338 11230 12350 11282
rect 12402 11230 12414 11282
rect 19058 11230 19070 11282
rect 19122 11230 19134 11282
rect 31378 11230 31390 11282
rect 31442 11230 31454 11282
rect 21758 11218 21810 11230
rect 34974 11218 35026 11230
rect 49198 11282 49250 11294
rect 49198 11218 49250 11230
rect 55022 11282 55074 11294
rect 55022 11218 55074 11230
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 3390 10834 3442 10846
rect 3390 10770 3442 10782
rect 7422 10834 7474 10846
rect 7422 10770 7474 10782
rect 8990 10834 9042 10846
rect 8990 10770 9042 10782
rect 10558 10834 10610 10846
rect 10558 10770 10610 10782
rect 13022 10834 13074 10846
rect 13022 10770 13074 10782
rect 14590 10834 14642 10846
rect 14590 10770 14642 10782
rect 18510 10834 18562 10846
rect 18510 10770 18562 10782
rect 49646 10834 49698 10846
rect 49646 10770 49698 10782
rect 51214 10834 51266 10846
rect 51214 10770 51266 10782
rect 52558 10834 52610 10846
rect 52558 10770 52610 10782
rect 48190 10722 48242 10734
rect 2146 10670 2158 10722
rect 2210 10670 2222 10722
rect 6066 10670 6078 10722
rect 6130 10670 6142 10722
rect 16930 10670 16942 10722
rect 16994 10670 17006 10722
rect 19618 10670 19630 10722
rect 19682 10670 19694 10722
rect 21858 10670 21870 10722
rect 21922 10670 21934 10722
rect 48190 10658 48242 10670
rect 54574 10722 54626 10734
rect 54574 10658 54626 10670
rect 56142 10722 56194 10734
rect 56142 10658 56194 10670
rect 41358 10610 41410 10622
rect 4386 10558 4398 10610
rect 4450 10558 4462 10610
rect 8194 10558 8206 10610
rect 8258 10558 8270 10610
rect 21074 10558 21086 10610
rect 21138 10558 21150 10610
rect 41358 10546 41410 10558
rect 42254 10610 42306 10622
rect 42254 10546 42306 10558
rect 42814 10610 42866 10622
rect 42814 10546 42866 10558
rect 47630 10610 47682 10622
rect 48850 10558 48862 10610
rect 48914 10558 48926 10610
rect 52098 10558 52110 10610
rect 52162 10558 52174 10610
rect 55346 10558 55358 10610
rect 55410 10558 55422 10610
rect 47630 10546 47682 10558
rect 36990 10498 37042 10510
rect 2818 10446 2830 10498
rect 2882 10446 2894 10498
rect 6850 10446 6862 10498
rect 6914 10446 6926 10498
rect 9986 10446 9998 10498
rect 10050 10446 10062 10498
rect 11554 10446 11566 10498
rect 11618 10446 11630 10498
rect 14018 10446 14030 10498
rect 14082 10446 14094 10498
rect 15586 10446 15598 10498
rect 15650 10446 15662 10498
rect 16146 10446 16158 10498
rect 16210 10446 16222 10498
rect 17938 10446 17950 10498
rect 18002 10446 18014 10498
rect 36990 10434 37042 10446
rect 41918 10498 41970 10510
rect 50194 10446 50206 10498
rect 50258 10446 50270 10498
rect 53554 10446 53566 10498
rect 53618 10446 53630 10498
rect 41918 10434 41970 10446
rect 20078 10386 20130 10398
rect 20078 10322 20130 10334
rect 37550 10386 37602 10398
rect 37550 10322 37602 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 17390 10050 17442 10062
rect 17390 9986 17442 9998
rect 26126 10050 26178 10062
rect 26126 9986 26178 9998
rect 9438 9938 9490 9950
rect 1474 9886 1486 9938
rect 1538 9886 1550 9938
rect 5282 9886 5294 9938
rect 5346 9886 5358 9938
rect 9438 9874 9490 9886
rect 16830 9938 16882 9950
rect 16830 9874 16882 9886
rect 23438 9938 23490 9950
rect 23438 9874 23490 9886
rect 23998 9938 24050 9950
rect 23998 9874 24050 9886
rect 25566 9938 25618 9950
rect 25566 9874 25618 9886
rect 36654 9938 36706 9950
rect 36654 9874 36706 9886
rect 6302 9826 6354 9838
rect 1250 9774 1262 9826
rect 1314 9774 1326 9826
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 6302 9762 6354 9774
rect 9998 9826 10050 9838
rect 9998 9762 10050 9774
rect 10894 9826 10946 9838
rect 10894 9762 10946 9774
rect 20862 9826 20914 9838
rect 20862 9762 20914 9774
rect 36094 9826 36146 9838
rect 36094 9762 36146 9774
rect 41470 9826 41522 9838
rect 41470 9762 41522 9774
rect 42590 9826 42642 9838
rect 48526 9826 48578 9838
rect 44706 9774 44718 9826
rect 44770 9774 44782 9826
rect 49634 9774 49646 9826
rect 49698 9774 49710 9826
rect 50194 9774 50206 9826
rect 50258 9774 50270 9826
rect 51090 9774 51102 9826
rect 51154 9774 51166 9826
rect 52546 9774 52558 9826
rect 52610 9774 52622 9826
rect 54226 9774 54238 9826
rect 54290 9774 54302 9826
rect 42590 9762 42642 9774
rect 48526 9762 48578 9774
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 4286 9714 4338 9726
rect 20302 9714 20354 9726
rect 43150 9714 43202 9726
rect 5842 9662 5854 9714
rect 5906 9662 5918 9714
rect 10434 9662 10446 9714
rect 10498 9662 10510 9714
rect 41906 9662 41918 9714
rect 41970 9662 41982 9714
rect 4286 9650 4338 9662
rect 20302 9650 20354 9662
rect 43150 9650 43202 9662
rect 45166 9714 45218 9726
rect 45166 9650 45218 9662
rect 49086 9714 49138 9726
rect 49086 9650 49138 9662
rect 51998 9714 52050 9726
rect 51998 9650 52050 9662
rect 53566 9714 53618 9726
rect 53566 9650 53618 9662
rect 55134 9602 55186 9614
rect 55134 9538 55186 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 51214 9266 51266 9278
rect 51214 9202 51266 9214
rect 53006 9266 53058 9278
rect 53006 9202 53058 9214
rect 2942 9154 2994 9166
rect 1698 9102 1710 9154
rect 1762 9102 1774 9154
rect 2942 9090 2994 9102
rect 5966 9154 6018 9166
rect 5966 9090 6018 9102
rect 3502 9042 3554 9054
rect 49746 8990 49758 9042
rect 49810 8990 49822 9042
rect 52098 8990 52110 9042
rect 52162 8990 52174 9042
rect 55234 8990 55246 9042
rect 55298 8990 55310 9042
rect 3502 8978 3554 8990
rect 10334 8930 10386 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 10334 8866 10386 8878
rect 22430 8930 22482 8942
rect 22430 8866 22482 8878
rect 47630 8930 47682 8942
rect 47630 8866 47682 8878
rect 49310 8930 49362 8942
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 55906 8878 55918 8930
rect 55970 8878 55982 8930
rect 49310 8866 49362 8878
rect 6526 8818 6578 8830
rect 6526 8754 6578 8766
rect 10894 8818 10946 8830
rect 10894 8754 10946 8766
rect 22990 8818 23042 8830
rect 22990 8754 23042 8766
rect 47070 8818 47122 8830
rect 47070 8754 47122 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 20526 8482 20578 8494
rect 20526 8418 20578 8430
rect 34638 8482 34690 8494
rect 34638 8418 34690 8430
rect 53330 8318 53342 8370
rect 53394 8318 53406 8370
rect 9438 8258 9490 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 5842 8206 5854 8258
rect 5906 8206 5918 8258
rect 9438 8194 9490 8206
rect 21534 8258 21586 8270
rect 21534 8194 21586 8206
rect 22094 8258 22146 8270
rect 48414 8258 48466 8270
rect 40338 8206 40350 8258
rect 40402 8206 40414 8258
rect 22094 8194 22146 8206
rect 48414 8194 48466 8206
rect 48974 8258 49026 8270
rect 48974 8194 49026 8206
rect 50094 8258 50146 8270
rect 50978 8206 50990 8258
rect 51042 8206 51054 8258
rect 52546 8206 52558 8258
rect 52610 8206 52622 8258
rect 54114 8206 54126 8258
rect 54178 8206 54190 8258
rect 50094 8194 50146 8206
rect 6302 8146 6354 8158
rect 19966 8146 20018 8158
rect 55134 8146 55186 8158
rect 1362 8094 1374 8146
rect 1426 8094 1438 8146
rect 8978 8094 8990 8146
rect 9042 8094 9054 8146
rect 35074 8094 35086 8146
rect 35138 8094 35150 8146
rect 40674 8094 40686 8146
rect 40738 8094 40750 8146
rect 50530 8094 50542 8146
rect 50594 8094 50606 8146
rect 51874 8094 51886 8146
rect 51938 8094 51950 8146
rect 6302 8082 6354 8094
rect 19966 8082 20018 8094
rect 55134 8082 55186 8094
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 53006 7698 53058 7710
rect 53006 7634 53058 7646
rect 56142 7698 56194 7710
rect 56142 7634 56194 7646
rect 10558 7586 10610 7598
rect 10558 7522 10610 7534
rect 18958 7586 19010 7598
rect 18958 7522 19010 7534
rect 54574 7586 54626 7598
rect 54574 7522 54626 7534
rect 30606 7474 30658 7486
rect 10098 7422 10110 7474
rect 10162 7422 10174 7474
rect 19394 7422 19406 7474
rect 19458 7422 19470 7474
rect 30606 7410 30658 7422
rect 50878 7474 50930 7486
rect 50878 7410 50930 7422
rect 51438 7474 51490 7486
rect 52098 7422 52110 7474
rect 52162 7422 52174 7474
rect 51438 7410 51490 7422
rect 31166 7362 31218 7374
rect 53554 7310 53566 7362
rect 53618 7310 53630 7362
rect 55122 7310 55134 7362
rect 55186 7310 55198 7362
rect 31166 7298 31218 7310
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 41582 6914 41634 6926
rect 41582 6850 41634 6862
rect 39230 6802 39282 6814
rect 39230 6738 39282 6750
rect 3502 6690 3554 6702
rect 3502 6626 3554 6638
rect 4062 6690 4114 6702
rect 4062 6626 4114 6638
rect 21198 6690 21250 6702
rect 23998 6690 24050 6702
rect 23538 6638 23550 6690
rect 23602 6638 23614 6690
rect 21198 6626 21250 6638
rect 23998 6626 24050 6638
rect 37550 6690 37602 6702
rect 37550 6626 37602 6638
rect 38670 6690 38722 6702
rect 52658 6638 52670 6690
rect 52722 6638 52734 6690
rect 54114 6638 54126 6690
rect 54178 6638 54190 6690
rect 38670 6626 38722 6638
rect 53566 6578 53618 6590
rect 20738 6526 20750 6578
rect 20802 6526 20814 6578
rect 37986 6526 37998 6578
rect 38050 6526 38062 6578
rect 42018 6526 42030 6578
rect 42082 6526 42094 6578
rect 53566 6514 53618 6526
rect 55134 6466 55186 6478
rect 55134 6402 55186 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 53006 6130 53058 6142
rect 53006 6066 53058 6078
rect 56142 6130 56194 6142
rect 56142 6066 56194 6078
rect 30942 6018 30994 6030
rect 13458 5966 13470 6018
rect 13522 5966 13534 6018
rect 14354 5966 14366 6018
rect 14418 5966 14430 6018
rect 19618 5966 19630 6018
rect 19682 5966 19694 6018
rect 30942 5954 30994 5966
rect 54574 6018 54626 6030
rect 54574 5954 54626 5966
rect 14814 5906 14866 5918
rect 14814 5842 14866 5854
rect 30382 5906 30434 5918
rect 52098 5854 52110 5906
rect 52162 5854 52174 5906
rect 30382 5842 30434 5854
rect 15710 5794 15762 5806
rect 15710 5730 15762 5742
rect 31726 5794 31778 5806
rect 53554 5742 53566 5794
rect 53618 5742 53630 5794
rect 55122 5742 55134 5794
rect 55186 5742 55198 5794
rect 31726 5730 31778 5742
rect 13918 5682 13970 5694
rect 13918 5618 13970 5630
rect 15150 5682 15202 5694
rect 15150 5618 15202 5630
rect 20078 5682 20130 5694
rect 20078 5618 20130 5630
rect 32286 5682 32338 5694
rect 32286 5618 32338 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 7310 5346 7362 5358
rect 7310 5282 7362 5294
rect 13134 5346 13186 5358
rect 13134 5282 13186 5294
rect 14142 5346 14194 5358
rect 14142 5282 14194 5294
rect 28478 5346 28530 5358
rect 28478 5282 28530 5294
rect 2046 5234 2098 5246
rect 2046 5170 2098 5182
rect 2606 5234 2658 5246
rect 2606 5170 2658 5182
rect 3950 5234 4002 5246
rect 3950 5170 4002 5182
rect 4510 5234 4562 5246
rect 4510 5170 4562 5182
rect 6750 5234 6802 5246
rect 6750 5170 6802 5182
rect 12574 5234 12626 5246
rect 12574 5170 12626 5182
rect 47518 5234 47570 5246
rect 47518 5170 47570 5182
rect 51998 5234 52050 5246
rect 51998 5170 52050 5182
rect 52894 5234 52946 5246
rect 54114 5182 54126 5234
rect 54178 5182 54190 5234
rect 52894 5170 52946 5182
rect 46958 5122 47010 5134
rect 46958 5058 47010 5070
rect 51438 5122 51490 5134
rect 51438 5058 51490 5070
rect 52334 5122 52386 5134
rect 52334 5058 52386 5070
rect 53230 5122 53282 5134
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 53230 5058 53282 5070
rect 27918 5010 27970 5022
rect 13682 4958 13694 5010
rect 13746 4958 13758 5010
rect 53666 4958 53678 5010
rect 53730 4958 53742 5010
rect 27918 4946 27970 4958
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 54574 4562 54626 4574
rect 54574 4498 54626 4510
rect 56142 4562 56194 4574
rect 56142 4498 56194 4510
rect 5742 4450 5794 4462
rect 39902 4450 39954 4462
rect 36978 4398 36990 4450
rect 37042 4398 37054 4450
rect 5742 4386 5794 4398
rect 39902 4386 39954 4398
rect 49870 4450 49922 4462
rect 52658 4398 52670 4450
rect 52722 4398 52734 4450
rect 49870 4386 49922 4398
rect 5182 4338 5234 4350
rect 5182 4274 5234 4286
rect 39342 4338 39394 4350
rect 39342 4274 39394 4286
rect 41694 4338 41746 4350
rect 41694 4274 41746 4286
rect 52222 4338 52274 4350
rect 52222 4274 52274 4286
rect 42254 4226 42306 4238
rect 53554 4174 53566 4226
rect 53618 4174 53630 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 42254 4162 42306 4174
rect 36542 4114 36594 4126
rect 36542 4050 36594 4062
rect 49310 4114 49362 4126
rect 49310 4050 49362 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 32958 3778 33010 3790
rect 32958 3714 33010 3726
rect 43934 3778 43986 3790
rect 43934 3714 43986 3726
rect 54798 3778 54850 3790
rect 54798 3714 54850 3726
rect 8878 3666 8930 3678
rect 8878 3602 8930 3614
rect 11006 3666 11058 3678
rect 11006 3602 11058 3614
rect 15598 3666 15650 3678
rect 15598 3602 15650 3614
rect 34750 3666 34802 3678
rect 34750 3602 34802 3614
rect 37102 3666 37154 3678
rect 37102 3602 37154 3614
rect 50542 3666 50594 3678
rect 50542 3602 50594 3614
rect 52222 3666 52274 3678
rect 52546 3614 52558 3666
rect 52610 3614 52622 3666
rect 52222 3602 52274 3614
rect 9438 3554 9490 3566
rect 9438 3490 9490 3502
rect 10446 3554 10498 3566
rect 18622 3554 18674 3566
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 10446 3490 10498 3502
rect 18622 3490 18674 3502
rect 19182 3554 19234 3566
rect 36542 3554 36594 3566
rect 35186 3502 35198 3554
rect 35250 3502 35262 3554
rect 19182 3490 19234 3502
rect 36542 3490 36594 3502
rect 49982 3554 50034 3566
rect 49982 3490 50034 3502
rect 51662 3554 51714 3566
rect 55122 3502 55134 3554
rect 55186 3502 55198 3554
rect 51662 3490 51714 3502
rect 32398 3442 32450 3454
rect 53566 3442 53618 3454
rect 44370 3390 44382 3442
rect 44434 3390 44446 3442
rect 32398 3378 32450 3390
rect 53566 3378 53618 3390
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 54574 2994 54626 3006
rect 54574 2930 54626 2942
rect 56142 2994 56194 3006
rect 56142 2930 56194 2942
rect 22094 2882 22146 2894
rect 32846 2882 32898 2894
rect 3938 2830 3950 2882
rect 4002 2830 4014 2882
rect 28578 2830 28590 2882
rect 28642 2830 28654 2882
rect 22094 2818 22146 2830
rect 32846 2818 32898 2830
rect 25454 2770 25506 2782
rect 4274 2718 4286 2770
rect 4338 2718 4350 2770
rect 25454 2706 25506 2718
rect 32286 2770 32338 2782
rect 32286 2706 32338 2718
rect 37886 2770 37938 2782
rect 52098 2718 52110 2770
rect 52162 2718 52174 2770
rect 53554 2718 53566 2770
rect 53618 2718 53630 2770
rect 55122 2718 55134 2770
rect 55186 2718 55198 2770
rect 37886 2706 37938 2718
rect 21534 2658 21586 2670
rect 21534 2594 21586 2606
rect 24894 2658 24946 2670
rect 24894 2594 24946 2606
rect 38446 2658 38498 2670
rect 52770 2606 52782 2658
rect 52834 2606 52846 2658
rect 38446 2594 38498 2606
rect 29038 2546 29090 2558
rect 29038 2482 29090 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 2494 2210 2546 2222
rect 2494 2146 2546 2158
rect 6974 2210 7026 2222
rect 6974 2146 7026 2158
rect 14254 2210 14306 2222
rect 14254 2146 14306 2158
rect 21310 2210 21362 2222
rect 21310 2146 21362 2158
rect 24558 2210 24610 2222
rect 24558 2146 24610 2158
rect 28926 2210 28978 2222
rect 28926 2146 28978 2158
rect 1934 2098 1986 2110
rect 1934 2034 1986 2046
rect 6414 2098 6466 2110
rect 6414 2034 6466 2046
rect 13694 2098 13746 2110
rect 13694 2034 13746 2046
rect 25118 2098 25170 2110
rect 25118 2034 25170 2046
rect 29486 2098 29538 2110
rect 52546 2046 52558 2098
rect 52610 2046 52622 2098
rect 54114 2046 54126 2098
rect 54178 2046 54190 2098
rect 54898 2046 54910 2098
rect 54962 2046 54974 2098
rect 29486 2034 29538 2046
rect 17838 1986 17890 1998
rect 3266 1934 3278 1986
rect 3330 1934 3342 1986
rect 17838 1922 17890 1934
rect 30942 1986 30994 1998
rect 51762 1934 51774 1986
rect 51826 1934 51838 1986
rect 30942 1922 30994 1934
rect 20750 1874 20802 1886
rect 53566 1874 53618 1886
rect 2930 1822 2942 1874
rect 2994 1822 3006 1874
rect 17378 1822 17390 1874
rect 17442 1822 17454 1874
rect 30482 1822 30494 1874
rect 30546 1822 30558 1874
rect 52098 1822 52110 1874
rect 52162 1822 52174 1874
rect 20750 1810 20802 1822
rect 53566 1810 53618 1822
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 53566 1426 53618 1438
rect 53566 1362 53618 1374
rect 56142 1426 56194 1438
rect 56142 1362 56194 1374
rect 51998 1314 52050 1326
rect 51998 1250 52050 1262
rect 50978 1150 50990 1202
rect 51042 1150 51054 1202
rect 52546 1150 52558 1202
rect 52610 1150 52622 1202
rect 55122 1150 55134 1202
rect 55186 1150 55198 1202
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 2158 13134 2210 13186
rect 3726 13134 3778 13186
rect 5966 13134 6018 13186
rect 7534 13134 7586 13186
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 21198 13134 21250 13186
rect 22654 13134 22706 13186
rect 25454 13134 25506 13186
rect 48974 13134 49026 13186
rect 51102 13134 51154 13186
rect 54910 13134 54962 13186
rect 14926 13022 14978 13074
rect 17502 13022 17554 13074
rect 52894 13022 52946 13074
rect 2606 12910 2658 12962
rect 4286 12910 4338 12962
rect 6526 12910 6578 12962
rect 8094 12910 8146 12962
rect 10334 12910 10386 12962
rect 11902 12910 11954 12962
rect 12910 12910 12962 12962
rect 15598 12910 15650 12962
rect 16942 12910 16994 12962
rect 18286 12910 18338 12962
rect 21758 12910 21810 12962
rect 22094 12910 22146 12962
rect 25118 12910 25170 12962
rect 44942 12910 44994 12962
rect 46846 12910 46898 12962
rect 48414 12910 48466 12962
rect 50542 12910 50594 12962
rect 52334 12910 52386 12962
rect 54350 12910 54402 12962
rect 13918 12798 13970 12850
rect 19294 12798 19346 12850
rect 24110 12798 24162 12850
rect 45950 12798 46002 12850
rect 47854 12798 47906 12850
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 2270 12350 2322 12402
rect 6974 12350 7026 12402
rect 8542 12350 8594 12402
rect 10110 12350 10162 12402
rect 11678 12350 11730 12402
rect 14814 12350 14866 12402
rect 16718 12350 16770 12402
rect 22318 12350 22370 12402
rect 23886 12350 23938 12402
rect 49422 12350 49474 12402
rect 52558 12350 52610 12402
rect 54126 12350 54178 12402
rect 55694 12350 55746 12402
rect 3614 12238 3666 12290
rect 5406 12238 5458 12290
rect 18174 12238 18226 12290
rect 19518 12238 19570 12290
rect 21086 12238 21138 12290
rect 27918 12238 27970 12290
rect 28590 12238 28642 12290
rect 38110 12238 38162 12290
rect 2718 12126 2770 12178
rect 5854 12126 5906 12178
rect 18846 12126 18898 12178
rect 20638 12126 20690 12178
rect 21982 12126 22034 12178
rect 23326 12126 23378 12178
rect 36878 12126 36930 12178
rect 44718 12126 44770 12178
rect 46398 12126 46450 12178
rect 52222 12126 52274 12178
rect 4398 12014 4450 12066
rect 7534 12014 7586 12066
rect 9102 12014 9154 12066
rect 10670 12014 10722 12066
rect 12238 12014 12290 12066
rect 12798 12014 12850 12066
rect 15374 12014 15426 12066
rect 15710 12014 15762 12066
rect 17278 12014 17330 12066
rect 29038 12014 29090 12066
rect 36318 12014 36370 12066
rect 45278 12014 45330 12066
rect 46958 12014 47010 12066
rect 48526 12014 48578 12066
rect 48862 12014 48914 12066
rect 50990 12014 51042 12066
rect 53566 12014 53618 12066
rect 55134 12014 55186 12066
rect 13358 11902 13410 11954
rect 27358 11902 27410 11954
rect 37662 11902 37714 11954
rect 47966 11902 48018 11954
rect 50430 11902 50482 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 4622 11566 4674 11618
rect 6190 11566 6242 11618
rect 7758 11566 7810 11618
rect 10894 11566 10946 11618
rect 13918 11566 13970 11618
rect 15486 11566 15538 11618
rect 17390 11566 17442 11618
rect 20526 11566 20578 11618
rect 30942 11566 30994 11618
rect 47182 11566 47234 11618
rect 47518 11566 47570 11618
rect 50318 11566 50370 11618
rect 51886 11566 51938 11618
rect 53454 11566 53506 11618
rect 2830 11454 2882 11506
rect 8318 11454 8370 11506
rect 25118 11454 25170 11506
rect 1934 11342 1986 11394
rect 3614 11342 3666 11394
rect 5182 11342 5234 11394
rect 6638 11342 6690 11394
rect 11454 11342 11506 11394
rect 13022 11342 13074 11394
rect 13582 11342 13634 11394
rect 14926 11342 14978 11394
rect 16830 11342 16882 11394
rect 18622 11342 18674 11394
rect 19966 11342 20018 11394
rect 22766 11342 22818 11394
rect 24558 11342 24610 11394
rect 34414 11342 34466 11394
rect 48302 11342 48354 11394
rect 49758 11342 49810 11394
rect 51326 11342 51378 11394
rect 52894 11342 52946 11394
rect 54462 11342 54514 11394
rect 1598 11230 1650 11282
rect 12350 11230 12402 11282
rect 19070 11230 19122 11282
rect 21758 11230 21810 11282
rect 31390 11230 31442 11282
rect 34974 11230 35026 11282
rect 49198 11230 49250 11282
rect 55022 11230 55074 11282
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 3390 10782 3442 10834
rect 7422 10782 7474 10834
rect 8990 10782 9042 10834
rect 10558 10782 10610 10834
rect 13022 10782 13074 10834
rect 14590 10782 14642 10834
rect 18510 10782 18562 10834
rect 49646 10782 49698 10834
rect 51214 10782 51266 10834
rect 52558 10782 52610 10834
rect 2158 10670 2210 10722
rect 6078 10670 6130 10722
rect 16942 10670 16994 10722
rect 19630 10670 19682 10722
rect 21870 10670 21922 10722
rect 48190 10670 48242 10722
rect 54574 10670 54626 10722
rect 56142 10670 56194 10722
rect 4398 10558 4450 10610
rect 8206 10558 8258 10610
rect 21086 10558 21138 10610
rect 41358 10558 41410 10610
rect 42254 10558 42306 10610
rect 42814 10558 42866 10610
rect 47630 10558 47682 10610
rect 48862 10558 48914 10610
rect 52110 10558 52162 10610
rect 55358 10558 55410 10610
rect 2830 10446 2882 10498
rect 6862 10446 6914 10498
rect 9998 10446 10050 10498
rect 11566 10446 11618 10498
rect 14030 10446 14082 10498
rect 15598 10446 15650 10498
rect 16158 10446 16210 10498
rect 17950 10446 18002 10498
rect 36990 10446 37042 10498
rect 41918 10446 41970 10498
rect 50206 10446 50258 10498
rect 53566 10446 53618 10498
rect 20078 10334 20130 10386
rect 37550 10334 37602 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 17390 9998 17442 10050
rect 26126 9998 26178 10050
rect 1486 9886 1538 9938
rect 5294 9886 5346 9938
rect 9438 9886 9490 9938
rect 16830 9886 16882 9938
rect 23438 9886 23490 9938
rect 23998 9886 24050 9938
rect 25566 9886 25618 9938
rect 36654 9886 36706 9938
rect 1262 9774 1314 9826
rect 3054 9774 3106 9826
rect 6302 9774 6354 9826
rect 9998 9774 10050 9826
rect 10894 9774 10946 9826
rect 20862 9774 20914 9826
rect 36094 9774 36146 9826
rect 41470 9774 41522 9826
rect 42590 9774 42642 9826
rect 44718 9774 44770 9826
rect 48526 9774 48578 9826
rect 49646 9774 49698 9826
rect 50206 9774 50258 9826
rect 51102 9774 51154 9826
rect 52558 9774 52610 9826
rect 54238 9774 54290 9826
rect 2046 9662 2098 9714
rect 4286 9662 4338 9714
rect 5854 9662 5906 9714
rect 10446 9662 10498 9714
rect 20302 9662 20354 9714
rect 41918 9662 41970 9714
rect 43150 9662 43202 9714
rect 45166 9662 45218 9714
rect 49086 9662 49138 9714
rect 51998 9662 52050 9714
rect 53566 9662 53618 9714
rect 55134 9550 55186 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 51214 9214 51266 9266
rect 53006 9214 53058 9266
rect 1710 9102 1762 9154
rect 2942 9102 2994 9154
rect 5966 9102 6018 9154
rect 3502 8990 3554 9042
rect 49758 8990 49810 9042
rect 52110 8990 52162 9042
rect 55246 8990 55298 9042
rect 2606 8878 2658 8930
rect 10334 8878 10386 8930
rect 22430 8878 22482 8930
rect 47630 8878 47682 8930
rect 49310 8878 49362 8930
rect 50206 8878 50258 8930
rect 53566 8878 53618 8930
rect 54350 8878 54402 8930
rect 55918 8878 55970 8930
rect 6526 8766 6578 8818
rect 10894 8766 10946 8818
rect 22990 8766 23042 8818
rect 47070 8766 47122 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 20526 8430 20578 8482
rect 34638 8430 34690 8482
rect 53342 8318 53394 8370
rect 2270 8206 2322 8258
rect 5854 8206 5906 8258
rect 9438 8206 9490 8258
rect 21534 8206 21586 8258
rect 22094 8206 22146 8258
rect 40350 8206 40402 8258
rect 48414 8206 48466 8258
rect 48974 8206 49026 8258
rect 50094 8206 50146 8258
rect 50990 8206 51042 8258
rect 52558 8206 52610 8258
rect 54126 8206 54178 8258
rect 1374 8094 1426 8146
rect 6302 8094 6354 8146
rect 8990 8094 9042 8146
rect 19966 8094 20018 8146
rect 35086 8094 35138 8146
rect 40686 8094 40738 8146
rect 50542 8094 50594 8146
rect 51886 8094 51938 8146
rect 55134 8094 55186 8146
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 53006 7646 53058 7698
rect 56142 7646 56194 7698
rect 10558 7534 10610 7586
rect 18958 7534 19010 7586
rect 54574 7534 54626 7586
rect 10110 7422 10162 7474
rect 19406 7422 19458 7474
rect 30606 7422 30658 7474
rect 50878 7422 50930 7474
rect 51438 7422 51490 7474
rect 52110 7422 52162 7474
rect 31166 7310 31218 7362
rect 53566 7310 53618 7362
rect 55134 7310 55186 7362
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 41582 6862 41634 6914
rect 39230 6750 39282 6802
rect 3502 6638 3554 6690
rect 4062 6638 4114 6690
rect 21198 6638 21250 6690
rect 23550 6638 23602 6690
rect 23998 6638 24050 6690
rect 37550 6638 37602 6690
rect 38670 6638 38722 6690
rect 52670 6638 52722 6690
rect 54126 6638 54178 6690
rect 20750 6526 20802 6578
rect 37998 6526 38050 6578
rect 42030 6526 42082 6578
rect 53566 6526 53618 6578
rect 55134 6414 55186 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 53006 6078 53058 6130
rect 56142 6078 56194 6130
rect 13470 5966 13522 6018
rect 14366 5966 14418 6018
rect 19630 5966 19682 6018
rect 30942 5966 30994 6018
rect 54574 5966 54626 6018
rect 14814 5854 14866 5906
rect 30382 5854 30434 5906
rect 52110 5854 52162 5906
rect 15710 5742 15762 5794
rect 31726 5742 31778 5794
rect 53566 5742 53618 5794
rect 55134 5742 55186 5794
rect 13918 5630 13970 5682
rect 15150 5630 15202 5682
rect 20078 5630 20130 5682
rect 32286 5630 32338 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 7310 5294 7362 5346
rect 13134 5294 13186 5346
rect 14142 5294 14194 5346
rect 28478 5294 28530 5346
rect 2046 5182 2098 5234
rect 2606 5182 2658 5234
rect 3950 5182 4002 5234
rect 4510 5182 4562 5234
rect 6750 5182 6802 5234
rect 12574 5182 12626 5234
rect 47518 5182 47570 5234
rect 51998 5182 52050 5234
rect 52894 5182 52946 5234
rect 54126 5182 54178 5234
rect 46958 5070 47010 5122
rect 51438 5070 51490 5122
rect 52334 5070 52386 5122
rect 53230 5070 53282 5122
rect 54910 5070 54962 5122
rect 13694 4958 13746 5010
rect 27918 4958 27970 5010
rect 53678 4958 53730 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 54574 4510 54626 4562
rect 56142 4510 56194 4562
rect 5742 4398 5794 4450
rect 36990 4398 37042 4450
rect 39902 4398 39954 4450
rect 49870 4398 49922 4450
rect 52670 4398 52722 4450
rect 5182 4286 5234 4338
rect 39342 4286 39394 4338
rect 41694 4286 41746 4338
rect 52222 4286 52274 4338
rect 42254 4174 42306 4226
rect 53566 4174 53618 4226
rect 55134 4174 55186 4226
rect 36542 4062 36594 4114
rect 49310 4062 49362 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 32958 3726 33010 3778
rect 43934 3726 43986 3778
rect 54798 3726 54850 3778
rect 8878 3614 8930 3666
rect 11006 3614 11058 3666
rect 15598 3614 15650 3666
rect 34750 3614 34802 3666
rect 37102 3614 37154 3666
rect 50542 3614 50594 3666
rect 52222 3614 52274 3666
rect 52558 3614 52610 3666
rect 9438 3502 9490 3554
rect 10446 3502 10498 3554
rect 15150 3502 15202 3554
rect 18622 3502 18674 3554
rect 19182 3502 19234 3554
rect 35198 3502 35250 3554
rect 36542 3502 36594 3554
rect 49982 3502 50034 3554
rect 51662 3502 51714 3554
rect 55134 3502 55186 3554
rect 32398 3390 32450 3442
rect 44382 3390 44434 3442
rect 53566 3390 53618 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 54574 2942 54626 2994
rect 56142 2942 56194 2994
rect 3950 2830 4002 2882
rect 22094 2830 22146 2882
rect 28590 2830 28642 2882
rect 32846 2830 32898 2882
rect 4286 2718 4338 2770
rect 25454 2718 25506 2770
rect 32286 2718 32338 2770
rect 37886 2718 37938 2770
rect 52110 2718 52162 2770
rect 53566 2718 53618 2770
rect 55134 2718 55186 2770
rect 21534 2606 21586 2658
rect 24894 2606 24946 2658
rect 38446 2606 38498 2658
rect 52782 2606 52834 2658
rect 29038 2494 29090 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 2494 2158 2546 2210
rect 6974 2158 7026 2210
rect 14254 2158 14306 2210
rect 21310 2158 21362 2210
rect 24558 2158 24610 2210
rect 28926 2158 28978 2210
rect 1934 2046 1986 2098
rect 6414 2046 6466 2098
rect 13694 2046 13746 2098
rect 25118 2046 25170 2098
rect 29486 2046 29538 2098
rect 52558 2046 52610 2098
rect 54126 2046 54178 2098
rect 54910 2046 54962 2098
rect 3278 1934 3330 1986
rect 17838 1934 17890 1986
rect 30942 1934 30994 1986
rect 51774 1934 51826 1986
rect 2942 1822 2994 1874
rect 17390 1822 17442 1874
rect 20750 1822 20802 1874
rect 30494 1822 30546 1874
rect 52110 1822 52162 1874
rect 53566 1822 53618 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 53566 1374 53618 1426
rect 56142 1374 56194 1426
rect 51998 1262 52050 1314
rect 50990 1150 51042 1202
rect 52558 1150 52610 1202
rect 55134 1150 55186 1202
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 672 14112 784 14224
rect 1120 14112 1232 14224
rect 1568 14112 1680 14224
rect 2016 14112 2128 14224
rect 2464 14112 2576 14224
rect 2912 14112 3024 14224
rect 3360 14112 3472 14224
rect 3808 14112 3920 14224
rect 4256 14112 4368 14224
rect 4704 14112 4816 14224
rect 5152 14112 5264 14224
rect 5600 14112 5712 14224
rect 6048 14112 6160 14224
rect 6496 14112 6608 14224
rect 6944 14112 7056 14224
rect 7392 14112 7504 14224
rect 7840 14112 7952 14224
rect 8288 14112 8400 14224
rect 8736 14112 8848 14224
rect 9184 14112 9296 14224
rect 9632 14112 9744 14224
rect 10080 14112 10192 14224
rect 10528 14112 10640 14224
rect 10976 14112 11088 14224
rect 11424 14112 11536 14224
rect 11872 14112 11984 14224
rect 12320 14112 12432 14224
rect 12768 14112 12880 14224
rect 13216 14112 13328 14224
rect 13664 14112 13776 14224
rect 14112 14112 14224 14224
rect 14560 14112 14672 14224
rect 15008 14112 15120 14224
rect 15456 14112 15568 14224
rect 15904 14112 16016 14224
rect 16352 14112 16464 14224
rect 16800 14112 16912 14224
rect 17248 14112 17360 14224
rect 17696 14112 17808 14224
rect 18144 14112 18256 14224
rect 18592 14112 18704 14224
rect 19040 14112 19152 14224
rect 19488 14112 19600 14224
rect 19936 14112 20048 14224
rect 20384 14112 20496 14224
rect 20832 14112 20944 14224
rect 21280 14112 21392 14224
rect 21728 14112 21840 14224
rect 22176 14112 22288 14224
rect 22624 14112 22736 14224
rect 23072 14112 23184 14224
rect 23520 14112 23632 14224
rect 23968 14112 24080 14224
rect 24416 14112 24528 14224
rect 24864 14112 24976 14224
rect 25312 14112 25424 14224
rect 25760 14112 25872 14224
rect 26208 14112 26320 14224
rect 26656 14112 26768 14224
rect 27104 14112 27216 14224
rect 27552 14112 27664 14224
rect 28000 14112 28112 14224
rect 28448 14112 28560 14224
rect 28896 14112 29008 14224
rect 29344 14112 29456 14224
rect 29792 14112 29904 14224
rect 30240 14112 30352 14224
rect 30688 14112 30800 14224
rect 31136 14112 31248 14224
rect 31584 14112 31696 14224
rect 32032 14112 32144 14224
rect 32480 14112 32592 14224
rect 32928 14112 33040 14224
rect 33376 14112 33488 14224
rect 33824 14112 33936 14224
rect 34272 14112 34384 14224
rect 34720 14112 34832 14224
rect 35168 14112 35280 14224
rect 35616 14112 35728 14224
rect 36064 14112 36176 14224
rect 36512 14112 36624 14224
rect 36960 14112 37072 14224
rect 37408 14112 37520 14224
rect 37856 14112 37968 14224
rect 38304 14112 38416 14224
rect 38752 14112 38864 14224
rect 39200 14112 39312 14224
rect 39648 14112 39760 14224
rect 40096 14112 40208 14224
rect 40544 14112 40656 14224
rect 40992 14112 41104 14224
rect 41440 14112 41552 14224
rect 41888 14112 42000 14224
rect 42336 14112 42448 14224
rect 42784 14112 42896 14224
rect 43232 14112 43344 14224
rect 43680 14112 43792 14224
rect 44128 14112 44240 14224
rect 44576 14112 44688 14224
rect 45024 14112 45136 14224
rect 45472 14112 45584 14224
rect 45920 14112 46032 14224
rect 46368 14112 46480 14224
rect 46816 14112 46928 14224
rect 47264 14112 47376 14224
rect 47712 14112 47824 14224
rect 48160 14112 48272 14224
rect 48608 14112 48720 14224
rect 49056 14112 49168 14224
rect 49504 14112 49616 14224
rect 49952 14112 50064 14224
rect 50400 14112 50512 14224
rect 50848 14112 50960 14224
rect 51296 14112 51408 14224
rect 51744 14112 51856 14224
rect 52192 14112 52304 14224
rect 52640 14112 52752 14224
rect 53088 14112 53200 14224
rect 53536 14112 53648 14224
rect 53984 14112 54096 14224
rect 54432 14112 54544 14224
rect 54880 14112 54992 14224
rect 55328 14112 55440 14224
rect 55776 14112 55888 14224
rect 56224 14112 56336 14224
rect 56672 14112 56784 14224
rect 364 13076 420 13086
rect 140 10612 196 10622
rect 140 9940 196 10556
rect 364 10052 420 13020
rect 476 12628 532 12638
rect 476 11396 532 12572
rect 476 11330 532 11340
rect 588 12180 644 12190
rect 364 9986 420 9996
rect 140 9874 196 9884
rect 588 9716 644 12124
rect 700 11284 756 14112
rect 1036 13524 1092 13534
rect 1036 11508 1092 13468
rect 1148 11844 1204 14112
rect 1596 11956 1652 14112
rect 1596 11900 1764 11956
rect 1148 11788 1652 11844
rect 1596 11620 1652 11788
rect 1708 11732 1764 11900
rect 2044 11844 2100 14112
rect 2156 13300 2212 13310
rect 2156 13186 2212 13244
rect 2156 13134 2158 13186
rect 2210 13134 2212 13186
rect 2156 13122 2212 13134
rect 2492 13188 2548 14112
rect 2492 13132 2884 13188
rect 2604 12964 2660 12974
rect 2380 12962 2660 12964
rect 2380 12910 2606 12962
rect 2658 12910 2660 12962
rect 2380 12908 2660 12910
rect 2268 12404 2324 12414
rect 2268 12310 2324 12348
rect 2268 11844 2324 11854
rect 2044 11788 2212 11844
rect 1708 11676 2100 11732
rect 1596 11564 1764 11620
rect 1036 11442 1092 11452
rect 1596 11284 1652 11294
rect 700 11228 1428 11284
rect 588 9650 644 9660
rect 924 11060 980 11070
rect 924 8372 980 11004
rect 1260 9828 1316 9838
rect 1260 9734 1316 9772
rect 812 8316 980 8372
rect 1148 9492 1204 9502
rect 812 6468 868 8316
rect 812 6402 868 6412
rect 1036 7028 1092 7038
rect 1036 1876 1092 6972
rect 1148 6692 1204 9436
rect 1148 6626 1204 6636
rect 1260 8596 1316 8606
rect 1260 4340 1316 8540
rect 1372 8146 1428 11228
rect 1596 11190 1652 11228
rect 1596 10836 1652 10846
rect 1372 8094 1374 8146
rect 1426 8094 1428 8146
rect 1372 8082 1428 8094
rect 1484 9938 1540 9950
rect 1484 9886 1486 9938
rect 1538 9886 1540 9938
rect 1372 7700 1428 7710
rect 1372 6356 1428 7644
rect 1372 6290 1428 6300
rect 1372 5796 1428 5806
rect 1372 4564 1428 5740
rect 1484 5124 1540 9886
rect 1596 8932 1652 10780
rect 1708 9154 1764 11564
rect 1932 11394 1988 11406
rect 1932 11342 1934 11394
rect 1986 11342 1988 11394
rect 1708 9102 1710 9154
rect 1762 9102 1764 9154
rect 1708 9090 1764 9102
rect 1820 9828 1876 9838
rect 1596 8876 1764 8932
rect 1596 8372 1652 8382
rect 1596 7252 1652 8316
rect 1708 7476 1764 8876
rect 1708 7410 1764 7420
rect 1596 7186 1652 7196
rect 1596 6132 1652 6142
rect 1596 5460 1652 6076
rect 1596 5394 1652 5404
rect 1484 5058 1540 5068
rect 1372 4498 1428 4508
rect 1260 4274 1316 4284
rect 1596 3780 1652 3790
rect 1596 3220 1652 3724
rect 1596 3154 1652 3164
rect 1036 1810 1092 1820
rect 1148 1988 1204 1998
rect 924 1764 980 1774
rect 924 980 980 1708
rect 924 914 980 924
rect 1148 84 1204 1932
rect 1820 112 1876 9772
rect 1932 4564 1988 11342
rect 2044 9714 2100 11676
rect 2156 10722 2212 11788
rect 2156 10670 2158 10722
rect 2210 10670 2212 10722
rect 2156 10658 2212 10670
rect 2044 9662 2046 9714
rect 2098 9662 2100 9714
rect 2044 9650 2100 9662
rect 2268 8428 2324 11788
rect 2044 8372 2324 8428
rect 2380 8428 2436 12908
rect 2604 12898 2660 12908
rect 2716 12178 2772 12190
rect 2716 12126 2718 12178
rect 2770 12126 2772 12178
rect 2492 10052 2548 10062
rect 2492 8708 2548 9996
rect 2604 8932 2660 8942
rect 2604 8838 2660 8876
rect 2492 8642 2548 8652
rect 2380 8372 2548 8428
rect 2044 5234 2100 8372
rect 2268 8260 2324 8270
rect 2268 8166 2324 8204
rect 2044 5182 2046 5234
rect 2098 5182 2100 5234
rect 2044 5170 2100 5182
rect 2380 7252 2436 7262
rect 1932 4508 2100 4564
rect 1932 4228 1988 4238
rect 1932 2098 1988 4172
rect 1932 2046 1934 2098
rect 1986 2046 1988 2098
rect 1932 2034 1988 2046
rect 2044 644 2100 4508
rect 2044 578 2100 588
rect 2380 532 2436 7196
rect 2492 4788 2548 8372
rect 2604 5236 2660 5246
rect 2604 5142 2660 5180
rect 2492 4732 2660 4788
rect 2492 2212 2548 2222
rect 2492 2118 2548 2156
rect 2604 980 2660 4732
rect 2716 3556 2772 12126
rect 2828 11506 2884 13132
rect 2940 11956 2996 14112
rect 3388 12404 3444 14112
rect 3388 12338 3444 12348
rect 3612 13524 3668 13534
rect 3612 12290 3668 13468
rect 3724 13188 3780 13198
rect 3724 13094 3780 13132
rect 3836 12740 3892 14112
rect 4284 13300 4340 14112
rect 4732 13524 4788 14112
rect 4732 13458 4788 13468
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4284 13234 4340 13244
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 3836 12684 4340 12740
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 3612 12238 3614 12290
rect 3666 12238 3668 12290
rect 3612 12226 3668 12238
rect 2940 11890 2996 11900
rect 3388 11956 3444 11966
rect 2828 11454 2830 11506
rect 2882 11454 2884 11506
rect 2828 11442 2884 11454
rect 3276 10836 3332 10846
rect 3164 10724 3220 10734
rect 2828 10500 2884 10510
rect 2828 10406 2884 10444
rect 2828 10276 2884 10286
rect 2828 8932 2884 10220
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 2940 9604 2996 9614
rect 2940 9154 2996 9548
rect 3052 9268 3108 9774
rect 3052 9202 3108 9212
rect 2940 9102 2942 9154
rect 2994 9102 2996 9154
rect 2940 9090 2996 9102
rect 2828 8876 2996 8932
rect 2716 3490 2772 3500
rect 2828 8708 2884 8718
rect 2828 1764 2884 8652
rect 2940 7140 2996 8876
rect 2940 7074 2996 7084
rect 3052 7588 3108 7598
rect 3052 4900 3108 7532
rect 3164 7028 3220 10668
rect 3276 8148 3332 10780
rect 3388 10834 3444 11900
rect 4172 11732 4228 11742
rect 3388 10782 3390 10834
rect 3442 10782 3444 10834
rect 3388 10770 3444 10782
rect 3612 11394 3668 11406
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3500 9604 3556 9614
rect 3500 9042 3556 9548
rect 3500 8990 3502 9042
rect 3554 8990 3556 9042
rect 3500 8978 3556 8990
rect 3276 8082 3332 8092
rect 3164 6962 3220 6972
rect 3500 7364 3556 7374
rect 3276 6916 3332 6926
rect 3276 5908 3332 6860
rect 3500 6690 3556 7308
rect 3500 6638 3502 6690
rect 3554 6638 3556 6690
rect 3500 6626 3556 6638
rect 3276 5842 3332 5852
rect 3052 4834 3108 4844
rect 3276 5684 3332 5694
rect 3276 4116 3332 5628
rect 3276 4050 3332 4060
rect 3612 3388 3668 11342
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4172 8260 4228 11676
rect 4284 9714 4340 12684
rect 4396 12068 4452 12078
rect 4396 11974 4452 12012
rect 5068 12068 5124 12078
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4620 11620 4676 11630
rect 4620 11526 4676 11564
rect 4956 11396 5012 11406
rect 4396 11060 4452 11070
rect 4396 10610 4452 11004
rect 4396 10558 4398 10610
rect 4450 10558 4452 10610
rect 4396 10546 4452 10558
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4284 9662 4286 9714
rect 4338 9662 4340 9714
rect 4284 9650 4340 9662
rect 4956 9492 5012 11340
rect 4956 9426 5012 9436
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 4172 8194 4228 8204
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 5068 7700 5124 12012
rect 5180 11620 5236 14112
rect 5404 13636 5460 13646
rect 5180 11554 5236 11564
rect 5292 13076 5348 13086
rect 5180 11394 5236 11406
rect 5180 11342 5182 11394
rect 5234 11342 5236 11394
rect 5180 10948 5236 11342
rect 5180 10882 5236 10892
rect 5292 10276 5348 13020
rect 5404 12290 5460 13580
rect 5628 13188 5684 14112
rect 5628 13122 5684 13132
rect 5964 13300 6020 13310
rect 5964 13186 6020 13244
rect 5964 13134 5966 13186
rect 6018 13134 6020 13186
rect 5964 13122 6020 13134
rect 5404 12238 5406 12290
rect 5458 12238 5460 12290
rect 5404 12226 5460 12238
rect 5964 12516 6020 12526
rect 5852 12180 5908 12190
rect 5180 10220 5348 10276
rect 5516 12178 5908 12180
rect 5516 12126 5854 12178
rect 5906 12126 5908 12178
rect 5516 12124 5908 12126
rect 5180 9044 5236 10220
rect 5292 10052 5348 10062
rect 5292 9938 5348 9996
rect 5292 9886 5294 9938
rect 5346 9886 5348 9938
rect 5292 9874 5348 9886
rect 5180 8978 5236 8988
rect 5068 7644 5348 7700
rect 4284 7140 4340 7150
rect 4060 6692 4116 6702
rect 4060 6690 4228 6692
rect 4060 6638 4062 6690
rect 4114 6638 4228 6690
rect 4060 6636 4228 6638
rect 4060 6626 4116 6636
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3724 5908 3780 5918
rect 3724 5684 3780 5852
rect 3724 5618 3780 5628
rect 3948 5684 4004 5694
rect 3948 5234 4004 5628
rect 3948 5182 3950 5234
rect 4002 5182 4004 5234
rect 3948 5170 4004 5182
rect 4172 4788 4228 6636
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4172 4722 4228 4732
rect 3804 4666 4068 4676
rect 4284 4676 4340 7084
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4508 5236 4564 5246
rect 4508 5142 4564 5180
rect 4284 4610 4340 4620
rect 5068 5124 5124 5134
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 3500 3332 3668 3388
rect 3500 3266 3556 3276
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3948 2884 4004 2894
rect 3948 2882 4228 2884
rect 3948 2830 3950 2882
rect 4002 2830 4228 2882
rect 3948 2828 4228 2830
rect 3948 2818 4004 2828
rect 3276 1986 3332 1998
rect 3276 1934 3278 1986
rect 3330 1934 3332 1986
rect 2940 1876 2996 1886
rect 2940 1782 2996 1820
rect 2828 1698 2884 1708
rect 3276 1428 3332 1934
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 3276 1362 3332 1372
rect 4172 1092 4228 2828
rect 4284 2770 4340 2782
rect 4284 2718 4286 2770
rect 4338 2718 4340 2770
rect 4284 1764 4340 2718
rect 5068 2548 5124 5068
rect 5180 4340 5236 4350
rect 5180 4246 5236 4284
rect 5292 3108 5348 7644
rect 5292 3042 5348 3052
rect 5404 4900 5460 4910
rect 5068 2482 5124 2492
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 5404 2100 5460 4844
rect 5404 2034 5460 2044
rect 4284 1698 4340 1708
rect 5516 1316 5572 12124
rect 5852 12114 5908 12124
rect 5964 11060 6020 12460
rect 5852 11004 6020 11060
rect 5852 9714 5908 11004
rect 6076 10722 6132 14112
rect 6524 13188 6580 14112
rect 6748 14084 6804 14094
rect 6748 13972 6804 14028
rect 6188 13132 6580 13188
rect 6636 13916 6804 13972
rect 6188 11618 6244 13132
rect 6188 11566 6190 11618
rect 6242 11566 6244 11618
rect 6188 11554 6244 11566
rect 6412 12964 6468 12974
rect 6076 10670 6078 10722
rect 6130 10670 6132 10722
rect 6076 10658 6132 10670
rect 5852 9662 5854 9714
rect 5906 9662 5908 9714
rect 5852 9650 5908 9662
rect 5964 10612 6020 10622
rect 5964 9154 6020 10556
rect 6188 10164 6244 10174
rect 6188 9716 6244 10108
rect 6188 9650 6244 9660
rect 6300 9826 6356 9838
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 5964 9102 5966 9154
rect 6018 9102 6020 9154
rect 5964 9090 6020 9102
rect 6300 8372 6356 9774
rect 6412 9716 6468 12908
rect 6524 12964 6580 12974
rect 6636 12964 6692 13916
rect 6524 12962 6692 12964
rect 6524 12910 6526 12962
rect 6578 12910 6692 12962
rect 6524 12908 6692 12910
rect 6524 12898 6580 12908
rect 6748 12852 6804 12862
rect 6412 9650 6468 9660
rect 6636 11394 6692 11406
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6300 8306 6356 8316
rect 6524 8818 6580 8830
rect 6524 8766 6526 8818
rect 6578 8766 6580 8818
rect 5852 8258 5908 8270
rect 5852 8206 5854 8258
rect 5906 8206 5908 8258
rect 5740 4452 5796 4462
rect 5740 4358 5796 4396
rect 5516 1250 5572 1260
rect 4172 1026 4228 1036
rect 2604 914 2660 924
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 2380 466 2436 476
rect 4508 420 4564 430
rect 4508 112 4564 364
rect 5852 420 5908 8206
rect 6300 8148 6356 8158
rect 6300 8054 6356 8092
rect 6300 7812 6356 7822
rect 6300 1988 6356 7756
rect 6524 5572 6580 8766
rect 6636 8036 6692 11342
rect 6636 7970 6692 7980
rect 6524 5506 6580 5516
rect 6748 5234 6804 12796
rect 6972 12628 7028 14112
rect 7420 13300 7476 14112
rect 7420 13234 7476 13244
rect 7532 13188 7588 13198
rect 7532 13094 7588 13132
rect 6972 12572 7476 12628
rect 6972 12404 7028 12414
rect 6972 12310 7028 12348
rect 7420 10834 7476 12572
rect 7868 12404 7924 14112
rect 8316 13188 8372 14112
rect 7868 12338 7924 12348
rect 7980 13132 8372 13188
rect 7980 12180 8036 13132
rect 7756 12124 8036 12180
rect 8092 12962 8148 12974
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 7420 10782 7422 10834
rect 7474 10782 7476 10834
rect 7420 10770 7476 10782
rect 7532 12066 7588 12078
rect 7532 12014 7534 12066
rect 7586 12014 7588 12066
rect 6860 10498 6916 10510
rect 6860 10446 6862 10498
rect 6914 10446 6916 10498
rect 6860 9044 6916 10446
rect 6860 8978 6916 8988
rect 7084 8372 7140 8382
rect 6748 5182 6750 5234
rect 6802 5182 6804 5234
rect 6748 5170 6804 5182
rect 6860 7700 6916 7710
rect 6748 4676 6804 4686
rect 6412 3444 6468 3454
rect 6412 2098 6468 3388
rect 6412 2046 6414 2098
rect 6466 2046 6468 2098
rect 6412 2034 6468 2046
rect 6300 1922 6356 1932
rect 6748 1540 6804 4620
rect 6860 3388 6916 7644
rect 6972 6692 7028 6702
rect 6972 4116 7028 6636
rect 6972 4050 7028 4060
rect 6860 3332 7028 3388
rect 6972 2210 7028 3332
rect 7084 2436 7140 8316
rect 7308 6692 7364 6702
rect 7308 5346 7364 6636
rect 7532 6580 7588 12014
rect 7756 11618 7812 12124
rect 7756 11566 7758 11618
rect 7810 11566 7812 11618
rect 7756 11554 7812 11566
rect 7756 10388 7812 10398
rect 7532 6514 7588 6524
rect 7644 8260 7700 8270
rect 7308 5294 7310 5346
rect 7362 5294 7364 5346
rect 7308 5282 7364 5294
rect 7644 3388 7700 8204
rect 7756 7364 7812 10332
rect 8092 10276 8148 12910
rect 8540 12404 8596 12414
rect 8540 12310 8596 12348
rect 8428 12292 8484 12302
rect 8316 11732 8372 11742
rect 8316 11506 8372 11676
rect 8316 11454 8318 11506
rect 8370 11454 8372 11506
rect 8316 11442 8372 11454
rect 8316 10724 8372 10734
rect 8092 10210 8148 10220
rect 8204 10610 8260 10622
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 7756 7298 7812 7308
rect 8092 9492 8148 9502
rect 8092 4004 8148 9436
rect 8092 3938 8148 3948
rect 8204 3388 8260 10558
rect 8316 10052 8372 10668
rect 8428 10388 8484 12236
rect 8428 10322 8484 10332
rect 8652 11508 8708 11518
rect 8652 10388 8708 11452
rect 8764 10836 8820 14112
rect 9212 13188 9268 14112
rect 9212 13122 9268 13132
rect 9436 12964 9492 12974
rect 9100 12068 9156 12078
rect 9100 12066 9268 12068
rect 9100 12014 9102 12066
rect 9154 12014 9268 12066
rect 9100 12012 9268 12014
rect 9100 12002 9156 12012
rect 8988 10836 9044 10846
rect 8764 10834 9044 10836
rect 8764 10782 8990 10834
rect 9042 10782 9044 10834
rect 8764 10780 9044 10782
rect 8988 10770 9044 10780
rect 8652 10322 8708 10332
rect 9100 10724 9156 10734
rect 8316 9996 8596 10052
rect 8316 9828 8372 9838
rect 8316 8428 8372 9772
rect 8540 9828 8596 9996
rect 8540 9762 8596 9772
rect 8316 8372 8484 8428
rect 8316 8148 8372 8158
rect 8316 4676 8372 8092
rect 8428 7140 8484 8372
rect 8876 8148 8932 8158
rect 8876 7924 8932 8092
rect 8988 8148 9044 8158
rect 9100 8148 9156 10668
rect 8988 8146 9156 8148
rect 8988 8094 8990 8146
rect 9042 8094 9156 8146
rect 8988 8092 9156 8094
rect 8988 8082 9044 8092
rect 8876 7858 8932 7868
rect 9212 7924 9268 12012
rect 9436 9938 9492 12908
rect 9660 12404 9716 14112
rect 9772 13188 9828 13198
rect 9772 13094 9828 13132
rect 10108 12628 10164 14112
rect 9660 12338 9716 12348
rect 9996 12572 10164 12628
rect 10332 12962 10388 12974
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 10332 12628 10388 12910
rect 9884 12180 9940 12190
rect 9996 12180 10052 12572
rect 10332 12562 10388 12572
rect 10108 12404 10164 12414
rect 10556 12404 10612 14112
rect 10108 12402 10612 12404
rect 10108 12350 10110 12402
rect 10162 12350 10612 12402
rect 10108 12348 10612 12350
rect 10108 12338 10164 12348
rect 9996 12124 10612 12180
rect 9548 11844 9604 11854
rect 9548 10500 9604 11788
rect 9884 11060 9940 12124
rect 9884 10994 9940 11004
rect 10444 11172 10500 11182
rect 9548 10434 9604 10444
rect 9660 10948 9716 10958
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 9212 7858 9268 7868
rect 9436 8258 9492 8270
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 8428 7084 8596 7140
rect 8428 6916 8484 6926
rect 8428 6244 8484 6860
rect 8428 6178 8484 6188
rect 8428 5796 8484 5806
rect 8428 4900 8484 5740
rect 8428 4834 8484 4844
rect 8316 4610 8372 4620
rect 7084 2370 7140 2380
rect 7420 3332 7700 3388
rect 8092 3332 8260 3388
rect 8540 3444 8596 7084
rect 9436 6468 9492 8206
rect 9436 6402 9492 6412
rect 8540 3378 8596 3388
rect 8764 6020 8820 6030
rect 8764 3332 8820 5964
rect 8876 5460 8932 5470
rect 8876 3666 8932 5404
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 8876 3602 8932 3614
rect 9660 3668 9716 10892
rect 9772 10500 9828 10510
rect 9772 9604 9828 10444
rect 9996 10498 10052 10510
rect 9996 10446 9998 10498
rect 10050 10446 10052 10498
rect 9996 10052 10052 10446
rect 10444 10164 10500 11116
rect 10556 10834 10612 12124
rect 10668 12068 10724 12078
rect 10668 12066 10836 12068
rect 10668 12014 10670 12066
rect 10722 12014 10836 12066
rect 10668 12012 10836 12014
rect 10668 12002 10724 12012
rect 10556 10782 10558 10834
rect 10610 10782 10612 10834
rect 10556 10770 10612 10782
rect 10444 10098 10500 10108
rect 9996 9996 10276 10052
rect 9772 9538 9828 9548
rect 9996 9826 10052 9838
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 9884 9492 9940 9502
rect 9772 7028 9828 7038
rect 9772 5236 9828 6972
rect 9884 6692 9940 9436
rect 9996 8820 10052 9774
rect 9996 8754 10052 8764
rect 9884 6626 9940 6636
rect 9996 8596 10052 8606
rect 9772 5170 9828 5180
rect 9996 5236 10052 8540
rect 10108 7476 10164 7486
rect 10108 7382 10164 7420
rect 10108 6916 10164 6926
rect 10108 5684 10164 6860
rect 10220 5796 10276 9996
rect 10444 9714 10500 9726
rect 10444 9662 10446 9714
rect 10498 9662 10500 9714
rect 10332 8932 10388 8942
rect 10332 8838 10388 8876
rect 10444 8596 10500 9662
rect 10444 8530 10500 8540
rect 10556 8484 10612 8494
rect 10332 8260 10388 8270
rect 10332 7476 10388 8204
rect 10556 7586 10612 8428
rect 10780 7700 10836 12012
rect 10892 11620 10948 11630
rect 11004 11620 11060 14112
rect 11340 13412 11396 13422
rect 11340 13186 11396 13356
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 11452 13188 11508 14112
rect 11900 13412 11956 14112
rect 11452 13122 11508 13132
rect 11676 13356 11956 13412
rect 12012 13860 12068 13870
rect 10892 11618 11060 11620
rect 10892 11566 10894 11618
rect 10946 11566 11060 11618
rect 10892 11564 11060 11566
rect 11116 12628 11172 12638
rect 10892 11554 10948 11564
rect 11116 11060 11172 12572
rect 11676 12402 11732 13356
rect 11676 12350 11678 12402
rect 11730 12350 11732 12402
rect 11676 12338 11732 12350
rect 11788 13188 11844 13198
rect 11116 10994 11172 11004
rect 11228 12292 11284 12302
rect 11228 9940 11284 12236
rect 11788 11732 11844 13132
rect 11900 12962 11956 12974
rect 11900 12910 11902 12962
rect 11954 12910 11956 12962
rect 11900 12068 11956 12910
rect 11900 12002 11956 12012
rect 11788 11666 11844 11676
rect 12012 11620 12068 13804
rect 12012 11554 12068 11564
rect 12124 13748 12180 13758
rect 11452 11396 11508 11406
rect 11452 11302 11508 11340
rect 11228 9874 11284 9884
rect 11452 10836 11508 10846
rect 10892 9828 10948 9838
rect 10892 9734 10948 9772
rect 10892 8820 10948 8830
rect 10892 8818 11396 8820
rect 10892 8766 10894 8818
rect 10946 8766 11396 8818
rect 10892 8764 11396 8766
rect 10892 8754 10948 8764
rect 10780 7644 11284 7700
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 10556 7522 10612 7534
rect 10332 7410 10388 7420
rect 10332 7252 10388 7262
rect 10332 6692 10388 7196
rect 10332 6626 10388 6636
rect 10444 6804 10500 6814
rect 10444 6356 10500 6748
rect 10444 6290 10500 6300
rect 10220 5730 10276 5740
rect 10332 6020 10388 6030
rect 10108 5618 10164 5628
rect 10332 5684 10388 5964
rect 10332 5618 10388 5628
rect 11116 5908 11172 5918
rect 9996 5170 10052 5180
rect 9660 3602 9716 3612
rect 9996 4564 10052 4574
rect 6972 2158 6974 2210
rect 7026 2158 7028 2210
rect 6972 2146 7028 2158
rect 6748 1474 6804 1484
rect 7196 1652 7252 1662
rect 5852 354 5908 364
rect 7196 112 7252 1596
rect 7420 1204 7476 3332
rect 8092 1652 8148 3332
rect 8764 3266 8820 3276
rect 9436 3554 9492 3566
rect 9436 3502 9438 3554
rect 9490 3502 9492 3554
rect 8092 1586 8148 1596
rect 8316 2884 8372 2894
rect 8316 1316 8372 2828
rect 8540 2772 8596 2782
rect 8540 1428 8596 2716
rect 9436 1876 9492 3502
rect 9436 1810 9492 1820
rect 9884 3556 9940 3566
rect 8540 1362 8596 1372
rect 8316 1250 8372 1260
rect 7420 1138 7476 1148
rect 9884 112 9940 3500
rect 9996 3220 10052 4508
rect 11004 3668 11060 3678
rect 11004 3574 11060 3612
rect 10444 3556 10500 3566
rect 10444 3462 10500 3500
rect 9996 3154 10052 3164
rect 10108 3332 10164 3342
rect 10108 2660 10164 3276
rect 10108 2594 10164 2604
rect 11116 2324 11172 5852
rect 11116 2258 11172 2268
rect 11228 1988 11284 7644
rect 11340 6020 11396 8764
rect 11452 8148 11508 10780
rect 12124 10836 12180 13692
rect 12124 10770 12180 10780
rect 12236 12066 12292 12078
rect 12236 12014 12238 12066
rect 12290 12014 12292 12066
rect 11788 10724 11844 10734
rect 11564 10498 11620 10510
rect 11564 10446 11566 10498
rect 11618 10446 11620 10498
rect 11564 9380 11620 10446
rect 11788 9828 11844 10668
rect 12236 10276 12292 12014
rect 12348 11282 12404 14112
rect 12796 12292 12852 14112
rect 13244 13412 13300 14112
rect 13244 13346 13300 13356
rect 13580 13412 13636 13422
rect 13468 13300 13524 13310
rect 12908 12964 12964 12974
rect 12908 12870 12964 12908
rect 12796 12236 12964 12292
rect 12796 12066 12852 12078
rect 12796 12014 12798 12066
rect 12850 12014 12852 12066
rect 12796 11844 12852 12014
rect 12796 11778 12852 11788
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 11218 12404 11230
rect 12236 10210 12292 10220
rect 12684 11060 12740 11070
rect 11564 9314 11620 9324
rect 11676 9772 11844 9828
rect 11676 9044 11732 9772
rect 11452 8082 11508 8092
rect 11564 8988 11732 9044
rect 11788 9604 11844 9614
rect 11564 7812 11620 8988
rect 11676 8820 11732 8830
rect 11676 8260 11732 8764
rect 11676 8194 11732 8204
rect 11564 7746 11620 7756
rect 11788 7700 11844 9548
rect 12684 9044 12740 11004
rect 12908 10836 12964 12236
rect 13356 11956 13412 11966
rect 13356 11862 13412 11900
rect 13020 11394 13076 11406
rect 13020 11342 13022 11394
rect 13074 11342 13076 11394
rect 13020 11060 13076 11342
rect 13020 10994 13076 11004
rect 13020 10836 13076 10846
rect 12908 10834 13076 10836
rect 12908 10782 13022 10834
rect 13074 10782 13076 10834
rect 12908 10780 13076 10782
rect 13020 10770 13076 10780
rect 12684 8978 12740 8988
rect 13356 9492 13412 9502
rect 12124 8932 12180 8942
rect 11788 7634 11844 7644
rect 12012 7700 12068 7710
rect 11900 7252 11956 7262
rect 11340 5954 11396 5964
rect 11452 6244 11508 6254
rect 11452 2884 11508 6188
rect 11788 6132 11844 6142
rect 11788 3444 11844 6076
rect 11900 5460 11956 7196
rect 11900 5394 11956 5404
rect 12012 4228 12068 7644
rect 12012 4162 12068 4172
rect 11788 3378 11844 3388
rect 11452 2818 11508 2828
rect 12124 2772 12180 8876
rect 13356 8820 13412 9436
rect 13356 8754 13412 8764
rect 13468 8372 13524 13244
rect 13580 11732 13636 13356
rect 13580 11666 13636 11676
rect 13692 11620 13748 14112
rect 13916 12852 13972 12862
rect 13916 12758 13972 12796
rect 13916 11620 13972 11630
rect 13692 11618 13972 11620
rect 13692 11566 13918 11618
rect 13970 11566 13972 11618
rect 13692 11564 13972 11566
rect 13916 11554 13972 11564
rect 13468 8306 13524 8316
rect 13580 11394 13636 11406
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 13468 6020 13524 6030
rect 13580 6020 13636 11342
rect 14140 10836 14196 14112
rect 14364 14084 14420 14094
rect 14364 11508 14420 14028
rect 14588 12852 14644 14112
rect 14924 13076 14980 13086
rect 14924 12982 14980 13020
rect 14588 12786 14644 12796
rect 14812 12404 14868 12414
rect 15036 12404 15092 14112
rect 14812 12402 15092 12404
rect 14812 12350 14814 12402
rect 14866 12350 15092 12402
rect 14812 12348 15092 12350
rect 14812 12338 14868 12348
rect 14588 12180 14644 12190
rect 15036 12180 15092 12190
rect 14644 12124 15036 12180
rect 14588 12114 14644 12124
rect 15036 12114 15092 12124
rect 14140 10770 14196 10780
rect 14252 11452 14420 11508
rect 15372 12066 15428 12078
rect 15372 12014 15374 12066
rect 15426 12014 15428 12066
rect 14028 10498 14084 10510
rect 14028 10446 14030 10498
rect 14082 10446 14084 10498
rect 14028 7588 14084 10446
rect 14140 7588 14196 7598
rect 14028 7532 14140 7588
rect 14140 7522 14196 7532
rect 14252 7476 14308 11452
rect 14924 11396 14980 11406
rect 14252 7410 14308 7420
rect 14364 11394 14980 11396
rect 14364 11342 14926 11394
rect 14978 11342 14980 11394
rect 14364 11340 14980 11342
rect 13468 6018 13636 6020
rect 13468 5966 13470 6018
rect 13522 5966 13636 6018
rect 13468 5964 13636 5966
rect 13804 6804 13860 6814
rect 13468 5954 13524 5964
rect 13132 5460 13188 5470
rect 13132 5346 13188 5404
rect 13132 5294 13134 5346
rect 13186 5294 13188 5346
rect 13132 5282 13188 5294
rect 12572 5236 12628 5246
rect 12572 5142 12628 5180
rect 12124 2706 12180 2716
rect 12684 5124 12740 5134
rect 11228 1922 11284 1932
rect 11788 2212 11844 2222
rect 11788 1204 11844 2156
rect 12684 1764 12740 5068
rect 13468 5124 13524 5134
rect 13468 4900 13524 5068
rect 13468 4834 13524 4844
rect 13692 5010 13748 5022
rect 13692 4958 13694 5010
rect 13746 4958 13748 5010
rect 13244 4676 13300 4686
rect 13244 3220 13300 4620
rect 13692 4676 13748 4958
rect 13692 4610 13748 4620
rect 13804 4340 13860 6748
rect 14364 6018 14420 11340
rect 14924 11330 14980 11340
rect 15148 11060 15204 11070
rect 15204 11004 15316 11060
rect 15148 10994 15204 11004
rect 14588 10836 14644 10846
rect 14588 10742 14644 10780
rect 15260 10276 15316 11004
rect 15260 10210 15316 10220
rect 15372 9940 15428 12014
rect 15484 11618 15540 14112
rect 15484 11566 15486 11618
rect 15538 11566 15540 11618
rect 15484 11554 15540 11566
rect 15596 12962 15652 12974
rect 15596 12910 15598 12962
rect 15650 12910 15652 12962
rect 15596 10724 15652 12910
rect 15820 12628 15876 12638
rect 15596 10658 15652 10668
rect 15708 12066 15764 12078
rect 15708 12014 15710 12066
rect 15762 12014 15764 12066
rect 15372 9874 15428 9884
rect 15596 10498 15652 10510
rect 15596 10446 15598 10498
rect 15650 10446 15652 10498
rect 15484 9604 15540 9614
rect 14700 9492 14756 9502
rect 14700 7140 14756 9436
rect 14924 8484 14980 8494
rect 14700 7074 14756 7084
rect 14812 8372 14868 8382
rect 14924 8372 15204 8428
rect 14364 5966 14366 6018
rect 14418 5966 14420 6018
rect 14364 5954 14420 5966
rect 14812 5906 14868 8316
rect 15148 6132 15204 8372
rect 15484 8260 15540 9548
rect 15596 8484 15652 10446
rect 15596 8418 15652 8428
rect 15484 8194 15540 8204
rect 15708 6916 15764 12014
rect 15820 11508 15876 12572
rect 15932 12292 15988 14112
rect 16380 13076 16436 14112
rect 16380 13010 16436 13020
rect 15932 12226 15988 12236
rect 16044 12628 16100 12638
rect 15820 11442 15876 11452
rect 16044 9044 16100 12572
rect 16716 12404 16772 12414
rect 16828 12404 16884 14112
rect 16940 12962 16996 12974
rect 16940 12910 16942 12962
rect 16994 12910 16996 12962
rect 16940 12516 16996 12910
rect 17276 12964 17332 14112
rect 17612 13748 17668 13758
rect 17500 13076 17556 13086
rect 17500 12982 17556 13020
rect 17276 12908 17444 12964
rect 16940 12450 16996 12460
rect 16156 12348 16660 12404
rect 16156 12180 16212 12348
rect 16156 12114 16212 12124
rect 16492 12180 16548 12190
rect 16268 12068 16324 12078
rect 16044 8978 16100 8988
rect 16156 10498 16212 10510
rect 16156 10446 16158 10498
rect 16210 10446 16212 10498
rect 15708 6850 15764 6860
rect 15820 7028 15876 7038
rect 15148 6066 15204 6076
rect 14812 5854 14814 5906
rect 14866 5854 14868 5906
rect 14812 5842 14868 5854
rect 15036 6020 15092 6030
rect 15036 5908 15092 5964
rect 15036 5852 15316 5908
rect 14140 5796 14196 5806
rect 13804 4274 13860 4284
rect 13916 5682 13972 5694
rect 13916 5630 13918 5682
rect 13970 5630 13972 5682
rect 13244 3154 13300 3164
rect 13916 3108 13972 5630
rect 14140 5346 14196 5740
rect 15148 5682 15204 5694
rect 15148 5630 15150 5682
rect 15202 5630 15204 5682
rect 15148 5572 15204 5630
rect 14140 5294 14142 5346
rect 14194 5294 14196 5346
rect 14140 5282 14196 5294
rect 14924 5516 15204 5572
rect 14924 5124 14980 5516
rect 14812 5068 14980 5124
rect 13916 3042 13972 3052
rect 14476 4452 14532 4462
rect 14476 2772 14532 4396
rect 14252 2716 14532 2772
rect 12684 1698 12740 1708
rect 13132 2436 13188 2446
rect 13132 1540 13188 2380
rect 14252 2210 14308 2716
rect 14812 2436 14868 5068
rect 15092 5012 15148 5022
rect 14252 2158 14254 2210
rect 14306 2158 14308 2210
rect 14252 2146 14308 2158
rect 14364 2380 14868 2436
rect 14924 4956 15092 5012
rect 13692 2100 13748 2110
rect 13692 2006 13748 2044
rect 13132 1474 13188 1484
rect 11788 1138 11844 1148
rect 12572 980 12628 990
rect 12572 112 12628 924
rect 14364 980 14420 2380
rect 14700 2212 14756 2222
rect 14924 2212 14980 4956
rect 15092 4946 15148 4956
rect 15260 3780 15316 5852
rect 15708 5794 15764 5806
rect 15708 5742 15710 5794
rect 15762 5742 15764 5794
rect 15484 5684 15540 5694
rect 15484 5236 15540 5628
rect 15484 5170 15540 5180
rect 15708 5236 15764 5742
rect 15708 5170 15764 5180
rect 15036 3724 15316 3780
rect 15596 4228 15652 4238
rect 15036 3332 15092 3724
rect 15596 3666 15652 4172
rect 15596 3614 15598 3666
rect 15650 3614 15652 3666
rect 15596 3602 15652 3614
rect 15148 3556 15204 3566
rect 15148 3554 15316 3556
rect 15148 3502 15150 3554
rect 15202 3502 15316 3554
rect 15148 3500 15316 3502
rect 15148 3490 15204 3500
rect 15036 3276 15204 3332
rect 14756 2156 14980 2212
rect 14700 2146 14756 2156
rect 15036 1876 15092 1886
rect 14700 1820 15036 1876
rect 14364 914 14420 924
rect 14588 1764 14644 1774
rect 14588 868 14644 1708
rect 14700 1652 14756 1820
rect 15036 1810 15092 1820
rect 14700 1586 14756 1596
rect 15148 1204 15204 3276
rect 15148 1138 15204 1148
rect 14588 802 14644 812
rect 15260 112 15316 3500
rect 15820 3388 15876 6972
rect 16156 5684 16212 10446
rect 16268 6804 16324 12012
rect 16268 6738 16324 6748
rect 16380 11172 16436 11182
rect 16380 6132 16436 11116
rect 16492 10164 16548 12124
rect 16492 10098 16548 10108
rect 16380 6066 16436 6076
rect 16492 9828 16548 9838
rect 16604 9828 16660 12348
rect 16716 12402 16884 12404
rect 16716 12350 16718 12402
rect 16770 12350 16884 12402
rect 16716 12348 16884 12350
rect 16716 12338 16772 12348
rect 16940 12292 16996 12302
rect 16716 11844 16772 11854
rect 16716 11284 16772 11788
rect 16716 11218 16772 11228
rect 16828 11394 16884 11406
rect 16828 11342 16830 11394
rect 16882 11342 16884 11394
rect 16828 10612 16884 11342
rect 16940 10722 16996 12236
rect 17276 12068 17332 12078
rect 17276 11974 17332 12012
rect 17388 11618 17444 12908
rect 17388 11566 17390 11618
rect 17442 11566 17444 11618
rect 17388 11554 17444 11566
rect 16940 10670 16942 10722
rect 16994 10670 16996 10722
rect 16940 10658 16996 10670
rect 17164 10836 17220 10846
rect 16828 10546 16884 10556
rect 17052 10612 17108 10622
rect 17052 10500 17108 10556
rect 16940 10444 17108 10500
rect 16940 10388 16996 10444
rect 16828 10332 16996 10388
rect 16828 10276 16884 10332
rect 16828 10210 16884 10220
rect 17052 10276 17108 10286
rect 16940 10164 16996 10174
rect 16828 9940 16884 9950
rect 16828 9846 16884 9884
rect 16716 9828 16772 9838
rect 16604 9772 16716 9828
rect 16156 5618 16212 5628
rect 15932 5348 15988 5358
rect 15932 4788 15988 5292
rect 15932 4722 15988 4732
rect 16492 3668 16548 9772
rect 16716 9762 16772 9772
rect 16604 8708 16660 8718
rect 16604 6132 16660 8652
rect 16828 7476 16884 7486
rect 16828 7252 16884 7420
rect 16828 7186 16884 7196
rect 16940 6692 16996 10108
rect 16604 6066 16660 6076
rect 16716 6636 16996 6692
rect 16492 3602 16548 3612
rect 15708 3332 15876 3388
rect 15484 2324 15540 2334
rect 15484 868 15540 2268
rect 15708 1540 15764 3332
rect 16716 2100 16772 6636
rect 17052 6580 17108 10220
rect 17164 7252 17220 10780
rect 17388 10052 17444 10062
rect 17612 10052 17668 13692
rect 17724 12404 17780 14112
rect 17724 12338 17780 12348
rect 17836 13188 17892 13198
rect 17836 12068 17892 13132
rect 17836 12002 17892 12012
rect 18060 13188 18116 13198
rect 17388 10050 17668 10052
rect 17388 9998 17390 10050
rect 17442 9998 17668 10050
rect 17388 9996 17668 9998
rect 17948 10498 18004 10510
rect 17948 10446 17950 10498
rect 18002 10446 18004 10498
rect 17388 9986 17444 9996
rect 17948 8036 18004 10446
rect 17948 7970 18004 7980
rect 18060 7476 18116 13132
rect 18172 12290 18228 14112
rect 18396 13972 18452 13982
rect 18284 12964 18340 12974
rect 18284 12870 18340 12908
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18396 11620 18452 13916
rect 18620 13076 18676 14112
rect 18620 13010 18676 13020
rect 18844 13636 18900 13646
rect 18620 12740 18676 12750
rect 18396 11554 18452 11564
rect 18508 12404 18564 12414
rect 18508 10834 18564 12348
rect 18620 11394 18676 12684
rect 18844 12178 18900 13580
rect 18844 12126 18846 12178
rect 18898 12126 18900 12178
rect 18844 12114 18900 12126
rect 18620 11342 18622 11394
rect 18674 11342 18676 11394
rect 18620 11330 18676 11342
rect 19068 11282 19124 14112
rect 19292 12852 19348 12862
rect 19292 12758 19348 12796
rect 19516 12290 19572 14112
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 12226 19572 12238
rect 19628 13636 19684 13646
rect 19068 11230 19070 11282
rect 19122 11230 19124 11282
rect 19068 11218 19124 11230
rect 19404 12180 19460 12190
rect 18508 10782 18510 10834
rect 18562 10782 18564 10834
rect 18508 10770 18564 10782
rect 18620 10836 18676 10846
rect 18060 7410 18116 7420
rect 18284 10612 18340 10622
rect 17164 7186 17220 7196
rect 17052 6514 17108 6524
rect 17836 7140 17892 7150
rect 17836 6580 17892 7084
rect 17836 6514 17892 6524
rect 18060 7140 18116 7150
rect 16716 2034 16772 2044
rect 16940 6020 16996 6030
rect 15708 1474 15764 1484
rect 15484 802 15540 812
rect 16940 644 16996 5964
rect 17948 3668 18004 3678
rect 17836 1986 17892 1998
rect 17836 1934 17838 1986
rect 17890 1934 17892 1986
rect 17388 1874 17444 1886
rect 17388 1822 17390 1874
rect 17442 1822 17444 1874
rect 17388 1540 17444 1822
rect 17388 1474 17444 1484
rect 16940 578 16996 588
rect 17836 308 17892 1934
rect 17836 242 17892 252
rect 17948 112 18004 3612
rect 18060 3556 18116 7084
rect 18284 6020 18340 10556
rect 18396 9716 18452 9726
rect 18396 8036 18452 9660
rect 18396 7970 18452 7980
rect 18620 7700 18676 10780
rect 19068 9940 19124 9950
rect 18732 9716 18788 9726
rect 18732 9492 18788 9660
rect 18732 9426 18788 9436
rect 18396 7644 18676 7700
rect 18396 6356 18452 7644
rect 18956 7588 19012 7598
rect 18956 7494 19012 7532
rect 18396 6290 18452 6300
rect 18508 7476 18564 7486
rect 18284 5954 18340 5964
rect 18508 5572 18564 7420
rect 18172 5516 18564 5572
rect 18844 6804 18900 6814
rect 18172 4228 18228 5516
rect 18396 5348 18452 5358
rect 18172 4162 18228 4172
rect 18284 5124 18340 5134
rect 18060 3490 18116 3500
rect 18284 2884 18340 5068
rect 18396 4564 18452 5292
rect 18396 4498 18452 4508
rect 18732 5236 18788 5246
rect 18620 4228 18676 4238
rect 18508 4172 18620 4228
rect 18508 2996 18564 4172
rect 18620 4162 18676 4172
rect 18620 3554 18676 3566
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 3332 18676 3502
rect 18620 3266 18676 3276
rect 18508 2930 18564 2940
rect 18284 2818 18340 2828
rect 18396 1764 18452 1774
rect 18396 1092 18452 1708
rect 18396 1026 18452 1036
rect 18732 980 18788 5180
rect 18844 3220 18900 6748
rect 18844 3154 18900 3164
rect 18956 4788 19012 4798
rect 18844 980 18900 990
rect 18732 924 18844 980
rect 18844 914 18900 924
rect 18956 868 19012 4732
rect 18956 802 19012 812
rect 19068 532 19124 9884
rect 19404 7474 19460 12124
rect 19516 11732 19572 11742
rect 19516 7812 19572 11676
rect 19628 10722 19684 13580
rect 19964 12852 20020 14112
rect 19964 12786 20020 12796
rect 20188 13300 20244 13310
rect 20188 12068 20244 13244
rect 20188 12002 20244 12012
rect 20300 12628 20356 12638
rect 20076 11956 20132 11966
rect 20076 11732 20132 11900
rect 20076 11666 20132 11676
rect 19964 11394 20020 11406
rect 19964 11342 19966 11394
rect 20018 11342 20020 11394
rect 19852 11172 19908 11182
rect 19628 10670 19630 10722
rect 19682 10670 19684 10722
rect 19628 10658 19684 10670
rect 19740 10724 19796 10734
rect 19516 7746 19572 7756
rect 19628 8484 19684 8494
rect 19404 7422 19406 7474
rect 19458 7422 19460 7474
rect 19404 7410 19460 7422
rect 19628 6018 19684 8428
rect 19740 8260 19796 10668
rect 19852 10052 19908 11116
rect 19964 10164 20020 11342
rect 20300 11284 20356 12572
rect 20412 11620 20468 14112
rect 20636 13412 20692 13422
rect 20524 12292 20580 12302
rect 20524 11956 20580 12236
rect 20636 12178 20692 13356
rect 20860 12292 20916 14112
rect 21196 13188 21252 13198
rect 21196 13094 21252 13132
rect 20860 12226 20916 12236
rect 21084 12290 21140 12302
rect 21084 12238 21086 12290
rect 21138 12238 21140 12290
rect 20636 12126 20638 12178
rect 20690 12126 20692 12178
rect 20636 12114 20692 12126
rect 20524 11900 20692 11956
rect 20524 11620 20580 11630
rect 20412 11618 20580 11620
rect 20412 11566 20526 11618
rect 20578 11566 20580 11618
rect 20412 11564 20580 11566
rect 20524 11554 20580 11564
rect 20300 11218 20356 11228
rect 19964 10098 20020 10108
rect 20076 10386 20132 10398
rect 20076 10334 20078 10386
rect 20130 10334 20132 10386
rect 19852 9986 19908 9996
rect 19740 8194 19796 8204
rect 19964 8146 20020 8158
rect 19964 8094 19966 8146
rect 20018 8094 20020 8146
rect 19964 7924 20020 8094
rect 19964 7858 20020 7868
rect 19628 5966 19630 6018
rect 19682 5966 19684 6018
rect 19628 5954 19684 5966
rect 19740 7252 19796 7262
rect 19180 5684 19236 5694
rect 19180 4788 19236 5628
rect 19180 4722 19236 4732
rect 19180 3556 19236 3566
rect 19180 3462 19236 3500
rect 19740 1092 19796 7196
rect 20076 6916 20132 10334
rect 20524 10052 20580 10062
rect 20300 9714 20356 9726
rect 20300 9662 20302 9714
rect 20354 9662 20356 9714
rect 20300 9380 20356 9662
rect 20300 9314 20356 9324
rect 20524 8482 20580 9996
rect 20524 8430 20526 8482
rect 20578 8430 20580 8482
rect 20524 8418 20580 8430
rect 20636 8372 20692 11900
rect 21084 11284 21140 12238
rect 21084 11218 21140 11228
rect 21196 11844 21252 11854
rect 21084 10948 21140 10958
rect 20748 10612 20804 10622
rect 20804 10556 21028 10612
rect 20748 10546 20804 10556
rect 20860 9826 20916 9838
rect 20860 9774 20862 9826
rect 20914 9774 20916 9826
rect 20860 9156 20916 9774
rect 20972 9268 21028 10556
rect 21084 10610 21140 10892
rect 21084 10558 21086 10610
rect 21138 10558 21140 10610
rect 21084 10546 21140 10558
rect 21196 9940 21252 11788
rect 21308 11284 21364 14112
rect 21756 13188 21812 14112
rect 21756 13122 21812 13132
rect 21980 13860 22036 13870
rect 21756 12962 21812 12974
rect 21756 12910 21758 12962
rect 21810 12910 21812 12962
rect 21756 12852 21812 12910
rect 21756 12786 21812 12796
rect 21868 12740 21924 12750
rect 21868 12516 21924 12684
rect 21756 12460 21924 12516
rect 21756 11732 21812 12460
rect 21756 11666 21812 11676
rect 21868 12292 21924 12302
rect 21756 11284 21812 11294
rect 21308 11282 21812 11284
rect 21308 11230 21758 11282
rect 21810 11230 21812 11282
rect 21308 11228 21812 11230
rect 21756 11218 21812 11228
rect 21868 10722 21924 12236
rect 21980 12178 22036 13804
rect 22092 12964 22148 12974
rect 22092 12870 22148 12908
rect 22204 12404 22260 14112
rect 22652 13186 22708 14112
rect 22652 13134 22654 13186
rect 22706 13134 22708 13186
rect 22652 13122 22708 13134
rect 22316 12404 22372 12414
rect 22204 12402 22372 12404
rect 22204 12350 22318 12402
rect 22370 12350 22372 12402
rect 22204 12348 22372 12350
rect 22316 12338 22372 12348
rect 23100 12404 23156 14112
rect 23548 13524 23604 14112
rect 23548 13458 23604 13468
rect 23996 13188 24052 14112
rect 23996 13122 24052 13132
rect 24108 13524 24164 13534
rect 24108 12850 24164 13468
rect 24444 13524 24500 14112
rect 24444 13458 24500 13468
rect 24892 13412 24948 14112
rect 24464 13356 24728 13366
rect 24332 13300 24388 13310
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24892 13346 24948 13356
rect 24464 13290 24728 13300
rect 25004 13300 25060 13310
rect 24332 13188 24388 13244
rect 25004 13188 25060 13244
rect 24332 13132 25060 13188
rect 25228 13076 25284 13086
rect 25116 12964 25172 12974
rect 25116 12870 25172 12908
rect 24108 12798 24110 12850
rect 24162 12798 24164 12850
rect 24108 12786 24164 12798
rect 23100 12338 23156 12348
rect 23324 12628 23380 12638
rect 21980 12126 21982 12178
rect 22034 12126 22036 12178
rect 21980 12114 22036 12126
rect 23324 12178 23380 12572
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 23884 12404 23940 12414
rect 23884 12310 23940 12348
rect 24556 12180 24612 12190
rect 23324 12126 23326 12178
rect 23378 12126 23380 12178
rect 23324 12114 23380 12126
rect 23660 12124 24556 12180
rect 21868 10670 21870 10722
rect 21922 10670 21924 10722
rect 21868 10658 21924 10670
rect 22092 11508 22148 11518
rect 21196 9874 21252 9884
rect 22092 9716 22148 11452
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 10388 22820 11342
rect 22764 10322 22820 10332
rect 23324 11284 23380 11294
rect 22092 9650 22148 9660
rect 20972 9202 21028 9212
rect 22316 9604 22372 9614
rect 20860 9090 20916 9100
rect 21980 8708 22036 8718
rect 21196 8372 21252 8382
rect 20636 8316 21196 8372
rect 21196 8306 21252 8316
rect 21532 8260 21588 8270
rect 21532 8166 21588 8204
rect 19740 1026 19796 1036
rect 19964 6860 20132 6916
rect 20972 7588 21028 7598
rect 19068 466 19124 476
rect 19964 196 20020 6860
rect 20748 6692 20804 6702
rect 20748 6578 20804 6636
rect 20748 6526 20750 6578
rect 20802 6526 20804 6578
rect 20748 6514 20804 6526
rect 20972 6244 21028 7532
rect 21868 7252 21924 7262
rect 20972 6178 21028 6188
rect 21196 6690 21252 6702
rect 21196 6638 21198 6690
rect 21250 6638 21252 6690
rect 20076 5684 20132 5694
rect 20076 5682 20356 5684
rect 20076 5630 20078 5682
rect 20130 5630 20356 5682
rect 20076 5628 20356 5630
rect 20076 5618 20132 5628
rect 20076 3332 20132 3342
rect 20076 1428 20132 3276
rect 20188 2884 20244 2894
rect 20188 1540 20244 2828
rect 20188 1474 20244 1484
rect 20076 1362 20132 1372
rect 20300 1428 20356 5628
rect 21196 5236 21252 6638
rect 21868 6468 21924 7196
rect 21980 7140 22036 8652
rect 21980 7074 22036 7084
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 21868 6402 21924 6412
rect 22092 6020 22148 8206
rect 22316 6244 22372 9548
rect 22540 9268 22596 9278
rect 22428 8932 22484 8942
rect 22428 8838 22484 8876
rect 22540 7140 22596 9212
rect 23324 9268 23380 11228
rect 23436 9940 23492 9950
rect 23436 9846 23492 9884
rect 23660 9716 23716 12124
rect 24556 12114 24612 12124
rect 24332 11844 24388 11854
rect 24332 11620 24388 11788
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24332 11564 24724 11620
rect 24444 11396 24500 11406
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 24444 10948 24500 11340
rect 24444 10882 24500 10892
rect 24556 11394 24612 11406
rect 24556 11342 24558 11394
rect 24610 11342 24612 11394
rect 24556 10388 24612 11342
rect 24668 10500 24724 11564
rect 25116 11508 25172 11518
rect 25228 11508 25284 13020
rect 25116 11506 25284 11508
rect 25116 11454 25118 11506
rect 25170 11454 25284 11506
rect 25116 11452 25284 11454
rect 25116 11442 25172 11452
rect 24668 10434 24724 10444
rect 25228 10836 25284 10846
rect 24332 10332 24612 10388
rect 24332 10276 24388 10332
rect 24892 10276 24948 10286
rect 24332 10210 24388 10220
rect 24464 10220 24728 10230
rect 24108 10164 24164 10174
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 24108 10052 24164 10108
rect 24892 10052 24948 10220
rect 24108 9996 24948 10052
rect 23996 9940 24052 9950
rect 23996 9846 24052 9884
rect 23324 9202 23380 9212
rect 23548 9660 23716 9716
rect 24892 9828 24948 9838
rect 22988 8818 23044 8830
rect 22988 8766 22990 8818
rect 23042 8766 23044 8818
rect 22988 8484 23044 8766
rect 23548 8596 23604 9660
rect 23660 9492 23716 9502
rect 23660 9268 23716 9436
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24220 9380 24276 9390
rect 24220 9268 24276 9324
rect 23660 9212 24276 9268
rect 23548 8530 23604 8540
rect 24332 8708 24388 8718
rect 22988 8418 23044 8428
rect 24332 8398 24388 8652
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24892 8596 24948 9772
rect 25228 9492 25284 10780
rect 25340 10500 25396 14112
rect 25452 13188 25508 13198
rect 25452 13094 25508 13132
rect 25564 12964 25620 12974
rect 25452 12068 25508 12078
rect 25452 10836 25508 12012
rect 25452 10770 25508 10780
rect 25340 10444 25508 10500
rect 25228 9426 25284 9436
rect 25340 9828 25396 9838
rect 25228 9044 25284 9054
rect 24892 8530 24948 8540
rect 25004 8708 25060 8718
rect 25004 8398 25060 8652
rect 24332 8342 25060 8398
rect 23548 7980 24388 8036
rect 23548 7924 23604 7980
rect 24332 7924 24388 7980
rect 23548 7858 23604 7868
rect 23804 7868 24068 7878
rect 23660 7812 23716 7822
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24332 7858 24388 7868
rect 23804 7802 24068 7812
rect 24220 7812 24276 7822
rect 23660 7700 23716 7756
rect 24220 7700 24276 7756
rect 23660 7644 24276 7700
rect 24780 7700 24836 7710
rect 24836 7644 24948 7700
rect 24780 7634 24836 7644
rect 22540 7074 22596 7084
rect 23660 7364 23716 7374
rect 23660 7028 23716 7308
rect 23660 6962 23716 6972
rect 24332 7140 24388 7150
rect 24892 7140 24948 7644
rect 25116 7140 25172 7150
rect 22092 5954 22148 5964
rect 22204 6188 22372 6244
rect 23548 6690 23604 6702
rect 23548 6638 23550 6690
rect 23602 6638 23604 6690
rect 22204 5796 22260 6188
rect 21868 5740 22260 5796
rect 21196 5170 21252 5180
rect 21644 5348 21700 5358
rect 21532 4564 21588 4574
rect 21532 3780 21588 4508
rect 21532 3714 21588 3724
rect 21420 3220 21476 3230
rect 21420 2996 21476 3164
rect 21644 3220 21700 5292
rect 21756 4340 21812 4350
rect 21756 3780 21812 4284
rect 21756 3714 21812 3724
rect 21644 3154 21700 3164
rect 21420 2930 21476 2940
rect 21868 2884 21924 5740
rect 21868 2818 21924 2828
rect 21980 5348 22036 5358
rect 21532 2660 21588 2670
rect 21532 2566 21588 2604
rect 21756 2660 21812 2670
rect 21756 2458 21812 2604
rect 21420 2402 21812 2458
rect 21308 2212 21364 2222
rect 21420 2212 21476 2402
rect 21980 2324 22036 5292
rect 22204 5348 22260 5358
rect 22092 4340 22148 4350
rect 22092 2882 22148 4284
rect 22092 2830 22094 2882
rect 22146 2830 22148 2882
rect 22092 2818 22148 2830
rect 22204 2324 22260 5292
rect 23548 4452 23604 6638
rect 23996 6692 24052 6702
rect 23996 6598 24052 6636
rect 23804 6300 24068 6310
rect 23660 6244 23716 6254
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24220 6244 24276 6254
rect 23660 5124 23716 6188
rect 24220 5460 24276 6188
rect 24332 5908 24388 7084
rect 24464 7084 24728 7094
rect 24892 7084 25116 7140
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 25116 7074 25172 7084
rect 24464 7018 24728 7028
rect 25228 6468 25284 8988
rect 25228 6402 25284 6412
rect 24332 5842 24388 5852
rect 25116 6020 25172 6030
rect 24332 5628 24948 5684
rect 24332 5572 24388 5628
rect 24892 5572 24948 5628
rect 24332 5506 24388 5516
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24892 5506 24948 5516
rect 24464 5450 24728 5460
rect 24220 5394 24276 5404
rect 23660 5068 24388 5124
rect 23660 4788 23716 4798
rect 24332 4788 24388 5068
rect 23660 4452 23716 4732
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24332 4722 24388 4732
rect 25116 4788 25172 5964
rect 25116 4722 25172 4732
rect 25228 5908 25284 5918
rect 23804 4666 24068 4676
rect 24220 4676 24276 4686
rect 23772 4452 23828 4462
rect 23660 4396 23772 4452
rect 23548 4386 23604 4396
rect 23772 4386 23828 4396
rect 21980 2268 22148 2324
rect 21308 2210 21476 2212
rect 21308 2158 21310 2210
rect 21362 2158 21476 2210
rect 21308 2156 21476 2158
rect 21308 2146 21364 2156
rect 21980 2100 22036 2110
rect 20748 1876 20804 1886
rect 20748 1782 20804 1820
rect 20300 1362 20356 1372
rect 19964 130 20020 140
rect 20636 1204 20692 1214
rect 20636 112 20692 1148
rect 20860 1204 20916 1214
rect 20860 980 20916 1148
rect 20860 914 20916 924
rect 21980 420 22036 2044
rect 21980 354 22036 364
rect 1148 18 1204 28
rect 1792 0 1904 112
rect 4480 0 4592 112
rect 7168 0 7280 112
rect 9856 0 9968 112
rect 12544 0 12656 112
rect 15232 0 15344 112
rect 17920 0 18032 112
rect 20608 0 20720 112
rect 22092 84 22148 2268
rect 22204 2258 22260 2268
rect 23660 4116 23716 4126
rect 23660 2212 23716 4060
rect 23884 4116 23940 4126
rect 23884 3780 23940 4060
rect 24220 4004 24276 4620
rect 24220 3938 24276 3948
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 24220 3780 24276 3790
rect 23884 3714 23940 3724
rect 23996 3724 24220 3780
rect 23996 3668 24052 3724
rect 24220 3714 24276 3724
rect 23996 3602 24052 3612
rect 25228 3388 25284 5852
rect 25340 5012 25396 9772
rect 25340 4946 25396 4956
rect 25228 3332 25396 3388
rect 24332 3220 24388 3230
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24332 2996 24388 3164
rect 23884 2940 24388 2996
rect 24444 3108 24500 3118
rect 23884 2436 23940 2940
rect 24444 2884 24500 3052
rect 23996 2828 24500 2884
rect 24668 2884 24724 2894
rect 23996 2772 24052 2828
rect 23996 2706 24052 2716
rect 24668 2660 24724 2828
rect 24668 2594 24724 2604
rect 24892 2658 24948 2670
rect 24892 2606 24894 2658
rect 24946 2606 24948 2658
rect 23884 2370 23940 2380
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24892 2324 24948 2606
rect 25116 2436 25172 2446
rect 24892 2258 24948 2268
rect 25004 2380 25116 2436
rect 24556 2212 24612 2222
rect 23660 2210 24612 2212
rect 23660 2158 24558 2210
rect 24610 2158 24612 2210
rect 23660 2156 24612 2158
rect 24556 2146 24612 2156
rect 24780 2100 24836 2110
rect 24780 1652 24836 2044
rect 23804 1596 24068 1606
rect 23660 1540 23716 1550
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24780 1586 24836 1596
rect 23804 1530 24068 1540
rect 24332 1540 24388 1550
rect 23660 1428 23716 1484
rect 24332 1428 24388 1484
rect 25004 1540 25060 2380
rect 25116 2370 25172 2380
rect 25116 2100 25172 2110
rect 25116 2006 25172 2044
rect 25004 1474 25060 1484
rect 25228 1764 25284 1774
rect 25228 1540 25284 1708
rect 25228 1474 25284 1484
rect 23660 1372 24388 1428
rect 22988 1316 23044 1326
rect 22988 868 23044 1260
rect 22988 802 23044 812
rect 24464 812 24728 822
rect 23324 756 23380 766
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 23324 112 23380 700
rect 22092 18 22148 28
rect 23296 0 23408 112
rect 25340 84 25396 3332
rect 25452 2770 25508 10444
rect 25564 9938 25620 12908
rect 25788 12068 25844 14112
rect 25788 12002 25844 12012
rect 25900 13972 25956 13982
rect 25900 10612 25956 13916
rect 26012 13412 26068 13422
rect 26012 11620 26068 13356
rect 26124 12516 26180 12526
rect 26124 11844 26180 12460
rect 26124 11778 26180 11788
rect 26012 11554 26068 11564
rect 25900 10546 25956 10556
rect 26124 11508 26180 11518
rect 25564 9886 25566 9938
rect 25618 9886 25620 9938
rect 25564 9874 25620 9886
rect 25676 10500 25732 10510
rect 25564 9604 25620 9614
rect 25564 9044 25620 9548
rect 25564 8978 25620 8988
rect 25564 8484 25620 8494
rect 25564 8260 25620 8428
rect 25564 8194 25620 8204
rect 25564 7924 25620 7934
rect 25564 4004 25620 7868
rect 25564 3938 25620 3948
rect 25452 2718 25454 2770
rect 25506 2718 25508 2770
rect 25452 2706 25508 2718
rect 25564 3332 25620 3342
rect 25564 868 25620 3276
rect 25676 1988 25732 10444
rect 26124 10050 26180 11452
rect 26236 11284 26292 14112
rect 26684 13412 26740 14112
rect 26684 13346 26740 13356
rect 27132 13188 27188 14112
rect 27468 13860 27524 13870
rect 27244 13188 27300 13198
rect 27132 13132 27244 13188
rect 27244 13122 27300 13132
rect 27020 12628 27076 12638
rect 27020 12180 27076 12572
rect 27020 12114 27076 12124
rect 26236 11218 26292 11228
rect 27356 11954 27412 11966
rect 27356 11902 27358 11954
rect 27410 11902 27412 11954
rect 26796 10052 26852 10062
rect 26124 9998 26126 10050
rect 26178 9998 26180 10050
rect 26124 9986 26180 9998
rect 26460 9996 26796 10052
rect 26460 9716 26516 9996
rect 26796 9986 26852 9996
rect 26460 9650 26516 9660
rect 27356 9716 27412 11902
rect 27468 11732 27524 13804
rect 27580 12180 27636 14112
rect 27916 13412 27972 13422
rect 27916 12516 27972 13356
rect 27916 12450 27972 12460
rect 27916 12292 27972 12302
rect 27916 12198 27972 12236
rect 27580 12114 27636 12124
rect 28028 11844 28084 14112
rect 28028 11778 28084 11788
rect 28252 13300 28308 13310
rect 27468 11666 27524 11676
rect 27356 9650 27412 9660
rect 27804 11620 27860 11630
rect 27244 9604 27300 9614
rect 26908 9380 26964 9390
rect 26684 9324 26908 9380
rect 26684 8036 26740 9324
rect 26908 9314 26964 9324
rect 26684 7970 26740 7980
rect 26796 9156 26852 9166
rect 26796 7924 26852 9100
rect 26796 7858 26852 7868
rect 26908 8036 26964 8046
rect 26796 6580 26852 6590
rect 26796 5572 26852 6524
rect 26908 6132 26964 7980
rect 27132 7028 27188 7038
rect 27132 6356 27188 6972
rect 27132 6290 27188 6300
rect 26908 6066 26964 6076
rect 26796 5516 27188 5572
rect 25788 5236 25844 5246
rect 25788 2212 25844 5180
rect 26572 5236 26628 5246
rect 26572 4228 26628 5180
rect 26572 4162 26628 4172
rect 26012 4116 26068 4126
rect 25900 3668 25956 3678
rect 25900 2548 25956 3612
rect 26012 2772 26068 4060
rect 26012 2706 26068 2716
rect 27020 3556 27076 3566
rect 25900 2482 25956 2492
rect 26348 2548 26404 2558
rect 25788 2156 26292 2212
rect 25676 1932 26068 1988
rect 25900 1764 25956 1774
rect 25900 1092 25956 1708
rect 26012 1316 26068 1932
rect 26012 1250 26068 1260
rect 26236 1204 26292 2156
rect 26236 1138 26292 1148
rect 25900 1026 25956 1036
rect 25564 802 25620 812
rect 26348 644 26404 2492
rect 27020 2212 27076 3500
rect 27132 2436 27188 5516
rect 27244 4452 27300 9548
rect 27692 9492 27748 9502
rect 27692 6020 27748 9436
rect 27804 6580 27860 11564
rect 28028 11284 28084 11294
rect 27916 10724 27972 10734
rect 27916 7812 27972 10668
rect 27916 7746 27972 7756
rect 27804 6514 27860 6524
rect 27692 5954 27748 5964
rect 27916 5010 27972 5022
rect 27916 4958 27918 5010
rect 27970 4958 27972 5010
rect 27916 4900 27972 4958
rect 27916 4834 27972 4844
rect 27244 4386 27300 4396
rect 27804 4788 27860 4798
rect 27580 4116 27636 4126
rect 27580 3556 27636 4060
rect 27804 4116 27860 4732
rect 28028 4788 28084 11228
rect 28252 11284 28308 13244
rect 28364 12404 28420 12414
rect 28364 11396 28420 12348
rect 28364 11330 28420 11340
rect 28252 11218 28308 11228
rect 28476 10500 28532 14112
rect 28700 13412 28756 13422
rect 28588 12852 28644 12862
rect 28588 12290 28644 12796
rect 28588 12238 28590 12290
rect 28642 12238 28644 12290
rect 28588 12226 28644 12238
rect 28476 10434 28532 10444
rect 28588 11956 28644 11966
rect 28476 10276 28532 10286
rect 28364 10164 28420 10174
rect 28364 9940 28420 10108
rect 28364 9874 28420 9884
rect 28140 9380 28196 9390
rect 28140 5908 28196 9324
rect 28476 9044 28532 10220
rect 28476 8978 28532 8988
rect 28476 8820 28532 8830
rect 28140 5842 28196 5852
rect 28364 8484 28420 8494
rect 28364 5908 28420 8428
rect 28476 7476 28532 8764
rect 28476 7410 28532 7420
rect 28364 5842 28420 5852
rect 28476 5348 28532 5358
rect 28588 5348 28644 11900
rect 28700 10052 28756 13356
rect 28924 12852 28980 14112
rect 28924 12786 28980 12796
rect 29148 12628 29204 12638
rect 28812 12068 28868 12078
rect 28812 11060 28868 12012
rect 29036 12068 29092 12078
rect 29036 11974 29092 12012
rect 28924 11844 28980 11854
rect 28924 11620 28980 11788
rect 29148 11844 29204 12572
rect 29372 12628 29428 14112
rect 29372 12562 29428 12572
rect 29820 12404 29876 14112
rect 29820 12338 29876 12348
rect 30044 12516 30100 12526
rect 29148 11778 29204 11788
rect 29932 12292 29988 12302
rect 30044 12292 30100 12460
rect 30268 12516 30324 14112
rect 30716 14084 30772 14112
rect 30716 14018 30772 14028
rect 30268 12450 30324 12460
rect 31052 12852 31108 12862
rect 30156 12292 30212 12302
rect 30044 12236 30156 12292
rect 28924 11554 28980 11564
rect 28812 10994 28868 11004
rect 28700 9986 28756 9996
rect 28812 10500 28868 10510
rect 29036 10500 29092 10510
rect 28812 9940 28868 10444
rect 28812 9874 28868 9884
rect 28924 10444 29036 10500
rect 28700 9156 28756 9166
rect 28700 8372 28756 9100
rect 28700 8306 28756 8316
rect 28476 5346 28644 5348
rect 28476 5294 28478 5346
rect 28530 5294 28644 5346
rect 28476 5292 28644 5294
rect 28700 6244 28756 6254
rect 28476 5282 28532 5292
rect 28028 4722 28084 4732
rect 28700 4564 28756 6188
rect 28812 6132 28868 6142
rect 28924 6132 28980 10444
rect 29036 10434 29092 10444
rect 29820 10052 29876 10062
rect 29708 8820 29764 8830
rect 29708 7028 29764 8764
rect 29820 7812 29876 9996
rect 29820 7746 29876 7756
rect 29708 6962 29764 6972
rect 28868 6076 28980 6132
rect 28812 6066 28868 6076
rect 29932 6020 29988 12236
rect 30156 12226 30212 12236
rect 30268 12180 30324 12190
rect 30044 9492 30100 9502
rect 30044 8036 30100 9436
rect 30044 7970 30100 7980
rect 30156 8372 30212 8382
rect 29932 5954 29988 5964
rect 29260 5908 29316 5918
rect 29708 5908 29764 5918
rect 29316 5852 29708 5908
rect 29260 5842 29316 5852
rect 29708 5842 29764 5852
rect 29148 5796 29204 5806
rect 28700 4498 28756 4508
rect 29036 5684 29092 5694
rect 27804 4050 27860 4060
rect 27580 3490 27636 3500
rect 28700 3444 28756 3454
rect 28588 2882 28644 2894
rect 28588 2830 28590 2882
rect 28642 2830 28644 2882
rect 28588 2660 28644 2830
rect 28588 2594 28644 2604
rect 28700 2548 28756 3388
rect 28700 2482 28756 2492
rect 28924 3332 28980 3342
rect 27132 2370 27188 2380
rect 28476 2324 28532 2334
rect 27020 2156 27300 2212
rect 26348 578 26404 588
rect 26796 1428 26852 1438
rect 27132 1428 27188 1438
rect 26796 420 26852 1372
rect 26908 1372 27132 1428
rect 26908 756 26964 1372
rect 27132 1362 27188 1372
rect 26908 690 26964 700
rect 27244 756 27300 2156
rect 28476 1428 28532 2268
rect 28924 2210 28980 3276
rect 29036 3220 29092 5628
rect 29036 3154 29092 3164
rect 28924 2158 28926 2210
rect 28978 2158 28980 2210
rect 28924 2146 28980 2158
rect 29036 2546 29092 2558
rect 29036 2494 29038 2546
rect 29090 2494 29092 2546
rect 28476 1362 28532 1372
rect 29036 1428 29092 2494
rect 29036 1362 29092 1372
rect 27244 690 27300 700
rect 28924 1316 28980 1326
rect 26796 354 26852 364
rect 28924 420 28980 1260
rect 29148 1316 29204 5740
rect 29484 4788 29540 4798
rect 29484 3108 29540 4732
rect 29484 3042 29540 3052
rect 29372 2996 29428 3006
rect 29372 1652 29428 2940
rect 30156 2884 30212 8316
rect 30268 8260 30324 12124
rect 30828 11844 30884 11854
rect 30380 11732 30436 11742
rect 30436 11676 30660 11732
rect 30380 11666 30436 11676
rect 30492 10948 30548 10958
rect 30268 8194 30324 8204
rect 30380 9716 30436 9726
rect 30380 6804 30436 9660
rect 30492 9604 30548 10892
rect 30492 9538 30548 9548
rect 30380 6738 30436 6748
rect 30492 9156 30548 9166
rect 30492 6468 30548 9100
rect 30604 8484 30660 11676
rect 30604 8418 30660 8428
rect 30716 10948 30772 10958
rect 30604 7476 30660 7486
rect 30604 7382 30660 7420
rect 30716 7028 30772 10892
rect 30828 8820 30884 11788
rect 30940 11620 30996 11630
rect 30940 11526 30996 11564
rect 30828 8754 30884 8764
rect 30716 6962 30772 6972
rect 30828 7140 30884 7150
rect 30268 6412 30548 6468
rect 30604 6804 30660 6814
rect 30268 6356 30324 6412
rect 30604 6356 30660 6748
rect 30268 6290 30324 6300
rect 30380 6300 30660 6356
rect 30716 6580 30772 6590
rect 30380 6132 30436 6300
rect 30380 6066 30436 6076
rect 30604 6132 30660 6142
rect 30380 5908 30436 5918
rect 30380 5814 30436 5852
rect 30268 5236 30324 5246
rect 30268 4676 30324 5180
rect 30268 4610 30324 4620
rect 30156 2818 30212 2828
rect 30268 3668 30324 3678
rect 29484 2660 29540 2670
rect 29484 2098 29540 2604
rect 29484 2046 29486 2098
rect 29538 2046 29540 2098
rect 29484 2034 29540 2046
rect 30268 1876 30324 3612
rect 30268 1810 30324 1820
rect 30492 1874 30548 1886
rect 30492 1822 30494 1874
rect 30546 1822 30548 1874
rect 29372 1586 29428 1596
rect 29148 1250 29204 1260
rect 30268 644 30324 654
rect 30268 478 30324 588
rect 30492 644 30548 1822
rect 30604 1764 30660 6076
rect 30716 2548 30772 6524
rect 30716 2482 30772 2492
rect 30604 1698 30660 1708
rect 30828 1652 30884 7084
rect 30940 7028 30996 7038
rect 30940 6018 30996 6972
rect 30940 5966 30942 6018
rect 30994 5966 30996 6018
rect 30940 5954 30996 5966
rect 31052 4900 31108 12796
rect 31164 11956 31220 14112
rect 31164 11890 31220 11900
rect 31500 13188 31556 13198
rect 31388 11282 31444 11294
rect 31388 11230 31390 11282
rect 31442 11230 31444 11282
rect 31388 11172 31444 11230
rect 31388 11106 31444 11116
rect 31500 10052 31556 13132
rect 31612 11732 31668 14112
rect 31724 13860 31780 13870
rect 31724 13188 31780 13804
rect 31724 13122 31780 13132
rect 31612 11676 32004 11732
rect 31836 10612 31892 10622
rect 31500 9986 31556 9996
rect 31724 10276 31780 10286
rect 31724 9828 31780 10220
rect 31836 9940 31892 10556
rect 31836 9874 31892 9884
rect 31724 9762 31780 9772
rect 31948 9828 32004 11676
rect 31948 9762 32004 9772
rect 32060 8372 32116 14112
rect 32284 13636 32340 13646
rect 32284 11620 32340 13580
rect 32284 11554 32340 11564
rect 32396 12180 32452 12190
rect 32060 8306 32116 8316
rect 32172 9604 32228 9614
rect 31164 7364 31220 7402
rect 31164 7298 31220 7308
rect 31164 7140 31220 7150
rect 31164 6804 31220 7084
rect 31164 6738 31220 6748
rect 31836 6804 31892 6814
rect 31724 5796 31780 5806
rect 31724 5702 31780 5740
rect 31052 4834 31108 4844
rect 31612 5124 31668 5134
rect 31612 4676 31668 5068
rect 31612 4610 31668 4620
rect 31836 4116 31892 6748
rect 31836 4050 31892 4060
rect 32172 3388 32228 9548
rect 32284 8932 32340 8942
rect 32284 6580 32340 8876
rect 32396 8484 32452 12124
rect 32508 11844 32564 14112
rect 32508 11778 32564 11788
rect 32732 12180 32788 12190
rect 32732 10500 32788 12124
rect 32732 10434 32788 10444
rect 32620 8484 32676 8494
rect 32396 8428 32620 8484
rect 32620 8418 32676 8428
rect 32284 6514 32340 6524
rect 32620 8260 32676 8270
rect 32284 5682 32340 5694
rect 32284 5630 32286 5682
rect 32338 5630 32340 5682
rect 32284 4564 32340 5630
rect 32284 4498 32340 4508
rect 32396 3442 32452 3454
rect 32396 3390 32398 3442
rect 32450 3390 32452 3442
rect 32172 3332 32340 3388
rect 32284 2770 32340 3332
rect 32396 3332 32452 3390
rect 32620 3388 32676 8204
rect 32844 8036 32900 8046
rect 32732 7924 32788 7934
rect 32732 7140 32788 7868
rect 32732 7074 32788 7084
rect 32844 4900 32900 7980
rect 32956 7812 33012 14112
rect 32956 7746 33012 7756
rect 33180 12292 33236 12302
rect 33180 7476 33236 12236
rect 33404 10500 33460 14112
rect 32844 4834 32900 4844
rect 33068 7420 33236 7476
rect 33292 10444 33460 10500
rect 33628 12852 33684 12862
rect 32956 3780 33012 3790
rect 33068 3780 33124 7420
rect 33292 6804 33348 10444
rect 33628 10388 33684 12796
rect 33292 6738 33348 6748
rect 33404 10332 33684 10388
rect 33292 4116 33348 4126
rect 33292 3892 33348 4060
rect 33292 3826 33348 3836
rect 32956 3778 33124 3780
rect 32956 3726 32958 3778
rect 33010 3726 33124 3778
rect 32956 3724 33124 3726
rect 32956 3714 33012 3724
rect 33404 3556 33460 10332
rect 33628 10164 33684 10174
rect 33628 9604 33684 10108
rect 33628 9538 33684 9548
rect 33852 9156 33908 14112
rect 34300 10948 34356 14112
rect 34748 13748 34804 14112
rect 35196 13972 35252 14112
rect 35196 13906 35252 13916
rect 34748 13682 34804 13692
rect 35084 13300 35140 13310
rect 34860 12628 34916 12638
rect 34636 11844 34692 11854
rect 34300 10882 34356 10892
rect 34412 11394 34468 11406
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 34412 10836 34468 11342
rect 34412 10770 34468 10780
rect 34524 10948 34580 10958
rect 33852 9090 33908 9100
rect 34412 9268 34468 9278
rect 33516 8596 33572 8606
rect 33516 5796 33572 8540
rect 33628 8484 33684 8494
rect 33628 7700 33684 8428
rect 33852 8484 33908 8494
rect 33740 7700 33796 7710
rect 33628 7644 33740 7700
rect 33740 7634 33796 7644
rect 33516 5740 33796 5796
rect 33628 5572 33684 5582
rect 33628 5012 33684 5516
rect 33628 4946 33684 4956
rect 33404 3490 33460 3500
rect 33516 3892 33572 3902
rect 32620 3332 32788 3388
rect 32396 3266 32452 3276
rect 32732 3266 32788 3276
rect 32844 2884 32900 2894
rect 32844 2790 32900 2828
rect 32284 2718 32286 2770
rect 32338 2718 32340 2770
rect 32284 2706 32340 2718
rect 33516 2324 33572 3836
rect 33740 3220 33796 5740
rect 33852 4452 33908 8428
rect 33852 4386 33908 4396
rect 34412 4116 34468 9212
rect 34412 4050 34468 4060
rect 33740 3154 33796 3164
rect 34188 3556 34244 3566
rect 34188 3108 34244 3500
rect 34188 3042 34244 3052
rect 34412 3108 34468 3118
rect 33516 2258 33572 2268
rect 30940 1988 30996 1998
rect 30940 1894 30996 1932
rect 34076 1988 34132 1998
rect 30828 1586 30884 1596
rect 30940 1764 30996 1774
rect 30492 578 30548 588
rect 30940 478 30996 1708
rect 32620 1764 32676 1774
rect 32676 1708 33012 1764
rect 32620 1698 32676 1708
rect 32956 1540 33012 1708
rect 32956 1474 33012 1484
rect 30268 422 30996 478
rect 31388 1316 31444 1326
rect 28924 354 28980 364
rect 25676 252 26068 308
rect 25676 84 25732 252
rect 26012 112 26068 252
rect 28700 196 28756 206
rect 28700 112 28756 140
rect 31388 112 31444 1260
rect 31612 1316 31668 1326
rect 31612 196 31668 1260
rect 31612 130 31668 140
rect 33628 1204 33684 1214
rect 33628 196 33684 1148
rect 33628 130 33684 140
rect 34076 112 34132 1932
rect 34412 1092 34468 3052
rect 34524 1316 34580 10892
rect 34636 8482 34692 11788
rect 34860 11172 34916 12572
rect 35084 11396 35140 13244
rect 35532 13076 35588 13086
rect 35308 12068 35364 12078
rect 35084 11330 35140 11340
rect 35196 11956 35252 11966
rect 34860 11106 34916 11116
rect 34972 11282 35028 11294
rect 34972 11230 34974 11282
rect 35026 11230 35028 11282
rect 34748 10836 34804 10846
rect 34748 9268 34804 10780
rect 34972 10052 35028 11230
rect 34972 9986 35028 9996
rect 34748 9202 34804 9212
rect 34636 8430 34638 8482
rect 34690 8430 34692 8482
rect 34636 8418 34692 8430
rect 34748 9044 34804 9054
rect 34636 8260 34692 8270
rect 34636 2212 34692 8204
rect 34748 4452 34804 8988
rect 34972 9044 35028 9054
rect 34972 8708 35028 8988
rect 34972 8642 35028 8652
rect 35084 8148 35140 8158
rect 35084 8054 35140 8092
rect 35084 7924 35140 7934
rect 34972 6692 35028 6702
rect 34748 4386 34804 4396
rect 34860 5348 34916 5358
rect 34748 3780 34804 3790
rect 34748 3666 34804 3724
rect 34748 3614 34750 3666
rect 34802 3614 34804 3666
rect 34748 3602 34804 3614
rect 34860 2772 34916 5292
rect 34860 2706 34916 2716
rect 34972 2660 35028 6636
rect 35084 6132 35140 7868
rect 35084 6066 35140 6076
rect 35084 5796 35140 5806
rect 35084 4116 35140 5740
rect 35084 4050 35140 4060
rect 35196 3554 35252 11900
rect 35308 8148 35364 12012
rect 35532 11284 35588 13020
rect 35532 11218 35588 11228
rect 35308 8082 35364 8092
rect 35420 9268 35476 9278
rect 35420 7028 35476 9212
rect 35532 8596 35588 8606
rect 35532 8036 35588 8540
rect 35644 8260 35700 14112
rect 35868 13076 35924 13086
rect 35644 8194 35700 8204
rect 35756 12404 35812 12414
rect 35532 7980 35700 8036
rect 35532 7812 35588 7822
rect 35532 7252 35588 7756
rect 35532 7186 35588 7196
rect 35420 6962 35476 6972
rect 35420 6132 35476 6142
rect 35308 5236 35364 5246
rect 35308 5012 35364 5180
rect 35308 4946 35364 4956
rect 35308 4676 35364 4686
rect 35308 3780 35364 4620
rect 35308 3714 35364 3724
rect 35196 3502 35198 3554
rect 35250 3502 35252 3554
rect 35196 3490 35252 3502
rect 35308 3220 35364 3230
rect 34972 2594 35028 2604
rect 35196 2660 35252 2670
rect 34636 2146 34692 2156
rect 34524 1250 34580 1260
rect 34412 1026 34468 1036
rect 35196 756 35252 2604
rect 35308 1204 35364 3164
rect 35420 2884 35476 6076
rect 35532 5908 35588 5918
rect 35532 4676 35588 5852
rect 35532 4610 35588 4620
rect 35420 2818 35476 2828
rect 35308 1138 35364 1148
rect 35196 690 35252 700
rect 35644 756 35700 7980
rect 35756 7252 35812 12348
rect 35868 8260 35924 13020
rect 36092 10836 36148 14112
rect 36540 13972 36596 14112
rect 36540 13906 36596 13916
rect 36988 13300 37044 14112
rect 36988 13234 37044 13244
rect 36876 12740 36932 12750
rect 36876 12178 36932 12684
rect 37436 12628 37492 14112
rect 37436 12562 37492 12572
rect 36876 12126 36878 12178
rect 36930 12126 36932 12178
rect 36876 12114 36932 12126
rect 37324 12516 37380 12526
rect 36092 10770 36148 10780
rect 36316 12066 36372 12078
rect 36316 12014 36318 12066
rect 36370 12014 36372 12066
rect 36316 10388 36372 12014
rect 36988 10500 37044 10510
rect 36988 10406 37044 10444
rect 36316 10322 36372 10332
rect 36652 9940 36708 9950
rect 36652 9846 36708 9884
rect 36092 9828 36148 9838
rect 36092 9734 36148 9772
rect 36316 9828 36372 9838
rect 36316 9492 36372 9772
rect 36316 9426 36372 9436
rect 35868 8194 35924 8204
rect 36092 8596 36148 8606
rect 35756 7186 35812 7196
rect 36092 1316 36148 8540
rect 36988 8372 37044 8382
rect 36652 7700 36708 7710
rect 36540 4116 36596 4126
rect 36428 4114 36596 4116
rect 36428 4062 36542 4114
rect 36594 4062 36596 4114
rect 36428 4060 36596 4062
rect 36428 3332 36484 4060
rect 36540 4050 36596 4060
rect 36540 3556 36596 3566
rect 36540 3462 36596 3500
rect 36428 3266 36484 3276
rect 36652 3108 36708 7644
rect 36876 7700 36932 7710
rect 36652 3042 36708 3052
rect 36764 4564 36820 4574
rect 36092 1250 36148 1260
rect 35644 690 35700 700
rect 36764 112 36820 4508
rect 36876 1428 36932 7644
rect 36988 5348 37044 8316
rect 37100 8036 37156 8046
rect 37100 7028 37156 7980
rect 37100 6962 37156 6972
rect 37100 6804 37156 6814
rect 37100 5572 37156 6748
rect 37100 5506 37156 5516
rect 36988 5282 37044 5292
rect 36988 4452 37044 4462
rect 36988 4358 37044 4396
rect 37100 4004 37156 4014
rect 37100 3666 37156 3948
rect 37100 3614 37102 3666
rect 37154 3614 37156 3666
rect 37100 3602 37156 3614
rect 37324 3220 37380 12460
rect 37772 12292 37828 12302
rect 37660 11954 37716 11966
rect 37660 11902 37662 11954
rect 37714 11902 37716 11954
rect 37548 10386 37604 10398
rect 37548 10334 37550 10386
rect 37602 10334 37604 10386
rect 37548 9044 37604 10334
rect 37660 10164 37716 11902
rect 37660 10098 37716 10108
rect 37548 8978 37604 8988
rect 37772 8596 37828 12236
rect 37884 11956 37940 14112
rect 38220 13524 38276 13534
rect 38108 12852 38164 12862
rect 38108 12290 38164 12796
rect 38108 12238 38110 12290
rect 38162 12238 38164 12290
rect 38108 12226 38164 12238
rect 37884 11890 37940 11900
rect 38220 11732 38276 13468
rect 38332 13076 38388 14112
rect 38332 13010 38388 13020
rect 38556 14084 38612 14094
rect 38220 11666 38276 11676
rect 38332 12852 38388 12862
rect 37772 8530 37828 8540
rect 37324 3154 37380 3164
rect 37548 6690 37604 6702
rect 37548 6638 37550 6690
rect 37602 6638 37604 6690
rect 36876 1362 36932 1372
rect 36988 2884 37044 2894
rect 36988 980 37044 2828
rect 37548 2548 37604 6638
rect 37996 6578 38052 6590
rect 37996 6526 37998 6578
rect 38050 6526 38052 6578
rect 37996 6468 38052 6526
rect 37996 6402 38052 6412
rect 38220 6468 38276 6478
rect 38220 2996 38276 6412
rect 38332 6132 38388 12796
rect 38556 10836 38612 14028
rect 38780 13748 38836 14112
rect 38780 13682 38836 13692
rect 38556 10770 38612 10780
rect 38556 9156 38612 9166
rect 38556 8596 38612 9100
rect 38780 9156 38836 9166
rect 38780 8596 38836 9100
rect 38556 8540 38836 8596
rect 39228 7700 39284 14112
rect 39340 12964 39396 12974
rect 39340 8036 39396 12908
rect 39452 12180 39508 12190
rect 39452 10164 39508 12124
rect 39452 10098 39508 10108
rect 39564 11060 39620 11070
rect 39340 7970 39396 7980
rect 39228 7634 39284 7644
rect 38556 7476 38612 7486
rect 38556 7252 38612 7420
rect 38556 7186 38612 7196
rect 39228 7252 39284 7262
rect 39228 6802 39284 7196
rect 39228 6750 39230 6802
rect 39282 6750 39284 6802
rect 39228 6738 39284 6750
rect 38332 6066 38388 6076
rect 38668 6690 38724 6702
rect 38668 6638 38670 6690
rect 38722 6638 38724 6690
rect 38668 6020 38724 6638
rect 38444 5964 38724 6020
rect 39564 6020 39620 11004
rect 39676 7140 39732 14112
rect 40124 13524 40180 14112
rect 40124 13458 40180 13468
rect 40236 13860 40292 13870
rect 40124 12964 40180 12974
rect 39788 11732 39844 11742
rect 39788 11060 39844 11676
rect 39788 10994 39844 11004
rect 40012 11732 40068 11742
rect 39900 10836 39956 10846
rect 40012 10836 40068 11676
rect 40124 11396 40180 12908
rect 40236 12292 40292 13804
rect 40236 12236 40404 12292
rect 40124 11330 40180 11340
rect 40236 12068 40292 12078
rect 39956 10780 40068 10836
rect 40124 10836 40180 10846
rect 39900 10770 39956 10780
rect 40012 10276 40068 10286
rect 39676 7074 39732 7084
rect 39788 8372 39844 8382
rect 38444 5460 38500 5964
rect 39564 5954 39620 5964
rect 39788 5908 39844 8316
rect 39788 5842 39844 5852
rect 39900 6692 39956 6702
rect 38444 5394 38500 5404
rect 39340 5348 39396 5358
rect 38668 4452 38724 4462
rect 38668 3892 38724 4396
rect 39340 4338 39396 5292
rect 39900 4450 39956 6636
rect 40012 6580 40068 10220
rect 40124 9268 40180 10780
rect 40236 10724 40292 12012
rect 40348 11396 40404 12236
rect 40572 11508 40628 14112
rect 41020 12964 41076 14112
rect 41020 12898 41076 12908
rect 41468 12292 41524 14112
rect 41468 12226 41524 12236
rect 40572 11442 40628 11452
rect 41356 11956 41412 11966
rect 40348 11330 40404 11340
rect 40236 10658 40292 10668
rect 40460 10724 40516 10734
rect 40124 9202 40180 9212
rect 40236 9156 40292 9166
rect 40124 8036 40180 8046
rect 40124 6580 40180 7980
rect 40236 7812 40292 9100
rect 40460 8484 40516 10668
rect 41356 10610 41412 11900
rect 41356 10558 41358 10610
rect 41410 10558 41412 10610
rect 41356 10546 41412 10558
rect 41692 11956 41748 11966
rect 41692 10276 41748 11900
rect 41804 11732 41860 11742
rect 41804 11508 41860 11676
rect 41804 11442 41860 11452
rect 41692 10210 41748 10220
rect 41804 11284 41860 11294
rect 40460 8418 40516 8428
rect 40572 9940 40628 9950
rect 40236 7746 40292 7756
rect 40348 8258 40404 8270
rect 40348 8206 40350 8258
rect 40402 8206 40404 8258
rect 40348 7028 40404 8206
rect 40348 6962 40404 6972
rect 40460 7700 40516 7710
rect 40236 6580 40292 6590
rect 40124 6524 40236 6580
rect 40012 6514 40068 6524
rect 40236 6514 40292 6524
rect 40460 6356 40516 7644
rect 40460 6290 40516 6300
rect 39900 4398 39902 4450
rect 39954 4398 39956 4450
rect 39900 4386 39956 4398
rect 40124 6132 40180 6142
rect 39340 4286 39342 4338
rect 39394 4286 39396 4338
rect 39340 4274 39396 4286
rect 40124 4228 40180 6076
rect 40124 4162 40180 4172
rect 40236 5684 40292 5694
rect 38668 3826 38724 3836
rect 40236 3892 40292 5628
rect 40348 5012 40404 5022
rect 40348 4564 40404 4956
rect 40348 4498 40404 4508
rect 40236 3826 40292 3836
rect 39788 3780 39844 3790
rect 38892 3668 38948 3678
rect 39788 3668 39844 3724
rect 40572 3668 40628 9884
rect 41468 9826 41524 9838
rect 41468 9774 41470 9826
rect 41522 9774 41524 9826
rect 40684 8146 40740 8158
rect 40684 8094 40686 8146
rect 40738 8094 40740 8146
rect 40684 6244 40740 8094
rect 41468 7924 41524 9774
rect 41468 7858 41524 7868
rect 41692 9044 41748 9054
rect 41580 7476 41636 7486
rect 41580 6914 41636 7420
rect 41580 6862 41582 6914
rect 41634 6862 41636 6914
rect 41580 6850 41636 6862
rect 41692 6244 41748 8988
rect 41804 6580 41860 11228
rect 41916 10948 41972 14112
rect 41916 10882 41972 10892
rect 42252 10612 42308 10622
rect 42252 10518 42308 10556
rect 41916 10500 41972 10510
rect 41916 10498 42196 10500
rect 41916 10446 41918 10498
rect 41970 10446 42196 10498
rect 41916 10444 42196 10446
rect 41916 10434 41972 10444
rect 41916 9714 41972 9726
rect 41916 9662 41918 9714
rect 41970 9662 41972 9714
rect 41916 9044 41972 9662
rect 41916 8978 41972 8988
rect 42140 7476 42196 10444
rect 42364 8148 42420 14112
rect 42812 12740 42868 14112
rect 43260 13300 43316 14112
rect 43260 13234 43316 13244
rect 43596 13972 43652 13982
rect 42812 12674 42868 12684
rect 43036 12740 43092 12750
rect 42476 12628 42532 12638
rect 42476 9268 42532 12572
rect 42812 10612 42868 10622
rect 42812 10518 42868 10556
rect 42476 9202 42532 9212
rect 42588 9826 42644 9838
rect 42588 9774 42590 9826
rect 42642 9774 42644 9826
rect 42588 8932 42644 9774
rect 42588 8866 42644 8876
rect 42364 8082 42420 8092
rect 42140 7410 42196 7420
rect 42028 6580 42084 6590
rect 41804 6578 42084 6580
rect 41804 6526 42030 6578
rect 42082 6526 42084 6578
rect 41804 6524 42084 6526
rect 42028 6514 42084 6524
rect 42364 6580 42420 6590
rect 41692 6188 41972 6244
rect 40684 6178 40740 6188
rect 41804 6020 41860 6030
rect 41132 5908 41188 5918
rect 39788 3612 40628 3668
rect 40684 4676 40740 4686
rect 38220 2930 38276 2940
rect 38668 3444 38724 3454
rect 37884 2772 37940 2782
rect 37884 2678 37940 2716
rect 38668 2772 38724 3388
rect 38668 2706 38724 2716
rect 37548 2482 37604 2492
rect 38444 2658 38500 2670
rect 38444 2606 38446 2658
rect 38498 2606 38500 2658
rect 38444 2212 38500 2606
rect 38892 2660 38948 3612
rect 40684 3388 40740 4620
rect 41132 4340 41188 5852
rect 41244 5124 41300 5134
rect 41244 4564 41300 5068
rect 41244 4508 41748 4564
rect 41132 4274 41188 4284
rect 41692 4338 41748 4508
rect 41692 4286 41694 4338
rect 41746 4286 41748 4338
rect 41692 4274 41748 4286
rect 40460 3332 40740 3388
rect 41468 3332 41524 3342
rect 38892 2594 38948 2604
rect 40236 3220 40292 3230
rect 38444 2146 38500 2156
rect 36988 914 37044 924
rect 39340 1988 39396 1998
rect 39340 532 39396 1932
rect 39452 1764 39508 1774
rect 39452 1540 39508 1708
rect 39452 1474 39508 1484
rect 39340 466 39396 476
rect 39452 1316 39508 1326
rect 39452 112 39508 1260
rect 40236 1092 40292 3164
rect 40236 1026 40292 1036
rect 40460 420 40516 3332
rect 41468 532 41524 3276
rect 41804 3220 41860 5964
rect 41916 3388 41972 6188
rect 42252 4228 42308 4238
rect 42252 4134 42308 4172
rect 42252 3892 42308 3902
rect 41916 3332 42196 3388
rect 41804 3164 42084 3220
rect 41580 1652 41636 1662
rect 41580 980 41636 1596
rect 42028 1204 42084 3164
rect 42028 1138 42084 1148
rect 41580 914 41636 924
rect 41468 466 41524 476
rect 40460 354 40516 364
rect 42140 112 42196 3332
rect 42252 3332 42308 3836
rect 42252 3266 42308 3276
rect 42364 1764 42420 6524
rect 42588 5236 42644 5246
rect 42588 4676 42644 5180
rect 42588 4610 42644 4620
rect 42364 1698 42420 1708
rect 43036 868 43092 12684
rect 43596 11620 43652 13916
rect 43708 12740 43764 14112
rect 43708 12674 43764 12684
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 44156 11956 44212 14112
rect 44604 13524 44660 14112
rect 44604 13468 44884 13524
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 44716 13188 44772 13198
rect 44156 11890 44212 11900
rect 44268 12516 44324 12526
rect 43596 11564 44212 11620
rect 43372 11396 43428 11406
rect 43148 9714 43204 9726
rect 43148 9662 43150 9714
rect 43202 9662 43204 9714
rect 43148 8484 43204 9662
rect 43148 8418 43204 8428
rect 43372 8148 43428 11340
rect 43596 11060 43652 11070
rect 43596 9940 43652 11004
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44156 10948 44212 11564
rect 44268 11172 44324 12460
rect 44716 12178 44772 13132
rect 44716 12126 44718 12178
rect 44770 12126 44772 12178
rect 44716 12114 44772 12126
rect 44828 11956 44884 13468
rect 44940 12962 44996 12974
rect 44940 12910 44942 12962
rect 44994 12910 44996 12962
rect 44940 12180 44996 12910
rect 44940 12114 44996 12124
rect 44828 11900 44996 11956
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44268 11106 44324 11116
rect 44156 10892 44324 10948
rect 43596 9874 43652 9884
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 44268 9380 44324 10892
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44716 9828 44772 9838
rect 44716 9826 44884 9828
rect 44716 9774 44718 9826
rect 44770 9774 44884 9826
rect 44716 9772 44884 9774
rect 44716 9762 44772 9772
rect 44268 9314 44324 9324
rect 43372 8082 43428 8092
rect 44156 9268 44212 9278
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 43596 5572 43652 5582
rect 43596 3780 43652 5516
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 44156 4452 44212 9212
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44464 7084 44728 7094
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 44828 5236 44884 9772
rect 44828 5170 44884 5180
rect 44940 5012 44996 11900
rect 45052 5124 45108 14112
rect 45500 13076 45556 14112
rect 45948 13188 46004 14112
rect 46396 13636 46452 14112
rect 46396 13570 46452 13580
rect 46844 13524 46900 14112
rect 46844 13458 46900 13468
rect 45948 13122 46004 13132
rect 46396 13076 46452 13086
rect 45500 13020 45780 13076
rect 45500 12852 45556 12862
rect 45276 12066 45332 12078
rect 45276 12014 45278 12066
rect 45330 12014 45332 12066
rect 45276 11844 45332 12014
rect 45276 11778 45332 11788
rect 45388 12068 45444 12078
rect 45388 11396 45444 12012
rect 45388 11330 45444 11340
rect 45500 10052 45556 12796
rect 45500 9986 45556 9996
rect 45612 9940 45668 9950
rect 45164 9716 45220 9726
rect 45164 9622 45220 9660
rect 45388 9268 45444 9278
rect 45388 7588 45444 9212
rect 45612 8148 45668 9884
rect 45724 9156 45780 13020
rect 45948 12852 46004 12862
rect 45948 12758 46004 12796
rect 46396 12178 46452 13020
rect 46844 12964 46900 12974
rect 46396 12126 46398 12178
rect 46450 12126 46452 12178
rect 46396 12114 46452 12126
rect 46620 12962 46900 12964
rect 46620 12910 46846 12962
rect 46898 12910 46900 12962
rect 46620 12908 46900 12910
rect 46172 10836 46228 10846
rect 45724 9090 45780 9100
rect 45836 9380 45892 9390
rect 45612 8082 45668 8092
rect 45388 7522 45444 7532
rect 45500 7812 45556 7822
rect 45052 5058 45108 5068
rect 45388 6804 45444 6814
rect 44940 4946 44996 4956
rect 43596 3714 43652 3724
rect 43932 4396 44212 4452
rect 43932 3778 43988 4396
rect 45276 4340 45332 4350
rect 45388 4340 45444 6748
rect 45500 4676 45556 7756
rect 45836 7812 45892 9324
rect 45836 7746 45892 7756
rect 45612 7588 45668 7598
rect 45612 5684 45668 7532
rect 46172 6580 46228 10780
rect 46172 6514 46228 6524
rect 46284 10164 46340 10174
rect 45612 5618 45668 5628
rect 45500 4610 45556 4620
rect 45332 4284 45444 4340
rect 45276 4274 45332 4284
rect 45724 4004 45780 4014
rect 44464 3948 44728 3958
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 43932 3726 43934 3778
rect 43986 3726 43988 3778
rect 43932 3714 43988 3726
rect 44044 3780 44100 3790
rect 44044 3556 44100 3724
rect 44044 3490 44100 3500
rect 44380 3444 44436 3482
rect 44380 3378 44436 3388
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 45724 1988 45780 3948
rect 46284 2772 46340 10108
rect 46620 8148 46676 12908
rect 46844 12898 46900 12908
rect 46956 12068 47012 12078
rect 46732 12066 47012 12068
rect 46732 12014 46958 12066
rect 47010 12014 47012 12066
rect 46732 12012 47012 12014
rect 46732 9828 46788 12012
rect 46956 12002 47012 12012
rect 46956 11620 47012 11630
rect 47180 11620 47236 11630
rect 47012 11618 47236 11620
rect 47012 11566 47182 11618
rect 47234 11566 47236 11618
rect 47012 11564 47236 11566
rect 46956 11554 47012 11564
rect 47180 11554 47236 11564
rect 46732 9762 46788 9772
rect 47180 9156 47236 9166
rect 47068 8818 47124 8830
rect 47068 8766 47070 8818
rect 47122 8766 47124 8818
rect 47068 8596 47124 8766
rect 47068 8530 47124 8540
rect 47180 8260 47236 9100
rect 47180 8194 47236 8204
rect 46620 8092 46900 8148
rect 46284 2706 46340 2716
rect 46508 7476 46564 7486
rect 45724 1922 45780 1932
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 46508 1540 46564 7420
rect 46620 7252 46676 7262
rect 46620 3108 46676 7196
rect 46844 3388 46900 8092
rect 47068 8036 47124 8046
rect 47068 6132 47124 7980
rect 47068 6066 47124 6076
rect 47180 6244 47236 6254
rect 46620 3042 46676 3052
rect 46732 3332 46900 3388
rect 46956 5122 47012 5134
rect 46956 5070 46958 5122
rect 47010 5070 47012 5122
rect 46732 1652 46788 3332
rect 46732 1586 46788 1596
rect 46508 1474 46564 1484
rect 46956 1316 47012 5070
rect 47068 5124 47124 5134
rect 47068 3332 47124 5068
rect 47180 4116 47236 6188
rect 47180 4050 47236 4060
rect 47068 3266 47124 3276
rect 47292 2996 47348 14112
rect 47404 12404 47460 12414
rect 47404 9940 47460 12348
rect 47516 11620 47572 11630
rect 47740 11620 47796 14112
rect 47852 13636 47908 13646
rect 47852 12850 47908 13580
rect 48188 13188 48244 14112
rect 48188 13122 48244 13132
rect 48412 12964 48468 12974
rect 47852 12798 47854 12850
rect 47906 12798 47908 12850
rect 47852 12786 47908 12798
rect 48076 12962 48468 12964
rect 48076 12910 48414 12962
rect 48466 12910 48468 12962
rect 48076 12908 48468 12910
rect 47964 11956 48020 11966
rect 47964 11862 48020 11900
rect 47516 11618 47796 11620
rect 47516 11566 47518 11618
rect 47570 11566 47796 11618
rect 47516 11564 47796 11566
rect 47516 11554 47572 11564
rect 47628 10836 47684 10846
rect 47628 10610 47684 10780
rect 47628 10558 47630 10610
rect 47682 10558 47684 10610
rect 47628 10546 47684 10558
rect 47404 9874 47460 9884
rect 48076 9156 48132 12908
rect 48412 12898 48468 12908
rect 48636 12404 48692 14112
rect 49084 13524 49140 14112
rect 49084 13458 49140 13468
rect 48972 13188 49028 13198
rect 48972 13094 49028 13132
rect 48636 12338 48692 12348
rect 49420 12404 49476 12414
rect 49420 12310 49476 12348
rect 48524 12066 48580 12078
rect 48524 12014 48526 12066
rect 48578 12014 48580 12066
rect 48300 11394 48356 11406
rect 48300 11342 48302 11394
rect 48354 11342 48356 11394
rect 48188 11172 48244 11182
rect 48188 10722 48244 11116
rect 48188 10670 48190 10722
rect 48242 10670 48244 10722
rect 48188 10658 48244 10670
rect 48300 10388 48356 11342
rect 48300 10322 48356 10332
rect 48524 10052 48580 12014
rect 48860 12068 48916 12078
rect 48860 11974 48916 12012
rect 49420 11844 49476 11854
rect 49196 11732 49252 11742
rect 49084 11508 49140 11518
rect 49084 11060 49140 11452
rect 49196 11282 49252 11676
rect 49196 11230 49198 11282
rect 49250 11230 49252 11282
rect 49196 11218 49252 11230
rect 49084 11004 49252 11060
rect 48748 10612 48804 10622
rect 48524 9996 48692 10052
rect 48524 9826 48580 9838
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 47292 2930 47348 2940
rect 47404 9100 48132 9156
rect 48300 9716 48356 9726
rect 47404 1876 47460 9100
rect 47628 8930 47684 8942
rect 47628 8878 47630 8930
rect 47682 8878 47684 8930
rect 47516 8708 47572 8718
rect 47516 5234 47572 8652
rect 47516 5182 47518 5234
rect 47570 5182 47572 5234
rect 47516 5170 47572 5182
rect 47628 2100 47684 8878
rect 48076 8484 48132 8494
rect 48076 3220 48132 8428
rect 48076 3154 48132 3164
rect 47628 2034 47684 2044
rect 47404 1810 47460 1820
rect 47068 1764 47124 1774
rect 47068 1428 47124 1708
rect 47068 1362 47124 1372
rect 46956 1250 47012 1260
rect 44828 980 44884 990
rect 43036 802 43092 812
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 44828 112 44884 924
rect 48300 980 48356 9660
rect 48524 8372 48580 9774
rect 48524 8306 48580 8316
rect 48412 8258 48468 8270
rect 48412 8206 48414 8258
rect 48466 8206 48468 8258
rect 48412 4564 48468 8206
rect 48636 5236 48692 9996
rect 48748 6132 48804 10556
rect 48748 6066 48804 6076
rect 48860 10610 48916 10622
rect 48860 10558 48862 10610
rect 48914 10558 48916 10610
rect 48860 5908 48916 10558
rect 49084 9714 49140 9726
rect 49084 9662 49086 9714
rect 49138 9662 49140 9714
rect 48972 8260 49028 8270
rect 48972 8166 49028 8204
rect 49084 7700 49140 9662
rect 49084 7634 49140 7644
rect 49196 7140 49252 11004
rect 49420 10052 49476 11788
rect 49532 11620 49588 14112
rect 49980 13076 50036 14112
rect 49980 13010 50036 13020
rect 50428 12404 50484 14112
rect 50428 12338 50484 12348
rect 50540 12962 50596 12974
rect 50540 12910 50542 12962
rect 50594 12910 50596 12962
rect 50428 11954 50484 11966
rect 50428 11902 50430 11954
rect 50482 11902 50484 11954
rect 49532 11554 49588 11564
rect 49868 11844 49924 11854
rect 49756 11394 49812 11406
rect 49756 11342 49758 11394
rect 49810 11342 49812 11394
rect 49644 11060 49700 11070
rect 49644 10834 49700 11004
rect 49644 10782 49646 10834
rect 49698 10782 49700 10834
rect 49644 10770 49700 10782
rect 49756 10164 49812 11342
rect 49756 10098 49812 10108
rect 49644 10052 49700 10062
rect 49420 9996 49588 10052
rect 49420 9044 49476 9054
rect 49308 8932 49364 8942
rect 49308 8838 49364 8876
rect 49196 7074 49252 7084
rect 48860 5842 48916 5852
rect 48636 5170 48692 5180
rect 48412 4498 48468 4508
rect 49308 4114 49364 4126
rect 49308 4062 49310 4114
rect 49362 4062 49364 4114
rect 48412 3444 48468 3454
rect 48412 1204 48468 3388
rect 48412 1138 48468 1148
rect 48300 914 48356 924
rect 47516 644 47572 654
rect 47516 112 47572 588
rect 49308 532 49364 4062
rect 49420 2772 49476 8988
rect 49420 2706 49476 2716
rect 49532 1652 49588 9996
rect 49644 9826 49700 9996
rect 49644 9774 49646 9826
rect 49698 9774 49700 9826
rect 49644 9762 49700 9774
rect 49868 9156 49924 11788
rect 50316 11620 50372 11630
rect 50316 11526 50372 11564
rect 50204 10500 50260 10510
rect 50204 10406 50260 10444
rect 50316 10052 50372 10062
rect 50204 9828 50260 9838
rect 50204 9734 50260 9772
rect 49868 9090 49924 9100
rect 49756 9042 49812 9054
rect 49756 8990 49758 9042
rect 49810 8990 49812 9042
rect 49756 4228 49812 8990
rect 50204 8932 50260 8942
rect 49980 8930 50260 8932
rect 49980 8878 50206 8930
rect 50258 8878 50260 8930
rect 49980 8876 50260 8878
rect 49868 4452 49924 4462
rect 49980 4452 50036 8876
rect 50204 8866 50260 8876
rect 50092 8258 50148 8270
rect 50092 8206 50094 8258
rect 50146 8206 50148 8258
rect 50092 8148 50148 8206
rect 50092 8082 50148 8092
rect 50316 7588 50372 9996
rect 50428 10052 50484 11902
rect 50428 9986 50484 9996
rect 50540 8428 50596 12910
rect 50876 11620 50932 14112
rect 51100 13524 51156 13534
rect 51100 13186 51156 13468
rect 51100 13134 51102 13186
rect 51154 13134 51156 13186
rect 51100 13122 51156 13134
rect 51324 12292 51380 14112
rect 51772 13300 51828 14112
rect 51772 13234 51828 13244
rect 52220 13188 52276 14112
rect 52220 13122 52276 13132
rect 52332 12962 52388 12974
rect 52332 12910 52334 12962
rect 52386 12910 52388 12962
rect 51772 12516 51828 12526
rect 51324 12236 51492 12292
rect 50988 12066 51044 12078
rect 50988 12014 50990 12066
rect 51042 12014 51044 12066
rect 50988 11844 51044 12014
rect 50988 11778 51044 11788
rect 51212 11844 51268 11854
rect 50876 11554 50932 11564
rect 51212 10834 51268 11788
rect 51436 11508 51492 12236
rect 51436 11442 51492 11452
rect 51212 10782 51214 10834
rect 51266 10782 51268 10834
rect 51212 10770 51268 10782
rect 51324 11394 51380 11406
rect 51324 11342 51326 11394
rect 51378 11342 51380 11394
rect 51324 10836 51380 11342
rect 51324 10770 51380 10780
rect 51660 11172 51716 11182
rect 50316 7522 50372 7532
rect 50428 8372 50596 8428
rect 51100 9826 51156 9838
rect 51100 9774 51102 9826
rect 51154 9774 51156 9826
rect 49868 4450 50036 4452
rect 49868 4398 49870 4450
rect 49922 4398 50036 4450
rect 49868 4396 50036 4398
rect 49868 4386 49924 4396
rect 49756 4172 50260 4228
rect 49532 1586 49588 1596
rect 49980 3554 50036 3566
rect 49980 3502 49982 3554
rect 50034 3502 50036 3554
rect 49308 466 49364 476
rect 49980 420 50036 3502
rect 49980 354 50036 364
rect 50204 112 50260 4172
rect 50428 3556 50484 8372
rect 50988 8260 51044 8270
rect 50988 8166 51044 8204
rect 50540 8148 50596 8158
rect 50540 8054 50596 8092
rect 50876 7812 50932 7822
rect 50876 7474 50932 7756
rect 50876 7422 50878 7474
rect 50930 7422 50932 7474
rect 50876 7410 50932 7422
rect 50540 3892 50596 3902
rect 50540 3666 50596 3836
rect 50540 3614 50542 3666
rect 50594 3614 50596 3666
rect 50540 3602 50596 3614
rect 50428 3490 50484 3500
rect 51100 1764 51156 9774
rect 51212 9380 51268 9390
rect 51212 9266 51268 9324
rect 51212 9214 51214 9266
rect 51266 9214 51268 9266
rect 51212 9202 51268 9214
rect 51436 7476 51492 7486
rect 51436 7382 51492 7420
rect 51660 6468 51716 11116
rect 51660 6402 51716 6412
rect 51100 1698 51156 1708
rect 51436 5122 51492 5134
rect 51436 5070 51438 5122
rect 51490 5070 51492 5122
rect 50988 1204 51044 1214
rect 50988 1110 51044 1148
rect 51436 644 51492 5070
rect 51660 3554 51716 3566
rect 51660 3502 51662 3554
rect 51714 3502 51716 3554
rect 51660 1316 51716 3502
rect 51772 1986 51828 12460
rect 52220 12178 52276 12190
rect 52220 12126 52222 12178
rect 52274 12126 52276 12178
rect 51884 11620 51940 11630
rect 51884 11526 51940 11564
rect 51884 10612 51940 10622
rect 51884 8146 51940 10556
rect 52108 10610 52164 10622
rect 52108 10558 52110 10610
rect 52162 10558 52164 10610
rect 52108 10164 52164 10558
rect 52108 10098 52164 10108
rect 51996 9716 52052 9726
rect 51996 9622 52052 9660
rect 52220 9492 52276 12126
rect 52220 9426 52276 9436
rect 52332 9268 52388 12910
rect 52668 12964 52724 14112
rect 53116 13412 53172 14112
rect 53116 13346 53172 13356
rect 52892 13076 52948 13086
rect 52892 12982 52948 13020
rect 52668 12908 52836 12964
rect 52556 12404 52612 12414
rect 52556 12310 52612 12348
rect 52780 11620 52836 12908
rect 53564 12292 53620 14112
rect 53788 13076 53844 13086
rect 53564 12236 53732 12292
rect 53564 12066 53620 12078
rect 53564 12014 53566 12066
rect 53618 12014 53620 12066
rect 53452 11620 53508 11630
rect 52780 11618 53508 11620
rect 52780 11566 53454 11618
rect 53506 11566 53508 11618
rect 52780 11564 53508 11566
rect 53452 11554 53508 11564
rect 52556 11508 52612 11518
rect 52556 10834 52612 11452
rect 52556 10782 52558 10834
rect 52610 10782 52612 10834
rect 52556 10770 52612 10782
rect 52892 11394 52948 11406
rect 52892 11342 52894 11394
rect 52946 11342 52948 11394
rect 52892 9940 52948 11342
rect 53564 11396 53620 12014
rect 53564 11330 53620 11340
rect 53564 10500 53620 10510
rect 52892 9874 52948 9884
rect 53452 10498 53620 10500
rect 53452 10446 53566 10498
rect 53618 10446 53620 10498
rect 53452 10444 53620 10446
rect 52556 9828 52612 9838
rect 52332 9202 52388 9212
rect 52444 9826 52612 9828
rect 52444 9774 52558 9826
rect 52610 9774 52612 9826
rect 52444 9772 52612 9774
rect 52108 9042 52164 9054
rect 52108 8990 52110 9042
rect 52162 8990 52164 9042
rect 52108 8708 52164 8990
rect 52108 8642 52164 8652
rect 51884 8094 51886 8146
rect 51938 8094 51940 8146
rect 51884 8082 51940 8094
rect 52108 7474 52164 7486
rect 52108 7422 52110 7474
rect 52162 7422 52164 7474
rect 52108 6804 52164 7422
rect 52108 6738 52164 6748
rect 52220 7140 52276 7150
rect 52108 5906 52164 5918
rect 52108 5854 52110 5906
rect 52162 5854 52164 5906
rect 52108 5348 52164 5854
rect 52108 5282 52164 5292
rect 51996 5236 52052 5246
rect 51996 5142 52052 5180
rect 52220 4338 52276 7084
rect 52444 6244 52500 9772
rect 52556 9762 52612 9772
rect 53004 9268 53060 9278
rect 53004 9174 53060 9212
rect 52668 8932 52724 8942
rect 52556 8258 52612 8270
rect 52556 8206 52558 8258
rect 52610 8206 52612 8258
rect 52556 7028 52612 8206
rect 52556 6962 52612 6972
rect 52668 6690 52724 8876
rect 53452 8820 53508 10444
rect 53564 10434 53620 10444
rect 53564 9716 53620 9726
rect 53676 9716 53732 12236
rect 53564 9714 53732 9716
rect 53564 9662 53566 9714
rect 53618 9662 53732 9714
rect 53564 9660 53732 9662
rect 53564 9650 53620 9660
rect 53788 9604 53844 13020
rect 53676 9548 53844 9604
rect 53900 10500 53956 10510
rect 53452 8754 53508 8764
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 8428 53620 8878
rect 53340 8372 53396 8382
rect 53340 8278 53396 8316
rect 53452 8372 53620 8428
rect 53004 7924 53060 7934
rect 53004 7698 53060 7868
rect 53004 7646 53006 7698
rect 53058 7646 53060 7698
rect 53004 7634 53060 7646
rect 53452 7476 53508 8372
rect 52668 6638 52670 6690
rect 52722 6638 52724 6690
rect 52668 6626 52724 6638
rect 53340 7420 53508 7476
rect 52444 6178 52500 6188
rect 52556 6132 52612 6142
rect 52332 5122 52388 5134
rect 52332 5070 52334 5122
rect 52386 5070 52388 5122
rect 52332 4452 52388 5070
rect 52332 4386 52388 4396
rect 52220 4286 52222 4338
rect 52274 4286 52276 4338
rect 52220 4274 52276 4286
rect 52332 4116 52388 4126
rect 52220 3780 52276 3790
rect 52220 3666 52276 3724
rect 52220 3614 52222 3666
rect 52274 3614 52276 3666
rect 52220 3602 52276 3614
rect 52108 2772 52164 2782
rect 52108 2678 52164 2716
rect 51772 1934 51774 1986
rect 51826 1934 51828 1986
rect 51772 1922 51828 1934
rect 52108 1876 52164 1886
rect 52108 1782 52164 1820
rect 51660 1250 51716 1260
rect 51996 1314 52052 1326
rect 51996 1262 51998 1314
rect 52050 1262 52052 1314
rect 51996 980 52052 1262
rect 51996 914 52052 924
rect 52332 756 52388 4060
rect 52556 3666 52612 6076
rect 53004 6132 53060 6142
rect 53004 6038 53060 6076
rect 52892 5236 52948 5246
rect 52892 5142 52948 5180
rect 53228 5122 53284 5134
rect 53228 5070 53230 5122
rect 53282 5070 53284 5122
rect 52668 4564 52724 4574
rect 52668 4450 52724 4508
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 52556 3614 52558 3666
rect 52610 3614 52612 3666
rect 52556 3602 52612 3614
rect 53228 3444 53284 5070
rect 53340 5124 53396 7420
rect 53564 7364 53620 7374
rect 53340 5058 53396 5068
rect 53452 7362 53620 7364
rect 53452 7310 53566 7362
rect 53618 7310 53620 7362
rect 53452 7308 53620 7310
rect 53452 3892 53508 7308
rect 53564 7298 53620 7308
rect 53564 6580 53620 6590
rect 53676 6580 53732 9548
rect 53564 6578 53732 6580
rect 53564 6526 53566 6578
rect 53618 6526 53732 6578
rect 53564 6524 53732 6526
rect 53564 6514 53620 6524
rect 53900 6132 53956 10444
rect 54012 9268 54068 14112
rect 54124 13300 54180 13310
rect 54124 12402 54180 13244
rect 54348 12962 54404 12974
rect 54348 12910 54350 12962
rect 54402 12910 54404 12962
rect 54124 12350 54126 12402
rect 54178 12350 54180 12402
rect 54124 12338 54180 12350
rect 54236 12628 54292 12638
rect 54236 10612 54292 12572
rect 54348 11284 54404 12910
rect 54460 11844 54516 14112
rect 54908 13636 54964 14112
rect 54908 13570 54964 13580
rect 54460 11778 54516 11788
rect 54684 13524 54740 13534
rect 54348 11218 54404 11228
rect 54460 11394 54516 11406
rect 54460 11342 54462 11394
rect 54514 11342 54516 11394
rect 54236 10546 54292 10556
rect 54012 9202 54068 9212
rect 54236 9826 54292 9838
rect 54236 9774 54238 9826
rect 54290 9774 54292 9826
rect 54124 8258 54180 8270
rect 54124 8206 54126 8258
rect 54178 8206 54180 8258
rect 54124 7364 54180 8206
rect 54124 7298 54180 7308
rect 54124 6692 54180 6702
rect 54124 6598 54180 6636
rect 53900 6066 53956 6076
rect 54124 6468 54180 6478
rect 53564 5796 53620 5806
rect 53564 5702 53620 5740
rect 54124 5234 54180 6412
rect 54124 5182 54126 5234
rect 54178 5182 54180 5234
rect 54124 5170 54180 5182
rect 53676 5010 53732 5022
rect 53676 4958 53678 5010
rect 53730 4958 53732 5010
rect 53564 4228 53620 4238
rect 53564 4134 53620 4172
rect 53676 4004 53732 4958
rect 53676 3938 53732 3948
rect 53452 3826 53508 3836
rect 53228 3378 53284 3388
rect 53564 3444 53620 3454
rect 53564 3350 53620 3388
rect 53564 3220 53620 3230
rect 53564 2770 53620 3164
rect 53564 2718 53566 2770
rect 53618 2718 53620 2770
rect 53564 2706 53620 2718
rect 52780 2660 52836 2670
rect 52780 2566 52836 2604
rect 54124 2436 54180 2446
rect 52556 2100 52612 2110
rect 52556 2006 52612 2044
rect 54124 2098 54180 2380
rect 54236 2324 54292 9774
rect 54348 8930 54404 8942
rect 54348 8878 54350 8930
rect 54402 8878 54404 8930
rect 54348 8596 54404 8878
rect 54348 8530 54404 8540
rect 54460 4900 54516 11342
rect 54572 10722 54628 10734
rect 54572 10670 54574 10722
rect 54626 10670 54628 10722
rect 54572 10164 54628 10670
rect 54572 10098 54628 10108
rect 54684 9828 54740 13468
rect 54908 13188 54964 13198
rect 54908 13094 54964 13132
rect 55132 12068 55188 12078
rect 54684 9762 54740 9772
rect 54796 12066 55188 12068
rect 54796 12014 55134 12066
rect 55186 12014 55188 12066
rect 54796 12012 55188 12014
rect 54572 7586 54628 7598
rect 54572 7534 54574 7586
rect 54626 7534 54628 7586
rect 54572 7252 54628 7534
rect 54572 7186 54628 7196
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 5908 54628 5966
rect 54572 5842 54628 5852
rect 54460 4834 54516 4844
rect 54572 4564 54628 4574
rect 54572 4470 54628 4508
rect 54796 4116 54852 12012
rect 55132 12002 55188 12012
rect 55356 11956 55412 14112
rect 55692 13412 55748 13422
rect 55692 12402 55748 13356
rect 55804 13076 55860 14112
rect 55804 13010 55860 13020
rect 56252 12852 56308 14112
rect 56252 12786 56308 12796
rect 56364 13972 56420 13982
rect 55692 12350 55694 12402
rect 55746 12350 55748 12402
rect 55692 12338 55748 12350
rect 55356 11890 55412 11900
rect 55020 11282 55076 11294
rect 55020 11230 55022 11282
rect 55074 11230 55076 11282
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 54796 4050 54852 4060
rect 54796 3778 54852 3790
rect 54796 3726 54798 3778
rect 54850 3726 54852 3778
rect 54796 3668 54852 3726
rect 54796 3602 54852 3612
rect 55020 3556 55076 11230
rect 55692 11284 55748 11294
rect 55356 10610 55412 10622
rect 55356 10558 55358 10610
rect 55410 10558 55412 10610
rect 55132 9602 55188 9614
rect 55132 9550 55134 9602
rect 55186 9550 55188 9602
rect 55132 9492 55188 9550
rect 55132 9426 55188 9436
rect 55244 9604 55300 9614
rect 55244 9042 55300 9548
rect 55244 8990 55246 9042
rect 55298 8990 55300 9042
rect 55244 8978 55300 8990
rect 55132 8148 55188 8158
rect 55132 8054 55188 8092
rect 55132 7362 55188 7374
rect 55132 7310 55134 7362
rect 55186 7310 55188 7362
rect 55132 6916 55188 7310
rect 55132 6850 55188 6860
rect 55132 6466 55188 6478
rect 55132 6414 55134 6466
rect 55186 6414 55188 6466
rect 55132 6356 55188 6414
rect 55132 6290 55188 6300
rect 55132 5796 55188 5806
rect 55132 5702 55188 5740
rect 55356 5236 55412 10558
rect 55468 10388 55524 10398
rect 55468 8148 55524 10332
rect 55692 8372 55748 11228
rect 56140 10722 56196 10734
rect 56140 10670 56142 10722
rect 56194 10670 56196 10722
rect 56140 9044 56196 10670
rect 56364 9380 56420 13916
rect 56700 12964 56756 14112
rect 56588 12908 56756 12964
rect 56924 13076 56980 13086
rect 56588 10500 56644 12908
rect 56924 11060 56980 13020
rect 56924 10994 56980 11004
rect 57260 12180 57316 12190
rect 56588 10434 56644 10444
rect 56700 10836 56756 10846
rect 56700 9716 56756 10780
rect 56700 9650 56756 9660
rect 56364 9314 56420 9324
rect 56140 8978 56196 8988
rect 55692 8306 55748 8316
rect 55916 8930 55972 8942
rect 55916 8878 55918 8930
rect 55970 8878 55972 8930
rect 55468 8082 55524 8092
rect 55916 8148 55972 8878
rect 55916 8082 55972 8092
rect 57260 7924 57316 12124
rect 57260 7858 57316 7868
rect 56140 7700 56196 7710
rect 56140 7606 56196 7644
rect 56140 6804 56196 6814
rect 56140 6130 56196 6748
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 55356 5170 55412 5180
rect 56140 5460 56196 5470
rect 56140 4562 56196 5404
rect 56140 4510 56142 4562
rect 56194 4510 56196 4562
rect 56140 4498 56196 4510
rect 55132 4226 55188 4238
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 3780 55188 4174
rect 55132 3714 55188 3724
rect 56140 4116 56196 4126
rect 55132 3556 55188 3566
rect 55020 3554 55188 3556
rect 55020 3502 55134 3554
rect 55186 3502 55188 3554
rect 55020 3500 55188 3502
rect 55132 3490 55188 3500
rect 54572 3220 54628 3230
rect 54572 2994 54628 3164
rect 54572 2942 54574 2994
rect 54626 2942 54628 2994
rect 54572 2930 54628 2942
rect 55132 3108 55188 3118
rect 55132 2770 55188 3052
rect 56140 2994 56196 4060
rect 56140 2942 56142 2994
rect 56194 2942 56196 2994
rect 56140 2930 56196 2942
rect 56812 3444 56868 3454
rect 55132 2718 55134 2770
rect 55186 2718 55188 2770
rect 55132 2706 55188 2718
rect 56140 2772 56196 2782
rect 54236 2258 54292 2268
rect 54908 2324 54964 2334
rect 54124 2046 54126 2098
rect 54178 2046 54180 2098
rect 54124 2034 54180 2046
rect 54908 2098 54964 2268
rect 54908 2046 54910 2098
rect 54962 2046 54964 2098
rect 54908 2034 54964 2046
rect 53564 1876 53620 1886
rect 53564 1782 53620 1820
rect 55132 1652 55188 1662
rect 52556 1540 52612 1550
rect 52556 1202 52612 1484
rect 53564 1428 53620 1438
rect 53564 1334 53620 1372
rect 52556 1150 52558 1202
rect 52610 1150 52612 1202
rect 52556 1138 52612 1150
rect 55132 1202 55188 1596
rect 56140 1426 56196 2716
rect 56140 1374 56142 1426
rect 56194 1374 56196 1426
rect 56140 1362 56196 1374
rect 56476 2660 56532 2670
rect 55132 1150 55134 1202
rect 55186 1150 55188 1202
rect 55132 1138 55188 1150
rect 52332 690 52388 700
rect 51436 578 51492 588
rect 55580 308 55636 318
rect 52892 196 52948 206
rect 52892 112 52948 140
rect 55580 112 55636 252
rect 25340 28 25732 84
rect 25984 0 26096 112
rect 28672 0 28784 112
rect 31360 0 31472 112
rect 34048 0 34160 112
rect 36736 0 36848 112
rect 39424 0 39536 112
rect 42112 0 42224 112
rect 44800 0 44912 112
rect 47488 0 47600 112
rect 50176 0 50288 112
rect 52864 0 52976 112
rect 55552 0 55664 112
rect 56476 84 56532 2604
rect 56812 532 56868 3388
rect 56812 466 56868 476
rect 56476 18 56532 28
<< via2 >>
rect 364 13020 420 13076
rect 140 10556 196 10612
rect 476 12572 532 12628
rect 476 11340 532 11396
rect 588 12124 644 12180
rect 364 9996 420 10052
rect 140 9884 196 9940
rect 1036 13468 1092 13524
rect 2156 13244 2212 13300
rect 2268 12402 2324 12404
rect 2268 12350 2270 12402
rect 2270 12350 2322 12402
rect 2322 12350 2324 12402
rect 2268 12348 2324 12350
rect 1036 11452 1092 11508
rect 588 9660 644 9716
rect 924 11004 980 11060
rect 1260 9826 1316 9828
rect 1260 9774 1262 9826
rect 1262 9774 1314 9826
rect 1314 9774 1316 9826
rect 1260 9772 1316 9774
rect 1148 9436 1204 9492
rect 812 6412 868 6468
rect 1036 6972 1092 7028
rect 1148 6636 1204 6692
rect 1260 8540 1316 8596
rect 1596 11282 1652 11284
rect 1596 11230 1598 11282
rect 1598 11230 1650 11282
rect 1650 11230 1652 11282
rect 1596 11228 1652 11230
rect 1596 10780 1652 10836
rect 1372 7644 1428 7700
rect 1372 6300 1428 6356
rect 1372 5740 1428 5796
rect 1820 9772 1876 9828
rect 1596 8316 1652 8372
rect 1708 7420 1764 7476
rect 1596 7196 1652 7252
rect 1596 6076 1652 6132
rect 1596 5404 1652 5460
rect 1484 5068 1540 5124
rect 1372 4508 1428 4564
rect 1260 4284 1316 4340
rect 1596 3724 1652 3780
rect 1596 3164 1652 3220
rect 1036 1820 1092 1876
rect 1148 1932 1204 1988
rect 924 1708 980 1764
rect 924 924 980 980
rect 2268 11788 2324 11844
rect 2492 9996 2548 10052
rect 2604 8930 2660 8932
rect 2604 8878 2606 8930
rect 2606 8878 2658 8930
rect 2658 8878 2660 8930
rect 2604 8876 2660 8878
rect 2492 8652 2548 8708
rect 2268 8258 2324 8260
rect 2268 8206 2270 8258
rect 2270 8206 2322 8258
rect 2322 8206 2324 8258
rect 2268 8204 2324 8206
rect 2380 7196 2436 7252
rect 1932 4172 1988 4228
rect 2044 588 2100 644
rect 2604 5234 2660 5236
rect 2604 5182 2606 5234
rect 2606 5182 2658 5234
rect 2658 5182 2660 5234
rect 2604 5180 2660 5182
rect 2492 2210 2548 2212
rect 2492 2158 2494 2210
rect 2494 2158 2546 2210
rect 2546 2158 2548 2210
rect 2492 2156 2548 2158
rect 3388 12348 3444 12404
rect 3612 13468 3668 13524
rect 3724 13186 3780 13188
rect 3724 13134 3726 13186
rect 3726 13134 3778 13186
rect 3778 13134 3780 13186
rect 3724 13132 3780 13134
rect 4732 13468 4788 13524
rect 4284 13244 4340 13300
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 2940 11900 2996 11956
rect 3388 11900 3444 11956
rect 3276 10780 3332 10836
rect 3164 10668 3220 10724
rect 2828 10498 2884 10500
rect 2828 10446 2830 10498
rect 2830 10446 2882 10498
rect 2882 10446 2884 10498
rect 2828 10444 2884 10446
rect 2828 10220 2884 10276
rect 2940 9548 2996 9604
rect 3052 9212 3108 9268
rect 2716 3500 2772 3556
rect 2828 8652 2884 8708
rect 2940 7084 2996 7140
rect 3052 7532 3108 7588
rect 4172 11676 4228 11732
rect 3500 9548 3556 9604
rect 3276 8092 3332 8148
rect 3164 6972 3220 7028
rect 3500 7308 3556 7364
rect 3276 6860 3332 6916
rect 3276 5852 3332 5908
rect 3052 4844 3108 4900
rect 3276 5628 3332 5684
rect 3276 4060 3332 4116
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4396 12066 4452 12068
rect 4396 12014 4398 12066
rect 4398 12014 4450 12066
rect 4450 12014 4452 12066
rect 4396 12012 4452 12014
rect 5068 12012 5124 12068
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4620 11618 4676 11620
rect 4620 11566 4622 11618
rect 4622 11566 4674 11618
rect 4674 11566 4676 11618
rect 4620 11564 4676 11566
rect 4956 11340 5012 11396
rect 4396 11004 4452 11060
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4956 9436 5012 9492
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 4172 8204 4228 8260
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 5404 13580 5460 13636
rect 5180 11564 5236 11620
rect 5292 13020 5348 13076
rect 5180 10892 5236 10948
rect 5628 13132 5684 13188
rect 5964 13244 6020 13300
rect 5964 12460 6020 12516
rect 5292 9996 5348 10052
rect 5180 8988 5236 9044
rect 4284 7084 4340 7140
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3724 5852 3780 5908
rect 3724 5628 3780 5684
rect 3948 5628 4004 5684
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4172 4732 4228 4788
rect 4012 4676 4068 4678
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4508 5234 4564 5236
rect 4508 5182 4510 5234
rect 4510 5182 4562 5234
rect 4562 5182 4564 5234
rect 4508 5180 4564 5182
rect 4284 4620 4340 4676
rect 5068 5068 5124 5124
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 3500 3276 3556 3332
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 2940 1874 2996 1876
rect 2940 1822 2942 1874
rect 2942 1822 2994 1874
rect 2994 1822 2996 1874
rect 2940 1820 2996 1822
rect 2828 1708 2884 1764
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 3276 1372 3332 1428
rect 5180 4338 5236 4340
rect 5180 4286 5182 4338
rect 5182 4286 5234 4338
rect 5234 4286 5236 4338
rect 5180 4284 5236 4286
rect 5292 3052 5348 3108
rect 5404 4844 5460 4900
rect 5068 2492 5124 2548
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 5404 2044 5460 2100
rect 4284 1708 4340 1764
rect 6748 14028 6804 14084
rect 6412 12908 6468 12964
rect 5964 10556 6020 10612
rect 6188 10108 6244 10164
rect 6188 9660 6244 9716
rect 6748 12796 6804 12852
rect 6412 9660 6468 9716
rect 6300 8316 6356 8372
rect 5740 4450 5796 4452
rect 5740 4398 5742 4450
rect 5742 4398 5794 4450
rect 5794 4398 5796 4450
rect 5740 4396 5796 4398
rect 5516 1260 5572 1316
rect 4172 1036 4228 1092
rect 2604 924 2660 980
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 2380 476 2436 532
rect 4508 364 4564 420
rect 6300 8146 6356 8148
rect 6300 8094 6302 8146
rect 6302 8094 6354 8146
rect 6354 8094 6356 8146
rect 6300 8092 6356 8094
rect 6300 7756 6356 7812
rect 6636 7980 6692 8036
rect 6524 5516 6580 5572
rect 7420 13244 7476 13300
rect 7532 13186 7588 13188
rect 7532 13134 7534 13186
rect 7534 13134 7586 13186
rect 7586 13134 7588 13186
rect 7532 13132 7588 13134
rect 6972 12402 7028 12404
rect 6972 12350 6974 12402
rect 6974 12350 7026 12402
rect 7026 12350 7028 12402
rect 6972 12348 7028 12350
rect 7868 12348 7924 12404
rect 6860 8988 6916 9044
rect 7084 8316 7140 8372
rect 6860 7644 6916 7700
rect 6748 4620 6804 4676
rect 6412 3388 6468 3444
rect 6300 1932 6356 1988
rect 6972 6636 7028 6692
rect 6972 4060 7028 4116
rect 7308 6636 7364 6692
rect 7756 10332 7812 10388
rect 7532 6524 7588 6580
rect 7644 8204 7700 8260
rect 8540 12402 8596 12404
rect 8540 12350 8542 12402
rect 8542 12350 8594 12402
rect 8594 12350 8596 12402
rect 8540 12348 8596 12350
rect 8428 12236 8484 12292
rect 8316 11676 8372 11732
rect 8316 10668 8372 10724
rect 8092 10220 8148 10276
rect 7756 7308 7812 7364
rect 8092 9436 8148 9492
rect 8092 3948 8148 4004
rect 8428 10332 8484 10388
rect 8652 11452 8708 11508
rect 9212 13132 9268 13188
rect 9436 12908 9492 12964
rect 8652 10332 8708 10388
rect 9100 10668 9156 10724
rect 8316 9772 8372 9828
rect 8540 9772 8596 9828
rect 8316 8092 8372 8148
rect 8876 8092 8932 8148
rect 8876 7868 8932 7924
rect 9772 13186 9828 13188
rect 9772 13134 9774 13186
rect 9774 13134 9826 13186
rect 9826 13134 9828 13186
rect 9772 13132 9828 13134
rect 9660 12348 9716 12404
rect 10332 12572 10388 12628
rect 9884 12124 9940 12180
rect 9548 11788 9604 11844
rect 9884 11004 9940 11060
rect 10444 11116 10500 11172
rect 9548 10444 9604 10500
rect 9660 10892 9716 10948
rect 9212 7868 9268 7924
rect 8428 6860 8484 6916
rect 8428 6188 8484 6244
rect 8428 5740 8484 5796
rect 8428 4844 8484 4900
rect 8316 4620 8372 4676
rect 7084 2380 7140 2436
rect 9436 6412 9492 6468
rect 8540 3388 8596 3444
rect 8764 5964 8820 6020
rect 8876 5404 8932 5460
rect 9772 10444 9828 10500
rect 10444 10108 10500 10164
rect 9772 9548 9828 9604
rect 9884 9436 9940 9492
rect 9772 6972 9828 7028
rect 9996 8764 10052 8820
rect 9884 6636 9940 6692
rect 9996 8540 10052 8596
rect 9772 5180 9828 5236
rect 10108 7474 10164 7476
rect 10108 7422 10110 7474
rect 10110 7422 10162 7474
rect 10162 7422 10164 7474
rect 10108 7420 10164 7422
rect 10108 6860 10164 6916
rect 10332 8930 10388 8932
rect 10332 8878 10334 8930
rect 10334 8878 10386 8930
rect 10386 8878 10388 8930
rect 10332 8876 10388 8878
rect 10444 8540 10500 8596
rect 10556 8428 10612 8484
rect 10332 8204 10388 8260
rect 11340 13356 11396 13412
rect 11452 13132 11508 13188
rect 12012 13804 12068 13860
rect 11116 12572 11172 12628
rect 11788 13132 11844 13188
rect 11116 11004 11172 11060
rect 11228 12236 11284 12292
rect 11900 12012 11956 12068
rect 11788 11676 11844 11732
rect 12012 11564 12068 11620
rect 12124 13692 12180 13748
rect 11452 11394 11508 11396
rect 11452 11342 11454 11394
rect 11454 11342 11506 11394
rect 11506 11342 11508 11394
rect 11452 11340 11508 11342
rect 11228 9884 11284 9940
rect 11452 10780 11508 10836
rect 10892 9826 10948 9828
rect 10892 9774 10894 9826
rect 10894 9774 10946 9826
rect 10946 9774 10948 9826
rect 10892 9772 10948 9774
rect 10332 7420 10388 7476
rect 10332 7196 10388 7252
rect 10332 6636 10388 6692
rect 10444 6748 10500 6804
rect 10444 6300 10500 6356
rect 10220 5740 10276 5796
rect 10332 5964 10388 6020
rect 10108 5628 10164 5684
rect 10332 5628 10388 5684
rect 11116 5852 11172 5908
rect 9996 5180 10052 5236
rect 9660 3612 9716 3668
rect 9996 4508 10052 4564
rect 6748 1484 6804 1540
rect 7196 1596 7252 1652
rect 5852 364 5908 420
rect 8764 3276 8820 3332
rect 8092 1596 8148 1652
rect 8316 2828 8372 2884
rect 8540 2716 8596 2772
rect 9436 1820 9492 1876
rect 9884 3500 9940 3556
rect 8540 1372 8596 1428
rect 8316 1260 8372 1316
rect 7420 1148 7476 1204
rect 11004 3666 11060 3668
rect 11004 3614 11006 3666
rect 11006 3614 11058 3666
rect 11058 3614 11060 3666
rect 11004 3612 11060 3614
rect 10444 3554 10500 3556
rect 10444 3502 10446 3554
rect 10446 3502 10498 3554
rect 10498 3502 10500 3554
rect 10444 3500 10500 3502
rect 9996 3164 10052 3220
rect 10108 3276 10164 3332
rect 10108 2604 10164 2660
rect 11116 2268 11172 2324
rect 12124 10780 12180 10836
rect 11788 10668 11844 10724
rect 13244 13356 13300 13412
rect 13580 13356 13636 13412
rect 13468 13244 13524 13300
rect 12908 12962 12964 12964
rect 12908 12910 12910 12962
rect 12910 12910 12962 12962
rect 12962 12910 12964 12962
rect 12908 12908 12964 12910
rect 12796 11788 12852 11844
rect 12236 10220 12292 10276
rect 12684 11004 12740 11060
rect 11564 9324 11620 9380
rect 11452 8092 11508 8148
rect 11788 9548 11844 9604
rect 11676 8764 11732 8820
rect 11676 8204 11732 8260
rect 11564 7756 11620 7812
rect 13356 11954 13412 11956
rect 13356 11902 13358 11954
rect 13358 11902 13410 11954
rect 13410 11902 13412 11954
rect 13356 11900 13412 11902
rect 13020 11004 13076 11060
rect 12684 8988 12740 9044
rect 13356 9436 13412 9492
rect 12124 8876 12180 8932
rect 11788 7644 11844 7700
rect 12012 7644 12068 7700
rect 11900 7196 11956 7252
rect 11340 5964 11396 6020
rect 11452 6188 11508 6244
rect 11788 6076 11844 6132
rect 11900 5404 11956 5460
rect 12012 4172 12068 4228
rect 11788 3388 11844 3444
rect 11452 2828 11508 2884
rect 13356 8764 13412 8820
rect 13580 11676 13636 11732
rect 13916 12850 13972 12852
rect 13916 12798 13918 12850
rect 13918 12798 13970 12850
rect 13970 12798 13972 12850
rect 13916 12796 13972 12798
rect 13468 8316 13524 8372
rect 14364 14028 14420 14084
rect 14924 13074 14980 13076
rect 14924 13022 14926 13074
rect 14926 13022 14978 13074
rect 14978 13022 14980 13074
rect 14924 13020 14980 13022
rect 14588 12796 14644 12852
rect 14588 12124 14644 12180
rect 15036 12124 15092 12180
rect 14140 10780 14196 10836
rect 14140 7532 14196 7588
rect 14252 7420 14308 7476
rect 13804 6748 13860 6804
rect 13132 5404 13188 5460
rect 12572 5234 12628 5236
rect 12572 5182 12574 5234
rect 12574 5182 12626 5234
rect 12626 5182 12628 5234
rect 12572 5180 12628 5182
rect 12124 2716 12180 2772
rect 12684 5068 12740 5124
rect 11228 1932 11284 1988
rect 11788 2156 11844 2212
rect 13468 5068 13524 5124
rect 13468 4844 13524 4900
rect 13244 4620 13300 4676
rect 13692 4620 13748 4676
rect 15148 11004 15204 11060
rect 14588 10834 14644 10836
rect 14588 10782 14590 10834
rect 14590 10782 14642 10834
rect 14642 10782 14644 10834
rect 14588 10780 14644 10782
rect 15260 10220 15316 10276
rect 15820 12572 15876 12628
rect 15596 10668 15652 10724
rect 15372 9884 15428 9940
rect 15484 9548 15540 9604
rect 14700 9436 14756 9492
rect 14924 8428 14980 8484
rect 14700 7084 14756 7140
rect 14812 8316 14868 8372
rect 15596 8428 15652 8484
rect 15484 8204 15540 8260
rect 16380 13020 16436 13076
rect 15932 12236 15988 12292
rect 16044 12572 16100 12628
rect 15820 11452 15876 11508
rect 17612 13692 17668 13748
rect 17500 13074 17556 13076
rect 17500 13022 17502 13074
rect 17502 13022 17554 13074
rect 17554 13022 17556 13074
rect 17500 13020 17556 13022
rect 16940 12460 16996 12516
rect 16156 12124 16212 12180
rect 16492 12124 16548 12180
rect 16268 12012 16324 12068
rect 16044 8988 16100 9044
rect 15708 6860 15764 6916
rect 15820 6972 15876 7028
rect 15148 6076 15204 6132
rect 15036 5964 15092 6020
rect 14140 5740 14196 5796
rect 13804 4284 13860 4340
rect 13244 3164 13300 3220
rect 13916 3052 13972 3108
rect 14476 4396 14532 4452
rect 12684 1708 12740 1764
rect 13132 2380 13188 2436
rect 15092 4956 15148 5012
rect 13692 2098 13748 2100
rect 13692 2046 13694 2098
rect 13694 2046 13746 2098
rect 13746 2046 13748 2098
rect 13692 2044 13748 2046
rect 13132 1484 13188 1540
rect 11788 1148 11844 1204
rect 12572 924 12628 980
rect 15484 5628 15540 5684
rect 15484 5180 15540 5236
rect 15708 5180 15764 5236
rect 15596 4172 15652 4228
rect 14700 2156 14756 2212
rect 15036 1820 15092 1876
rect 14364 924 14420 980
rect 14588 1708 14644 1764
rect 14700 1596 14756 1652
rect 15148 1148 15204 1204
rect 14588 812 14644 868
rect 16268 6748 16324 6804
rect 16380 11116 16436 11172
rect 16492 10108 16548 10164
rect 16380 6076 16436 6132
rect 16492 9772 16548 9828
rect 16940 12236 16996 12292
rect 16716 11788 16772 11844
rect 16716 11228 16772 11284
rect 17276 12066 17332 12068
rect 17276 12014 17278 12066
rect 17278 12014 17330 12066
rect 17330 12014 17332 12066
rect 17276 12012 17332 12014
rect 17164 10780 17220 10836
rect 16828 10556 16884 10612
rect 17052 10556 17108 10612
rect 16828 10220 16884 10276
rect 17052 10220 17108 10276
rect 16940 10108 16996 10164
rect 16828 9938 16884 9940
rect 16828 9886 16830 9938
rect 16830 9886 16882 9938
rect 16882 9886 16884 9938
rect 16828 9884 16884 9886
rect 16716 9772 16772 9828
rect 16156 5628 16212 5684
rect 15932 5292 15988 5348
rect 15932 4732 15988 4788
rect 16604 8652 16660 8708
rect 16828 7420 16884 7476
rect 16828 7196 16884 7252
rect 16604 6076 16660 6132
rect 16492 3612 16548 3668
rect 15484 2268 15540 2324
rect 17724 12348 17780 12404
rect 17836 13132 17892 13188
rect 17836 12012 17892 12068
rect 18060 13132 18116 13188
rect 17948 7980 18004 8036
rect 18396 13916 18452 13972
rect 18284 12962 18340 12964
rect 18284 12910 18286 12962
rect 18286 12910 18338 12962
rect 18338 12910 18340 12962
rect 18284 12908 18340 12910
rect 18620 13020 18676 13076
rect 18844 13580 18900 13636
rect 18620 12684 18676 12740
rect 18396 11564 18452 11620
rect 18508 12348 18564 12404
rect 19292 12850 19348 12852
rect 19292 12798 19294 12850
rect 19294 12798 19346 12850
rect 19346 12798 19348 12850
rect 19292 12796 19348 12798
rect 19628 13580 19684 13636
rect 19404 12124 19460 12180
rect 18620 10780 18676 10836
rect 18060 7420 18116 7476
rect 18284 10556 18340 10612
rect 17164 7196 17220 7252
rect 17052 6524 17108 6580
rect 17836 7084 17892 7140
rect 17836 6524 17892 6580
rect 18060 7084 18116 7140
rect 16716 2044 16772 2100
rect 16940 5964 16996 6020
rect 15708 1484 15764 1540
rect 15484 812 15540 868
rect 17948 3612 18004 3668
rect 17388 1484 17444 1540
rect 16940 588 16996 644
rect 17836 252 17892 308
rect 18396 9660 18452 9716
rect 18396 7980 18452 8036
rect 19068 9884 19124 9940
rect 18732 9660 18788 9716
rect 18732 9436 18788 9492
rect 18956 7586 19012 7588
rect 18956 7534 18958 7586
rect 18958 7534 19010 7586
rect 19010 7534 19012 7586
rect 18956 7532 19012 7534
rect 18396 6300 18452 6356
rect 18508 7420 18564 7476
rect 18284 5964 18340 6020
rect 18844 6748 18900 6804
rect 18396 5292 18452 5348
rect 18172 4172 18228 4228
rect 18284 5068 18340 5124
rect 18060 3500 18116 3556
rect 18396 4508 18452 4564
rect 18732 5180 18788 5236
rect 18620 4172 18676 4228
rect 18620 3276 18676 3332
rect 18508 2940 18564 2996
rect 18284 2828 18340 2884
rect 18396 1708 18452 1764
rect 18396 1036 18452 1092
rect 18844 3164 18900 3220
rect 18956 4732 19012 4788
rect 18844 924 18900 980
rect 18956 812 19012 868
rect 19516 11676 19572 11732
rect 19964 12796 20020 12852
rect 20188 13244 20244 13300
rect 20188 12012 20244 12068
rect 20300 12572 20356 12628
rect 20076 11900 20132 11956
rect 20076 11676 20132 11732
rect 19852 11116 19908 11172
rect 19740 10668 19796 10724
rect 19516 7756 19572 7812
rect 19628 8428 19684 8484
rect 20636 13356 20692 13412
rect 20524 12236 20580 12292
rect 21196 13186 21252 13188
rect 21196 13134 21198 13186
rect 21198 13134 21250 13186
rect 21250 13134 21252 13186
rect 21196 13132 21252 13134
rect 20860 12236 20916 12292
rect 20300 11228 20356 11284
rect 19964 10108 20020 10164
rect 19852 9996 19908 10052
rect 19740 8204 19796 8260
rect 19964 7868 20020 7924
rect 19740 7196 19796 7252
rect 19180 5628 19236 5684
rect 19180 4732 19236 4788
rect 19180 3554 19236 3556
rect 19180 3502 19182 3554
rect 19182 3502 19234 3554
rect 19234 3502 19236 3554
rect 19180 3500 19236 3502
rect 20524 9996 20580 10052
rect 20300 9324 20356 9380
rect 21084 11228 21140 11284
rect 21196 11788 21252 11844
rect 21084 10892 21140 10948
rect 20748 10556 20804 10612
rect 21756 13132 21812 13188
rect 21980 13804 22036 13860
rect 21756 12796 21812 12852
rect 21868 12684 21924 12740
rect 21756 11676 21812 11732
rect 21868 12236 21924 12292
rect 22092 12962 22148 12964
rect 22092 12910 22094 12962
rect 22094 12910 22146 12962
rect 22146 12910 22148 12962
rect 22092 12908 22148 12910
rect 23548 13468 23604 13524
rect 23996 13132 24052 13188
rect 24108 13468 24164 13524
rect 24444 13468 24500 13524
rect 24464 13354 24520 13356
rect 24332 13244 24388 13300
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24892 13356 24948 13412
rect 24672 13300 24728 13302
rect 25004 13244 25060 13300
rect 25228 13020 25284 13076
rect 25116 12962 25172 12964
rect 25116 12910 25118 12962
rect 25118 12910 25170 12962
rect 25170 12910 25172 12962
rect 25116 12908 25172 12910
rect 23100 12348 23156 12404
rect 23324 12572 23380 12628
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 23884 12402 23940 12404
rect 23884 12350 23886 12402
rect 23886 12350 23938 12402
rect 23938 12350 23940 12402
rect 23884 12348 23940 12350
rect 24556 12124 24612 12180
rect 22092 11452 22148 11508
rect 21196 9884 21252 9940
rect 22764 10332 22820 10388
rect 23324 11228 23380 11284
rect 22092 9660 22148 9716
rect 20972 9212 21028 9268
rect 22316 9548 22372 9604
rect 20860 9100 20916 9156
rect 21980 8652 22036 8708
rect 21196 8316 21252 8372
rect 21532 8258 21588 8260
rect 21532 8206 21534 8258
rect 21534 8206 21586 8258
rect 21586 8206 21588 8258
rect 21532 8204 21588 8206
rect 19740 1036 19796 1092
rect 20972 7532 21028 7588
rect 19068 476 19124 532
rect 20748 6636 20804 6692
rect 21868 7196 21924 7252
rect 20972 6188 21028 6244
rect 20076 3276 20132 3332
rect 20188 2828 20244 2884
rect 20188 1484 20244 1540
rect 20076 1372 20132 1428
rect 21980 7084 22036 7140
rect 21868 6412 21924 6468
rect 22540 9212 22596 9268
rect 22428 8930 22484 8932
rect 22428 8878 22430 8930
rect 22430 8878 22482 8930
rect 22482 8878 22484 8930
rect 22428 8876 22484 8878
rect 23436 9938 23492 9940
rect 23436 9886 23438 9938
rect 23438 9886 23490 9938
rect 23490 9886 23492 9938
rect 23436 9884 23492 9886
rect 24332 11788 24388 11844
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 24444 11340 24500 11396
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 24444 10892 24500 10948
rect 24668 10444 24724 10500
rect 25228 10780 25284 10836
rect 24332 10220 24388 10276
rect 24464 10218 24520 10220
rect 24108 10108 24164 10164
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24892 10220 24948 10276
rect 23996 9938 24052 9940
rect 23996 9886 23998 9938
rect 23998 9886 24050 9938
rect 24050 9886 24052 9938
rect 23996 9884 24052 9886
rect 23324 9212 23380 9268
rect 24892 9772 24948 9828
rect 23660 9436 23716 9492
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24220 9324 24276 9380
rect 23548 8540 23604 8596
rect 24332 8652 24388 8708
rect 22988 8428 23044 8484
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 25452 13186 25508 13188
rect 25452 13134 25454 13186
rect 25454 13134 25506 13186
rect 25506 13134 25508 13186
rect 25452 13132 25508 13134
rect 25564 12908 25620 12964
rect 25452 12012 25508 12068
rect 25452 10780 25508 10836
rect 25228 9436 25284 9492
rect 25340 9772 25396 9828
rect 25228 8988 25284 9044
rect 24892 8540 24948 8596
rect 25004 8652 25060 8708
rect 23548 7868 23604 7924
rect 23804 7866 23860 7868
rect 23660 7756 23716 7812
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24332 7868 24388 7924
rect 24012 7812 24068 7814
rect 24220 7756 24276 7812
rect 24780 7644 24836 7700
rect 22540 7084 22596 7140
rect 23660 7308 23716 7364
rect 23660 6972 23716 7028
rect 24332 7084 24388 7140
rect 22092 5964 22148 6020
rect 21196 5180 21252 5236
rect 21644 5292 21700 5348
rect 21532 4508 21588 4564
rect 21532 3724 21588 3780
rect 21420 3164 21476 3220
rect 21756 4284 21812 4340
rect 21756 3724 21812 3780
rect 21644 3164 21700 3220
rect 21420 2940 21476 2996
rect 21868 2828 21924 2884
rect 21980 5292 22036 5348
rect 21532 2658 21588 2660
rect 21532 2606 21534 2658
rect 21534 2606 21586 2658
rect 21586 2606 21588 2658
rect 21532 2604 21588 2606
rect 21756 2604 21812 2660
rect 22204 5292 22260 5348
rect 22092 4284 22148 4340
rect 23996 6690 24052 6692
rect 23996 6638 23998 6690
rect 23998 6638 24050 6690
rect 24050 6638 24052 6690
rect 23996 6636 24052 6638
rect 23804 6298 23860 6300
rect 23660 6188 23716 6244
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24220 6188 24276 6244
rect 25116 7084 25172 7140
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 25228 6412 25284 6468
rect 24332 5852 24388 5908
rect 25116 5964 25172 6020
rect 24332 5516 24388 5572
rect 24464 5514 24520 5516
rect 24220 5404 24276 5460
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24892 5516 24948 5572
rect 24672 5460 24728 5462
rect 23548 4396 23604 4452
rect 23660 4732 23716 4788
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24332 4732 24388 4788
rect 25116 4732 25172 4788
rect 25228 5852 25284 5908
rect 24012 4676 24068 4678
rect 24220 4620 24276 4676
rect 23772 4396 23828 4452
rect 21980 2044 22036 2100
rect 20748 1874 20804 1876
rect 20748 1822 20750 1874
rect 20750 1822 20802 1874
rect 20802 1822 20804 1874
rect 20748 1820 20804 1822
rect 20300 1372 20356 1428
rect 19964 140 20020 196
rect 20636 1148 20692 1204
rect 20860 1148 20916 1204
rect 20860 924 20916 980
rect 21980 364 22036 420
rect 1148 28 1204 84
rect 22204 2268 22260 2324
rect 23660 4060 23716 4116
rect 23884 4060 23940 4116
rect 24220 3948 24276 4004
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 23884 3724 23940 3780
rect 24220 3724 24276 3780
rect 23996 3612 24052 3668
rect 25340 4956 25396 5012
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 24332 3164 24388 3220
rect 24444 3052 24500 3108
rect 24668 2828 24724 2884
rect 23996 2716 24052 2772
rect 24668 2604 24724 2660
rect 23884 2380 23940 2436
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24892 2268 24948 2324
rect 25116 2380 25172 2436
rect 24780 2044 24836 2100
rect 23804 1594 23860 1596
rect 23660 1484 23716 1540
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24780 1596 24836 1652
rect 24012 1540 24068 1542
rect 24332 1484 24388 1540
rect 25116 2098 25172 2100
rect 25116 2046 25118 2098
rect 25118 2046 25170 2098
rect 25170 2046 25172 2098
rect 25116 2044 25172 2046
rect 25004 1484 25060 1540
rect 25228 1708 25284 1764
rect 25228 1484 25284 1540
rect 22988 1260 23044 1316
rect 22988 812 23044 868
rect 24464 810 24520 812
rect 23324 700 23380 756
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 22092 28 22148 84
rect 25788 12012 25844 12068
rect 25900 13916 25956 13972
rect 26012 13356 26068 13412
rect 26124 12460 26180 12516
rect 26124 11788 26180 11844
rect 26012 11564 26068 11620
rect 25900 10556 25956 10612
rect 26124 11452 26180 11508
rect 25676 10444 25732 10500
rect 25564 9548 25620 9604
rect 25564 8988 25620 9044
rect 25564 8428 25620 8484
rect 25564 8204 25620 8260
rect 25564 7868 25620 7924
rect 25564 3948 25620 4004
rect 25564 3276 25620 3332
rect 26684 13356 26740 13412
rect 27468 13804 27524 13860
rect 27244 13132 27300 13188
rect 27020 12572 27076 12628
rect 27020 12124 27076 12180
rect 26236 11228 26292 11284
rect 26796 9996 26852 10052
rect 26460 9660 26516 9716
rect 27916 13356 27972 13412
rect 27916 12460 27972 12516
rect 27916 12290 27972 12292
rect 27916 12238 27918 12290
rect 27918 12238 27970 12290
rect 27970 12238 27972 12290
rect 27916 12236 27972 12238
rect 27580 12124 27636 12180
rect 28028 11788 28084 11844
rect 28252 13244 28308 13300
rect 27468 11676 27524 11732
rect 27356 9660 27412 9716
rect 27804 11564 27860 11620
rect 27244 9548 27300 9604
rect 26908 9324 26964 9380
rect 26684 7980 26740 8036
rect 26796 9100 26852 9156
rect 26796 7868 26852 7924
rect 26908 7980 26964 8036
rect 26796 6524 26852 6580
rect 27132 6972 27188 7028
rect 27132 6300 27188 6356
rect 26908 6076 26964 6132
rect 25788 5180 25844 5236
rect 26572 5180 26628 5236
rect 26572 4172 26628 4228
rect 26012 4060 26068 4116
rect 25900 3612 25956 3668
rect 26012 2716 26068 2772
rect 27020 3500 27076 3556
rect 25900 2492 25956 2548
rect 26348 2492 26404 2548
rect 25900 1708 25956 1764
rect 26012 1260 26068 1316
rect 26236 1148 26292 1204
rect 25900 1036 25956 1092
rect 25564 812 25620 868
rect 27692 9436 27748 9492
rect 28028 11228 28084 11284
rect 27916 10668 27972 10724
rect 27916 7756 27972 7812
rect 27804 6524 27860 6580
rect 27692 5964 27748 6020
rect 27916 4844 27972 4900
rect 27244 4396 27300 4452
rect 27804 4732 27860 4788
rect 27580 4060 27636 4116
rect 28364 12348 28420 12404
rect 28364 11340 28420 11396
rect 28252 11228 28308 11284
rect 28700 13356 28756 13412
rect 28588 12796 28644 12852
rect 28476 10444 28532 10500
rect 28588 11900 28644 11956
rect 28476 10220 28532 10276
rect 28364 10108 28420 10164
rect 28364 9884 28420 9940
rect 28140 9324 28196 9380
rect 28476 8988 28532 9044
rect 28476 8764 28532 8820
rect 28140 5852 28196 5908
rect 28364 8428 28420 8484
rect 28476 7420 28532 7476
rect 28364 5852 28420 5908
rect 28924 12796 28980 12852
rect 29148 12572 29204 12628
rect 28812 12012 28868 12068
rect 29036 12066 29092 12068
rect 29036 12014 29038 12066
rect 29038 12014 29090 12066
rect 29090 12014 29092 12066
rect 29036 12012 29092 12014
rect 28924 11788 28980 11844
rect 29372 12572 29428 12628
rect 29820 12348 29876 12404
rect 30044 12460 30100 12516
rect 29148 11788 29204 11844
rect 29932 12236 29988 12292
rect 30716 14028 30772 14084
rect 30268 12460 30324 12516
rect 31052 12796 31108 12852
rect 30156 12236 30212 12292
rect 28924 11564 28980 11620
rect 28812 11004 28868 11060
rect 28700 9996 28756 10052
rect 28812 10444 28868 10500
rect 28812 9884 28868 9940
rect 29036 10444 29092 10500
rect 28700 9100 28756 9156
rect 28700 8316 28756 8372
rect 28700 6188 28756 6244
rect 28028 4732 28084 4788
rect 29820 9996 29876 10052
rect 29708 8764 29764 8820
rect 29820 7756 29876 7812
rect 29708 6972 29764 7028
rect 28812 6076 28868 6132
rect 30268 12124 30324 12180
rect 30044 9436 30100 9492
rect 30044 7980 30100 8036
rect 30156 8316 30212 8372
rect 29932 5964 29988 6020
rect 29260 5852 29316 5908
rect 29708 5852 29764 5908
rect 29148 5740 29204 5796
rect 28700 4508 28756 4564
rect 29036 5628 29092 5684
rect 27804 4060 27860 4116
rect 27580 3500 27636 3556
rect 28700 3388 28756 3444
rect 28588 2604 28644 2660
rect 28700 2492 28756 2548
rect 28924 3276 28980 3332
rect 27132 2380 27188 2436
rect 28476 2268 28532 2324
rect 26348 588 26404 644
rect 26796 1372 26852 1428
rect 27132 1372 27188 1428
rect 26908 700 26964 756
rect 29036 3164 29092 3220
rect 28476 1372 28532 1428
rect 29036 1372 29092 1428
rect 27244 700 27300 756
rect 28924 1260 28980 1316
rect 26796 364 26852 420
rect 29484 4732 29540 4788
rect 29484 3052 29540 3108
rect 29372 2940 29428 2996
rect 30828 11788 30884 11844
rect 30380 11676 30436 11732
rect 30492 10892 30548 10948
rect 30268 8204 30324 8260
rect 30380 9660 30436 9716
rect 30492 9548 30548 9604
rect 30380 6748 30436 6804
rect 30492 9100 30548 9156
rect 30604 8428 30660 8484
rect 30716 10892 30772 10948
rect 30604 7474 30660 7476
rect 30604 7422 30606 7474
rect 30606 7422 30658 7474
rect 30658 7422 30660 7474
rect 30604 7420 30660 7422
rect 30940 11618 30996 11620
rect 30940 11566 30942 11618
rect 30942 11566 30994 11618
rect 30994 11566 30996 11618
rect 30940 11564 30996 11566
rect 30828 8764 30884 8820
rect 30716 6972 30772 7028
rect 30828 7084 30884 7140
rect 30604 6748 30660 6804
rect 30268 6300 30324 6356
rect 30716 6524 30772 6580
rect 30380 6076 30436 6132
rect 30604 6076 30660 6132
rect 30380 5906 30436 5908
rect 30380 5854 30382 5906
rect 30382 5854 30434 5906
rect 30434 5854 30436 5906
rect 30380 5852 30436 5854
rect 30268 5180 30324 5236
rect 30268 4620 30324 4676
rect 30156 2828 30212 2884
rect 30268 3612 30324 3668
rect 29484 2604 29540 2660
rect 30268 1820 30324 1876
rect 29372 1596 29428 1652
rect 29148 1260 29204 1316
rect 30268 588 30324 644
rect 30716 2492 30772 2548
rect 30604 1708 30660 1764
rect 30940 6972 30996 7028
rect 31164 11900 31220 11956
rect 31500 13132 31556 13188
rect 31388 11116 31444 11172
rect 31724 13804 31780 13860
rect 31724 13132 31780 13188
rect 31836 10556 31892 10612
rect 31500 9996 31556 10052
rect 31724 10220 31780 10276
rect 31836 9884 31892 9940
rect 31724 9772 31780 9828
rect 31948 9772 32004 9828
rect 32284 13580 32340 13636
rect 32284 11564 32340 11620
rect 32396 12124 32452 12180
rect 32060 8316 32116 8372
rect 32172 9548 32228 9604
rect 31164 7362 31220 7364
rect 31164 7310 31166 7362
rect 31166 7310 31218 7362
rect 31218 7310 31220 7362
rect 31164 7308 31220 7310
rect 31164 7084 31220 7140
rect 31164 6748 31220 6804
rect 31836 6748 31892 6804
rect 31724 5794 31780 5796
rect 31724 5742 31726 5794
rect 31726 5742 31778 5794
rect 31778 5742 31780 5794
rect 31724 5740 31780 5742
rect 31052 4844 31108 4900
rect 31612 5068 31668 5124
rect 31612 4620 31668 4676
rect 31836 4060 31892 4116
rect 32284 8876 32340 8932
rect 32508 11788 32564 11844
rect 32732 12124 32788 12180
rect 32732 10444 32788 10500
rect 32620 8428 32676 8484
rect 32284 6524 32340 6580
rect 32620 8204 32676 8260
rect 32284 4508 32340 4564
rect 32844 7980 32900 8036
rect 32732 7868 32788 7924
rect 32732 7084 32788 7140
rect 32956 7756 33012 7812
rect 33180 12236 33236 12292
rect 32844 4844 32900 4900
rect 33628 12796 33684 12852
rect 33292 6748 33348 6804
rect 33292 4060 33348 4116
rect 33292 3836 33348 3892
rect 33628 10108 33684 10164
rect 33628 9548 33684 9604
rect 35196 13916 35252 13972
rect 34748 13692 34804 13748
rect 35084 13244 35140 13300
rect 34860 12572 34916 12628
rect 34636 11788 34692 11844
rect 34300 10892 34356 10948
rect 34412 10780 34468 10836
rect 34524 10892 34580 10948
rect 33852 9100 33908 9156
rect 34412 9212 34468 9268
rect 33516 8540 33572 8596
rect 33628 8428 33684 8484
rect 33852 8428 33908 8484
rect 33740 7644 33796 7700
rect 33628 5516 33684 5572
rect 33628 4956 33684 5012
rect 33404 3500 33460 3556
rect 33516 3836 33572 3892
rect 32396 3276 32452 3332
rect 32732 3276 32788 3332
rect 32844 2882 32900 2884
rect 32844 2830 32846 2882
rect 32846 2830 32898 2882
rect 32898 2830 32900 2882
rect 32844 2828 32900 2830
rect 33852 4396 33908 4452
rect 34412 4060 34468 4116
rect 33740 3164 33796 3220
rect 34188 3500 34244 3556
rect 34188 3052 34244 3108
rect 34412 3052 34468 3108
rect 33516 2268 33572 2324
rect 30940 1986 30996 1988
rect 30940 1934 30942 1986
rect 30942 1934 30994 1986
rect 30994 1934 30996 1986
rect 30940 1932 30996 1934
rect 34076 1932 34132 1988
rect 30828 1596 30884 1652
rect 30940 1708 30996 1764
rect 30492 588 30548 644
rect 32620 1708 32676 1764
rect 32956 1484 33012 1540
rect 31388 1260 31444 1316
rect 28924 364 28980 420
rect 28700 140 28756 196
rect 31612 1260 31668 1316
rect 31612 140 31668 196
rect 33628 1148 33684 1204
rect 33628 140 33684 196
rect 35532 13020 35588 13076
rect 35308 12012 35364 12068
rect 35084 11340 35140 11396
rect 35196 11900 35252 11956
rect 34860 11116 34916 11172
rect 34748 10780 34804 10836
rect 34972 9996 35028 10052
rect 34748 9212 34804 9268
rect 34748 8988 34804 9044
rect 34636 8204 34692 8260
rect 34972 8988 35028 9044
rect 34972 8652 35028 8708
rect 35084 8146 35140 8148
rect 35084 8094 35086 8146
rect 35086 8094 35138 8146
rect 35138 8094 35140 8146
rect 35084 8092 35140 8094
rect 35084 7868 35140 7924
rect 34972 6636 35028 6692
rect 34748 4396 34804 4452
rect 34860 5292 34916 5348
rect 34748 3724 34804 3780
rect 34860 2716 34916 2772
rect 35084 6076 35140 6132
rect 35084 5740 35140 5796
rect 35084 4060 35140 4116
rect 35532 11228 35588 11284
rect 35308 8092 35364 8148
rect 35420 9212 35476 9268
rect 35532 8540 35588 8596
rect 35868 13020 35924 13076
rect 35644 8204 35700 8260
rect 35756 12348 35812 12404
rect 35532 7756 35588 7812
rect 35532 7196 35588 7252
rect 35420 6972 35476 7028
rect 35420 6076 35476 6132
rect 35308 5180 35364 5236
rect 35308 4956 35364 5012
rect 35308 4620 35364 4676
rect 35308 3724 35364 3780
rect 35308 3164 35364 3220
rect 34972 2604 35028 2660
rect 35196 2604 35252 2660
rect 34636 2156 34692 2212
rect 34524 1260 34580 1316
rect 34412 1036 34468 1092
rect 35532 5852 35588 5908
rect 35532 4620 35588 4676
rect 35420 2828 35476 2884
rect 35308 1148 35364 1204
rect 35196 700 35252 756
rect 36540 13916 36596 13972
rect 36988 13244 37044 13300
rect 36876 12684 36932 12740
rect 37436 12572 37492 12628
rect 37324 12460 37380 12516
rect 36092 10780 36148 10836
rect 36988 10498 37044 10500
rect 36988 10446 36990 10498
rect 36990 10446 37042 10498
rect 37042 10446 37044 10498
rect 36988 10444 37044 10446
rect 36316 10332 36372 10388
rect 36652 9938 36708 9940
rect 36652 9886 36654 9938
rect 36654 9886 36706 9938
rect 36706 9886 36708 9938
rect 36652 9884 36708 9886
rect 36092 9826 36148 9828
rect 36092 9774 36094 9826
rect 36094 9774 36146 9826
rect 36146 9774 36148 9826
rect 36092 9772 36148 9774
rect 36316 9772 36372 9828
rect 36316 9436 36372 9492
rect 35868 8204 35924 8260
rect 36092 8540 36148 8596
rect 35756 7196 35812 7252
rect 36988 8316 37044 8372
rect 36652 7644 36708 7700
rect 36540 3554 36596 3556
rect 36540 3502 36542 3554
rect 36542 3502 36594 3554
rect 36594 3502 36596 3554
rect 36540 3500 36596 3502
rect 36428 3276 36484 3332
rect 36876 7644 36932 7700
rect 36652 3052 36708 3108
rect 36764 4508 36820 4564
rect 36092 1260 36148 1316
rect 35644 700 35700 756
rect 37100 7980 37156 8036
rect 37100 6972 37156 7028
rect 37100 6748 37156 6804
rect 37100 5516 37156 5572
rect 36988 5292 37044 5348
rect 36988 4450 37044 4452
rect 36988 4398 36990 4450
rect 36990 4398 37042 4450
rect 37042 4398 37044 4450
rect 36988 4396 37044 4398
rect 37100 3948 37156 4004
rect 37772 12236 37828 12292
rect 37660 10108 37716 10164
rect 37548 8988 37604 9044
rect 38220 13468 38276 13524
rect 38108 12796 38164 12852
rect 37884 11900 37940 11956
rect 38332 13020 38388 13076
rect 38556 14028 38612 14084
rect 38220 11676 38276 11732
rect 38332 12796 38388 12852
rect 37772 8540 37828 8596
rect 37324 3164 37380 3220
rect 36876 1372 36932 1428
rect 36988 2828 37044 2884
rect 37996 6412 38052 6468
rect 38220 6412 38276 6468
rect 38780 13692 38836 13748
rect 38556 10780 38612 10836
rect 38556 9100 38612 9156
rect 38780 9100 38836 9156
rect 39340 12908 39396 12964
rect 39452 12124 39508 12180
rect 39452 10108 39508 10164
rect 39564 11004 39620 11060
rect 39340 7980 39396 8036
rect 39228 7644 39284 7700
rect 38556 7420 38612 7476
rect 38556 7196 38612 7252
rect 39228 7196 39284 7252
rect 38332 6076 38388 6132
rect 40124 13468 40180 13524
rect 40236 13804 40292 13860
rect 40124 12908 40180 12964
rect 39788 11676 39844 11732
rect 39788 11004 39844 11060
rect 40012 11676 40068 11732
rect 40124 11340 40180 11396
rect 40236 12012 40292 12068
rect 39900 10780 39956 10836
rect 40124 10780 40180 10836
rect 40012 10220 40068 10276
rect 39676 7084 39732 7140
rect 39788 8316 39844 8372
rect 39564 5964 39620 6020
rect 39788 5852 39844 5908
rect 39900 6636 39956 6692
rect 38444 5404 38500 5460
rect 39340 5292 39396 5348
rect 38668 4396 38724 4452
rect 41020 12908 41076 12964
rect 41468 12236 41524 12292
rect 40572 11452 40628 11508
rect 41356 11900 41412 11956
rect 40348 11340 40404 11396
rect 40236 10668 40292 10724
rect 40460 10668 40516 10724
rect 40124 9212 40180 9268
rect 40236 9100 40292 9156
rect 40012 6524 40068 6580
rect 40124 7980 40180 8036
rect 41692 11900 41748 11956
rect 41804 11676 41860 11732
rect 41804 11452 41860 11508
rect 41692 10220 41748 10276
rect 41804 11228 41860 11284
rect 40460 8428 40516 8484
rect 40572 9884 40628 9940
rect 40236 7756 40292 7812
rect 40348 6972 40404 7028
rect 40460 7644 40516 7700
rect 40236 6524 40292 6580
rect 40460 6300 40516 6356
rect 40124 6076 40180 6132
rect 40124 4172 40180 4228
rect 40236 5628 40292 5684
rect 38668 3836 38724 3892
rect 40348 4956 40404 5012
rect 40348 4508 40404 4564
rect 40236 3836 40292 3892
rect 39788 3724 39844 3780
rect 38892 3612 38948 3668
rect 41468 7868 41524 7924
rect 41692 8988 41748 9044
rect 41580 7420 41636 7476
rect 40684 6188 40740 6244
rect 41916 10892 41972 10948
rect 42252 10610 42308 10612
rect 42252 10558 42254 10610
rect 42254 10558 42306 10610
rect 42306 10558 42308 10610
rect 42252 10556 42308 10558
rect 41916 8988 41972 9044
rect 43260 13244 43316 13300
rect 43596 13916 43652 13972
rect 42812 12684 42868 12740
rect 43036 12684 43092 12740
rect 42476 12572 42532 12628
rect 42812 10610 42868 10612
rect 42812 10558 42814 10610
rect 42814 10558 42866 10610
rect 42866 10558 42868 10610
rect 42812 10556 42868 10558
rect 42476 9212 42532 9268
rect 42588 8876 42644 8932
rect 42364 8092 42420 8148
rect 42140 7420 42196 7476
rect 42364 6524 42420 6580
rect 41804 5964 41860 6020
rect 41132 5852 41188 5908
rect 40684 4620 40740 4676
rect 38220 2940 38276 2996
rect 38668 3388 38724 3444
rect 37884 2770 37940 2772
rect 37884 2718 37886 2770
rect 37886 2718 37938 2770
rect 37938 2718 37940 2770
rect 37884 2716 37940 2718
rect 38668 2716 38724 2772
rect 37548 2492 37604 2548
rect 41244 5068 41300 5124
rect 41132 4284 41188 4340
rect 38892 2604 38948 2660
rect 40236 3164 40292 3220
rect 38444 2156 38500 2212
rect 36988 924 37044 980
rect 39340 1932 39396 1988
rect 39452 1708 39508 1764
rect 39452 1484 39508 1540
rect 39340 476 39396 532
rect 39452 1260 39508 1316
rect 40236 1036 40292 1092
rect 41468 3276 41524 3332
rect 42252 4226 42308 4228
rect 42252 4174 42254 4226
rect 42254 4174 42306 4226
rect 42306 4174 42308 4226
rect 42252 4172 42308 4174
rect 42252 3836 42308 3892
rect 41580 1596 41636 1652
rect 42028 1148 42084 1204
rect 41580 924 41636 980
rect 41468 476 41524 532
rect 40460 364 40516 420
rect 42252 3276 42308 3332
rect 42588 5180 42644 5236
rect 42588 4620 42644 4676
rect 42364 1708 42420 1764
rect 43708 12684 43764 12740
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 44716 13132 44772 13188
rect 44156 11900 44212 11956
rect 44268 12460 44324 12516
rect 43372 11340 43428 11396
rect 43148 8428 43204 8484
rect 43596 11004 43652 11060
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 44940 12124 44996 12180
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44268 11116 44324 11172
rect 43596 9884 43652 9940
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 44268 9324 44324 9380
rect 43372 8092 43428 8148
rect 44156 9212 44212 9268
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 43596 5516 43652 5572
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 44464 7082 44520 7084
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 44828 5180 44884 5236
rect 46396 13580 46452 13636
rect 46844 13468 46900 13524
rect 45948 13132 46004 13188
rect 45500 12796 45556 12852
rect 45276 11788 45332 11844
rect 45388 12012 45444 12068
rect 45388 11340 45444 11396
rect 45500 9996 45556 10052
rect 45612 9884 45668 9940
rect 45164 9714 45220 9716
rect 45164 9662 45166 9714
rect 45166 9662 45218 9714
rect 45218 9662 45220 9714
rect 45164 9660 45220 9662
rect 45388 9212 45444 9268
rect 46396 13020 46452 13076
rect 45948 12850 46004 12852
rect 45948 12798 45950 12850
rect 45950 12798 46002 12850
rect 46002 12798 46004 12850
rect 45948 12796 46004 12798
rect 46172 10780 46228 10836
rect 45724 9100 45780 9156
rect 45836 9324 45892 9380
rect 45612 8092 45668 8148
rect 45388 7532 45444 7588
rect 45500 7756 45556 7812
rect 45052 5068 45108 5124
rect 45388 6748 45444 6804
rect 44940 4956 44996 5012
rect 43596 3724 43652 3780
rect 45836 7756 45892 7812
rect 45612 7532 45668 7588
rect 46172 6524 46228 6580
rect 46284 10108 46340 10164
rect 45612 5628 45668 5684
rect 45500 4620 45556 4676
rect 45276 4284 45332 4340
rect 44464 3946 44520 3948
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 45724 3948 45780 4004
rect 44044 3724 44100 3780
rect 44044 3500 44100 3556
rect 44380 3442 44436 3444
rect 44380 3390 44382 3442
rect 44382 3390 44434 3442
rect 44434 3390 44436 3442
rect 44380 3388 44436 3390
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 46956 11564 47012 11620
rect 46732 9772 46788 9828
rect 47180 9100 47236 9156
rect 47068 8540 47124 8596
rect 47180 8204 47236 8260
rect 46284 2716 46340 2772
rect 46508 7420 46564 7476
rect 45724 1932 45780 1988
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 46620 7196 46676 7252
rect 47068 7980 47124 8036
rect 47068 6076 47124 6132
rect 47180 6188 47236 6244
rect 46620 3052 46676 3108
rect 46732 1596 46788 1652
rect 46508 1484 46564 1540
rect 47068 5068 47124 5124
rect 47180 4060 47236 4116
rect 47068 3276 47124 3332
rect 47404 12348 47460 12404
rect 47852 13580 47908 13636
rect 48188 13132 48244 13188
rect 47964 11954 48020 11956
rect 47964 11902 47966 11954
rect 47966 11902 48018 11954
rect 48018 11902 48020 11954
rect 47964 11900 48020 11902
rect 47628 10780 47684 10836
rect 47404 9884 47460 9940
rect 49084 13468 49140 13524
rect 48972 13186 49028 13188
rect 48972 13134 48974 13186
rect 48974 13134 49026 13186
rect 49026 13134 49028 13186
rect 48972 13132 49028 13134
rect 48636 12348 48692 12404
rect 49420 12402 49476 12404
rect 49420 12350 49422 12402
rect 49422 12350 49474 12402
rect 49474 12350 49476 12402
rect 49420 12348 49476 12350
rect 48188 11116 48244 11172
rect 48300 10332 48356 10388
rect 48860 12066 48916 12068
rect 48860 12014 48862 12066
rect 48862 12014 48914 12066
rect 48914 12014 48916 12066
rect 48860 12012 48916 12014
rect 49420 11788 49476 11844
rect 49196 11676 49252 11732
rect 49084 11452 49140 11508
rect 48748 10556 48804 10612
rect 47292 2940 47348 2996
rect 48300 9660 48356 9716
rect 47516 8652 47572 8708
rect 48076 8428 48132 8484
rect 48076 3164 48132 3220
rect 47628 2044 47684 2100
rect 47404 1820 47460 1876
rect 47068 1708 47124 1764
rect 47068 1372 47124 1428
rect 46956 1260 47012 1316
rect 43036 812 43092 868
rect 44828 924 44884 980
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 48524 8316 48580 8372
rect 48748 6076 48804 6132
rect 48972 8258 49028 8260
rect 48972 8206 48974 8258
rect 48974 8206 49026 8258
rect 49026 8206 49028 8258
rect 48972 8204 49028 8206
rect 49084 7644 49140 7700
rect 49980 13020 50036 13076
rect 50428 12348 50484 12404
rect 49532 11564 49588 11620
rect 49868 11788 49924 11844
rect 49644 11004 49700 11060
rect 49756 10108 49812 10164
rect 49420 8988 49476 9044
rect 49308 8930 49364 8932
rect 49308 8878 49310 8930
rect 49310 8878 49362 8930
rect 49362 8878 49364 8930
rect 49308 8876 49364 8878
rect 49196 7084 49252 7140
rect 48860 5852 48916 5908
rect 48636 5180 48692 5236
rect 48412 4508 48468 4564
rect 48412 3388 48468 3444
rect 48412 1148 48468 1204
rect 48300 924 48356 980
rect 47516 588 47572 644
rect 49420 2716 49476 2772
rect 49644 9996 49700 10052
rect 50316 11618 50372 11620
rect 50316 11566 50318 11618
rect 50318 11566 50370 11618
rect 50370 11566 50372 11618
rect 50316 11564 50372 11566
rect 50204 10498 50260 10500
rect 50204 10446 50206 10498
rect 50206 10446 50258 10498
rect 50258 10446 50260 10498
rect 50204 10444 50260 10446
rect 50316 9996 50372 10052
rect 50204 9826 50260 9828
rect 50204 9774 50206 9826
rect 50206 9774 50258 9826
rect 50258 9774 50260 9826
rect 50204 9772 50260 9774
rect 49868 9100 49924 9156
rect 50092 8092 50148 8148
rect 50428 9996 50484 10052
rect 51100 13468 51156 13524
rect 51772 13244 51828 13300
rect 52220 13132 52276 13188
rect 51772 12460 51828 12516
rect 50988 11788 51044 11844
rect 51212 11788 51268 11844
rect 50876 11564 50932 11620
rect 51436 11452 51492 11508
rect 51324 10780 51380 10836
rect 51660 11116 51716 11172
rect 50316 7532 50372 7588
rect 49532 1596 49588 1652
rect 49308 476 49364 532
rect 49980 364 50036 420
rect 50988 8258 51044 8260
rect 50988 8206 50990 8258
rect 50990 8206 51042 8258
rect 51042 8206 51044 8258
rect 50988 8204 51044 8206
rect 50540 8146 50596 8148
rect 50540 8094 50542 8146
rect 50542 8094 50594 8146
rect 50594 8094 50596 8146
rect 50540 8092 50596 8094
rect 50876 7756 50932 7812
rect 50540 3836 50596 3892
rect 50428 3500 50484 3556
rect 51212 9324 51268 9380
rect 51436 7474 51492 7476
rect 51436 7422 51438 7474
rect 51438 7422 51490 7474
rect 51490 7422 51492 7474
rect 51436 7420 51492 7422
rect 51660 6412 51716 6468
rect 51100 1708 51156 1764
rect 50988 1202 51044 1204
rect 50988 1150 50990 1202
rect 50990 1150 51042 1202
rect 51042 1150 51044 1202
rect 50988 1148 51044 1150
rect 51884 11618 51940 11620
rect 51884 11566 51886 11618
rect 51886 11566 51938 11618
rect 51938 11566 51940 11618
rect 51884 11564 51940 11566
rect 51884 10556 51940 10612
rect 52108 10108 52164 10164
rect 51996 9714 52052 9716
rect 51996 9662 51998 9714
rect 51998 9662 52050 9714
rect 52050 9662 52052 9714
rect 51996 9660 52052 9662
rect 52220 9436 52276 9492
rect 53116 13356 53172 13412
rect 52892 13074 52948 13076
rect 52892 13022 52894 13074
rect 52894 13022 52946 13074
rect 52946 13022 52948 13074
rect 52892 13020 52948 13022
rect 52556 12402 52612 12404
rect 52556 12350 52558 12402
rect 52558 12350 52610 12402
rect 52610 12350 52612 12402
rect 52556 12348 52612 12350
rect 53788 13020 53844 13076
rect 52556 11452 52612 11508
rect 53564 11340 53620 11396
rect 52892 9884 52948 9940
rect 52332 9212 52388 9268
rect 52108 8652 52164 8708
rect 52108 6748 52164 6804
rect 52220 7084 52276 7140
rect 52108 5292 52164 5348
rect 51996 5234 52052 5236
rect 51996 5182 51998 5234
rect 51998 5182 52050 5234
rect 52050 5182 52052 5234
rect 51996 5180 52052 5182
rect 53004 9266 53060 9268
rect 53004 9214 53006 9266
rect 53006 9214 53058 9266
rect 53058 9214 53060 9266
rect 53004 9212 53060 9214
rect 52668 8876 52724 8932
rect 52556 6972 52612 7028
rect 53900 10444 53956 10500
rect 53452 8764 53508 8820
rect 53340 8370 53396 8372
rect 53340 8318 53342 8370
rect 53342 8318 53394 8370
rect 53394 8318 53396 8370
rect 53340 8316 53396 8318
rect 53004 7868 53060 7924
rect 52444 6188 52500 6244
rect 52556 6076 52612 6132
rect 52332 4396 52388 4452
rect 52332 4060 52388 4116
rect 52220 3724 52276 3780
rect 52108 2770 52164 2772
rect 52108 2718 52110 2770
rect 52110 2718 52162 2770
rect 52162 2718 52164 2770
rect 52108 2716 52164 2718
rect 52108 1874 52164 1876
rect 52108 1822 52110 1874
rect 52110 1822 52162 1874
rect 52162 1822 52164 1874
rect 52108 1820 52164 1822
rect 51660 1260 51716 1316
rect 51996 924 52052 980
rect 53004 6130 53060 6132
rect 53004 6078 53006 6130
rect 53006 6078 53058 6130
rect 53058 6078 53060 6130
rect 53004 6076 53060 6078
rect 52892 5234 52948 5236
rect 52892 5182 52894 5234
rect 52894 5182 52946 5234
rect 52946 5182 52948 5234
rect 52892 5180 52948 5182
rect 52668 4508 52724 4564
rect 53340 5068 53396 5124
rect 54124 13244 54180 13300
rect 54236 12572 54292 12628
rect 54908 13580 54964 13636
rect 54460 11788 54516 11844
rect 54684 13468 54740 13524
rect 54348 11228 54404 11284
rect 54236 10556 54292 10612
rect 54012 9212 54068 9268
rect 54124 7308 54180 7364
rect 54124 6690 54180 6692
rect 54124 6638 54126 6690
rect 54126 6638 54178 6690
rect 54178 6638 54180 6690
rect 54124 6636 54180 6638
rect 53900 6076 53956 6132
rect 54124 6412 54180 6468
rect 53564 5794 53620 5796
rect 53564 5742 53566 5794
rect 53566 5742 53618 5794
rect 53618 5742 53620 5794
rect 53564 5740 53620 5742
rect 53564 4226 53620 4228
rect 53564 4174 53566 4226
rect 53566 4174 53618 4226
rect 53618 4174 53620 4226
rect 53564 4172 53620 4174
rect 53676 3948 53732 4004
rect 53452 3836 53508 3892
rect 53228 3388 53284 3444
rect 53564 3442 53620 3444
rect 53564 3390 53566 3442
rect 53566 3390 53618 3442
rect 53618 3390 53620 3442
rect 53564 3388 53620 3390
rect 53564 3164 53620 3220
rect 52780 2658 52836 2660
rect 52780 2606 52782 2658
rect 52782 2606 52834 2658
rect 52834 2606 52836 2658
rect 52780 2604 52836 2606
rect 54124 2380 54180 2436
rect 52556 2098 52612 2100
rect 52556 2046 52558 2098
rect 52558 2046 52610 2098
rect 52610 2046 52612 2098
rect 52556 2044 52612 2046
rect 54348 8540 54404 8596
rect 54572 10108 54628 10164
rect 54908 13186 54964 13188
rect 54908 13134 54910 13186
rect 54910 13134 54962 13186
rect 54962 13134 54964 13186
rect 54908 13132 54964 13134
rect 54684 9772 54740 9828
rect 54572 7196 54628 7252
rect 54572 5852 54628 5908
rect 54460 4844 54516 4900
rect 54572 4562 54628 4564
rect 54572 4510 54574 4562
rect 54574 4510 54626 4562
rect 54626 4510 54628 4562
rect 54572 4508 54628 4510
rect 55692 13356 55748 13412
rect 55804 13020 55860 13076
rect 56252 12796 56308 12852
rect 56364 13916 56420 13972
rect 55356 11900 55412 11956
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 54796 4060 54852 4116
rect 54796 3612 54852 3668
rect 55692 11228 55748 11284
rect 55132 9436 55188 9492
rect 55244 9548 55300 9604
rect 55132 8146 55188 8148
rect 55132 8094 55134 8146
rect 55134 8094 55186 8146
rect 55186 8094 55188 8146
rect 55132 8092 55188 8094
rect 55132 6860 55188 6916
rect 55132 6300 55188 6356
rect 55132 5794 55188 5796
rect 55132 5742 55134 5794
rect 55134 5742 55186 5794
rect 55186 5742 55188 5794
rect 55132 5740 55188 5742
rect 55468 10332 55524 10388
rect 56924 13020 56980 13076
rect 56924 11004 56980 11060
rect 57260 12124 57316 12180
rect 56588 10444 56644 10500
rect 56700 10780 56756 10836
rect 56700 9660 56756 9716
rect 56364 9324 56420 9380
rect 56140 8988 56196 9044
rect 55692 8316 55748 8372
rect 55468 8092 55524 8148
rect 55916 8092 55972 8148
rect 57260 7868 57316 7924
rect 56140 7698 56196 7700
rect 56140 7646 56142 7698
rect 56142 7646 56194 7698
rect 56194 7646 56196 7698
rect 56140 7644 56196 7646
rect 56140 6748 56196 6804
rect 55356 5180 55412 5236
rect 56140 5404 56196 5460
rect 55132 3724 55188 3780
rect 56140 4060 56196 4116
rect 54572 3164 54628 3220
rect 55132 3052 55188 3108
rect 56812 3388 56868 3444
rect 56140 2716 56196 2772
rect 54236 2268 54292 2324
rect 54908 2268 54964 2324
rect 53564 1874 53620 1876
rect 53564 1822 53566 1874
rect 53566 1822 53618 1874
rect 53618 1822 53620 1874
rect 53564 1820 53620 1822
rect 55132 1596 55188 1652
rect 52556 1484 52612 1540
rect 53564 1426 53620 1428
rect 53564 1374 53566 1426
rect 53566 1374 53618 1426
rect 53618 1374 53620 1426
rect 53564 1372 53620 1374
rect 56476 2604 56532 2660
rect 52332 700 52388 756
rect 51436 588 51492 644
rect 55580 252 55636 308
rect 52892 140 52948 196
rect 56812 476 56868 532
rect 56476 28 56532 84
<< metal3 >>
rect 6748 14140 20524 14196
rect 20580 14140 20590 14196
rect 20748 14140 38108 14196
rect 38164 14140 38174 14196
rect 6748 14084 6804 14140
rect 20748 14084 20804 14140
rect 6738 14028 6748 14084
rect 6804 14028 6814 14084
rect 14354 14028 14364 14084
rect 14420 14028 20804 14084
rect 20962 14028 20972 14084
rect 21028 14028 28028 14084
rect 28084 14028 28094 14084
rect 28242 14028 28252 14084
rect 28308 14028 30492 14084
rect 30548 14028 30558 14084
rect 30706 14028 30716 14084
rect 30772 14028 38556 14084
rect 38612 14028 38622 14084
rect 0 13972 112 14000
rect 57344 13972 57456 14000
rect 0 13916 18396 13972
rect 18452 13916 18462 13972
rect 20514 13916 20524 13972
rect 20580 13916 25900 13972
rect 25956 13916 25966 13972
rect 26852 13916 35196 13972
rect 35252 13916 35262 13972
rect 36530 13916 36540 13972
rect 36596 13916 43596 13972
rect 43652 13916 43662 13972
rect 56354 13916 56364 13972
rect 56420 13916 57456 13972
rect 0 13888 112 13916
rect 26852 13860 26908 13916
rect 57344 13888 57456 13916
rect 12002 13804 12012 13860
rect 12068 13804 21980 13860
rect 22036 13804 22046 13860
rect 23650 13804 23660 13860
rect 23716 13804 26908 13860
rect 27458 13804 27468 13860
rect 27524 13804 31724 13860
rect 31780 13804 31790 13860
rect 31938 13804 31948 13860
rect 32004 13804 32508 13860
rect 32564 13804 32574 13860
rect 32722 13804 32732 13860
rect 32788 13804 40236 13860
rect 40292 13804 40302 13860
rect 12114 13692 12124 13748
rect 12180 13692 17388 13748
rect 17444 13692 17454 13748
rect 17602 13692 17612 13748
rect 17668 13692 34748 13748
rect 34804 13692 34814 13748
rect 36978 13692 36988 13748
rect 37044 13692 38780 13748
rect 38836 13692 38846 13748
rect 5394 13580 5404 13636
rect 5460 13580 18844 13636
rect 18900 13580 18910 13636
rect 19618 13580 19628 13636
rect 19684 13580 32284 13636
rect 32340 13580 32350 13636
rect 32498 13580 32508 13636
rect 32564 13580 38444 13636
rect 38500 13580 38510 13636
rect 38882 13580 38892 13636
rect 38948 13580 46396 13636
rect 46452 13580 46462 13636
rect 47842 13580 47852 13636
rect 47908 13580 54908 13636
rect 54964 13580 54974 13636
rect 0 13524 112 13552
rect 57344 13524 57456 13552
rect 0 13468 1036 13524
rect 1092 13468 1102 13524
rect 3602 13468 3612 13524
rect 3668 13468 4732 13524
rect 4788 13468 4798 13524
rect 6290 13468 6300 13524
rect 6356 13468 20972 13524
rect 21028 13468 21038 13524
rect 23538 13468 23548 13524
rect 23604 13468 24108 13524
rect 24164 13468 24174 13524
rect 24434 13468 24444 13524
rect 24500 13468 38220 13524
rect 38276 13468 38286 13524
rect 38444 13468 40124 13524
rect 40180 13468 40190 13524
rect 44268 13468 46844 13524
rect 46900 13468 46910 13524
rect 49074 13468 49084 13524
rect 49140 13468 51100 13524
rect 51156 13468 51166 13524
rect 54674 13468 54684 13524
rect 54740 13468 57456 13524
rect 0 13440 112 13468
rect 38444 13412 38500 13468
rect 44268 13412 44324 13468
rect 57344 13440 57456 13468
rect 11330 13356 11340 13412
rect 11396 13356 13244 13412
rect 13300 13356 13310 13412
rect 13570 13356 13580 13412
rect 13636 13356 20636 13412
rect 20692 13356 20702 13412
rect 24882 13356 24892 13412
rect 24948 13356 26012 13412
rect 26068 13356 26078 13412
rect 26674 13356 26684 13412
rect 26740 13356 27916 13412
rect 27972 13356 27982 13412
rect 28130 13356 28140 13412
rect 28196 13356 28532 13412
rect 28690 13356 28700 13412
rect 28756 13356 38500 13412
rect 38602 13356 38612 13412
rect 38668 13356 44324 13412
rect 53106 13356 53116 13412
rect 53172 13356 55692 13412
rect 55748 13356 55758 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 28476 13300 28532 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 2146 13244 2156 13300
rect 2212 13244 4284 13300
rect 4340 13244 4350 13300
rect 5954 13244 5964 13300
rect 6020 13244 7420 13300
rect 7476 13244 7486 13300
rect 13458 13244 13468 13300
rect 13524 13244 20188 13300
rect 20244 13244 20254 13300
rect 20962 13244 20972 13300
rect 21028 13244 24332 13300
rect 24388 13244 24398 13300
rect 24994 13244 25004 13300
rect 25060 13244 28252 13300
rect 28308 13244 28318 13300
rect 28476 13244 33740 13300
rect 33796 13244 33806 13300
rect 35074 13244 35084 13300
rect 35140 13244 36988 13300
rect 37044 13244 37054 13300
rect 37212 13244 43260 13300
rect 43316 13244 43326 13300
rect 51762 13244 51772 13300
rect 51828 13244 54124 13300
rect 54180 13244 54190 13300
rect 37212 13188 37268 13244
rect 3714 13132 3724 13188
rect 3780 13132 5628 13188
rect 5684 13132 5694 13188
rect 7522 13132 7532 13188
rect 7588 13132 9212 13188
rect 9268 13132 9278 13188
rect 9762 13132 9772 13188
rect 9828 13132 11452 13188
rect 11508 13132 11518 13188
rect 11778 13132 11788 13188
rect 11844 13132 15820 13188
rect 15876 13132 15886 13188
rect 16034 13132 16044 13188
rect 16100 13132 17836 13188
rect 17892 13132 17902 13188
rect 18050 13132 18060 13188
rect 18116 13132 18900 13188
rect 21186 13132 21196 13188
rect 21252 13132 21756 13188
rect 21812 13132 21822 13188
rect 23986 13132 23996 13188
rect 24052 13132 25452 13188
rect 25508 13132 25518 13188
rect 25666 13132 25676 13188
rect 25732 13132 27076 13188
rect 27234 13132 27244 13188
rect 27300 13132 31500 13188
rect 31556 13132 31566 13188
rect 31714 13132 31724 13188
rect 31780 13132 33852 13188
rect 33908 13132 33918 13188
rect 34066 13132 34076 13188
rect 34132 13132 37268 13188
rect 37324 13132 44716 13188
rect 44772 13132 44782 13188
rect 45910 13132 45948 13188
rect 46004 13132 46014 13188
rect 48178 13132 48188 13188
rect 48244 13132 48972 13188
rect 49028 13132 49038 13188
rect 52210 13132 52220 13188
rect 52276 13132 54908 13188
rect 54964 13132 54974 13188
rect 0 13076 112 13104
rect 18844 13076 18900 13132
rect 27020 13076 27076 13132
rect 37324 13076 37380 13132
rect 57344 13076 57456 13104
rect 0 13020 364 13076
rect 420 13020 430 13076
rect 5282 13020 5292 13076
rect 5348 13020 13188 13076
rect 14914 13020 14924 13076
rect 14980 13020 16380 13076
rect 16436 13020 16446 13076
rect 17490 13020 17500 13076
rect 17556 13020 18620 13076
rect 18676 13020 18686 13076
rect 18844 13020 22372 13076
rect 23538 13020 23548 13076
rect 23604 13020 25004 13076
rect 25060 13020 25070 13076
rect 25218 13020 25228 13076
rect 25284 13020 26908 13076
rect 27020 13020 35532 13076
rect 35588 13020 35598 13076
rect 35858 13020 35868 13076
rect 35924 13020 37380 13076
rect 38322 13020 38332 13076
rect 38388 13020 46396 13076
rect 46452 13020 46462 13076
rect 49970 13020 49980 13076
rect 50036 13020 52892 13076
rect 52948 13020 52958 13076
rect 53778 13020 53788 13076
rect 53844 13020 55804 13076
rect 55860 13020 55870 13076
rect 56914 13020 56924 13076
rect 56980 13020 57456 13076
rect 0 12992 112 13020
rect 13132 12964 13188 13020
rect 22316 12964 22372 13020
rect 26852 12964 26908 13020
rect 57344 12992 57456 13020
rect 4274 12908 4284 12964
rect 4340 12908 6412 12964
rect 6468 12908 6478 12964
rect 9426 12908 9436 12964
rect 9492 12908 12908 12964
rect 12964 12908 12974 12964
rect 13132 12908 18284 12964
rect 18340 12908 18350 12964
rect 18620 12908 22092 12964
rect 22148 12908 22158 12964
rect 22316 12908 24220 12964
rect 24276 12908 24286 12964
rect 25106 12908 25116 12964
rect 25172 12908 25564 12964
rect 25620 12908 25630 12964
rect 26852 12908 39340 12964
rect 39396 12908 39406 12964
rect 40114 12908 40124 12964
rect 40180 12908 41020 12964
rect 41076 12908 41086 12964
rect 18620 12852 18676 12908
rect 6738 12796 6748 12852
rect 6804 12796 13300 12852
rect 13906 12796 13916 12852
rect 13972 12796 14588 12852
rect 14644 12796 14654 12852
rect 14802 12796 14812 12852
rect 14868 12796 18676 12852
rect 19282 12796 19292 12852
rect 19348 12796 19964 12852
rect 20020 12796 20030 12852
rect 21746 12796 21756 12852
rect 21812 12796 28588 12852
rect 28644 12796 28654 12852
rect 28914 12796 28924 12852
rect 28980 12796 31052 12852
rect 31108 12796 31118 12852
rect 31266 12796 31276 12852
rect 31332 12796 33292 12852
rect 33348 12796 33358 12852
rect 33618 12796 33628 12852
rect 33684 12796 38108 12852
rect 38164 12796 38174 12852
rect 38322 12796 38332 12852
rect 38388 12796 45500 12852
rect 45556 12796 45566 12852
rect 45938 12796 45948 12852
rect 46004 12796 56252 12852
rect 56308 12796 56318 12852
rect 13244 12740 13300 12796
rect 13244 12684 18620 12740
rect 18676 12684 18686 12740
rect 18844 12684 20972 12740
rect 21028 12684 21038 12740
rect 21858 12684 21868 12740
rect 21924 12684 32732 12740
rect 32788 12684 32798 12740
rect 36866 12684 36876 12740
rect 36932 12684 42812 12740
rect 42868 12684 42878 12740
rect 43026 12684 43036 12740
rect 43092 12684 43708 12740
rect 43764 12684 43774 12740
rect 0 12628 112 12656
rect 18844 12628 18900 12684
rect 57344 12628 57456 12656
rect 0 12572 476 12628
rect 532 12572 542 12628
rect 10322 12572 10332 12628
rect 10388 12572 11116 12628
rect 11172 12572 11182 12628
rect 11778 12572 11788 12628
rect 11844 12572 15820 12628
rect 15876 12572 15886 12628
rect 16034 12572 16044 12628
rect 16100 12572 18900 12628
rect 20290 12572 20300 12628
rect 20356 12572 23324 12628
rect 23380 12572 23390 12628
rect 25218 12572 25228 12628
rect 25284 12572 26908 12628
rect 27010 12572 27020 12628
rect 27076 12572 29148 12628
rect 29204 12572 29214 12628
rect 29362 12572 29372 12628
rect 29428 12572 34860 12628
rect 34916 12572 34926 12628
rect 37426 12572 37436 12628
rect 37492 12572 42476 12628
rect 42532 12572 42542 12628
rect 54226 12572 54236 12628
rect 54292 12572 57456 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 26852 12516 26908 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 57344 12544 57456 12572
rect 5954 12460 5964 12516
rect 6020 12460 16940 12516
rect 16996 12460 17006 12516
rect 17164 12460 18284 12516
rect 18340 12460 18350 12516
rect 18498 12460 18508 12516
rect 18564 12460 21756 12516
rect 21812 12460 21822 12516
rect 24210 12460 24220 12516
rect 24276 12460 26124 12516
rect 26180 12460 26190 12516
rect 26852 12460 27692 12516
rect 27748 12460 27758 12516
rect 27906 12460 27916 12516
rect 27972 12460 30044 12516
rect 30100 12460 30110 12516
rect 30258 12460 30268 12516
rect 30324 12460 37324 12516
rect 37380 12460 37390 12516
rect 44258 12460 44268 12516
rect 44324 12460 51772 12516
rect 51828 12460 51838 12516
rect 17164 12404 17220 12460
rect 2258 12348 2268 12404
rect 2324 12348 3388 12404
rect 3444 12348 3454 12404
rect 6962 12348 6972 12404
rect 7028 12348 7868 12404
rect 7924 12348 7934 12404
rect 8530 12348 8540 12404
rect 8596 12348 9660 12404
rect 9716 12348 9726 12404
rect 9884 12348 14812 12404
rect 14868 12348 14878 12404
rect 15810 12348 15820 12404
rect 15876 12348 17220 12404
rect 17714 12348 17724 12404
rect 17780 12348 18508 12404
rect 18564 12348 18574 12404
rect 18732 12348 22260 12404
rect 23090 12348 23100 12404
rect 23156 12348 23884 12404
rect 23940 12348 23950 12404
rect 24332 12348 28364 12404
rect 28420 12348 28430 12404
rect 29810 12348 29820 12404
rect 29876 12348 35756 12404
rect 35812 12348 35822 12404
rect 39330 12348 39340 12404
rect 39396 12348 47404 12404
rect 47460 12348 47470 12404
rect 48626 12348 48636 12404
rect 48692 12348 49420 12404
rect 49476 12348 49486 12404
rect 50418 12348 50428 12404
rect 50484 12348 52556 12404
rect 52612 12348 52622 12404
rect 9884 12292 9940 12348
rect 18732 12292 18788 12348
rect 22204 12292 22260 12348
rect 8418 12236 8428 12292
rect 8484 12236 9940 12292
rect 11218 12236 11228 12292
rect 11284 12236 14868 12292
rect 15922 12236 15932 12292
rect 15988 12236 16940 12292
rect 16996 12236 17006 12292
rect 17164 12236 18788 12292
rect 18844 12236 20524 12292
rect 20580 12236 20590 12292
rect 20850 12236 20860 12292
rect 20916 12236 21868 12292
rect 21924 12236 21934 12292
rect 22204 12236 23548 12292
rect 23604 12236 23614 12292
rect 0 12180 112 12208
rect 0 12124 588 12180
rect 644 12124 654 12180
rect 9874 12124 9884 12180
rect 9940 12124 14588 12180
rect 14644 12124 14654 12180
rect 0 12096 112 12124
rect 14812 12068 14868 12236
rect 17164 12180 17220 12236
rect 18844 12180 18900 12236
rect 24332 12180 24388 12348
rect 27906 12236 27916 12292
rect 27972 12236 29932 12292
rect 29988 12236 29998 12292
rect 30146 12236 30156 12292
rect 30212 12236 32956 12292
rect 33012 12236 33022 12292
rect 33170 12236 33180 12292
rect 33236 12236 36988 12292
rect 37044 12236 37054 12292
rect 37762 12236 37772 12292
rect 37828 12236 41468 12292
rect 41524 12236 41534 12292
rect 57344 12180 57456 12208
rect 15026 12124 15036 12180
rect 15092 12124 16156 12180
rect 16212 12124 16222 12180
rect 16482 12124 16492 12180
rect 16548 12124 17220 12180
rect 17378 12124 17388 12180
rect 17444 12124 18900 12180
rect 19394 12124 19404 12180
rect 19460 12124 24388 12180
rect 24546 12124 24556 12180
rect 24612 12124 27020 12180
rect 27076 12124 27086 12180
rect 27570 12124 27580 12180
rect 27636 12124 30268 12180
rect 30324 12124 30334 12180
rect 30482 12124 30492 12180
rect 30548 12124 32396 12180
rect 32452 12124 32462 12180
rect 32722 12124 32732 12180
rect 32788 12124 37324 12180
rect 37380 12124 37390 12180
rect 38612 12124 39228 12180
rect 39284 12124 39294 12180
rect 39442 12124 39452 12180
rect 39508 12124 44940 12180
rect 44996 12124 45006 12180
rect 57250 12124 57260 12180
rect 57316 12124 57456 12180
rect 38612 12068 38668 12124
rect 57344 12096 57456 12124
rect 4386 12012 4396 12068
rect 4452 12012 5068 12068
rect 5124 12012 5134 12068
rect 11890 12012 11900 12068
rect 11956 12012 14644 12068
rect 14812 12012 16044 12068
rect 16100 12012 16110 12068
rect 16258 12012 16268 12068
rect 16324 12012 17276 12068
rect 17332 12012 17342 12068
rect 17826 12012 17836 12068
rect 17892 12012 19964 12068
rect 20020 12012 20030 12068
rect 20178 12012 20188 12068
rect 20244 12012 25452 12068
rect 25508 12012 25518 12068
rect 25778 12012 25788 12068
rect 25844 12012 28812 12068
rect 28868 12012 28878 12068
rect 29026 12012 29036 12068
rect 29092 12012 35308 12068
rect 35364 12012 35374 12068
rect 35522 12012 35532 12068
rect 35588 12012 38668 12068
rect 40226 12012 40236 12068
rect 40292 12012 45388 12068
rect 45444 12012 45454 12068
rect 48822 12012 48860 12068
rect 48916 12012 48926 12068
rect 2930 11900 2940 11956
rect 2996 11900 3388 11956
rect 3444 11900 3454 11956
rect 4284 11900 8148 11956
rect 13346 11900 13356 11956
rect 13412 11900 14252 11956
rect 14308 11900 14318 11956
rect 4284 11844 4340 11900
rect 2258 11788 2268 11844
rect 2324 11788 4340 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 0 11676 4172 11732
rect 4228 11676 4238 11732
rect 0 11648 112 11676
rect 8092 11620 8148 11900
rect 14588 11844 14644 12012
rect 14914 11900 14924 11956
rect 14980 11900 16268 11956
rect 16324 11900 16334 11956
rect 16492 11900 20076 11956
rect 20132 11900 20142 11956
rect 20290 11900 20300 11956
rect 20356 11900 21700 11956
rect 21858 11900 21868 11956
rect 21924 11900 28364 11956
rect 28420 11900 28430 11956
rect 28578 11900 28588 11956
rect 28644 11900 31164 11956
rect 31220 11900 31230 11956
rect 31388 11900 34972 11956
rect 35028 11900 35038 11956
rect 35186 11900 35196 11956
rect 35252 11900 37884 11956
rect 37940 11900 37950 11956
rect 38098 11900 38108 11956
rect 38164 11900 41356 11956
rect 41412 11900 41422 11956
rect 41682 11900 41692 11956
rect 41748 11900 44156 11956
rect 44212 11900 44222 11956
rect 47954 11900 47964 11956
rect 48020 11900 55356 11956
rect 55412 11900 55422 11956
rect 16492 11844 16548 11900
rect 21644 11844 21700 11900
rect 31388 11844 31444 11900
rect 9538 11788 9548 11844
rect 9604 11788 12068 11844
rect 12786 11788 12796 11844
rect 12852 11788 14420 11844
rect 14588 11788 16548 11844
rect 16706 11788 16716 11844
rect 16772 11788 21196 11844
rect 21252 11788 21262 11844
rect 21644 11788 22036 11844
rect 12012 11732 12068 11788
rect 14364 11732 14420 11788
rect 21980 11732 22036 11788
rect 22316 11788 24332 11844
rect 24388 11788 24398 11844
rect 26114 11788 26124 11844
rect 26180 11788 27860 11844
rect 28018 11788 28028 11844
rect 28084 11788 28924 11844
rect 28980 11788 28990 11844
rect 29138 11788 29148 11844
rect 29204 11788 30492 11844
rect 30548 11788 30558 11844
rect 30818 11788 30828 11844
rect 30884 11788 31444 11844
rect 32498 11788 32508 11844
rect 32564 11788 34636 11844
rect 34692 11788 34702 11844
rect 35308 11788 42196 11844
rect 45266 11788 45276 11844
rect 45332 11788 49420 11844
rect 49476 11788 49486 11844
rect 49858 11788 49868 11844
rect 49924 11788 50988 11844
rect 51044 11788 51054 11844
rect 51202 11788 51212 11844
rect 51268 11788 54460 11844
rect 54516 11788 54526 11844
rect 22316 11732 22372 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 27804 11732 27860 11788
rect 35308 11732 35364 11788
rect 42140 11732 42196 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 57344 11732 57456 11760
rect 8306 11676 8316 11732
rect 8372 11676 11788 11732
rect 11844 11676 11854 11732
rect 12012 11676 13580 11732
rect 13636 11676 13646 11732
rect 14364 11676 19516 11732
rect 19572 11676 19582 11732
rect 20066 11676 20076 11732
rect 20132 11676 21756 11732
rect 21812 11676 21822 11732
rect 21980 11676 22372 11732
rect 24892 11676 27468 11732
rect 27524 11676 27534 11732
rect 27804 11676 30380 11732
rect 30436 11676 30446 11732
rect 30706 11676 30716 11732
rect 30772 11676 35364 11732
rect 38210 11676 38220 11732
rect 38276 11676 39788 11732
rect 39844 11676 39854 11732
rect 40002 11676 40012 11732
rect 40068 11676 41804 11732
rect 41860 11676 41870 11732
rect 42140 11676 43876 11732
rect 49186 11676 49196 11732
rect 49252 11676 57456 11732
rect 24892 11620 24948 11676
rect 43820 11620 43876 11676
rect 57344 11648 57456 11676
rect 4610 11564 4620 11620
rect 4676 11564 5180 11620
rect 5236 11564 5246 11620
rect 8092 11564 12012 11620
rect 12068 11564 12078 11620
rect 15092 11564 17948 11620
rect 18004 11564 18014 11620
rect 18386 11564 18396 11620
rect 18452 11564 21756 11620
rect 21812 11564 21822 11620
rect 21970 11564 21980 11620
rect 22036 11564 24948 11620
rect 26002 11564 26012 11620
rect 26068 11564 27804 11620
rect 27860 11564 27870 11620
rect 28914 11564 28924 11620
rect 28980 11564 30940 11620
rect 30996 11564 31006 11620
rect 32274 11564 32284 11620
rect 32340 11564 43596 11620
rect 43652 11564 43662 11620
rect 43820 11564 46956 11620
rect 47012 11564 47022 11620
rect 49522 11564 49532 11620
rect 49588 11564 50316 11620
rect 50372 11564 50382 11620
rect 50866 11564 50876 11620
rect 50932 11564 51884 11620
rect 51940 11564 51950 11620
rect 15092 11508 15148 11564
rect 1026 11452 1036 11508
rect 1092 11452 8652 11508
rect 8708 11452 8718 11508
rect 9212 11452 15148 11508
rect 15810 11452 15820 11508
rect 15876 11452 22092 11508
rect 22148 11452 22158 11508
rect 26114 11452 26124 11508
rect 26180 11452 40572 11508
rect 40628 11452 40638 11508
rect 41794 11452 41804 11508
rect 41860 11452 49084 11508
rect 49140 11452 49150 11508
rect 51426 11452 51436 11508
rect 51492 11452 52556 11508
rect 52612 11452 52622 11508
rect 466 11340 476 11396
rect 532 11340 4956 11396
rect 5012 11340 5022 11396
rect 0 11284 112 11312
rect 0 11228 980 11284
rect 1586 11228 1596 11284
rect 1652 11228 6076 11284
rect 6132 11228 6142 11284
rect 0 11200 112 11228
rect 924 11060 980 11228
rect 9212 11172 9268 11452
rect 11442 11340 11452 11396
rect 11508 11340 13692 11396
rect 13748 11340 13758 11396
rect 13906 11340 13916 11396
rect 13972 11340 24444 11396
rect 24500 11340 24510 11396
rect 28354 11340 28364 11396
rect 28420 11340 35084 11396
rect 35140 11340 35150 11396
rect 35308 11340 40124 11396
rect 40180 11340 40190 11396
rect 40338 11340 40348 11396
rect 40404 11340 43372 11396
rect 43428 11340 43438 11396
rect 45378 11340 45388 11396
rect 45444 11340 53564 11396
rect 53620 11340 53630 11396
rect 35308 11284 35364 11340
rect 57344 11284 57456 11312
rect 2594 11116 2604 11172
rect 2660 11116 9268 11172
rect 10220 11228 16716 11284
rect 16772 11228 16782 11284
rect 16940 11228 20300 11284
rect 20356 11228 20366 11284
rect 21074 11228 21084 11284
rect 21140 11228 23324 11284
rect 23380 11228 23390 11284
rect 23538 11228 23548 11284
rect 23604 11228 26012 11284
rect 26068 11228 26078 11284
rect 26226 11228 26236 11284
rect 26292 11228 28028 11284
rect 28084 11228 28094 11284
rect 28242 11228 28252 11284
rect 28308 11228 35364 11284
rect 35522 11228 35532 11284
rect 35588 11228 41804 11284
rect 41860 11228 41870 11284
rect 43586 11228 43596 11284
rect 43652 11228 54348 11284
rect 54404 11228 54414 11284
rect 55682 11228 55692 11284
rect 55748 11228 57456 11284
rect 914 11004 924 11060
rect 980 11004 990 11060
rect 4386 11004 4396 11060
rect 4452 11004 9884 11060
rect 9940 11004 9950 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 5170 10892 5180 10948
rect 5236 10892 9660 10948
rect 9716 10892 9726 10948
rect 0 10836 112 10864
rect 10220 10836 10276 11228
rect 16940 11172 16996 11228
rect 57344 11200 57456 11228
rect 10434 11116 10444 11172
rect 10500 11116 15428 11172
rect 16370 11116 16380 11172
rect 16436 11116 16996 11172
rect 17154 11116 17164 11172
rect 17220 11116 19628 11172
rect 19684 11116 19694 11172
rect 19842 11116 19852 11172
rect 19908 11116 31388 11172
rect 31444 11116 31454 11172
rect 31602 11116 31612 11172
rect 31668 11116 34076 11172
rect 34132 11116 34142 11172
rect 34850 11116 34860 11172
rect 34916 11116 44268 11172
rect 44324 11116 44334 11172
rect 48178 11116 48188 11172
rect 48244 11116 51660 11172
rect 51716 11116 51726 11172
rect 15372 11060 15428 11116
rect 11106 11004 11116 11060
rect 11172 11004 12684 11060
rect 12740 11004 12750 11060
rect 13010 11004 13020 11060
rect 13076 11004 15148 11060
rect 15204 11004 15214 11060
rect 15372 11004 21980 11060
rect 22036 11004 22046 11060
rect 24210 11004 24220 11060
rect 24276 11004 28532 11060
rect 28802 11004 28812 11060
rect 28868 11004 39564 11060
rect 39620 11004 39630 11060
rect 39778 11004 39788 11060
rect 39844 11004 43596 11060
rect 43652 11004 43662 11060
rect 49634 11004 49644 11060
rect 49700 11004 56924 11060
rect 56980 11004 56990 11060
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 28476 10948 28532 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 0 10780 1596 10836
rect 1652 10780 1662 10836
rect 3266 10780 3276 10836
rect 3332 10780 10276 10836
rect 11004 10892 21084 10948
rect 21140 10892 21150 10948
rect 21298 10892 21308 10948
rect 21364 10892 23548 10948
rect 23604 10892 23614 10948
rect 24434 10892 24444 10948
rect 24500 10892 28252 10948
rect 28308 10892 28318 10948
rect 28476 10892 30492 10948
rect 30548 10892 30558 10948
rect 30706 10892 30716 10948
rect 30772 10892 34300 10948
rect 34356 10892 34366 10948
rect 34514 10892 34524 10948
rect 34580 10892 41916 10948
rect 41972 10892 41982 10948
rect 0 10752 112 10780
rect 11004 10724 11060 10892
rect 57344 10836 57456 10864
rect 11442 10780 11452 10836
rect 11508 10780 12124 10836
rect 12180 10780 12190 10836
rect 14130 10780 14140 10836
rect 14196 10780 14588 10836
rect 14644 10780 14654 10836
rect 15092 10780 17164 10836
rect 17220 10780 17230 10836
rect 18610 10780 18620 10836
rect 18676 10780 25228 10836
rect 25284 10780 25294 10836
rect 25442 10780 25452 10836
rect 25508 10780 34412 10836
rect 34468 10780 34478 10836
rect 34738 10780 34748 10836
rect 34804 10780 36092 10836
rect 36148 10780 36158 10836
rect 38546 10780 38556 10836
rect 38612 10780 39900 10836
rect 39956 10780 39966 10836
rect 40114 10780 40124 10836
rect 40180 10780 46172 10836
rect 46228 10780 46238 10836
rect 47590 10780 47628 10836
rect 47684 10780 47694 10836
rect 50372 10780 51324 10836
rect 51380 10780 51390 10836
rect 56690 10780 56700 10836
rect 56756 10780 57456 10836
rect 15092 10724 15148 10780
rect 50372 10724 50428 10780
rect 57344 10752 57456 10780
rect 3154 10668 3164 10724
rect 3220 10668 8316 10724
rect 8372 10668 8382 10724
rect 9090 10668 9100 10724
rect 9156 10668 11060 10724
rect 11778 10668 11788 10724
rect 11844 10668 15148 10724
rect 15586 10668 15596 10724
rect 15652 10668 19740 10724
rect 19796 10668 19806 10724
rect 20066 10668 20076 10724
rect 20132 10668 26572 10724
rect 26628 10668 26638 10724
rect 27906 10668 27916 10724
rect 27972 10668 40236 10724
rect 40292 10668 40302 10724
rect 40450 10668 40460 10724
rect 40516 10668 50428 10724
rect 130 10556 140 10612
rect 196 10556 3332 10612
rect 5954 10556 5964 10612
rect 6020 10556 16828 10612
rect 16884 10556 16894 10612
rect 17042 10556 17052 10612
rect 17108 10556 18284 10612
rect 18340 10556 18350 10612
rect 19618 10556 19628 10612
rect 19684 10556 20748 10612
rect 20804 10556 20814 10612
rect 20972 10556 25228 10612
rect 25284 10556 25294 10612
rect 25890 10556 25900 10612
rect 25956 10556 31836 10612
rect 31892 10556 31902 10612
rect 33618 10556 33628 10612
rect 33684 10556 42252 10612
rect 42308 10556 42318 10612
rect 42802 10556 42812 10612
rect 42868 10556 48748 10612
rect 48804 10556 48814 10612
rect 51874 10556 51884 10612
rect 51940 10556 54236 10612
rect 54292 10556 54302 10612
rect 3276 10500 3332 10556
rect 20972 10500 21028 10556
rect 2790 10444 2828 10500
rect 2884 10444 2894 10500
rect 3276 10444 9548 10500
rect 9604 10444 9614 10500
rect 9762 10444 9772 10500
rect 9828 10444 13916 10500
rect 13972 10444 13982 10500
rect 14130 10444 14140 10500
rect 14196 10444 21028 10500
rect 21980 10444 24220 10500
rect 24276 10444 24286 10500
rect 24658 10444 24668 10500
rect 24724 10444 25676 10500
rect 25732 10444 25742 10500
rect 28466 10444 28476 10500
rect 28532 10444 28812 10500
rect 28868 10444 28878 10500
rect 29026 10444 29036 10500
rect 29092 10444 30716 10500
rect 30772 10444 30782 10500
rect 31490 10444 31500 10500
rect 31556 10444 32732 10500
rect 32788 10444 32798 10500
rect 33506 10444 33516 10500
rect 33572 10444 36596 10500
rect 36978 10444 36988 10500
rect 37044 10444 50204 10500
rect 50260 10444 50270 10500
rect 53890 10444 53900 10500
rect 53956 10444 56588 10500
rect 56644 10444 56654 10500
rect 0 10388 112 10416
rect 21980 10388 22036 10444
rect 36540 10388 36596 10444
rect 57344 10388 57456 10416
rect 0 10332 2884 10388
rect 7746 10332 7756 10388
rect 7812 10332 8428 10388
rect 8484 10332 8494 10388
rect 8642 10332 8652 10388
rect 8708 10332 22036 10388
rect 22754 10332 22764 10388
rect 22820 10332 36316 10388
rect 36372 10332 36382 10388
rect 36540 10332 42028 10388
rect 42084 10332 42094 10388
rect 43484 10332 48300 10388
rect 48356 10332 48366 10388
rect 55458 10332 55468 10388
rect 55524 10332 57456 10388
rect 0 10304 112 10332
rect 2828 10276 2884 10332
rect 2818 10220 2828 10276
rect 2884 10220 2894 10276
rect 8082 10220 8092 10276
rect 8148 10220 11620 10276
rect 12226 10220 12236 10276
rect 12292 10220 15036 10276
rect 15092 10220 15102 10276
rect 15250 10220 15260 10276
rect 15316 10220 16828 10276
rect 16884 10220 16894 10276
rect 17042 10220 17052 10276
rect 17108 10220 24332 10276
rect 24388 10220 24398 10276
rect 24882 10220 24892 10276
rect 24948 10220 28476 10276
rect 28532 10220 28542 10276
rect 30258 10220 30268 10276
rect 30324 10220 31500 10276
rect 31556 10220 31566 10276
rect 31714 10220 31724 10276
rect 31780 10220 35196 10276
rect 35252 10220 35262 10276
rect 35410 10220 35420 10276
rect 35476 10220 38668 10276
rect 40002 10220 40012 10276
rect 40068 10220 41692 10276
rect 41748 10220 41758 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 11564 10164 11620 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 38612 10164 38668 10220
rect 43484 10164 43540 10332
rect 57344 10304 57456 10332
rect 45500 10220 50428 10276
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 45500 10164 45556 10220
rect 50372 10164 50428 10220
rect 6178 10108 6188 10164
rect 6244 10108 10444 10164
rect 10500 10108 10510 10164
rect 11564 10108 16492 10164
rect 16548 10108 16558 10164
rect 16930 10108 16940 10164
rect 16996 10108 19964 10164
rect 20020 10108 20030 10164
rect 20188 10108 24108 10164
rect 24164 10108 24174 10164
rect 26572 10108 27300 10164
rect 28354 10108 28364 10164
rect 28420 10108 33628 10164
rect 33684 10108 33694 10164
rect 34748 10108 37660 10164
rect 37716 10108 37726 10164
rect 38612 10108 39452 10164
rect 39508 10108 39518 10164
rect 41916 10108 43540 10164
rect 45276 10108 45556 10164
rect 46274 10108 46284 10164
rect 46340 10108 49756 10164
rect 49812 10108 49822 10164
rect 50372 10108 52108 10164
rect 52164 10108 52174 10164
rect 54562 10108 54572 10164
rect 54628 10108 55468 10164
rect 354 9996 364 10052
rect 420 9996 1764 10052
rect 2482 9996 2492 10052
rect 2548 9996 5124 10052
rect 5282 9996 5292 10052
rect 5348 9996 19852 10052
rect 19908 9996 19918 10052
rect 0 9940 112 9968
rect 1708 9940 1764 9996
rect 5068 9940 5124 9996
rect 20188 9940 20244 10108
rect 26572 10052 26628 10108
rect 27244 10052 27300 10108
rect 34748 10052 34804 10108
rect 41916 10052 41972 10108
rect 45276 10052 45332 10108
rect 20514 9996 20524 10052
rect 20580 9996 26628 10052
rect 26786 9996 26796 10052
rect 26908 9996 26928 10052
rect 27244 9996 28700 10052
rect 28756 9996 28766 10052
rect 29810 9996 29820 10052
rect 29876 9996 31276 10052
rect 31332 9996 31342 10052
rect 31490 9996 31500 10052
rect 31556 9996 34804 10052
rect 34962 9996 34972 10052
rect 35028 9996 41972 10052
rect 42028 9996 45332 10052
rect 45490 9996 45500 10052
rect 45556 9996 49644 10052
rect 49700 9996 49710 10052
rect 50306 9996 50316 10052
rect 50372 9996 50428 10052
rect 50484 9996 50494 10052
rect 42028 9940 42084 9996
rect 55412 9940 55468 10108
rect 57344 9940 57456 9968
rect 0 9884 140 9940
rect 196 9884 206 9940
rect 1708 9884 3388 9940
rect 5068 9884 11228 9940
rect 11284 9884 11294 9940
rect 11442 9884 11452 9940
rect 11508 9884 14700 9940
rect 14756 9884 14766 9940
rect 15362 9884 15372 9940
rect 15428 9884 16828 9940
rect 16884 9884 16894 9940
rect 19058 9884 19068 9940
rect 19124 9884 20244 9940
rect 21186 9884 21196 9940
rect 21252 9884 23436 9940
rect 23492 9884 23502 9940
rect 23986 9884 23996 9940
rect 24052 9884 28364 9940
rect 28420 9884 28430 9940
rect 28802 9884 28812 9940
rect 28868 9884 31612 9940
rect 31668 9884 31678 9940
rect 31826 9884 31836 9940
rect 31892 9884 36652 9940
rect 36708 9884 36718 9940
rect 40562 9884 40572 9940
rect 40628 9884 42084 9940
rect 43586 9884 43596 9940
rect 43652 9884 45612 9940
rect 45668 9884 45678 9940
rect 47394 9884 47404 9940
rect 47460 9884 52892 9940
rect 52948 9884 52958 9940
rect 55412 9884 57456 9940
rect 0 9856 112 9884
rect 3332 9828 3388 9884
rect 57344 9856 57456 9884
rect 1250 9772 1260 9828
rect 1316 9772 1820 9828
rect 1876 9772 1886 9828
rect 3332 9772 8316 9828
rect 8372 9772 8382 9828
rect 8530 9772 8540 9828
rect 8596 9772 10108 9828
rect 10164 9772 10174 9828
rect 10882 9772 10892 9828
rect 10948 9772 16492 9828
rect 16548 9772 16558 9828
rect 16706 9772 16716 9828
rect 16772 9772 21196 9828
rect 21252 9772 21262 9828
rect 21970 9772 21980 9828
rect 22036 9772 24892 9828
rect 24948 9772 24958 9828
rect 25330 9772 25340 9828
rect 25396 9772 26740 9828
rect 29362 9772 29372 9828
rect 29428 9772 31724 9828
rect 31780 9772 31790 9828
rect 31938 9772 31948 9828
rect 32004 9772 36092 9828
rect 36148 9772 36158 9828
rect 36306 9772 36316 9828
rect 36372 9772 46732 9828
rect 46788 9772 46798 9828
rect 50194 9772 50204 9828
rect 50260 9772 54684 9828
rect 54740 9772 54750 9828
rect 26684 9716 26740 9772
rect 578 9660 588 9716
rect 644 9660 6188 9716
rect 6244 9660 6254 9716
rect 6402 9660 6412 9716
rect 6468 9660 18396 9716
rect 18452 9660 18462 9716
rect 18722 9660 18732 9716
rect 18788 9660 21812 9716
rect 22082 9660 22092 9716
rect 22148 9660 26460 9716
rect 26516 9660 26526 9716
rect 26684 9660 27356 9716
rect 27412 9660 27422 9716
rect 30370 9660 30380 9716
rect 30436 9660 35420 9716
rect 35476 9660 35486 9716
rect 45154 9660 45164 9716
rect 45220 9660 48300 9716
rect 48356 9660 48366 9716
rect 51986 9660 51996 9716
rect 52052 9660 56700 9716
rect 56756 9660 56766 9716
rect 2930 9548 2940 9604
rect 2996 9548 3388 9604
rect 3490 9548 3500 9604
rect 3556 9548 9772 9604
rect 9828 9548 9838 9604
rect 10098 9548 10108 9604
rect 10164 9548 11452 9604
rect 11508 9548 11518 9604
rect 11778 9548 11788 9604
rect 11844 9548 13804 9604
rect 13860 9548 13870 9604
rect 14028 9548 15260 9604
rect 15316 9548 15326 9604
rect 15474 9548 15484 9604
rect 15540 9548 21028 9604
rect 0 9492 112 9520
rect 3332 9492 3388 9548
rect 14028 9492 14084 9548
rect 0 9436 1148 9492
rect 1204 9436 1214 9492
rect 3332 9436 3612 9492
rect 3668 9436 3678 9492
rect 4946 9436 4956 9492
rect 5012 9436 8092 9492
rect 8148 9436 8158 9492
rect 9874 9436 9884 9492
rect 9940 9436 13356 9492
rect 13412 9436 13422 9492
rect 13682 9436 13692 9492
rect 13748 9436 14084 9492
rect 14690 9436 14700 9492
rect 14756 9436 15148 9492
rect 15204 9436 15214 9492
rect 15362 9436 15372 9492
rect 15428 9436 18732 9492
rect 18788 9436 18798 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 20972 9380 21028 9548
rect 21756 9492 21812 9660
rect 22306 9548 22316 9604
rect 22372 9548 25564 9604
rect 25620 9548 25630 9604
rect 26898 9548 26908 9604
rect 26964 9548 27244 9604
rect 27300 9548 27310 9604
rect 27458 9548 27468 9604
rect 27524 9548 30156 9604
rect 30212 9548 30222 9604
rect 30482 9548 30492 9604
rect 30548 9548 32172 9604
rect 32228 9548 32238 9604
rect 32386 9548 32396 9604
rect 32452 9548 33404 9604
rect 33460 9548 33470 9604
rect 33618 9548 33628 9604
rect 33684 9548 55244 9604
rect 55300 9548 55310 9604
rect 57344 9492 57456 9520
rect 21756 9436 23660 9492
rect 23716 9436 23726 9492
rect 25218 9436 25228 9492
rect 25284 9436 27692 9492
rect 27748 9436 27758 9492
rect 27916 9436 29372 9492
rect 29428 9436 29438 9492
rect 30034 9436 30044 9492
rect 30100 9436 36316 9492
rect 36372 9436 36382 9492
rect 44258 9436 44268 9492
rect 44324 9436 52220 9492
rect 52276 9436 52286 9492
rect 55122 9436 55132 9492
rect 55188 9436 57456 9492
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 27916 9380 27972 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 57344 9408 57456 9436
rect 6066 9324 6076 9380
rect 6132 9324 9996 9380
rect 10052 9324 10062 9380
rect 11554 9324 11564 9380
rect 11620 9324 20300 9380
rect 20356 9324 20366 9380
rect 20972 9324 23660 9380
rect 23716 9324 23726 9380
rect 24210 9324 24220 9380
rect 24276 9324 26684 9380
rect 26740 9324 26750 9380
rect 26898 9324 26908 9380
rect 26964 9324 27972 9380
rect 28130 9324 28140 9380
rect 28196 9324 38780 9380
rect 38836 9324 38846 9380
rect 44258 9324 44268 9380
rect 44324 9324 45836 9380
rect 45892 9324 45902 9380
rect 51202 9324 51212 9380
rect 51268 9324 56364 9380
rect 56420 9324 56430 9380
rect 3042 9212 3052 9268
rect 3108 9212 20692 9268
rect 20962 9212 20972 9268
rect 21028 9212 22540 9268
rect 22596 9212 22606 9268
rect 23314 9212 23324 9268
rect 23380 9212 32956 9268
rect 33012 9212 33022 9268
rect 33730 9212 33740 9268
rect 33796 9212 34132 9268
rect 34402 9212 34412 9268
rect 34468 9212 34748 9268
rect 34804 9212 34814 9268
rect 35410 9212 35420 9268
rect 35476 9212 40124 9268
rect 40180 9212 40190 9268
rect 42466 9212 42476 9268
rect 42532 9212 44156 9268
rect 44212 9212 44222 9268
rect 45378 9212 45388 9268
rect 45444 9212 52332 9268
rect 52388 9212 52398 9268
rect 52994 9212 53004 9268
rect 53060 9212 54012 9268
rect 54068 9212 54078 9268
rect 1820 9100 20076 9156
rect 20132 9100 20142 9156
rect 0 9044 112 9072
rect 1820 9044 1876 9100
rect 20636 9044 20692 9212
rect 34076 9156 34132 9212
rect 20850 9100 20860 9156
rect 20916 9100 26796 9156
rect 26852 9100 26862 9156
rect 27132 9100 28700 9156
rect 28756 9100 28766 9156
rect 28914 9100 28924 9156
rect 28980 9100 30268 9156
rect 30324 9100 30334 9156
rect 30482 9100 30492 9156
rect 30548 9100 33852 9156
rect 33908 9100 33918 9156
rect 34076 9100 38556 9156
rect 38612 9100 38622 9156
rect 38770 9100 38780 9156
rect 38836 9100 38892 9156
rect 38948 9100 38958 9156
rect 40226 9100 40236 9156
rect 40292 9100 45724 9156
rect 45780 9100 45790 9156
rect 47170 9100 47180 9156
rect 47236 9100 49868 9156
rect 49924 9100 49934 9156
rect 27132 9044 27188 9100
rect 57344 9044 57456 9072
rect 0 8988 1876 9044
rect 3602 8988 3612 9044
rect 3668 8988 5180 9044
rect 5236 8988 5246 9044
rect 6850 8988 6860 9044
rect 6916 8988 12404 9044
rect 12674 8988 12684 9044
rect 12740 8988 13580 9044
rect 13636 8988 13646 9044
rect 13794 8988 13804 9044
rect 13860 8988 16044 9044
rect 16100 8988 16110 9044
rect 16258 8988 16268 9044
rect 16324 8988 19628 9044
rect 19684 8988 19694 9044
rect 20636 8988 25228 9044
rect 25284 8988 25294 9044
rect 25554 8988 25564 9044
rect 25620 8988 27188 9044
rect 28466 8988 28476 9044
rect 28532 8988 34748 9044
rect 34804 8988 34814 9044
rect 34962 8988 34972 9044
rect 35028 8988 36876 9044
rect 36932 8988 36942 9044
rect 37538 8988 37548 9044
rect 37604 8988 41692 9044
rect 41748 8988 41758 9044
rect 41906 8988 41916 9044
rect 41972 8988 49420 9044
rect 49476 8988 49486 9044
rect 56130 8988 56140 9044
rect 56196 8988 57456 9044
rect 0 8960 112 8988
rect 12348 8932 12404 8988
rect 57344 8960 57456 8988
rect 2594 8876 2604 8932
rect 2660 8876 4900 8932
rect 10322 8876 10332 8932
rect 10388 8876 12124 8932
rect 12180 8876 12190 8932
rect 12348 8876 22428 8932
rect 22484 8876 22494 8932
rect 23426 8876 23436 8932
rect 23492 8876 28028 8932
rect 28084 8876 28094 8932
rect 28242 8876 28252 8932
rect 28308 8876 32284 8932
rect 32340 8876 32350 8932
rect 32498 8876 32508 8932
rect 32564 8876 42588 8932
rect 42644 8876 42654 8932
rect 49298 8876 49308 8932
rect 49364 8876 52668 8932
rect 52724 8876 52734 8932
rect 2482 8652 2492 8708
rect 2548 8652 2828 8708
rect 2884 8652 2894 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 4844 8596 4900 8876
rect 9986 8764 9996 8820
rect 10052 8764 11676 8820
rect 11732 8764 11742 8820
rect 13346 8764 13356 8820
rect 13412 8764 15260 8820
rect 15316 8764 15326 8820
rect 15922 8764 15932 8820
rect 15988 8764 28476 8820
rect 28532 8764 28542 8820
rect 29698 8764 29708 8820
rect 29764 8764 30828 8820
rect 30884 8764 30894 8820
rect 31042 8764 31052 8820
rect 31108 8764 32564 8820
rect 32946 8764 32956 8820
rect 33012 8764 53452 8820
rect 53508 8764 53518 8820
rect 32508 8708 32564 8764
rect 10220 8652 13356 8708
rect 13412 8652 13422 8708
rect 13570 8652 13580 8708
rect 13636 8652 16604 8708
rect 16660 8652 16670 8708
rect 19506 8652 19516 8708
rect 19572 8652 20356 8708
rect 21970 8652 21980 8708
rect 22036 8652 24332 8708
rect 24388 8652 24398 8708
rect 24994 8652 25004 8708
rect 25060 8652 32284 8708
rect 32340 8652 32350 8708
rect 32508 8652 34972 8708
rect 35028 8652 35038 8708
rect 35186 8652 35196 8708
rect 35252 8652 44268 8708
rect 44324 8652 44334 8708
rect 47506 8652 47516 8708
rect 47572 8652 52108 8708
rect 52164 8652 52174 8708
rect 0 8540 1260 8596
rect 1316 8540 1326 8596
rect 4844 8540 9996 8596
rect 10052 8540 10062 8596
rect 0 8512 112 8540
rect 10220 8484 10276 8652
rect 20300 8596 20356 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 57344 8596 57456 8624
rect 10434 8540 10444 8596
rect 10500 8540 15148 8596
rect 15092 8484 15148 8540
rect 15372 8540 20076 8596
rect 20132 8540 20142 8596
rect 20300 8540 23548 8596
rect 23604 8540 23614 8596
rect 24882 8540 24892 8596
rect 24948 8540 32172 8596
rect 32228 8540 32238 8596
rect 32396 8540 33516 8596
rect 33572 8540 33582 8596
rect 33842 8540 33852 8596
rect 33908 8540 35532 8596
rect 35588 8540 35598 8596
rect 36082 8540 36092 8596
rect 36148 8540 37772 8596
rect 37828 8540 37838 8596
rect 38780 8540 44156 8596
rect 44212 8540 44222 8596
rect 45378 8540 45388 8596
rect 45444 8540 47068 8596
rect 47124 8540 47134 8596
rect 54338 8540 54348 8596
rect 54404 8540 57456 8596
rect 15372 8484 15428 8540
rect 32396 8484 32452 8540
rect 38780 8484 38836 8540
rect 57344 8512 57456 8540
rect 1596 8428 10276 8484
rect 10546 8428 10556 8484
rect 10612 8428 14924 8484
rect 14980 8428 14990 8484
rect 15092 8428 15428 8484
rect 15586 8428 15596 8484
rect 15652 8428 19628 8484
rect 19684 8428 19694 8484
rect 20972 8428 22820 8484
rect 22978 8428 22988 8484
rect 23044 8428 25564 8484
rect 25620 8428 25630 8484
rect 26852 8428 28364 8484
rect 28420 8428 28430 8484
rect 30594 8428 30604 8484
rect 30660 8428 32452 8484
rect 32610 8428 32620 8484
rect 32676 8428 33628 8484
rect 33684 8428 33694 8484
rect 33842 8428 33852 8484
rect 33908 8428 38276 8484
rect 38434 8428 38444 8484
rect 38500 8428 38836 8484
rect 38892 8428 40460 8484
rect 40516 8428 40526 8484
rect 43138 8428 43148 8484
rect 43204 8428 48076 8484
rect 48132 8428 48142 8484
rect 1596 8372 1652 8428
rect 20972 8372 21028 8428
rect 22764 8372 22820 8428
rect 26852 8372 26908 8428
rect 38220 8372 38276 8428
rect 38892 8372 38948 8428
rect 1586 8316 1596 8372
rect 1652 8316 1662 8372
rect 6290 8316 6300 8372
rect 6356 8316 7084 8372
rect 7140 8316 7150 8372
rect 7308 8316 13468 8372
rect 13524 8316 13534 8372
rect 14802 8316 14812 8372
rect 14868 8316 21028 8372
rect 21186 8316 21196 8372
rect 21252 8316 21812 8372
rect 22764 8316 24892 8372
rect 24948 8316 24958 8372
rect 25116 8316 26908 8372
rect 28690 8316 28700 8372
rect 28756 8316 29932 8372
rect 29988 8316 29998 8372
rect 30146 8316 30156 8372
rect 30212 8316 32060 8372
rect 32116 8316 32126 8372
rect 32274 8316 32284 8372
rect 32340 8316 36988 8372
rect 37044 8316 37054 8372
rect 38220 8316 38948 8372
rect 39778 8316 39788 8372
rect 39844 8316 48524 8372
rect 48580 8316 48590 8372
rect 53330 8316 53340 8372
rect 53396 8316 55692 8372
rect 55748 8316 55758 8372
rect 7308 8260 7364 8316
rect 21756 8260 21812 8316
rect 25116 8260 25172 8316
rect 2230 8204 2268 8260
rect 2324 8204 2334 8260
rect 4162 8204 4172 8260
rect 4228 8204 7364 8260
rect 7634 8204 7644 8260
rect 7700 8204 10332 8260
rect 10388 8204 10398 8260
rect 11666 8204 11676 8260
rect 11732 8204 15484 8260
rect 15540 8204 15550 8260
rect 15698 8204 15708 8260
rect 15764 8204 19516 8260
rect 19572 8204 19582 8260
rect 19730 8204 19740 8260
rect 19796 8204 21532 8260
rect 21588 8204 21598 8260
rect 21756 8204 25172 8260
rect 25554 8204 25564 8260
rect 25620 8204 30044 8260
rect 30100 8204 30110 8260
rect 30258 8204 30268 8260
rect 30324 8204 32620 8260
rect 32676 8204 32686 8260
rect 34626 8204 34636 8260
rect 34692 8204 35644 8260
rect 35700 8204 35710 8260
rect 35858 8204 35868 8260
rect 35924 8204 35962 8260
rect 38770 8204 38780 8260
rect 38836 8204 47180 8260
rect 47236 8204 47246 8260
rect 48962 8204 48972 8260
rect 49028 8204 50988 8260
rect 51044 8204 51054 8260
rect 0 8148 112 8176
rect 57344 8148 57456 8176
rect 0 8092 3276 8148
rect 3332 8092 3342 8148
rect 6290 8092 6300 8148
rect 6356 8092 8316 8148
rect 8372 8092 8382 8148
rect 8866 8092 8876 8148
rect 8932 8092 11452 8148
rect 11508 8092 11518 8148
rect 13468 8092 35084 8148
rect 35140 8092 35150 8148
rect 35298 8092 35308 8148
rect 35364 8092 42364 8148
rect 42420 8092 42430 8148
rect 43362 8092 43372 8148
rect 43428 8092 44660 8148
rect 45602 8092 45612 8148
rect 45668 8092 50092 8148
rect 50148 8092 50158 8148
rect 50372 8092 50540 8148
rect 50596 8092 50606 8148
rect 55122 8092 55132 8148
rect 55188 8092 55468 8148
rect 55524 8092 55534 8148
rect 55906 8092 55916 8148
rect 55972 8092 57456 8148
rect 0 8064 112 8092
rect 13468 8036 13524 8092
rect 44604 8036 44660 8092
rect 50372 8036 50428 8092
rect 57344 8064 57456 8092
rect 6626 7980 6636 8036
rect 6692 7980 13524 8036
rect 13682 7980 13692 8036
rect 13748 7980 17948 8036
rect 18004 7980 18014 8036
rect 18386 7980 18396 8036
rect 18452 7980 19852 8036
rect 19908 7980 19918 8036
rect 20066 7980 20076 8036
rect 20132 7980 26684 8036
rect 26740 7980 26750 8036
rect 26898 7980 26908 8036
rect 26964 7980 30044 8036
rect 30100 7980 30110 8036
rect 30258 7980 30268 8036
rect 30324 7980 32844 8036
rect 32900 7980 32910 8036
rect 33058 7980 33068 8036
rect 33124 7980 37100 8036
rect 37156 7980 37166 8036
rect 39330 7980 39340 8036
rect 39396 7980 40124 8036
rect 40180 7980 40190 8036
rect 44604 7980 46732 8036
rect 46788 7980 46798 8036
rect 47058 7980 47068 8036
rect 47124 7980 50428 8036
rect 6076 7868 8876 7924
rect 8932 7868 8942 7924
rect 9202 7868 9212 7924
rect 9268 7868 19964 7924
rect 20020 7868 20030 7924
rect 20178 7868 20188 7924
rect 20244 7868 23548 7924
rect 23604 7868 23614 7924
rect 24322 7868 24332 7924
rect 24388 7868 25564 7924
rect 25620 7868 25630 7924
rect 26786 7868 26796 7924
rect 26852 7868 32732 7924
rect 32788 7868 32798 7924
rect 32946 7868 32956 7924
rect 33012 7868 33236 7924
rect 33394 7868 33404 7924
rect 33460 7868 34860 7924
rect 34916 7868 34926 7924
rect 35074 7868 35084 7924
rect 35140 7868 41468 7924
rect 41524 7868 41534 7924
rect 52994 7868 53004 7924
rect 53060 7868 57260 7924
rect 57316 7868 57326 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 0 7700 112 7728
rect 6076 7700 6132 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 33180 7812 33236 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 6290 7756 6300 7812
rect 6356 7756 11564 7812
rect 11620 7756 11630 7812
rect 13346 7756 13356 7812
rect 13412 7756 18508 7812
rect 18564 7756 18574 7812
rect 19506 7756 19516 7812
rect 19572 7756 23660 7812
rect 23716 7756 23726 7812
rect 24210 7756 24220 7812
rect 24276 7756 27916 7812
rect 27972 7756 27982 7812
rect 28242 7756 28252 7812
rect 28308 7756 29820 7812
rect 29876 7756 29886 7812
rect 30034 7756 30044 7812
rect 30100 7756 32956 7812
rect 33012 7756 33022 7812
rect 33180 7756 35308 7812
rect 35364 7756 35374 7812
rect 35522 7756 35532 7812
rect 35588 7756 40236 7812
rect 40292 7756 40302 7812
rect 44146 7756 44156 7812
rect 44212 7756 45500 7812
rect 45556 7756 45566 7812
rect 45826 7756 45836 7812
rect 45892 7756 50876 7812
rect 50932 7756 50942 7812
rect 57344 7700 57456 7728
rect 0 7644 1204 7700
rect 1362 7644 1372 7700
rect 1428 7644 6132 7700
rect 6850 7644 6860 7700
rect 6916 7644 11788 7700
rect 11844 7644 11854 7700
rect 12002 7644 12012 7700
rect 12068 7644 13692 7700
rect 13748 7644 13758 7700
rect 13916 7644 24780 7700
rect 24836 7644 24846 7700
rect 25004 7644 33516 7700
rect 33572 7644 33582 7700
rect 33730 7644 33740 7700
rect 33796 7644 36652 7700
rect 36708 7644 36718 7700
rect 36866 7644 36876 7700
rect 36932 7644 39228 7700
rect 39284 7644 39294 7700
rect 40450 7644 40460 7700
rect 40516 7644 49084 7700
rect 49140 7644 49150 7700
rect 56130 7644 56140 7700
rect 56196 7644 57456 7700
rect 0 7616 112 7644
rect 1148 7588 1204 7644
rect 13916 7588 13972 7644
rect 25004 7588 25060 7644
rect 57344 7616 57456 7644
rect 1148 7532 3052 7588
rect 3108 7532 3118 7588
rect 6738 7532 6748 7588
rect 6804 7532 13972 7588
rect 14130 7532 14140 7588
rect 14196 7532 18956 7588
rect 19012 7532 19022 7588
rect 20962 7532 20972 7588
rect 21028 7532 25060 7588
rect 25116 7532 45388 7588
rect 45444 7532 45454 7588
rect 45602 7532 45612 7588
rect 45668 7532 50316 7588
rect 50372 7532 50382 7588
rect 25116 7476 25172 7532
rect 1698 7420 1708 7476
rect 1764 7420 10108 7476
rect 10164 7420 10174 7476
rect 10322 7420 10332 7476
rect 10388 7420 14252 7476
rect 14308 7420 14318 7476
rect 15138 7420 15148 7476
rect 15204 7420 16268 7476
rect 16324 7420 16334 7476
rect 16818 7420 16828 7476
rect 16884 7420 18060 7476
rect 18116 7420 18126 7476
rect 18498 7420 18508 7476
rect 18564 7420 25172 7476
rect 26898 7420 26908 7476
rect 26964 7420 28252 7476
rect 28308 7420 28318 7476
rect 28466 7420 28476 7476
rect 28532 7420 30604 7476
rect 30660 7420 30670 7476
rect 30828 7420 38332 7476
rect 38388 7420 38398 7476
rect 38546 7420 38556 7476
rect 38612 7420 41580 7476
rect 41636 7420 41646 7476
rect 42130 7420 42140 7476
rect 42196 7420 46508 7476
rect 46564 7420 46574 7476
rect 46722 7420 46732 7476
rect 46788 7420 51436 7476
rect 51492 7420 51502 7476
rect 30828 7364 30884 7420
rect 3490 7308 3500 7364
rect 3556 7308 7756 7364
rect 7812 7308 7822 7364
rect 9986 7308 9996 7364
rect 10052 7308 23436 7364
rect 23492 7308 23502 7364
rect 23650 7308 23660 7364
rect 23716 7308 25060 7364
rect 25218 7308 25228 7364
rect 25284 7308 29932 7364
rect 29988 7308 29998 7364
rect 30146 7308 30156 7364
rect 30212 7308 30884 7364
rect 31154 7308 31164 7364
rect 31220 7308 54124 7364
rect 54180 7308 54190 7364
rect 0 7252 112 7280
rect 25004 7252 25060 7308
rect 57344 7252 57456 7280
rect 0 7196 1596 7252
rect 1652 7196 1662 7252
rect 2370 7196 2380 7252
rect 2436 7196 10332 7252
rect 10388 7196 10398 7252
rect 10546 7196 10556 7252
rect 10612 7196 11676 7252
rect 11732 7196 11742 7252
rect 11890 7196 11900 7252
rect 11956 7196 16828 7252
rect 16884 7196 16894 7252
rect 17154 7196 17164 7252
rect 17220 7196 19740 7252
rect 19796 7196 19806 7252
rect 20178 7196 20188 7252
rect 20244 7196 21308 7252
rect 21364 7196 21374 7252
rect 21858 7196 21868 7252
rect 21924 7196 24948 7252
rect 25004 7196 35532 7252
rect 35588 7196 35598 7252
rect 35746 7196 35756 7252
rect 35812 7196 38556 7252
rect 38612 7196 38622 7252
rect 39218 7196 39228 7252
rect 39284 7196 46620 7252
rect 46676 7196 46686 7252
rect 54562 7196 54572 7252
rect 54628 7196 57456 7252
rect 0 7168 112 7196
rect 2930 7084 2940 7140
rect 2996 7084 4284 7140
rect 4340 7084 4350 7140
rect 7970 7084 7980 7140
rect 8036 7084 9772 7140
rect 9828 7084 9838 7140
rect 10658 7084 10668 7140
rect 10724 7084 14700 7140
rect 14756 7084 14766 7140
rect 15250 7084 15260 7140
rect 15316 7084 17836 7140
rect 17892 7084 17902 7140
rect 18050 7084 18060 7140
rect 18116 7084 21980 7140
rect 22036 7084 22046 7140
rect 22530 7084 22540 7140
rect 22596 7084 24332 7140
rect 24388 7084 24398 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 24892 7028 24948 7196
rect 57344 7168 57456 7196
rect 25106 7084 25116 7140
rect 25172 7084 30828 7140
rect 30884 7084 30894 7140
rect 31154 7084 31164 7140
rect 31220 7084 32508 7140
rect 32564 7084 32574 7140
rect 32722 7084 32732 7140
rect 32788 7084 39676 7140
rect 39732 7084 39742 7140
rect 49186 7084 49196 7140
rect 49252 7084 52220 7140
rect 52276 7084 52286 7140
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 1026 6972 1036 7028
rect 1092 6972 3164 7028
rect 3220 6972 3230 7028
rect 9762 6972 9772 7028
rect 9828 6972 15596 7028
rect 15652 6972 15662 7028
rect 15810 6972 15820 7028
rect 15876 6972 23660 7028
rect 23716 6972 23726 7028
rect 24892 6972 26908 7028
rect 26964 6972 26974 7028
rect 27122 6972 27132 7028
rect 27188 6972 29708 7028
rect 29764 6972 29774 7028
rect 29922 6972 29932 7028
rect 29988 6972 30716 7028
rect 30772 6972 30782 7028
rect 30930 6972 30940 7028
rect 30996 6972 35420 7028
rect 35476 6972 35486 7028
rect 37090 6972 37100 7028
rect 37156 6972 40348 7028
rect 40404 6972 40414 7028
rect 44828 6972 52556 7028
rect 52612 6972 52622 7028
rect 44828 6916 44884 6972
rect 3266 6860 3276 6916
rect 3332 6860 8428 6916
rect 8484 6860 8494 6916
rect 10098 6860 10108 6916
rect 10164 6860 15708 6916
rect 15764 6860 15774 6916
rect 18620 6860 33404 6916
rect 33460 6860 33470 6916
rect 33628 6860 44884 6916
rect 44940 6860 55132 6916
rect 55188 6860 55198 6916
rect 0 6804 112 6832
rect 0 6748 10164 6804
rect 10434 6748 10444 6804
rect 10500 6748 13804 6804
rect 13860 6748 13870 6804
rect 14018 6748 14028 6804
rect 14084 6748 16268 6804
rect 16324 6748 16334 6804
rect 0 6720 112 6748
rect 1138 6636 1148 6692
rect 1204 6636 6972 6692
rect 7028 6636 7038 6692
rect 7298 6636 7308 6692
rect 7364 6636 9884 6692
rect 9940 6636 9950 6692
rect 10108 6580 10164 6748
rect 18620 6692 18676 6860
rect 18834 6748 18844 6804
rect 18900 6748 20188 6804
rect 20244 6748 20254 6804
rect 20748 6748 30380 6804
rect 30436 6748 30446 6804
rect 30594 6748 30604 6804
rect 30660 6748 31164 6804
rect 31220 6748 31230 6804
rect 31826 6748 31836 6804
rect 31892 6748 33292 6804
rect 33348 6748 33358 6804
rect 20748 6692 20804 6748
rect 33628 6692 33684 6860
rect 44940 6804 44996 6860
rect 57344 6804 57456 6832
rect 33954 6748 33964 6804
rect 34020 6748 37100 6804
rect 37156 6748 37166 6804
rect 38780 6748 44996 6804
rect 45378 6748 45388 6804
rect 45444 6748 47628 6804
rect 47684 6748 47694 6804
rect 48748 6748 52108 6804
rect 52164 6748 52174 6804
rect 56130 6748 56140 6804
rect 56196 6748 57456 6804
rect 38780 6692 38836 6748
rect 48748 6692 48804 6748
rect 57344 6720 57456 6748
rect 10322 6636 10332 6692
rect 10388 6636 18676 6692
rect 20738 6636 20748 6692
rect 20804 6636 20814 6692
rect 23986 6636 23996 6692
rect 24052 6636 33684 6692
rect 34962 6636 34972 6692
rect 35028 6636 38836 6692
rect 39890 6636 39900 6692
rect 39956 6636 48804 6692
rect 50372 6636 54124 6692
rect 54180 6636 54190 6692
rect 50372 6580 50428 6636
rect 7522 6524 7532 6580
rect 7588 6524 9884 6580
rect 9940 6524 9950 6580
rect 10108 6524 17052 6580
rect 17108 6524 17118 6580
rect 17826 6524 17836 6580
rect 17892 6524 26796 6580
rect 26852 6524 26862 6580
rect 27794 6524 27804 6580
rect 27860 6524 30716 6580
rect 30772 6524 30782 6580
rect 32274 6524 32284 6580
rect 32340 6524 40012 6580
rect 40068 6524 40078 6580
rect 40226 6524 40236 6580
rect 40292 6524 42140 6580
rect 42196 6524 42206 6580
rect 42354 6524 42364 6580
rect 42420 6524 45948 6580
rect 46004 6524 46014 6580
rect 46162 6524 46172 6580
rect 46228 6524 50428 6580
rect 802 6412 812 6468
rect 868 6412 9268 6468
rect 9426 6412 9436 6468
rect 9492 6412 21868 6468
rect 21924 6412 21934 6468
rect 22092 6412 24276 6468
rect 25218 6412 25228 6468
rect 25284 6412 37996 6468
rect 38052 6412 38062 6468
rect 38210 6412 38220 6468
rect 38276 6412 45388 6468
rect 45444 6412 45454 6468
rect 51650 6412 51660 6468
rect 51716 6412 54124 6468
rect 54180 6412 54190 6468
rect 0 6356 112 6384
rect 9212 6356 9268 6412
rect 22092 6356 22148 6412
rect 0 6300 1372 6356
rect 1428 6300 1438 6356
rect 9212 6300 10444 6356
rect 10500 6300 10510 6356
rect 10658 6300 10668 6356
rect 10724 6300 12740 6356
rect 15586 6300 15596 6356
rect 15652 6300 18396 6356
rect 18452 6300 18462 6356
rect 18610 6300 18620 6356
rect 18676 6300 21364 6356
rect 21746 6300 21756 6356
rect 21812 6300 22148 6356
rect 24220 6356 24276 6412
rect 57344 6356 57456 6384
rect 24220 6300 27132 6356
rect 27188 6300 27198 6356
rect 28364 6300 30268 6356
rect 30324 6300 30334 6356
rect 32722 6300 32732 6356
rect 32788 6300 40460 6356
rect 40516 6300 40526 6356
rect 55122 6300 55132 6356
rect 55188 6300 57456 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 8418 6188 8428 6244
rect 8484 6188 11452 6244
rect 11508 6188 11518 6244
rect 12684 6132 12740 6300
rect 21308 6244 21364 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 28364 6244 28420 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 57344 6272 57456 6300
rect 13458 6188 13468 6244
rect 13524 6188 20972 6244
rect 21028 6188 21038 6244
rect 21308 6188 23660 6244
rect 23716 6188 23726 6244
rect 24210 6188 24220 6244
rect 24276 6188 28420 6244
rect 28690 6188 28700 6244
rect 28756 6188 40684 6244
rect 40740 6188 40750 6244
rect 47170 6188 47180 6244
rect 47236 6188 52444 6244
rect 52500 6188 52510 6244
rect 1586 6076 1596 6132
rect 1652 6076 11788 6132
rect 11844 6076 11854 6132
rect 12684 6076 13692 6132
rect 13748 6076 13758 6132
rect 15138 6076 15148 6132
rect 15204 6076 15316 6132
rect 15474 6076 15484 6132
rect 15540 6076 16380 6132
rect 16436 6076 16446 6132
rect 16594 6076 16604 6132
rect 16660 6076 26908 6132
rect 26964 6076 26974 6132
rect 27132 6076 28812 6132
rect 28868 6076 28878 6132
rect 29026 6076 29036 6132
rect 29092 6076 30380 6132
rect 30436 6076 30446 6132
rect 30594 6076 30604 6132
rect 30660 6076 35084 6132
rect 35140 6076 35150 6132
rect 35410 6076 35420 6132
rect 35476 6076 38332 6132
rect 38388 6076 38398 6132
rect 40114 6076 40124 6132
rect 40180 6076 47068 6132
rect 47124 6076 47134 6132
rect 48738 6076 48748 6132
rect 48804 6076 52556 6132
rect 52612 6076 52622 6132
rect 52994 6076 53004 6132
rect 53060 6076 53900 6132
rect 53956 6076 53966 6132
rect 15260 6020 15316 6076
rect 27132 6020 27188 6076
rect 8754 5964 8764 6020
rect 8820 5964 10332 6020
rect 10388 5964 10398 6020
rect 11330 5964 11340 6020
rect 11396 5964 15036 6020
rect 15092 5964 15102 6020
rect 15260 5964 16940 6020
rect 16996 5964 17006 6020
rect 18274 5964 18284 6020
rect 18340 5964 21868 6020
rect 21924 5964 21934 6020
rect 22082 5964 22092 6020
rect 22148 5964 25116 6020
rect 25172 5964 25182 6020
rect 25778 5964 25788 6020
rect 25844 5964 27188 6020
rect 27682 5964 27692 6020
rect 27748 5964 29540 6020
rect 29922 5964 29932 6020
rect 29988 5964 35308 6020
rect 35364 5964 35374 6020
rect 36978 5964 36988 6020
rect 37044 5964 38556 6020
rect 38612 5964 38622 6020
rect 39554 5964 39564 6020
rect 39620 5964 41804 6020
rect 41860 5964 41870 6020
rect 42130 5964 42140 6020
rect 42196 5964 50428 6020
rect 0 5908 112 5936
rect 0 5852 3276 5908
rect 3332 5852 3342 5908
rect 3714 5852 3724 5908
rect 3780 5852 11116 5908
rect 11172 5852 11182 5908
rect 12572 5852 22988 5908
rect 23044 5852 23054 5908
rect 24322 5852 24332 5908
rect 24388 5852 25228 5908
rect 25284 5852 25294 5908
rect 25666 5852 25676 5908
rect 25732 5852 28140 5908
rect 28196 5852 28206 5908
rect 28354 5852 28364 5908
rect 28420 5852 29260 5908
rect 29316 5852 29326 5908
rect 0 5824 112 5852
rect 12572 5796 12628 5852
rect 29484 5796 29540 5964
rect 50372 5908 50428 5964
rect 57344 5908 57456 5936
rect 29698 5852 29708 5908
rect 29764 5852 30380 5908
rect 30436 5852 30446 5908
rect 30604 5852 35532 5908
rect 35588 5852 35598 5908
rect 35746 5852 35756 5908
rect 35812 5852 39788 5908
rect 39844 5852 39854 5908
rect 41122 5852 41132 5908
rect 41188 5852 48860 5908
rect 48916 5852 48926 5908
rect 50372 5852 53844 5908
rect 54562 5852 54572 5908
rect 54628 5852 57456 5908
rect 30604 5796 30660 5852
rect 53788 5796 53844 5852
rect 57344 5824 57456 5852
rect 1362 5740 1372 5796
rect 1428 5740 8428 5796
rect 8484 5740 8494 5796
rect 10210 5740 10220 5796
rect 10276 5740 12628 5796
rect 14130 5740 14140 5796
rect 14196 5740 29148 5796
rect 29204 5740 29214 5796
rect 29484 5740 30660 5796
rect 31714 5740 31724 5796
rect 31780 5740 35084 5796
rect 35140 5740 35150 5796
rect 35298 5740 35308 5796
rect 35364 5740 53564 5796
rect 53620 5740 53630 5796
rect 53788 5740 55132 5796
rect 55188 5740 55198 5796
rect 3266 5628 3276 5684
rect 3332 5628 3724 5684
rect 3780 5628 3790 5684
rect 3938 5628 3948 5684
rect 4004 5628 10108 5684
rect 10164 5628 10174 5684
rect 10322 5628 10332 5684
rect 10388 5628 15260 5684
rect 15316 5628 15326 5684
rect 15474 5628 15484 5684
rect 15540 5628 16156 5684
rect 16212 5628 16222 5684
rect 16370 5628 16380 5684
rect 16436 5628 19180 5684
rect 19236 5628 19246 5684
rect 20972 5628 27580 5684
rect 27636 5628 27646 5684
rect 29026 5628 29036 5684
rect 29092 5628 40236 5684
rect 40292 5628 40302 5684
rect 43820 5628 45612 5684
rect 45668 5628 45678 5684
rect 20972 5572 21028 5628
rect 6514 5516 6524 5572
rect 6580 5516 21028 5572
rect 21186 5516 21196 5572
rect 21252 5516 24332 5572
rect 24388 5516 24398 5572
rect 24882 5516 24892 5572
rect 24948 5516 32732 5572
rect 32788 5516 32798 5572
rect 33618 5516 33628 5572
rect 33684 5516 35756 5572
rect 35812 5516 35822 5572
rect 37090 5516 37100 5572
rect 37156 5516 40796 5572
rect 40852 5516 40862 5572
rect 41458 5516 41468 5572
rect 41524 5516 43596 5572
rect 43652 5516 43662 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 43820 5460 43876 5628
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 57344 5460 57456 5488
rect 0 5404 1596 5460
rect 1652 5404 1662 5460
rect 8866 5404 8876 5460
rect 8932 5404 11900 5460
rect 11956 5404 11966 5460
rect 13122 5404 13132 5460
rect 13188 5404 24220 5460
rect 24276 5404 24286 5460
rect 25228 5404 38444 5460
rect 38500 5404 38510 5460
rect 41356 5404 43876 5460
rect 56130 5404 56140 5460
rect 56196 5404 57456 5460
rect 0 5376 112 5404
rect 25228 5348 25284 5404
rect 3332 5292 15932 5348
rect 15988 5292 15998 5348
rect 18386 5292 18396 5348
rect 18452 5292 21644 5348
rect 21700 5292 21710 5348
rect 21858 5292 21868 5348
rect 21924 5292 21980 5348
rect 22036 5292 22046 5348
rect 22194 5292 22204 5348
rect 22260 5292 25284 5348
rect 26852 5292 34860 5348
rect 34916 5292 34926 5348
rect 35074 5292 35084 5348
rect 35140 5292 35588 5348
rect 36978 5292 36988 5348
rect 37044 5292 39340 5348
rect 39396 5292 39406 5348
rect 3332 5236 3388 5292
rect 26852 5236 26908 5292
rect 35532 5236 35588 5292
rect 41356 5236 41412 5404
rect 57344 5376 57456 5404
rect 42028 5292 52108 5348
rect 52164 5292 52174 5348
rect 42028 5236 42084 5292
rect 2594 5180 2604 5236
rect 2660 5180 3388 5236
rect 4498 5180 4508 5236
rect 4564 5180 9772 5236
rect 9828 5180 9838 5236
rect 9986 5180 9996 5236
rect 10052 5180 11956 5236
rect 12562 5180 12572 5236
rect 12628 5180 15484 5236
rect 15540 5180 15550 5236
rect 15698 5180 15708 5236
rect 15764 5180 18732 5236
rect 18788 5180 18798 5236
rect 21186 5180 21196 5236
rect 21252 5180 25788 5236
rect 25844 5180 25854 5236
rect 26562 5180 26572 5236
rect 26628 5180 26908 5236
rect 30258 5180 30268 5236
rect 30324 5180 35308 5236
rect 35364 5180 35374 5236
rect 35532 5180 41412 5236
rect 41468 5180 42084 5236
rect 42578 5180 42588 5236
rect 42644 5180 44828 5236
rect 44884 5180 44894 5236
rect 48626 5180 48636 5236
rect 48692 5180 51996 5236
rect 52052 5180 52062 5236
rect 52882 5180 52892 5236
rect 52948 5180 55356 5236
rect 55412 5180 55422 5236
rect 11900 5124 11956 5180
rect 1474 5068 1484 5124
rect 1540 5068 5068 5124
rect 5124 5068 5134 5124
rect 5404 5068 11844 5124
rect 11900 5068 12684 5124
rect 12740 5068 12750 5124
rect 13458 5068 13468 5124
rect 13524 5068 16884 5124
rect 18274 5068 18284 5124
rect 18340 5068 18452 5124
rect 18610 5068 18620 5124
rect 18676 5068 28532 5124
rect 28690 5068 28700 5124
rect 28756 5068 31612 5124
rect 31668 5068 31678 5124
rect 31836 5068 41244 5124
rect 41300 5068 41310 5124
rect 0 5012 112 5040
rect 5404 5012 5460 5068
rect 0 4956 5460 5012
rect 11788 5012 11844 5068
rect 16828 5012 16884 5068
rect 18396 5012 18452 5068
rect 28476 5012 28532 5068
rect 31836 5012 31892 5068
rect 41468 5012 41524 5180
rect 41682 5068 41692 5124
rect 41748 5068 45052 5124
rect 45108 5068 45118 5124
rect 47058 5068 47068 5124
rect 47124 5068 53340 5124
rect 53396 5068 53406 5124
rect 54898 5068 54908 5124
rect 54964 5068 55468 5124
rect 55412 5012 55468 5068
rect 57344 5012 57456 5040
rect 11788 4956 14924 5012
rect 14980 4956 14990 5012
rect 15082 4956 15092 5012
rect 15148 4956 15484 5012
rect 15540 4956 15550 5012
rect 16828 4956 18060 5012
rect 18116 4956 18126 5012
rect 18396 4956 25340 5012
rect 25396 4956 25406 5012
rect 25554 4956 25564 5012
rect 25620 4956 28420 5012
rect 28476 4956 31892 5012
rect 31948 4956 33628 5012
rect 33684 4956 33694 5012
rect 35298 4956 35308 5012
rect 35364 4956 40348 5012
rect 40404 4956 40414 5012
rect 40684 4956 41524 5012
rect 43362 4956 43372 5012
rect 43428 4956 44940 5012
rect 44996 4956 45006 5012
rect 55412 4956 57456 5012
rect 0 4928 112 4956
rect 28364 4900 28420 4956
rect 31948 4900 32004 4956
rect 40684 4900 40740 4956
rect 57344 4928 57456 4956
rect 3042 4844 3052 4900
rect 3108 4844 5404 4900
rect 5460 4844 5470 4900
rect 8418 4844 8428 4900
rect 8484 4844 13468 4900
rect 13524 4844 13534 4900
rect 13682 4844 13692 4900
rect 13748 4844 27916 4900
rect 27972 4844 27982 4900
rect 28364 4844 30156 4900
rect 30212 4844 30222 4900
rect 31042 4844 31052 4900
rect 31108 4844 32004 4900
rect 32834 4844 32844 4900
rect 32900 4844 40740 4900
rect 40796 4844 54460 4900
rect 54516 4844 54526 4900
rect 40796 4788 40852 4844
rect 4162 4732 4172 4788
rect 4228 4732 15652 4788
rect 15922 4732 15932 4788
rect 15988 4732 18956 4788
rect 19012 4732 19022 4788
rect 19170 4732 19180 4788
rect 19236 4732 23660 4788
rect 23716 4732 23726 4788
rect 24322 4732 24332 4788
rect 24388 4732 24892 4788
rect 24948 4732 24958 4788
rect 25106 4732 25116 4788
rect 25172 4732 27804 4788
rect 27860 4732 27870 4788
rect 28018 4732 28028 4788
rect 28084 4732 29484 4788
rect 29540 4732 29550 4788
rect 30492 4732 37156 4788
rect 37314 4732 37324 4788
rect 37380 4732 40852 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 4274 4620 4284 4676
rect 4340 4620 6748 4676
rect 6804 4620 6814 4676
rect 8306 4620 8316 4676
rect 8372 4620 13244 4676
rect 13300 4620 13310 4676
rect 13682 4620 13692 4676
rect 13748 4620 15372 4676
rect 15428 4620 15438 4676
rect 0 4564 112 4592
rect 15596 4564 15652 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 15810 4620 15820 4676
rect 15876 4620 21756 4676
rect 21812 4620 21822 4676
rect 24210 4620 24220 4676
rect 24276 4620 30268 4676
rect 30324 4620 30334 4676
rect 0 4508 1372 4564
rect 1428 4508 1438 4564
rect 9986 4508 9996 4564
rect 10052 4508 13468 4564
rect 13524 4508 13534 4564
rect 15596 4508 18396 4564
rect 18452 4508 18462 4564
rect 21522 4508 21532 4564
rect 21588 4508 28700 4564
rect 28756 4508 28766 4564
rect 0 4480 112 4508
rect 30492 4452 30548 4732
rect 37100 4676 37156 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 31602 4620 31612 4676
rect 31668 4620 35308 4676
rect 35364 4620 35374 4676
rect 35522 4620 35532 4676
rect 35588 4620 37044 4676
rect 37100 4620 39060 4676
rect 40674 4620 40684 4676
rect 40740 4620 42588 4676
rect 42644 4620 42654 4676
rect 45490 4620 45500 4676
rect 45556 4620 50428 4676
rect 36988 4564 37044 4620
rect 32274 4508 32284 4564
rect 32340 4508 36764 4564
rect 36820 4508 36830 4564
rect 36988 4508 38668 4564
rect 5730 4396 5740 4452
rect 5796 4396 9772 4452
rect 9828 4396 9838 4452
rect 14466 4396 14476 4452
rect 14532 4396 18844 4452
rect 18900 4396 18910 4452
rect 19292 4396 23548 4452
rect 23604 4396 23614 4452
rect 23762 4396 23772 4452
rect 23828 4396 25116 4452
rect 25172 4396 25182 4452
rect 27234 4396 27244 4452
rect 27300 4396 30548 4452
rect 30706 4396 30716 4452
rect 30772 4396 33852 4452
rect 33908 4396 33918 4452
rect 34738 4396 34748 4452
rect 34804 4396 36988 4452
rect 37044 4396 37054 4452
rect 38612 4396 38668 4508
rect 39004 4452 39060 4620
rect 50372 4564 50428 4620
rect 57344 4564 57456 4592
rect 40338 4508 40348 4564
rect 40404 4508 48412 4564
rect 48468 4508 48478 4564
rect 50372 4508 52668 4564
rect 52724 4508 52734 4564
rect 54562 4508 54572 4564
rect 54628 4508 57456 4564
rect 57344 4480 57456 4508
rect 38724 4396 38734 4452
rect 39004 4396 42196 4452
rect 42354 4396 42364 4452
rect 42420 4396 52332 4452
rect 52388 4396 52398 4452
rect 19292 4340 19348 4396
rect 42140 4340 42196 4396
rect 1250 4284 1260 4340
rect 1316 4284 5180 4340
rect 5236 4284 5246 4340
rect 13794 4284 13804 4340
rect 13860 4284 19348 4340
rect 19618 4284 19628 4340
rect 19684 4284 21756 4340
rect 21812 4284 21822 4340
rect 22082 4284 22092 4340
rect 22148 4284 41132 4340
rect 41188 4284 41198 4340
rect 42140 4284 45276 4340
rect 45332 4284 45342 4340
rect 1922 4172 1932 4228
rect 1988 4172 12012 4228
rect 12068 4172 12078 4228
rect 12898 4172 12908 4228
rect 12964 4172 15372 4228
rect 15428 4172 15438 4228
rect 15586 4172 15596 4228
rect 15652 4172 18172 4228
rect 18228 4172 18238 4228
rect 18610 4172 18620 4228
rect 18676 4172 26572 4228
rect 26628 4172 26638 4228
rect 26786 4172 26796 4228
rect 26852 4172 40124 4228
rect 40180 4172 40190 4228
rect 42242 4172 42252 4228
rect 42308 4172 53564 4228
rect 53620 4172 53630 4228
rect 0 4116 112 4144
rect 57344 4116 57456 4144
rect 0 4060 3276 4116
rect 3332 4060 3342 4116
rect 6962 4060 6972 4116
rect 7028 4060 23660 4116
rect 23716 4060 23726 4116
rect 23874 4060 23884 4116
rect 23940 4060 25788 4116
rect 25844 4060 25854 4116
rect 26002 4060 26012 4116
rect 26068 4060 27580 4116
rect 27636 4060 27646 4116
rect 27794 4060 27804 4116
rect 27860 4060 31836 4116
rect 31892 4060 31902 4116
rect 33282 4060 33292 4116
rect 33348 4060 34412 4116
rect 34468 4060 34478 4116
rect 35074 4060 35084 4116
rect 35140 4060 47180 4116
rect 47236 4060 47246 4116
rect 52322 4060 52332 4116
rect 52388 4060 54796 4116
rect 54852 4060 54862 4116
rect 56130 4060 56140 4116
rect 56196 4060 57456 4116
rect 0 4032 112 4060
rect 57344 4032 57456 4060
rect 8082 3948 8092 4004
rect 8148 3948 24220 4004
rect 24276 3948 24286 4004
rect 25554 3948 25564 4004
rect 25620 3948 37100 4004
rect 37156 3948 37166 4004
rect 37324 3948 44324 4004
rect 45714 3948 45724 4004
rect 45780 3948 53676 4004
rect 53732 3948 53742 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 37324 3892 37380 3948
rect 9212 3836 15708 3892
rect 15764 3836 15774 3892
rect 15932 3836 24220 3892
rect 24276 3836 24286 3892
rect 24892 3836 29148 3892
rect 29204 3836 29214 3892
rect 29810 3836 29820 3892
rect 29876 3836 33292 3892
rect 33348 3836 33358 3892
rect 33506 3836 33516 3892
rect 33572 3836 37380 3892
rect 38658 3836 38668 3892
rect 38724 3836 40068 3892
rect 40226 3836 40236 3892
rect 40292 3836 42252 3892
rect 42308 3836 42318 3892
rect 9212 3780 9268 3836
rect 15932 3780 15988 3836
rect 24892 3780 24948 3836
rect 40012 3780 40068 3836
rect 44268 3780 44324 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 50530 3836 50540 3892
rect 50596 3836 53452 3892
rect 53508 3836 53518 3892
rect 1586 3724 1596 3780
rect 1652 3724 9268 3780
rect 9324 3724 15988 3780
rect 16146 3724 16156 3780
rect 16212 3724 21532 3780
rect 21588 3724 21598 3780
rect 21746 3724 21756 3780
rect 21812 3724 23548 3780
rect 23650 3724 23660 3780
rect 23716 3724 23884 3780
rect 23940 3724 23950 3780
rect 24210 3724 24220 3780
rect 24276 3724 24948 3780
rect 25106 3724 25116 3780
rect 25172 3724 34748 3780
rect 34804 3724 34814 3780
rect 35298 3724 35308 3780
rect 35364 3724 39788 3780
rect 39844 3724 39854 3780
rect 40012 3724 43372 3780
rect 43428 3724 43438 3780
rect 43586 3724 43596 3780
rect 43652 3724 44044 3780
rect 44100 3724 44110 3780
rect 44268 3724 52220 3780
rect 52276 3724 52286 3780
rect 52444 3724 55132 3780
rect 55188 3724 55198 3780
rect 0 3668 112 3696
rect 0 3612 7980 3668
rect 8036 3612 8046 3668
rect 0 3584 112 3612
rect 9324 3556 9380 3724
rect 23492 3668 23548 3724
rect 52444 3668 52500 3724
rect 57344 3668 57456 3696
rect 9650 3612 9660 3668
rect 9716 3612 10836 3668
rect 10994 3612 11004 3668
rect 11060 3612 14140 3668
rect 14196 3612 14206 3668
rect 15092 3612 15484 3668
rect 15540 3612 15550 3668
rect 16482 3612 16492 3668
rect 16548 3612 17948 3668
rect 18004 3612 18014 3668
rect 18834 3612 18844 3668
rect 18900 3612 22764 3668
rect 22820 3612 22830 3668
rect 23492 3612 23996 3668
rect 24052 3612 24062 3668
rect 24210 3612 24220 3668
rect 24276 3612 25676 3668
rect 25732 3612 25742 3668
rect 25890 3612 25900 3668
rect 25956 3612 30100 3668
rect 30258 3612 30268 3668
rect 30324 3612 38556 3668
rect 38612 3612 38622 3668
rect 38882 3612 38892 3668
rect 38948 3612 52500 3668
rect 54786 3612 54796 3668
rect 54852 3612 57456 3668
rect 10780 3556 10836 3612
rect 15092 3556 15148 3612
rect 30044 3556 30100 3612
rect 57344 3584 57456 3612
rect 2706 3500 2716 3556
rect 2772 3500 9380 3556
rect 9874 3500 9884 3556
rect 9940 3500 10444 3556
rect 10500 3500 10510 3556
rect 10780 3500 15148 3556
rect 15698 3500 15708 3556
rect 15764 3500 18060 3556
rect 18116 3500 18126 3556
rect 18274 3500 18284 3556
rect 18340 3500 19012 3556
rect 19170 3500 19180 3556
rect 19236 3500 27020 3556
rect 27076 3500 27086 3556
rect 27570 3500 27580 3556
rect 27636 3500 29820 3556
rect 29876 3500 29886 3556
rect 30044 3500 33404 3556
rect 33460 3500 33470 3556
rect 34178 3500 34188 3556
rect 34244 3500 36540 3556
rect 36596 3500 36606 3556
rect 37090 3500 37100 3556
rect 37156 3500 42364 3556
rect 42420 3500 42430 3556
rect 44034 3500 44044 3556
rect 44100 3500 50428 3556
rect 50484 3500 50494 3556
rect 18956 3444 19012 3500
rect 6402 3388 6412 3444
rect 6468 3388 8428 3444
rect 8530 3388 8540 3444
rect 8596 3388 10164 3444
rect 11778 3388 11788 3444
rect 11844 3388 15988 3444
rect 17938 3388 17948 3444
rect 18004 3388 18900 3444
rect 18956 3388 26964 3444
rect 28690 3388 28700 3444
rect 28756 3388 36820 3444
rect 38658 3388 38668 3444
rect 38724 3388 44380 3444
rect 44436 3388 44446 3444
rect 48402 3388 48412 3444
rect 48468 3388 53228 3444
rect 53284 3388 53294 3444
rect 53554 3388 53564 3444
rect 53620 3388 56812 3444
rect 56868 3388 56878 3444
rect 8372 3332 8428 3388
rect 10108 3332 10164 3388
rect 15932 3332 15988 3388
rect 18844 3332 18900 3388
rect 26908 3332 26964 3388
rect 36764 3332 36820 3388
rect 2818 3276 2828 3332
rect 2884 3276 3388 3332
rect 3490 3276 3500 3332
rect 3556 3276 4564 3332
rect 8372 3276 8764 3332
rect 8820 3276 8830 3332
rect 10098 3276 10108 3332
rect 10164 3276 10174 3332
rect 10332 3276 15036 3332
rect 15092 3276 15102 3332
rect 15932 3276 18620 3332
rect 18676 3276 18686 3332
rect 18844 3276 19124 3332
rect 20066 3276 20076 3332
rect 20132 3276 22596 3332
rect 22754 3276 22764 3332
rect 22820 3276 25564 3332
rect 25620 3276 25630 3332
rect 26908 3276 28924 3332
rect 28980 3276 28990 3332
rect 29138 3276 29148 3332
rect 29204 3276 32396 3332
rect 32452 3276 32462 3332
rect 32722 3276 32732 3332
rect 32788 3276 36428 3332
rect 36484 3276 36494 3332
rect 36764 3276 37660 3332
rect 37716 3276 37726 3332
rect 38658 3276 38668 3332
rect 38724 3276 41468 3332
rect 41524 3276 41534 3332
rect 42242 3276 42252 3332
rect 42308 3276 47068 3332
rect 47124 3276 47134 3332
rect 0 3220 112 3248
rect 3332 3220 3388 3276
rect 4508 3220 4564 3276
rect 0 3164 1596 3220
rect 1652 3164 1662 3220
rect 3332 3164 3612 3220
rect 3668 3164 3678 3220
rect 4508 3164 9996 3220
rect 10052 3164 10062 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 10332 3108 10388 3276
rect 19068 3220 19124 3276
rect 22540 3220 22596 3276
rect 57344 3220 57456 3248
rect 13234 3164 13244 3220
rect 13300 3164 18844 3220
rect 18900 3164 18910 3220
rect 19068 3164 21420 3220
rect 21476 3164 21486 3220
rect 21634 3164 21644 3220
rect 21700 3164 22204 3220
rect 22260 3164 22270 3220
rect 22540 3164 23660 3220
rect 23716 3164 23726 3220
rect 24322 3164 24332 3220
rect 24388 3164 29036 3220
rect 29092 3164 29102 3220
rect 29260 3164 30716 3220
rect 30772 3164 30782 3220
rect 33730 3164 33740 3220
rect 33796 3164 35308 3220
rect 35364 3164 35374 3220
rect 36428 3164 37100 3220
rect 37156 3164 37166 3220
rect 37314 3164 37324 3220
rect 37380 3164 40236 3220
rect 40292 3164 40302 3220
rect 48066 3164 48076 3220
rect 48132 3164 53564 3220
rect 53620 3164 53630 3220
rect 54562 3164 54572 3220
rect 54628 3164 57456 3220
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 29260 3108 29316 3164
rect 36428 3108 36484 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 57344 3136 57456 3164
rect 924 3052 2604 3108
rect 2660 3052 2670 3108
rect 5282 3052 5292 3108
rect 5348 3052 10388 3108
rect 10546 3052 10556 3108
rect 10612 3052 13692 3108
rect 13748 3052 13758 3108
rect 13906 3052 13916 3108
rect 13972 3052 19012 3108
rect 0 2772 112 2800
rect 924 2772 980 3052
rect 18956 2996 19012 3052
rect 19180 3052 21756 3108
rect 21812 3052 21822 3108
rect 24434 3052 24444 3108
rect 24500 3052 29316 3108
rect 29474 3052 29484 3108
rect 29540 3052 34188 3108
rect 34244 3052 34254 3108
rect 34402 3052 34412 3108
rect 34468 3052 36484 3108
rect 36642 3052 36652 3108
rect 36708 3052 43204 3108
rect 46610 3052 46620 3108
rect 46676 3052 55132 3108
rect 55188 3052 55198 3108
rect 19180 2996 19236 3052
rect 43148 2996 43204 3052
rect 0 2716 980 2772
rect 1036 2940 18508 2996
rect 18564 2940 18574 2996
rect 18956 2940 19236 2996
rect 21410 2940 21420 2996
rect 21476 2940 29036 2996
rect 29092 2940 29102 2996
rect 29362 2940 29372 2996
rect 29428 2940 38220 2996
rect 38276 2940 38286 2996
rect 43148 2940 47292 2996
rect 47348 2940 47358 2996
rect 0 2688 112 2716
rect 0 2324 112 2352
rect 1036 2324 1092 2940
rect 2258 2828 2268 2884
rect 2324 2828 8316 2884
rect 8372 2828 8382 2884
rect 11442 2828 11452 2884
rect 11508 2828 18284 2884
rect 18340 2828 18350 2884
rect 20178 2828 20188 2884
rect 20244 2828 21868 2884
rect 21924 2828 21934 2884
rect 22082 2828 22092 2884
rect 22148 2828 24276 2884
rect 24658 2828 24668 2884
rect 24724 2828 30156 2884
rect 30212 2828 30222 2884
rect 32834 2828 32844 2884
rect 32900 2828 35420 2884
rect 35476 2828 35486 2884
rect 36978 2828 36988 2884
rect 37044 2828 42532 2884
rect 24220 2772 24276 2828
rect 42476 2772 42532 2828
rect 57344 2772 57456 2800
rect 3602 2716 3612 2772
rect 3668 2716 8540 2772
rect 8596 2716 8606 2772
rect 12114 2716 12124 2772
rect 12180 2716 23996 2772
rect 24052 2716 24062 2772
rect 24220 2716 26012 2772
rect 26068 2716 26078 2772
rect 34850 2716 34860 2772
rect 34916 2716 37884 2772
rect 37940 2716 37950 2772
rect 38098 2716 38108 2772
rect 38164 2716 38668 2772
rect 38724 2716 38734 2772
rect 42476 2716 46284 2772
rect 46340 2716 46350 2772
rect 49410 2716 49420 2772
rect 49476 2716 52108 2772
rect 52164 2716 52174 2772
rect 56130 2716 56140 2772
rect 56196 2716 57456 2772
rect 57344 2688 57456 2716
rect 10098 2604 10108 2660
rect 10164 2604 21532 2660
rect 21588 2604 21598 2660
rect 21746 2604 21756 2660
rect 21812 2604 24668 2660
rect 24724 2604 24734 2660
rect 24994 2604 25004 2660
rect 25060 2604 28588 2660
rect 28644 2604 28654 2660
rect 29474 2604 29484 2660
rect 29540 2604 34972 2660
rect 35028 2604 35038 2660
rect 35186 2604 35196 2660
rect 35252 2604 38892 2660
rect 38948 2604 38958 2660
rect 41804 2604 48860 2660
rect 48916 2604 48926 2660
rect 52770 2604 52780 2660
rect 52836 2604 56476 2660
rect 56532 2604 56542 2660
rect 41804 2548 41860 2604
rect 5058 2492 5068 2548
rect 5124 2492 23548 2548
rect 23604 2492 23614 2548
rect 24332 2492 25900 2548
rect 25956 2492 25966 2548
rect 26338 2492 26348 2548
rect 26404 2492 28700 2548
rect 28756 2492 28766 2548
rect 30706 2492 30716 2548
rect 30772 2492 37548 2548
rect 37604 2492 37614 2548
rect 38546 2492 38556 2548
rect 38612 2492 41860 2548
rect 42018 2492 42028 2548
rect 42084 2492 47628 2548
rect 47684 2492 47694 2548
rect 7074 2380 7084 2436
rect 7140 2380 13132 2436
rect 13188 2380 13198 2436
rect 13458 2380 13468 2436
rect 13524 2380 16044 2436
rect 16100 2380 16110 2436
rect 16258 2380 16268 2436
rect 16324 2380 23884 2436
rect 23940 2380 23950 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24332 2324 24388 2492
rect 25106 2380 25116 2436
rect 25172 2380 26796 2436
rect 26852 2380 26862 2436
rect 27122 2380 27132 2436
rect 27188 2380 41692 2436
rect 41748 2380 41758 2436
rect 44828 2380 54124 2436
rect 54180 2380 54190 2436
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 0 2268 1092 2324
rect 11106 2268 11116 2324
rect 11172 2268 14812 2324
rect 14868 2268 14878 2324
rect 15474 2268 15484 2324
rect 15540 2268 18732 2324
rect 18788 2268 18798 2324
rect 18956 2268 22204 2324
rect 22260 2268 22270 2324
rect 23650 2268 23660 2324
rect 23716 2268 24388 2324
rect 24882 2268 24892 2324
rect 24948 2268 24958 2324
rect 28466 2268 28476 2324
rect 28532 2268 33516 2324
rect 33572 2268 33582 2324
rect 33730 2268 33740 2324
rect 33796 2268 38108 2324
rect 38164 2268 38174 2324
rect 0 2240 112 2268
rect 2482 2156 2492 2212
rect 2548 2156 6300 2212
rect 6356 2156 6366 2212
rect 11778 2156 11788 2212
rect 11844 2156 14700 2212
rect 14756 2156 14766 2212
rect 16034 2156 16044 2212
rect 16100 2156 18284 2212
rect 18340 2156 18350 2212
rect 18956 2100 19012 2268
rect 24892 2212 24948 2268
rect 44828 2212 44884 2380
rect 57344 2324 57456 2352
rect 19170 2156 19180 2212
rect 19236 2156 24948 2212
rect 25330 2156 25340 2212
rect 25396 2156 34636 2212
rect 34692 2156 34702 2212
rect 38434 2156 38444 2212
rect 38500 2156 44884 2212
rect 44940 2268 54236 2324
rect 54292 2268 54302 2324
rect 54898 2268 54908 2324
rect 54964 2268 57456 2324
rect 44940 2100 44996 2268
rect 57344 2240 57456 2268
rect 5394 2044 5404 2100
rect 5460 2044 13468 2100
rect 13524 2044 13534 2100
rect 13682 2044 13692 2100
rect 13748 2044 16716 2100
rect 16772 2044 16782 2100
rect 17154 2044 17164 2100
rect 17220 2044 19012 2100
rect 21970 2044 21980 2100
rect 22036 2044 24780 2100
rect 24836 2044 24846 2100
rect 25106 2044 25116 2100
rect 25172 2044 44996 2100
rect 47618 2044 47628 2100
rect 47684 2044 52556 2100
rect 52612 2044 52622 2100
rect 1138 1932 1148 1988
rect 1204 1932 6300 1988
rect 6356 1932 6366 1988
rect 8876 1932 10556 1988
rect 10612 1932 10622 1988
rect 11218 1932 11228 1988
rect 11284 1932 25004 1988
rect 25060 1932 25070 1988
rect 26002 1932 26012 1988
rect 26068 1932 30548 1988
rect 30930 1932 30940 1988
rect 30996 1932 34076 1988
rect 34132 1932 34142 1988
rect 39330 1932 39340 1988
rect 39396 1932 45724 1988
rect 45780 1932 45790 1988
rect 0 1876 112 1904
rect 8876 1876 8932 1932
rect 30492 1876 30548 1932
rect 57344 1876 57456 1904
rect 0 1820 1036 1876
rect 1092 1820 1102 1876
rect 2930 1820 2940 1876
rect 2996 1820 8932 1876
rect 9426 1820 9436 1876
rect 9492 1820 14588 1876
rect 14644 1820 14654 1876
rect 14802 1820 14812 1876
rect 14868 1820 14878 1876
rect 15026 1820 15036 1876
rect 15092 1820 20748 1876
rect 20804 1820 20814 1876
rect 20972 1820 30268 1876
rect 30324 1820 30334 1876
rect 30492 1820 47404 1876
rect 47460 1820 47470 1876
rect 47618 1820 47628 1876
rect 47684 1820 52108 1876
rect 52164 1820 52174 1876
rect 53554 1820 53564 1876
rect 53620 1820 57456 1876
rect 0 1792 112 1820
rect 14812 1764 14868 1820
rect 20972 1764 21028 1820
rect 57344 1792 57456 1820
rect 914 1708 924 1764
rect 980 1708 2828 1764
rect 2884 1708 2894 1764
rect 4274 1708 4284 1764
rect 4340 1708 6692 1764
rect 12674 1708 12684 1764
rect 12740 1708 14588 1764
rect 14644 1708 14654 1764
rect 14812 1708 17164 1764
rect 17220 1708 17230 1764
rect 18386 1708 18396 1764
rect 18452 1708 21028 1764
rect 21868 1708 25228 1764
rect 25284 1708 25294 1764
rect 25890 1708 25900 1764
rect 25956 1708 30604 1764
rect 30660 1708 30670 1764
rect 30930 1708 30940 1764
rect 30996 1708 32620 1764
rect 32676 1708 32686 1764
rect 32834 1708 32844 1764
rect 32900 1708 38668 1764
rect 39442 1708 39452 1764
rect 39508 1708 42364 1764
rect 42420 1708 42430 1764
rect 43596 1708 44212 1764
rect 47058 1708 47068 1764
rect 47124 1708 51100 1764
rect 51156 1708 51166 1764
rect 6636 1652 6692 1708
rect 21868 1652 21924 1708
rect 38612 1652 38668 1708
rect 43596 1652 43652 1708
rect 6636 1596 7196 1652
rect 7252 1596 7262 1652
rect 8082 1596 8092 1652
rect 8148 1596 14700 1652
rect 14756 1596 14766 1652
rect 15026 1596 15036 1652
rect 15092 1596 21924 1652
rect 24770 1596 24780 1652
rect 24836 1596 29372 1652
rect 29428 1596 29438 1652
rect 30818 1596 30828 1652
rect 30884 1596 33964 1652
rect 34020 1596 34030 1652
rect 38612 1596 41580 1652
rect 41636 1596 41646 1652
rect 41794 1596 41804 1652
rect 41860 1596 43652 1652
rect 44156 1652 44212 1708
rect 44156 1596 46732 1652
rect 46788 1596 46798 1652
rect 49522 1596 49532 1652
rect 49588 1596 55132 1652
rect 55188 1596 55198 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 6738 1484 6748 1540
rect 6804 1484 12908 1540
rect 12964 1484 12974 1540
rect 13122 1484 13132 1540
rect 13188 1484 15708 1540
rect 15764 1484 15774 1540
rect 17378 1484 17388 1540
rect 17444 1484 20188 1540
rect 20244 1484 20254 1540
rect 20402 1484 20412 1540
rect 20468 1484 23660 1540
rect 23716 1484 23726 1540
rect 24322 1484 24332 1540
rect 24388 1484 25004 1540
rect 25060 1484 25070 1540
rect 25218 1484 25228 1540
rect 25284 1484 32732 1540
rect 32788 1484 32798 1540
rect 32946 1484 32956 1540
rect 33012 1484 33852 1540
rect 33908 1484 33918 1540
rect 34402 1484 34412 1540
rect 34468 1484 39452 1540
rect 39508 1484 39518 1540
rect 46498 1484 46508 1540
rect 46564 1484 52556 1540
rect 52612 1484 52622 1540
rect 0 1428 112 1456
rect 57344 1428 57456 1456
rect 0 1372 2548 1428
rect 3266 1372 3276 1428
rect 3332 1372 6748 1428
rect 6804 1372 6814 1428
rect 8530 1372 8540 1428
rect 8596 1372 15148 1428
rect 15204 1372 15214 1428
rect 15362 1372 15372 1428
rect 15428 1372 20076 1428
rect 20132 1372 20142 1428
rect 20290 1372 20300 1428
rect 20356 1372 25340 1428
rect 25396 1372 25406 1428
rect 25564 1372 26796 1428
rect 26852 1372 26862 1428
rect 27122 1372 27132 1428
rect 27188 1372 28476 1428
rect 28532 1372 28542 1428
rect 29026 1372 29036 1428
rect 29092 1372 36876 1428
rect 36932 1372 36942 1428
rect 37650 1372 37660 1428
rect 37716 1372 47068 1428
rect 47124 1372 47134 1428
rect 53554 1372 53564 1428
rect 53620 1372 57456 1428
rect 0 1344 112 1372
rect 2492 1204 2548 1372
rect 25564 1316 25620 1372
rect 57344 1344 57456 1372
rect 5506 1260 5516 1316
rect 5572 1260 7700 1316
rect 8306 1260 8316 1316
rect 8372 1260 21980 1316
rect 22036 1260 22046 1316
rect 22978 1260 22988 1316
rect 23044 1260 25620 1316
rect 26002 1260 26012 1316
rect 26068 1260 28924 1316
rect 28980 1260 28990 1316
rect 29138 1260 29148 1316
rect 29204 1260 31388 1316
rect 31444 1260 31454 1316
rect 31602 1260 31612 1316
rect 31668 1260 34524 1316
rect 34580 1260 34590 1316
rect 34748 1260 36092 1316
rect 36148 1260 36158 1316
rect 39442 1260 39452 1316
rect 39508 1260 46956 1316
rect 47012 1260 47022 1316
rect 48972 1260 51660 1316
rect 51716 1260 51726 1316
rect 7644 1204 7700 1260
rect 34748 1204 34804 1260
rect 2492 1148 7420 1204
rect 7476 1148 7486 1204
rect 7644 1148 11788 1204
rect 11844 1148 11854 1204
rect 15138 1148 15148 1204
rect 15204 1148 20636 1204
rect 20692 1148 20702 1204
rect 20850 1148 20860 1204
rect 20916 1148 25116 1204
rect 25172 1148 25182 1204
rect 26226 1148 26236 1204
rect 26292 1148 33628 1204
rect 33684 1148 33694 1204
rect 33842 1148 33852 1204
rect 33908 1148 34804 1204
rect 35298 1148 35308 1204
rect 35364 1148 41804 1204
rect 41860 1148 41870 1204
rect 42018 1148 42028 1204
rect 42084 1148 48412 1204
rect 48468 1148 48478 1204
rect 48972 1092 49028 1260
rect 4162 1036 4172 1092
rect 4228 1036 18396 1092
rect 18452 1036 18462 1092
rect 18620 1036 19516 1092
rect 19572 1036 19582 1092
rect 19730 1036 19740 1092
rect 19796 1036 25900 1092
rect 25956 1036 25966 1092
rect 26898 1036 26908 1092
rect 26964 1036 34412 1092
rect 34468 1036 34478 1092
rect 40226 1036 40236 1092
rect 40292 1036 49028 1092
rect 50372 1148 50988 1204
rect 51044 1148 51054 1204
rect 0 980 112 1008
rect 18620 980 18676 1036
rect 50372 980 50428 1148
rect 57344 980 57456 1008
rect 0 924 924 980
rect 980 924 990 980
rect 2594 924 2604 980
rect 2660 924 9212 980
rect 9268 924 9278 980
rect 12562 924 12572 980
rect 12628 924 14364 980
rect 14420 924 14430 980
rect 15138 924 15148 980
rect 15204 924 18676 980
rect 18834 924 18844 980
rect 18900 924 20860 980
rect 20916 924 20926 980
rect 22978 924 22988 980
rect 23044 924 24948 980
rect 25106 924 25116 980
rect 25172 924 36988 980
rect 37044 924 37054 980
rect 41570 924 41580 980
rect 41636 924 44828 980
rect 44884 924 44894 980
rect 48290 924 48300 980
rect 48356 924 50428 980
rect 51986 924 51996 980
rect 52052 924 57456 980
rect 0 896 112 924
rect 14578 812 14588 868
rect 14644 812 15484 868
rect 15540 812 15550 868
rect 18946 812 18956 868
rect 19012 812 22988 868
rect 23044 812 23054 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 24892 756 24948 924
rect 57344 896 57456 924
rect 25554 812 25564 868
rect 25620 812 43036 868
rect 43092 812 43102 868
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 8652 700 23324 756
rect 23380 700 23390 756
rect 24892 700 26908 756
rect 26964 700 26974 756
rect 27234 700 27244 756
rect 27300 700 35196 756
rect 35252 700 35262 756
rect 35634 700 35644 756
rect 35700 700 40684 756
rect 40740 700 40750 756
rect 40908 700 41412 756
rect 2034 588 2044 644
rect 2100 588 2660 644
rect 0 532 112 560
rect 2604 532 2660 588
rect 8652 532 8708 700
rect 9202 588 9212 644
rect 9268 588 16772 644
rect 16930 588 16940 644
rect 16996 588 26348 644
rect 26404 588 26414 644
rect 26572 588 30268 644
rect 30324 588 30334 644
rect 30482 588 30492 644
rect 30548 588 40628 644
rect 0 476 2380 532
rect 2436 476 2446 532
rect 2604 476 8708 532
rect 16716 532 16772 588
rect 16716 476 19068 532
rect 19124 476 19134 532
rect 21970 476 21980 532
rect 22036 476 26124 532
rect 26180 476 26190 532
rect 0 448 112 476
rect 26572 420 26628 588
rect 40572 532 40628 588
rect 40908 532 40964 700
rect 41356 644 41412 700
rect 44828 700 52332 756
rect 52388 700 52398 756
rect 44828 644 44884 700
rect 41356 588 44884 644
rect 47506 588 47516 644
rect 47572 588 51436 644
rect 51492 588 51502 644
rect 57344 532 57456 560
rect 26786 476 26796 532
rect 26852 476 39340 532
rect 39396 476 39406 532
rect 40572 476 40964 532
rect 41458 476 41468 532
rect 41524 476 49308 532
rect 49364 476 49374 532
rect 56802 476 56812 532
rect 56868 476 57456 532
rect 57344 448 57456 476
rect 4498 364 4508 420
rect 4564 364 5852 420
rect 5908 364 5918 420
rect 14466 364 14476 420
rect 14532 364 21980 420
rect 22036 364 22046 420
rect 22194 364 22204 420
rect 22260 364 26628 420
rect 26786 364 26796 420
rect 26852 364 28700 420
rect 28756 364 28766 420
rect 28914 364 28924 420
rect 28980 364 40460 420
rect 40516 364 40526 420
rect 40674 364 40684 420
rect 40740 364 49980 420
rect 50036 364 50046 420
rect 17826 252 17836 308
rect 17892 252 55580 308
rect 55636 252 55646 308
rect 19954 140 19964 196
rect 20020 140 28700 196
rect 28756 140 28766 196
rect 28914 140 28924 196
rect 28980 140 31612 196
rect 31668 140 31678 196
rect 33618 140 33628 196
rect 33684 140 52892 196
rect 52948 140 52958 196
rect 0 84 112 112
rect 57344 84 57456 112
rect 0 28 1148 84
rect 1204 28 1214 84
rect 22082 28 22092 84
rect 22148 28 33740 84
rect 33796 28 33806 84
rect 56466 28 56476 84
rect 56532 28 57456 84
rect 0 0 112 28
rect 57344 0 57456 28
<< via3 >>
rect 20524 14140 20580 14196
rect 38108 14140 38164 14196
rect 20972 14028 21028 14084
rect 28028 14028 28084 14084
rect 28252 14028 28308 14084
rect 30492 14028 30548 14084
rect 20524 13916 20580 13972
rect 23660 13804 23716 13860
rect 31948 13804 32004 13860
rect 32508 13804 32564 13860
rect 32732 13804 32788 13860
rect 17388 13692 17444 13748
rect 36988 13692 37044 13748
rect 32508 13580 32564 13636
rect 38444 13580 38500 13636
rect 38892 13580 38948 13636
rect 6300 13468 6356 13524
rect 20972 13468 21028 13524
rect 28140 13356 28196 13412
rect 38612 13356 38668 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 20972 13244 21028 13300
rect 33740 13244 33796 13300
rect 15820 13132 15876 13188
rect 16044 13132 16100 13188
rect 25676 13132 25732 13188
rect 33852 13132 33908 13188
rect 34076 13132 34132 13188
rect 45948 13132 46004 13188
rect 23548 13020 23604 13076
rect 25004 13020 25060 13076
rect 24220 12908 24276 12964
rect 14812 12796 14868 12852
rect 31276 12796 31332 12852
rect 33292 12796 33348 12852
rect 20972 12684 21028 12740
rect 32732 12684 32788 12740
rect 11788 12572 11844 12628
rect 25228 12572 25284 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 18284 12460 18340 12516
rect 18508 12460 18564 12516
rect 21756 12460 21812 12516
rect 24220 12460 24276 12516
rect 27692 12460 27748 12516
rect 14812 12348 14868 12404
rect 15820 12348 15876 12404
rect 39340 12348 39396 12404
rect 23548 12236 23604 12292
rect 32956 12236 33012 12292
rect 36988 12236 37044 12292
rect 17388 12124 17444 12180
rect 30492 12124 30548 12180
rect 37324 12124 37380 12180
rect 39228 12124 39284 12180
rect 16044 12012 16100 12068
rect 19964 12012 20020 12068
rect 35532 12012 35588 12068
rect 48860 12012 48916 12068
rect 14252 11900 14308 11956
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 14924 11900 14980 11956
rect 16268 11900 16324 11956
rect 20300 11900 20356 11956
rect 21868 11900 21924 11956
rect 28364 11900 28420 11956
rect 34972 11900 35028 11956
rect 38108 11900 38164 11956
rect 30492 11788 30548 11844
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 30716 11676 30772 11732
rect 17948 11564 18004 11620
rect 21756 11564 21812 11620
rect 21980 11564 22036 11620
rect 43596 11564 43652 11620
rect 6076 11228 6132 11284
rect 13692 11340 13748 11396
rect 13916 11340 13972 11396
rect 2604 11116 2660 11172
rect 23548 11228 23604 11284
rect 26012 11228 26068 11284
rect 43596 11228 43652 11284
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 17164 11116 17220 11172
rect 19628 11116 19684 11172
rect 31612 11116 31668 11172
rect 34076 11116 34132 11172
rect 21980 11004 22036 11060
rect 24220 11004 24276 11060
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 21308 10892 21364 10948
rect 23548 10892 23604 10948
rect 28252 10892 28308 10948
rect 47628 10780 47684 10836
rect 20076 10668 20132 10724
rect 26572 10668 26628 10724
rect 19628 10556 19684 10612
rect 25228 10556 25284 10612
rect 33628 10556 33684 10612
rect 2828 10444 2884 10500
rect 13916 10444 13972 10500
rect 14140 10444 14196 10500
rect 24220 10444 24276 10500
rect 30716 10444 30772 10500
rect 31500 10444 31556 10500
rect 33516 10444 33572 10500
rect 42028 10332 42084 10388
rect 15036 10220 15092 10276
rect 30268 10220 30324 10276
rect 31500 10220 31556 10276
rect 35196 10220 35252 10276
rect 35420 10220 35476 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 26852 9996 26908 10052
rect 31276 9996 31332 10052
rect 11452 9884 11508 9940
rect 14700 9884 14756 9940
rect 31612 9884 31668 9940
rect 10108 9772 10164 9828
rect 21196 9772 21252 9828
rect 21980 9772 22036 9828
rect 29372 9772 29428 9828
rect 35420 9660 35476 9716
rect 10108 9548 10164 9604
rect 11452 9548 11508 9604
rect 13804 9548 13860 9604
rect 15260 9548 15316 9604
rect 3612 9436 3668 9492
rect 13692 9436 13748 9492
rect 15148 9436 15204 9492
rect 15372 9436 15428 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 26908 9548 26964 9604
rect 27468 9548 27524 9604
rect 30156 9548 30212 9604
rect 32396 9548 32452 9604
rect 33404 9548 33460 9604
rect 29372 9436 29428 9492
rect 44268 9436 44324 9492
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 6076 9324 6132 9380
rect 9996 9324 10052 9380
rect 23660 9324 23716 9380
rect 26684 9324 26740 9380
rect 38780 9324 38836 9380
rect 32956 9212 33012 9268
rect 33740 9212 33796 9268
rect 20076 9100 20132 9156
rect 28924 9100 28980 9156
rect 30268 9100 30324 9156
rect 38892 9100 38948 9156
rect 3612 8988 3668 9044
rect 13580 8988 13636 9044
rect 13804 8988 13860 9044
rect 16268 8988 16324 9044
rect 19628 8988 19684 9044
rect 36876 8988 36932 9044
rect 23436 8876 23492 8932
rect 28028 8876 28084 8932
rect 28252 8876 28308 8932
rect 32508 8876 32564 8932
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 15260 8764 15316 8820
rect 15932 8764 15988 8820
rect 31052 8764 31108 8820
rect 32956 8764 33012 8820
rect 13356 8652 13412 8708
rect 13580 8652 13636 8708
rect 19516 8652 19572 8708
rect 32284 8652 32340 8708
rect 35196 8652 35252 8708
rect 44268 8652 44324 8708
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 20076 8540 20132 8596
rect 32172 8540 32228 8596
rect 33852 8540 33908 8596
rect 44156 8540 44212 8596
rect 45388 8540 45444 8596
rect 38444 8428 38500 8484
rect 24892 8316 24948 8372
rect 29932 8316 29988 8372
rect 32284 8316 32340 8372
rect 2268 8204 2324 8260
rect 15708 8204 15764 8260
rect 19516 8204 19572 8260
rect 30044 8204 30100 8260
rect 35868 8204 35924 8260
rect 38780 8204 38836 8260
rect 13692 7980 13748 8036
rect 19852 7980 19908 8036
rect 20076 7980 20132 8036
rect 30268 7980 30324 8036
rect 33068 7980 33124 8036
rect 46732 7980 46788 8036
rect 20188 7868 20244 7924
rect 32956 7868 33012 7924
rect 33404 7868 33460 7924
rect 34860 7868 34916 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 13356 7756 13412 7812
rect 18508 7756 18564 7812
rect 28252 7756 28308 7812
rect 30044 7756 30100 7812
rect 35308 7756 35364 7812
rect 44156 7756 44212 7812
rect 13692 7644 13748 7700
rect 33516 7644 33572 7700
rect 6748 7532 6804 7588
rect 15148 7420 15204 7476
rect 16268 7420 16324 7476
rect 26908 7420 26964 7476
rect 28252 7420 28308 7476
rect 38332 7420 38388 7476
rect 46732 7420 46788 7476
rect 9996 7308 10052 7364
rect 23436 7308 23492 7364
rect 25228 7308 25284 7364
rect 29932 7308 29988 7364
rect 30156 7308 30212 7364
rect 10556 7196 10612 7252
rect 11676 7196 11732 7252
rect 20188 7196 20244 7252
rect 21308 7196 21364 7252
rect 7980 7084 8036 7140
rect 9772 7084 9828 7140
rect 10668 7084 10724 7140
rect 15260 7084 15316 7140
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 32508 7084 32564 7140
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 15596 6972 15652 7028
rect 26908 6972 26964 7028
rect 29932 6972 29988 7028
rect 33404 6860 33460 6916
rect 14028 6748 14084 6804
rect 20188 6748 20244 6804
rect 33964 6748 34020 6804
rect 47628 6748 47684 6804
rect 9884 6524 9940 6580
rect 42140 6524 42196 6580
rect 45948 6524 46004 6580
rect 45388 6412 45444 6468
rect 10668 6300 10724 6356
rect 15596 6300 15652 6356
rect 18620 6300 18676 6356
rect 21756 6300 21812 6356
rect 32732 6300 32788 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 13468 6188 13524 6244
rect 13692 6076 13748 6132
rect 15484 6076 15540 6132
rect 29036 6076 29092 6132
rect 21868 5964 21924 6020
rect 25788 5964 25844 6020
rect 35308 5964 35364 6020
rect 36988 5964 37044 6020
rect 38556 5964 38612 6020
rect 42140 5964 42196 6020
rect 22988 5852 23044 5908
rect 25676 5852 25732 5908
rect 35756 5852 35812 5908
rect 35308 5740 35364 5796
rect 15260 5628 15316 5684
rect 16380 5628 16436 5684
rect 27580 5628 27636 5684
rect 21196 5516 21252 5572
rect 32732 5516 32788 5572
rect 35756 5516 35812 5572
rect 40796 5516 40852 5572
rect 41468 5516 41524 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 21868 5292 21924 5348
rect 35084 5292 35140 5348
rect 18620 5068 18676 5124
rect 28700 5068 28756 5124
rect 41692 5068 41748 5124
rect 14924 4956 14980 5012
rect 15484 4956 15540 5012
rect 18060 4956 18116 5012
rect 25564 4956 25620 5012
rect 43372 4956 43428 5012
rect 13692 4844 13748 4900
rect 30156 4844 30212 4900
rect 24892 4732 24948 4788
rect 37324 4732 37380 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 15372 4620 15428 4676
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 15820 4620 15876 4676
rect 21756 4620 21812 4676
rect 13468 4508 13524 4564
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 9772 4396 9828 4452
rect 18844 4396 18900 4452
rect 25116 4396 25172 4452
rect 30716 4396 30772 4452
rect 42364 4396 42420 4452
rect 19628 4284 19684 4340
rect 12908 4172 12964 4228
rect 15372 4172 15428 4228
rect 26796 4172 26852 4228
rect 25788 4060 25844 4116
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 15708 3836 15764 3892
rect 24220 3836 24276 3892
rect 29148 3836 29204 3892
rect 29820 3836 29876 3892
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 16156 3724 16212 3780
rect 23660 3724 23716 3780
rect 25116 3724 25172 3780
rect 43372 3724 43428 3780
rect 7980 3612 8036 3668
rect 14140 3612 14196 3668
rect 15484 3612 15540 3668
rect 18844 3612 18900 3668
rect 22764 3612 22820 3668
rect 24220 3612 24276 3668
rect 25676 3612 25732 3668
rect 38556 3612 38612 3668
rect 15708 3500 15764 3556
rect 18284 3500 18340 3556
rect 29820 3500 29876 3556
rect 37100 3500 37156 3556
rect 42364 3500 42420 3556
rect 17948 3388 18004 3444
rect 2828 3276 2884 3332
rect 15036 3276 15092 3332
rect 22764 3276 22820 3332
rect 29148 3276 29204 3332
rect 37660 3276 37716 3332
rect 38668 3276 38724 3332
rect 3612 3164 3668 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 22204 3164 22260 3220
rect 23660 3164 23716 3220
rect 30716 3164 30772 3220
rect 37100 3164 37156 3220
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 2604 3052 2660 3108
rect 10556 3052 10612 3108
rect 13692 3052 13748 3108
rect 21756 3052 21812 3108
rect 29036 2940 29092 2996
rect 2268 2828 2324 2884
rect 22092 2828 22148 2884
rect 3612 2716 3668 2772
rect 38108 2716 38164 2772
rect 25004 2604 25060 2660
rect 48860 2604 48916 2660
rect 23548 2492 23604 2548
rect 38556 2492 38612 2548
rect 42028 2492 42084 2548
rect 47628 2492 47684 2548
rect 13468 2380 13524 2436
rect 16044 2380 16100 2436
rect 16268 2380 16324 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 26796 2380 26852 2436
rect 41692 2380 41748 2436
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 14812 2268 14868 2324
rect 18732 2268 18788 2324
rect 23660 2268 23716 2324
rect 33740 2268 33796 2324
rect 38108 2268 38164 2324
rect 6300 2156 6356 2212
rect 16044 2156 16100 2212
rect 18284 2156 18340 2212
rect 19180 2156 19236 2212
rect 25340 2156 25396 2212
rect 13468 2044 13524 2100
rect 17164 2044 17220 2100
rect 10556 1932 10612 1988
rect 25004 1932 25060 1988
rect 26012 1932 26068 1988
rect 14588 1820 14644 1876
rect 14812 1820 14868 1876
rect 47628 1820 47684 1876
rect 17164 1708 17220 1764
rect 32844 1708 32900 1764
rect 15036 1596 15092 1652
rect 33964 1596 34020 1652
rect 41804 1596 41860 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 12908 1484 12964 1540
rect 20412 1484 20468 1540
rect 32732 1484 32788 1540
rect 33852 1484 33908 1540
rect 34412 1484 34468 1540
rect 6748 1372 6804 1428
rect 15148 1372 15204 1428
rect 15372 1372 15428 1428
rect 25340 1372 25396 1428
rect 37660 1372 37716 1428
rect 21980 1260 22036 1316
rect 25116 1148 25172 1204
rect 33852 1148 33908 1204
rect 41804 1148 41860 1204
rect 19516 1036 19572 1092
rect 26908 1036 26964 1092
rect 9212 924 9268 980
rect 15148 924 15204 980
rect 22988 924 23044 980
rect 25116 924 25172 980
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 40684 700 40740 756
rect 9212 588 9268 644
rect 21980 476 22036 532
rect 26124 476 26180 532
rect 26796 476 26852 532
rect 14476 364 14532 420
rect 22204 364 22260 420
rect 28700 364 28756 420
rect 40684 364 40740 420
rect 28924 140 28980 196
rect 33740 28 33796 84
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 2604 11172 2660 11182
rect 2268 8260 2324 8270
rect 2268 2884 2324 8204
rect 2604 3108 2660 11116
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 2828 10500 2884 10510
rect 2828 3332 2884 10444
rect 3612 9492 3668 9502
rect 3612 9044 3668 9436
rect 3612 8978 3668 8988
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 2828 3266 2884 3276
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 2604 3042 2660 3052
rect 3612 3220 3668 3230
rect 2268 2818 2324 2828
rect 3612 2772 3668 3164
rect 3612 2706 3668 2716
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14224
rect 20524 14196 20580 14206
rect 20524 13972 20580 14140
rect 20524 13906 20580 13916
rect 20972 14084 21028 14094
rect 17388 13748 17444 13758
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 6300 13524 6356 13534
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 6076 11284 6132 11294
rect 6076 9380 6132 11228
rect 6076 9314 6132 9324
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 6300 2212 6356 13468
rect 15820 13188 15876 13198
rect 14812 12852 14868 12862
rect 11788 12628 11844 12638
rect 11452 9940 11508 9950
rect 10108 9828 10164 9838
rect 10108 9604 10164 9772
rect 10108 9538 10164 9548
rect 11452 9604 11508 9884
rect 11452 9538 11508 9548
rect 9996 9380 10052 9390
rect 6300 2146 6356 2156
rect 6748 7588 6804 7598
rect 6748 1428 6804 7532
rect 9996 7364 10052 9324
rect 11788 7318 11844 12572
rect 14812 12404 14868 12796
rect 14812 12338 14868 12348
rect 15820 12404 15876 13132
rect 15820 12338 15876 12348
rect 16044 13188 16100 13198
rect 16044 12068 16100 13132
rect 17388 12180 17444 13692
rect 20972 13524 21028 14028
rect 20972 13458 21028 13468
rect 23660 13860 23716 13870
rect 20972 13300 21028 13310
rect 20972 12740 21028 13244
rect 20972 12674 21028 12684
rect 23548 13076 23604 13086
rect 17388 12114 17444 12124
rect 18284 12516 18340 12526
rect 16044 12002 16100 12012
rect 14252 11956 14980 11998
rect 14308 11942 14924 11956
rect 14252 11890 14308 11900
rect 14924 11890 14980 11900
rect 16268 11956 16324 11966
rect 13692 11396 13748 11406
rect 13692 9492 13748 11340
rect 13916 11396 13972 11406
rect 13916 10500 13972 11340
rect 16268 11278 16324 11900
rect 17948 11620 18004 11630
rect 16268 11222 17220 11278
rect 17164 11172 17220 11222
rect 17164 11106 17220 11116
rect 13916 10434 13972 10444
rect 14140 10500 14196 10510
rect 13692 9426 13748 9436
rect 13804 9604 13860 9614
rect 13580 9044 13636 9054
rect 13356 8708 13412 8718
rect 13356 7812 13412 8652
rect 13580 8708 13636 8988
rect 13804 9044 13860 9548
rect 13804 8978 13860 8988
rect 13580 8642 13636 8652
rect 13356 7746 13412 7756
rect 13692 8036 13748 8046
rect 13692 7700 13748 7980
rect 13692 7634 13748 7644
rect 9996 7298 10052 7308
rect 11676 7262 11844 7318
rect 10556 7252 10612 7262
rect 7980 7140 8036 7150
rect 7980 3668 8036 7084
rect 9772 7140 9828 7150
rect 10556 7138 10612 7196
rect 11676 7252 11732 7262
rect 11676 7186 11732 7196
rect 9828 7084 10612 7138
rect 9772 7082 10612 7084
rect 10668 7140 10724 7150
rect 9772 7074 9828 7082
rect 10668 6958 10724 7084
rect 9772 6902 10724 6958
rect 9772 4452 9828 6902
rect 14028 6804 14084 6814
rect 9884 6580 9940 6590
rect 9884 6418 9940 6524
rect 9884 6362 10724 6418
rect 10668 6356 10724 6362
rect 10668 6290 10724 6300
rect 13468 6244 13524 6254
rect 13468 4564 13524 6188
rect 13692 6132 13748 6142
rect 13692 4900 13748 6076
rect 13692 4834 13748 4844
rect 13468 4498 13524 4508
rect 9772 4386 9828 4396
rect 7980 3602 8036 3612
rect 12908 4228 12964 4238
rect 10556 3108 10612 3118
rect 10556 1988 10612 3052
rect 10556 1922 10612 1932
rect 12908 1540 12964 4172
rect 14028 3358 14084 6748
rect 14140 3668 14196 10444
rect 15036 10276 15092 10286
rect 15036 10018 15092 10220
rect 15036 9962 16436 10018
rect 14140 3602 14196 3612
rect 14700 9940 14756 9950
rect 13692 3302 14084 3358
rect 13692 3108 13748 3302
rect 13692 3042 13748 3052
rect 13468 2436 13524 2446
rect 13468 2100 13524 2380
rect 14700 2098 14756 9884
rect 15260 9604 16324 9658
rect 15316 9602 16324 9604
rect 15260 9538 15316 9548
rect 15148 9492 15204 9502
rect 15148 7476 15204 9436
rect 15372 9492 15428 9502
rect 15148 7410 15204 7420
rect 15260 8820 15316 8830
rect 15260 7140 15316 8764
rect 15260 7074 15316 7084
rect 15372 6238 15428 9436
rect 16268 9044 16324 9602
rect 16268 8978 16324 8988
rect 15932 8820 15988 8830
rect 15708 8260 15764 8270
rect 15708 7138 15764 8204
rect 15596 7082 15764 7138
rect 15596 7028 15652 7082
rect 15596 6962 15652 6972
rect 15148 6182 15428 6238
rect 15596 6356 15652 6366
rect 14924 5012 14980 5022
rect 14924 4618 14980 4956
rect 15148 4618 15204 6182
rect 15484 6132 15540 6142
rect 15484 6058 15540 6076
rect 15260 6002 15540 6058
rect 15260 5684 15316 6002
rect 15596 5878 15652 6300
rect 15260 5618 15316 5628
rect 15484 5822 15652 5878
rect 15484 5012 15540 5822
rect 15484 4946 15540 4956
rect 14924 4562 15204 4618
rect 15372 4676 15428 4686
rect 15372 4618 15428 4620
rect 15820 4676 15876 4686
rect 15820 4618 15876 4620
rect 15372 4562 15876 4618
rect 15932 4258 15988 8764
rect 15372 4228 15988 4258
rect 15428 4202 15988 4228
rect 16268 7476 16324 7486
rect 15372 4162 15428 4172
rect 15708 3892 15764 3902
rect 15484 3668 15540 3678
rect 15484 3358 15540 3612
rect 15708 3556 15764 3836
rect 15708 3490 15764 3500
rect 16156 3780 16212 3790
rect 16156 3358 16212 3724
rect 15036 3332 15092 3342
rect 15484 3302 16212 3358
rect 15036 2458 15092 3276
rect 15036 2402 15428 2458
rect 13468 2034 13524 2044
rect 14476 2042 14756 2098
rect 14812 2324 14868 2334
rect 12908 1474 12964 1484
rect 6748 1362 6804 1372
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 9212 980 9268 990
rect 9212 644 9268 924
rect 9212 578 9268 588
rect 14476 420 14532 2042
rect 14588 1876 14644 1886
rect 14588 1738 14644 1820
rect 14812 1876 14868 2268
rect 14812 1810 14868 1820
rect 14588 1682 15092 1738
rect 15036 1652 15092 1682
rect 15036 1586 15092 1596
rect 15148 1428 15204 1438
rect 15148 980 15204 1372
rect 15372 1428 15428 2402
rect 16044 2436 16100 2446
rect 16044 2212 16100 2380
rect 16268 2436 16324 7420
rect 16380 5684 16436 9962
rect 16380 5618 16436 5628
rect 17948 3444 18004 11564
rect 18284 6778 18340 12460
rect 18508 12516 18564 12526
rect 18508 7812 18564 12460
rect 21756 12516 21812 12526
rect 21756 12178 21812 12460
rect 23548 12292 23604 13020
rect 23548 12226 23604 12236
rect 21756 12122 22036 12178
rect 19964 12068 20020 12078
rect 19964 11998 20020 12012
rect 19964 11956 20356 11998
rect 19964 11942 20300 11956
rect 20300 11890 20356 11900
rect 21868 11956 21924 11966
rect 21868 11638 21924 11900
rect 21756 11620 21924 11638
rect 21812 11582 21924 11620
rect 21980 11620 22036 12122
rect 21756 11554 21812 11564
rect 21980 11554 22036 11564
rect 23548 11284 23604 11294
rect 19628 11172 19684 11182
rect 19628 10612 19684 11116
rect 21980 11060 22036 11070
rect 21308 10948 21364 10958
rect 19628 10546 19684 10556
rect 20076 10724 20132 10734
rect 20076 9156 20132 10668
rect 20076 9090 20132 9100
rect 21196 9828 21252 9838
rect 19628 9044 19684 9054
rect 19516 8708 19572 8718
rect 19516 8260 19572 8652
rect 19516 8194 19572 8204
rect 18508 7746 18564 7756
rect 18284 6722 18676 6778
rect 18620 6356 18676 6722
rect 18620 6290 18676 6300
rect 18620 5124 18676 5134
rect 18060 5012 18116 5022
rect 18620 4978 18676 5068
rect 18116 4956 18676 4978
rect 18060 4922 18676 4956
rect 18844 4452 18900 4462
rect 18844 3668 18900 4396
rect 19628 4340 19684 8988
rect 20076 8596 20132 8606
rect 19852 8036 19908 8046
rect 19852 7858 19908 7980
rect 20076 8036 20132 8540
rect 20076 7970 20132 7980
rect 20188 7924 20244 7934
rect 20188 7858 20244 7868
rect 19852 7802 20244 7858
rect 20188 7252 20244 7262
rect 20188 6804 20244 7196
rect 20188 6738 20244 6748
rect 21196 5572 21252 9772
rect 21308 7252 21364 10892
rect 21980 9828 22036 11004
rect 23548 10948 23604 11228
rect 23548 10882 23604 10892
rect 21980 9762 22036 9772
rect 23660 9380 23716 13804
rect 23660 9314 23716 9324
rect 23776 12572 24096 14224
rect 24436 13356 24756 14224
rect 38108 14196 38164 14206
rect 28028 14084 28084 14094
rect 28028 13978 28084 14028
rect 28252 14084 28308 14094
rect 28028 13922 28196 13978
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 28140 13412 28196 13922
rect 28140 13346 28196 13356
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 24220 12964 24276 12974
rect 24220 12516 24276 12908
rect 24220 12450 24276 12460
rect 24436 11788 24756 13300
rect 25676 13188 25732 13198
rect 25004 13078 25060 13086
rect 25676 13078 25732 13132
rect 25004 13076 25732 13078
rect 25060 13022 25732 13076
rect 25004 13010 25060 13020
rect 28252 12898 28308 14028
rect 30492 14084 30548 14094
rect 30492 13978 30548 14028
rect 30492 13922 32004 13978
rect 31948 13860 32004 13922
rect 31948 13794 32004 13804
rect 32508 13860 32564 13870
rect 32508 13636 32564 13804
rect 32508 13570 32564 13580
rect 32732 13860 32788 13870
rect 27580 12842 28308 12898
rect 31276 12852 31332 12862
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 24220 11060 24276 11070
rect 24220 10500 24276 11004
rect 24220 10434 24276 10444
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23436 8932 23492 8942
rect 23436 7364 23492 8876
rect 23436 7298 23492 7308
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 21308 7186 21364 7196
rect 21196 5506 21252 5516
rect 21756 6356 21812 6366
rect 21756 4676 21812 6300
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 21868 6020 21924 6030
rect 21868 5348 21924 5964
rect 21868 5282 21924 5292
rect 22988 5908 23044 5918
rect 21756 4610 21812 4620
rect 19628 4274 19684 4284
rect 18844 3602 18900 3612
rect 22764 3668 22820 3678
rect 17948 3378 18004 3388
rect 18284 3556 18340 3566
rect 16268 2370 16324 2380
rect 16044 2146 16100 2156
rect 18284 2212 18340 3500
rect 22764 3332 22820 3612
rect 22764 3266 22820 3276
rect 22204 3220 22260 3230
rect 21756 3108 21812 3118
rect 21756 2998 21812 3052
rect 21756 2942 22148 2998
rect 22092 2884 22148 2942
rect 22092 2818 22148 2828
rect 18732 2324 18788 2334
rect 18788 2268 19236 2278
rect 18732 2222 19236 2268
rect 18284 2146 18340 2156
rect 19180 2212 19236 2222
rect 19180 2146 19236 2156
rect 17164 2100 17220 2110
rect 17164 1764 17220 2044
rect 17164 1698 17220 1708
rect 20412 1540 20468 1550
rect 20412 1378 20468 1484
rect 15372 1362 15428 1372
rect 19516 1322 20468 1378
rect 19516 1092 19572 1322
rect 19516 1026 19572 1036
rect 21980 1316 22036 1326
rect 15148 914 15204 924
rect 21980 532 22036 1260
rect 21980 466 22036 476
rect 14476 354 14532 364
rect 22204 420 22260 3164
rect 22988 980 23044 5852
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23660 3780 23716 3790
rect 23660 3358 23716 3724
rect 23548 3302 23716 3358
rect 23548 2548 23604 3302
rect 23548 2482 23604 2492
rect 23660 3220 23716 3230
rect 23660 2324 23716 3164
rect 23660 2258 23716 2268
rect 23776 3164 24096 4676
rect 24436 10220 24756 11732
rect 25228 12628 25284 12638
rect 25228 10612 25284 12572
rect 25228 10546 25284 10556
rect 26012 11284 26068 11294
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 24892 8372 24948 8382
rect 24892 7678 24948 8316
rect 24892 7622 25284 7678
rect 25228 7364 25284 7622
rect 25228 7298 25284 7308
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 25788 6020 25844 6030
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 25676 5908 25732 5918
rect 25564 5012 25620 5022
rect 24892 4956 25564 4978
rect 24892 4922 25620 4956
rect 24892 4788 24948 4922
rect 24892 4722 24948 4732
rect 24220 3892 24276 3902
rect 24220 3668 24276 3836
rect 24220 3602 24276 3612
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 22988 914 23044 924
rect 23776 1596 24096 3108
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 22204 354 22260 364
rect 23776 0 24096 1540
rect 24436 2380 24756 3892
rect 25116 4452 25172 4462
rect 25116 3780 25172 4396
rect 25116 3714 25172 3724
rect 25676 3668 25732 5852
rect 25788 4116 25844 5964
rect 25788 4050 25844 4060
rect 25676 3602 25732 3612
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 25004 2660 25060 2670
rect 25004 1988 25060 2604
rect 25004 1922 25060 1932
rect 25340 2212 25396 2222
rect 25340 1428 25396 2156
rect 26012 1988 26068 11228
rect 26572 10724 26628 10734
rect 26572 5158 26628 10668
rect 26852 10052 26908 10062
rect 26908 9996 27524 10018
rect 26852 9962 27524 9996
rect 26684 9782 26964 9838
rect 26684 9380 26740 9782
rect 26908 9604 26964 9782
rect 26908 9538 26964 9548
rect 27468 9604 27524 9962
rect 27468 9538 27524 9548
rect 26684 9314 26740 9324
rect 26908 7476 26964 7486
rect 26908 7028 26964 7420
rect 26908 6962 26964 6972
rect 27580 5684 27636 12842
rect 31276 12718 31332 12796
rect 27692 12662 31332 12718
rect 32732 12740 32788 13804
rect 36988 13748 37044 13758
rect 33740 13300 33796 13310
rect 32732 12674 32788 12684
rect 33292 12852 33348 12862
rect 27692 12516 27748 12662
rect 27692 12450 27748 12460
rect 32956 12292 33012 12302
rect 30492 12180 30548 12190
rect 28364 11956 28644 11998
rect 28420 11942 28644 11956
rect 28364 11890 28420 11900
rect 28252 10948 28308 10958
rect 28028 8932 28084 8942
rect 28028 8758 28084 8876
rect 28252 8932 28308 10892
rect 28588 10378 28644 11942
rect 30492 11844 30548 12124
rect 30492 11778 30548 11788
rect 30716 11732 30772 11742
rect 30716 10500 30772 11676
rect 32956 11458 33012 12236
rect 32956 11402 33124 11458
rect 31612 11172 31668 11182
rect 31612 11098 31668 11116
rect 30716 10434 30772 10444
rect 31276 11042 31668 11098
rect 28588 10322 28980 10378
rect 28924 9156 28980 10322
rect 30268 10276 30324 10286
rect 29372 9828 29428 9838
rect 29372 9492 29428 9772
rect 30268 9658 30324 10220
rect 31276 10052 31332 11042
rect 31500 10500 31556 10510
rect 31500 10276 31556 10444
rect 31500 10210 31556 10220
rect 31276 9986 31332 9996
rect 31612 9940 31668 9950
rect 31612 9838 31668 9884
rect 31612 9782 32452 9838
rect 30156 9604 30324 9658
rect 30212 9602 30324 9604
rect 32396 9604 32452 9782
rect 30156 9538 30212 9548
rect 32396 9538 32452 9548
rect 29372 9426 29428 9436
rect 32956 9268 33012 9278
rect 28924 9090 28980 9100
rect 30268 9156 30324 9166
rect 30324 9100 31108 9118
rect 30268 9062 31108 9100
rect 28252 8866 28308 8876
rect 31052 8820 31108 9062
rect 28028 8702 28756 8758
rect 31052 8754 31108 8764
rect 32508 8932 32564 8942
rect 32508 8758 32564 8876
rect 28252 7812 28308 7822
rect 28252 7476 28308 7756
rect 28252 7410 28308 7420
rect 27580 5618 27636 5628
rect 26572 5102 26964 5158
rect 26796 4228 26852 4238
rect 26796 2436 26852 4172
rect 26796 2370 26852 2380
rect 26012 1922 26068 1932
rect 25340 1362 25396 1372
rect 25116 1204 25172 1214
rect 25116 980 25172 1148
rect 26908 1092 26964 5102
rect 28700 5124 28756 8702
rect 32284 8708 32564 8758
rect 32956 8820 33012 9212
rect 32956 8754 33012 8764
rect 32340 8702 32564 8708
rect 32284 8642 32340 8652
rect 32172 8596 32228 8606
rect 32228 8540 32340 8578
rect 32172 8522 32340 8540
rect 29932 8372 30212 8398
rect 29988 8342 30212 8372
rect 29932 8306 29988 8316
rect 30044 8260 30100 8270
rect 30044 7812 30100 8204
rect 30156 8218 30212 8342
rect 32284 8372 32340 8522
rect 32284 8306 32340 8316
rect 30156 8162 30324 8218
rect 30268 8036 30324 8162
rect 30268 7970 30324 7980
rect 33068 8036 33124 11402
rect 33068 7970 33124 7980
rect 32956 7924 33012 7934
rect 32956 7858 33012 7868
rect 30044 7746 30100 7756
rect 32508 7802 33012 7858
rect 29932 7364 29988 7374
rect 29932 7028 29988 7308
rect 29932 6962 29988 6972
rect 30156 7364 30212 7374
rect 28700 5058 28756 5068
rect 29036 6132 29092 6142
rect 29036 2996 29092 6076
rect 30156 4900 30212 7308
rect 32508 7140 32564 7802
rect 32508 7074 32564 7084
rect 33292 6778 33348 12796
rect 33628 10612 33684 10622
rect 33516 10500 33572 10510
rect 33404 9604 33460 9614
rect 33404 7924 33460 9548
rect 33404 7858 33460 7868
rect 33516 7700 33572 10444
rect 33516 7634 33572 7644
rect 33628 6958 33684 10556
rect 33740 9268 33796 13244
rect 33740 9202 33796 9212
rect 33852 13188 33908 13198
rect 33852 8596 33908 13132
rect 34076 13188 34132 13198
rect 34076 11172 34132 13132
rect 36988 12292 37044 13692
rect 36988 12226 37044 12236
rect 37324 12180 37380 12190
rect 35532 12068 35588 12078
rect 35532 11998 35588 12012
rect 34972 11956 35588 11998
rect 35028 11942 35588 11956
rect 34972 11890 35028 11900
rect 34076 11106 34132 11116
rect 35196 10276 35252 10286
rect 35196 8708 35252 10220
rect 35420 10276 35476 10286
rect 35420 9716 35476 10220
rect 35420 9650 35476 9660
rect 36876 9044 36932 9054
rect 36876 8938 36932 8988
rect 36876 8882 37044 8938
rect 35196 8642 35252 8652
rect 33852 8530 33908 8540
rect 35868 8260 35924 8270
rect 35308 8204 35868 8218
rect 35308 8162 35924 8204
rect 34860 7924 34916 7934
rect 34860 7858 34916 7868
rect 34860 7802 35140 7858
rect 33404 6916 33684 6958
rect 33460 6902 33684 6916
rect 33740 6902 34020 6958
rect 33404 6850 33460 6860
rect 33740 6778 33796 6902
rect 33292 6722 33796 6778
rect 33964 6804 34020 6902
rect 33964 6738 34020 6748
rect 32732 6356 32788 6366
rect 32732 5572 32788 6300
rect 32732 5506 32788 5516
rect 35084 5348 35140 7802
rect 35308 7812 35364 8162
rect 35308 7746 35364 7756
rect 35308 6020 35364 6030
rect 35308 5796 35364 5964
rect 36988 6020 37044 8882
rect 36988 5954 37044 5964
rect 35308 5730 35364 5740
rect 35756 5908 35812 5918
rect 35756 5572 35812 5852
rect 35756 5506 35812 5516
rect 35084 5282 35140 5292
rect 30156 4834 30212 4844
rect 37324 4788 37380 12124
rect 38108 11956 38164 14140
rect 38444 13636 38500 13646
rect 38444 13438 38500 13580
rect 38892 13636 38948 13646
rect 38444 13412 38668 13438
rect 38444 13382 38612 13412
rect 38612 13346 38668 13356
rect 38108 11890 38164 11900
rect 38780 9380 38836 9390
rect 38444 8484 38500 8494
rect 38444 7498 38500 8428
rect 38780 8260 38836 9324
rect 38892 9156 38948 13580
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 39340 12404 39396 12414
rect 39228 12348 39340 12358
rect 39228 12302 39396 12348
rect 39228 12180 39284 12302
rect 39228 12114 39284 12124
rect 43596 11620 43652 11630
rect 43596 11284 43652 11564
rect 43596 11218 43652 11228
rect 43776 11004 44096 12516
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 38892 9090 38948 9100
rect 42028 10388 42084 10398
rect 38780 8194 38836 8204
rect 38332 7476 38500 7498
rect 38388 7442 38500 7476
rect 38332 7410 38388 7420
rect 38556 6020 38612 6030
rect 38556 5158 38612 5964
rect 40796 5572 40852 5582
rect 41468 5572 41524 5582
rect 40852 5516 41468 5518
rect 40796 5462 41524 5516
rect 38556 5102 38724 5158
rect 37324 4722 37380 4732
rect 30716 4452 30772 4462
rect 29148 3892 29204 3902
rect 29148 3332 29204 3836
rect 29820 3892 29876 3902
rect 29820 3556 29876 3836
rect 29820 3490 29876 3500
rect 29148 3266 29204 3276
rect 30716 3220 30772 4396
rect 38556 3668 38612 3678
rect 30716 3154 30772 3164
rect 37100 3556 37156 3566
rect 37100 3220 37156 3500
rect 37100 3154 37156 3164
rect 37660 3332 37716 3342
rect 29036 2930 29092 2940
rect 33740 2324 33796 2334
rect 32844 1764 32900 1774
rect 32844 1558 32900 1708
rect 32732 1540 32900 1558
rect 32788 1502 32900 1540
rect 32732 1474 32788 1484
rect 26908 1026 26964 1036
rect 25116 914 25172 924
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 26124 532 26180 542
rect 26796 532 26852 542
rect 26180 476 26796 478
rect 26124 422 26852 476
rect 28700 420 28756 430
rect 28700 298 28756 364
rect 28700 242 28980 298
rect 28924 196 28980 242
rect 28924 130 28980 140
rect 33740 84 33796 2268
rect 33964 1652 34020 1662
rect 33964 1558 34020 1596
rect 33852 1540 33908 1550
rect 33964 1540 34468 1558
rect 33964 1502 34412 1540
rect 33852 1204 33908 1484
rect 34412 1474 34468 1484
rect 37660 1428 37716 3276
rect 38108 2772 38164 2782
rect 38108 2324 38164 2716
rect 38556 2548 38612 3612
rect 38668 3332 38724 5102
rect 38668 3266 38724 3276
rect 41692 5124 41748 5134
rect 38556 2482 38612 2492
rect 41692 2436 41748 5068
rect 42028 2548 42084 10332
rect 43776 9436 44096 10948
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 43776 7868 44096 9380
rect 44268 9492 44324 9502
rect 44268 8708 44324 9436
rect 44268 8642 44324 8652
rect 44436 8652 44756 10164
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 42140 6580 42196 6590
rect 42140 6020 42196 6524
rect 42140 5954 42196 5964
rect 43776 6300 44096 7812
rect 44156 8596 44212 8606
rect 44156 7812 44212 8540
rect 44156 7746 44212 7756
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 45948 13188 46004 13198
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 43372 5012 43428 5022
rect 42364 4452 42420 4462
rect 42364 3556 42420 4396
rect 43372 3780 43428 4956
rect 43372 3714 43428 3724
rect 43776 4732 44096 6244
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 42364 3490 42420 3500
rect 42028 2482 42084 2492
rect 43776 3164 44096 4676
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 41692 2370 41748 2380
rect 38108 2258 38164 2268
rect 37660 1362 37716 1372
rect 41804 1652 41860 1662
rect 33852 1138 33908 1148
rect 41804 1204 41860 1596
rect 41804 1138 41860 1148
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 40684 756 40740 766
rect 40684 420 40740 700
rect 40684 354 40740 364
rect 33740 18 33796 28
rect 43776 0 44096 1540
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 45388 8596 45444 8606
rect 45388 6468 45444 8540
rect 45948 6580 46004 13132
rect 48860 12068 48916 12078
rect 47628 10836 47684 10846
rect 46732 8036 46788 8046
rect 46732 7476 46788 7980
rect 46732 7410 46788 7420
rect 47628 6804 47684 10780
rect 47628 6738 47684 6748
rect 45948 6514 46004 6524
rect 45388 6402 45444 6412
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44436 3948 44756 5460
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 48860 2660 48916 12012
rect 48860 2594 48916 2604
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 47628 2548 47684 2558
rect 47628 1876 47684 2492
rect 47628 1810 47684 1820
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 41328 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 42112 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 44464 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 41216 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 46928 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 37744 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 44576 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 42448 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 54320 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 38528 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 41552 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 47488 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 18480 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 27216 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 30240 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 49840 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 28784 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 23296 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 5040 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 52192 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 30464 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 9856 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 23296 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 34272 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 39200 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 48272 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 21392 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 32144 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 49168 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 5600 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 4592 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 10304 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 14896 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 11088 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 11088 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 2240 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 13552 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 14336 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 31136 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 32480 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform 1 0 46816 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 37744 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 9632 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform 1 0 51296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 50064 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 21392 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 18032 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform -1 0 25648 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 37408 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 49952 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform 1 0 51520 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 50288 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 30800 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 36400 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 37520 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 36400 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform -1 0 23184 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 34496 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform -1 0 21504 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 35952 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform -1 0 28672 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 52080 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 51520 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform 1 0 41440 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform -1 0 20720 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform -1 0 21056 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform -1 0 29232 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 33152 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 46256 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 35504 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 43792 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 19712 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 50736 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 14112 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform -1 0 20272 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 10192 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 17584 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 13328 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform -1 0 22288 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform -1 0 4704 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 6720 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 2688 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 3584 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 6496 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 7504 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 6160 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 3696 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 14448 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 9632 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 37072 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 29232 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 2800 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 4256 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 7168 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _104_
timestamp 1486834041
transform -1 0 26320 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1486834041
transform 1 0 1008 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_444
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 54656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 54880 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_26
timestamp 1486834041
transform 1 0 3584 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_42
timestamp 1486834041
transform 1 0 5376 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_58
timestamp 1486834041
transform 1 0 7168 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1486834041
transform 1 0 12320 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1486834041
transform 1 0 13216 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_114
timestamp 1486834041
transform 1 0 13440 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_123
timestamp 1486834041
transform 1 0 14448 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_146
timestamp 1486834041
transform 1 0 17024 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_155
timestamp 1486834041
transform 1 0 18032 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_171
timestamp 1486834041
transform 1 0 19824 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_175
timestamp 1486834041
transform 1 0 20272 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_177
timestamp 1486834041
transform 1 0 20496 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_186
timestamp 1486834041
transform 1 0 21504 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_202
timestamp 1486834041
transform 1 0 23296 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_220
timestamp 1486834041
transform 1 0 25312 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_236
timestamp 1486834041
transform 1 0 27104 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_244
timestamp 1486834041
transform 1 0 28000 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_248
timestamp 1486834041
transform 1 0 28448 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_250
timestamp 1486834041
transform 1 0 28672 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_259
timestamp 1486834041
transform 1 0 29680 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_263
timestamp 1486834041
transform 1 0 30128 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_272
timestamp 1486834041
transform 1 0 31136 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_282
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_346
timestamp 1486834041
transform 1 0 39424 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_416
timestamp 1486834041
transform 1 0 47264 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 55776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 56224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_18
timestamp 1486834041
transform 1 0 2688 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_26
timestamp 1486834041
transform 1 0 3584 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_193
timestamp 1486834041
transform 1 0 22288 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_213
timestamp 1486834041
transform 1 0 24528 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_223
timestamp 1486834041
transform 1 0 25648 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_239
timestamp 1486834041
transform 1 0 27440 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_243
timestamp 1486834041
transform 1 0 27888 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_255
timestamp 1486834041
transform 1 0 29232 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_271
timestamp 1486834041
transform 1 0 31024 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_279
timestamp 1486834041
transform 1 0 31920 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_289
timestamp 1486834041
transform 1 0 33040 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_305
timestamp 1486834041
transform 1 0 34832 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_313
timestamp 1486834041
transform 1 0 35728 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_325
timestamp 1486834041
transform 1 0 37072 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_329
timestamp 1486834041
transform 1 0 37520 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_339
timestamp 1486834041
transform 1 0 38640 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_371
timestamp 1486834041
transform 1 0 42224 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_379
timestamp 1486834041
transform 1 0 43120 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_383
timestamp 1486834041
transform 1 0 43568 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 51184 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_80
timestamp 1486834041
transform 1 0 9632 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_84
timestamp 1486834041
transform 1 0 10080 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_94
timestamp 1486834041
transform 1 0 11200 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_126
timestamp 1486834041
transform 1 0 14784 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_135
timestamp 1486834041
transform 1 0 15792 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1486834041
transform 1 0 16240 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_158
timestamp 1486834041
transform 1 0 18368 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_167
timestamp 1486834041
transform 1 0 19376 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_199
timestamp 1486834041
transform 1 0 22960 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_207
timestamp 1486834041
transform 1 0 23856 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_276
timestamp 1486834041
transform 1 0 31584 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_290
timestamp 1486834041
transform 1 0 33152 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_298
timestamp 1486834041
transform 1 0 34048 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_302
timestamp 1486834041
transform 1 0 34496 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_311
timestamp 1486834041
transform 1 0 35504 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_327
timestamp 1486834041
transform 1 0 37296 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_343
timestamp 1486834041
transform 1 0 39088 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_347
timestamp 1486834041
transform 1 0 39536 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 39760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_384
timestamp 1486834041
transform 1 0 43680 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_393
timestamp 1486834041
transform 1 0 44688 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_409
timestamp 1486834041
transform 1 0 46480 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1486834041
transform 1 0 47376 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1486834041
transform 1 0 47600 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_438
timestamp 1486834041
transform 1 0 49728 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_447
timestamp 1486834041
transform 1 0 50736 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_451
timestamp 1486834041
transform 1 0 51184 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_453
timestamp 1486834041
transform 1 0 51408 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 56224 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 56448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_47
timestamp 1486834041
transform 1 0 5936 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_79
timestamp 1486834041
transform 1 0 9520 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_95
timestamp 1486834041
transform 1 0 11312 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1486834041
transform 1 0 12208 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 27664 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 35504 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_317
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_327
timestamp 1486834041
transform 1 0 37296 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_343
timestamp 1486834041
transform 1 0 39088 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_352
timestamp 1486834041
transform 1 0 40096 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_360
timestamp 1486834041
transform 1 0 40992 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_364
timestamp 1486834041
transform 1 0 41440 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_373
timestamp 1486834041
transform 1 0 42448 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_381
timestamp 1486834041
transform 1 0 43344 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_387
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_419
timestamp 1486834041
transform 1 0 47600 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_427
timestamp 1486834041
transform 1 0 48496 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_431
timestamp 1486834041
transform 1 0 48944 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_441
timestamp 1486834041
transform 1 0 50064 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_449
timestamp 1486834041
transform 1 0 50960 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_453
timestamp 1486834041
transform 1 0 51408 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_457
timestamp 1486834041
transform 1 0 51856 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_467
timestamp 1486834041
transform 1 0 52976 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_10
timestamp 1486834041
transform 1 0 1792 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_19
timestamp 1486834041
transform 1 0 2800 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_27
timestamp 1486834041
transform 1 0 3696 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_36
timestamp 1486834041
transform 1 0 4704 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_52
timestamp 1486834041
transform 1 0 6496 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_61
timestamp 1486834041
transform 1 0 7504 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_69
timestamp 1486834041
transform 1 0 8400 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_104
timestamp 1486834041
transform 1 0 12320 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_113
timestamp 1486834041
transform 1 0 13328 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_122
timestamp 1486834041
transform 1 0 14336 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_138
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 27104 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_240
timestamp 1486834041
transform 1 0 27552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_250
timestamp 1486834041
transform 1 0 28672 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_266
timestamp 1486834041
transform 1 0 30464 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_274
timestamp 1486834041
transform 1 0 31360 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_278
timestamp 1486834041
transform 1 0 31808 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_346
timestamp 1486834041
transform 1 0 39424 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_384
timestamp 1486834041
transform 1 0 43680 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_400
timestamp 1486834041
transform 1 0 45472 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_408
timestamp 1486834041
transform 1 0 46368 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_438
timestamp 1486834041
transform 1 0 49728 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_446
timestamp 1486834041
transform 1 0 50624 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_450
timestamp 1486834041
transform 1 0 51072 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 55776 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 56224 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 11984 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_111
timestamp 1486834041
transform 1 0 13104 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_136
timestamp 1486834041
transform 1 0 15904 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_152
timestamp 1486834041
transform 1 0 17696 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_160
timestamp 1486834041
transform 1 0 18592 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_164
timestamp 1486834041
transform 1 0 19040 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_166
timestamp 1486834041
transform 1 0 19264 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1486834041
transform 1 0 27664 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_263
timestamp 1486834041
transform 1 0 30128 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_272
timestamp 1486834041
transform 1 0 31136 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_284
timestamp 1486834041
transform 1 0 32480 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_300
timestamp 1486834041
transform 1 0 34272 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_308
timestamp 1486834041
transform 1 0 35168 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_312
timestamp 1486834041
transform 1 0 35616 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 35840 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_381
timestamp 1486834041
transform 1 0 43344 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_451
timestamp 1486834041
transform 1 0 51184 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_18
timestamp 1486834041
transform 1 0 2688 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_22
timestamp 1486834041
transform 1 0 3136 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_32
timestamp 1486834041
transform 1 0 4256 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_64
timestamp 1486834041
transform 1 0 7840 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1486834041
transform 1 0 8288 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1486834041
transform 1 0 15904 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_174
timestamp 1486834041
transform 1 0 20160 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_176
timestamp 1486834041
transform 1 0 20384 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_185
timestamp 1486834041
transform 1 0 21392 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_201
timestamp 1486834041
transform 1 0 23184 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_276
timestamp 1486834041
transform 1 0 31584 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_314
timestamp 1486834041
transform 1 0 35840 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_322
timestamp 1486834041
transform 1 0 36736 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_326
timestamp 1486834041
transform 1 0 37184 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_336
timestamp 1486834041
transform 1 0 38304 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_360
timestamp 1486834041
transform 1 0 40992 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_372
timestamp 1486834041
transform 1 0 42336 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_404
timestamp 1486834041
transform 1 0 45920 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_454
timestamp 1486834041
transform 1 0 51520 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 55776 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 56224 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1486834041
transform 1 0 9296 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_81
timestamp 1486834041
transform 1 0 9744 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_90
timestamp 1486834041
transform 1 0 10752 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_98
timestamp 1486834041
transform 1 0 11648 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_102
timestamp 1486834041
transform 1 0 12096 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_104
timestamp 1486834041
transform 1 0 12320 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_139
timestamp 1486834041
transform 1 0 16240 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_159
timestamp 1486834041
transform 1 0 18480 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_161
timestamp 1486834041
transform 1 0 18704 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_170
timestamp 1486834041
transform 1 0 19712 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 20160 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_263
timestamp 1486834041
transform 1 0 30128 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_265
timestamp 1486834041
transform 1 0 30352 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_274
timestamp 1486834041
transform 1 0 31360 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_306
timestamp 1486834041
transform 1 0 34944 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 35840 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_435
timestamp 1486834041
transform 1 0 49392 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_443
timestamp 1486834041
transform 1 0 50288 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_16
timestamp 1486834041
transform 1 0 2464 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_32
timestamp 1486834041
transform 1 0 4256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_40
timestamp 1486834041
transform 1 0 5152 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_52
timestamp 1486834041
transform 1 0 6496 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_68
timestamp 1486834041
transform 1 0 8288 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_80
timestamp 1486834041
transform 1 0 9632 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_112
timestamp 1486834041
transform 1 0 13216 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_128
timestamp 1486834041
transform 1 0 15008 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 15904 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_158
timestamp 1486834041
transform 1 0 18368 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_170
timestamp 1486834041
transform 1 0 19712 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_179
timestamp 1486834041
transform 1 0 20720 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_183
timestamp 1486834041
transform 1 0 21168 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_193
timestamp 1486834041
transform 1 0 22288 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_276
timestamp 1486834041
transform 1 0 31584 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_282
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_298
timestamp 1486834041
transform 1 0 34048 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_310
timestamp 1486834041
transform 1 0 35392 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_342
timestamp 1486834041
transform 1 0 38976 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_360
timestamp 1486834041
transform 1 0 40992 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_392
timestamp 1486834041
transform 1 0 44576 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_408
timestamp 1486834041
transform 1 0 46368 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 47264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_424
timestamp 1486834041
transform 1 0 48160 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_433
timestamp 1486834041
transform 1 0 49168 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_437
timestamp 1486834041
transform 1 0 49616 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_439
timestamp 1486834041
transform 1 0 49840 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 56224 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 56448 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1486834041
transform 1 0 1120 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_27
timestamp 1486834041
transform 1 0 3696 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_45
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_54
timestamp 1486834041
transform 1 0 6720 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_70
timestamp 1486834041
transform 1 0 8512 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_78
timestamp 1486834041
transform 1 0 9408 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_82
timestamp 1486834041
transform 1 0 9856 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_84
timestamp 1486834041
transform 1 0 10080 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_93
timestamp 1486834041
transform 1 0 11088 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 11984 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 19824 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_201
timestamp 1486834041
transform 1 0 23184 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_233
timestamp 1486834041
transform 1 0 26768 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1486834041
transform 1 0 27664 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_381
timestamp 1486834041
transform 1 0 43344 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_403
timestamp 1486834041
transform 1 0 45808 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_411
timestamp 1486834041
transform 1 0 46704 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_421
timestamp 1486834041
transform 1 0 47824 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_429
timestamp 1486834041
transform 1 0 48720 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_23
timestamp 1486834041
transform 1 0 3248 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_27
timestamp 1486834041
transform 1 0 3696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_52
timestamp 1486834041
transform 1 0 6496 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_68
timestamp 1486834041
transform 1 0 8288 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_76
timestamp 1486834041
transform 1 0 9184 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_93
timestamp 1486834041
transform 1 0 11088 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_125
timestamp 1486834041
transform 1 0 14672 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_133
timestamp 1486834041
transform 1 0 15568 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_137
timestamp 1486834041
transform 1 0 16016 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_151
timestamp 1486834041
transform 1 0 17584 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_167
timestamp 1486834041
transform 1 0 19376 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_171
timestamp 1486834041
transform 1 0 19824 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_173
timestamp 1486834041
transform 1 0 20048 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_182
timestamp 1486834041
transform 1 0 21056 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_198
timestamp 1486834041
transform 1 0 22848 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_220
timestamp 1486834041
transform 1 0 25312 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_229
timestamp 1486834041
transform 1 0 26320 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_261
timestamp 1486834041
transform 1 0 29904 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_277
timestamp 1486834041
transform 1 0 31696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_314
timestamp 1486834041
transform 1 0 35840 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_323
timestamp 1486834041
transform 1 0 36848 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_339
timestamp 1486834041
transform 1 0 38640 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_347
timestamp 1486834041
transform 1 0 39536 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_349
timestamp 1486834041
transform 1 0 39760 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_360
timestamp 1486834041
transform 1 0 40992 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_362
timestamp 1486834041
transform 1 0 41216 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_371
timestamp 1486834041
transform 1 0 42224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_381
timestamp 1486834041
transform 1 0 43344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_389
timestamp 1486834041
transform 1 0 44240 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_399
timestamp 1486834041
transform 1 0 45360 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_415
timestamp 1486834041
transform 1 0 47152 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 56224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 56448 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_41
timestamp 1486834041
transform 1 0 5264 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_99
timestamp 1486834041
transform 1 0 11760 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_103
timestamp 1486834041
transform 1 0 12208 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_135
timestamp 1486834041
transform 1 0 15792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_151
timestamp 1486834041
transform 1 0 17584 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_195
timestamp 1486834041
transform 1 0 22512 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_227
timestamp 1486834041
transform 1 0 26096 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1486834041
transform 1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 35504 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_321
timestamp 1486834041
transform 1 0 36624 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_331
timestamp 1486834041
transform 1 0 37744 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_347
timestamp 1486834041
transform 1 0 39536 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_355
timestamp 1486834041
transform 1 0 40432 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_359
timestamp 1486834041
transform 1 0 40880 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_361
timestamp 1486834041
transform 1 0 41104 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_378
timestamp 1486834041
transform 1 0 43008 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_382
timestamp 1486834041
transform 1 0 43456 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 43680 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_403
timestamp 1486834041
transform 1 0 45808 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_411
timestamp 1486834041
transform 1 0 46704 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_415
timestamp 1486834041
transform 1 0 47152 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_417
timestamp 1486834041
transform 1 0 47376 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_426
timestamp 1486834041
transform 1 0 48384 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_207
timestamp 1486834041
transform 1 0 23856 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_209
timestamp 1486834041
transform 1 0 24080 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_252
timestamp 1486834041
transform 1 0 28896 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_268
timestamp 1486834041
transform 1 0 30688 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_277
timestamp 1486834041
transform 1 0 31696 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 31920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_298
timestamp 1486834041
transform 1 0 34048 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_308
timestamp 1486834041
transform 1 0 35168 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_340
timestamp 1486834041
transform 1 0 38752 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_348
timestamp 1486834041
transform 1 0 39648 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_384
timestamp 1486834041
transform 1 0 43680 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_400
timestamp 1486834041
transform 1 0 45472 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_408
timestamp 1486834041
transform 1 0 46368 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_412
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_487
timestamp 1486834041
transform 1 0 55216 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 55440 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 56224 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 56448 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_115
timestamp 1486834041
transform 1 0 13552 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_185
timestamp 1486834041
transform 1 0 21392 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_215
timestamp 1486834041
transform 1 0 24752 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_231
timestamp 1486834041
transform 1 0 26544 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_235
timestamp 1486834041
transform 1 0 26992 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_255
timestamp 1486834041
transform 1 0 29232 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_287
timestamp 1486834041
transform 1 0 32816 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_303
timestamp 1486834041
transform 1 0 34608 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_311
timestamp 1486834041
transform 1 0 35504 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_325
timestamp 1486834041
transform 1 0 37072 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_337
timestamp 1486834041
transform 1 0 38416 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_369
timestamp 1486834041
transform 1 0 42000 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_391
timestamp 1486834041
transform 1 0 44464 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_400
timestamp 1486834041
transform 1 0 45472 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_404
timestamp 1486834041
transform 1 0 45920 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_406
timestamp 1486834041
transform 1 0 46144 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 51184 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_224
timestamp 1486834041
transform 1 0 25760 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_232
timestamp 1486834041
transform 1 0 26656 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_236
timestamp 1486834041
transform 1 0 27104 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_342
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_376
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_392
timestamp 1486834041
transform 1 0 44576 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_439
timestamp 1486834041
transform 1 0 49840 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 50064 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_472
timestamp 1486834041
transform 1 0 53536 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1486834041
transform 1 0 55776 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_496
timestamp 1486834041
transform 1 0 56224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_498
timestamp 1486834041
transform 1 0 56448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 53424 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 53984 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 54992 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 53424 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 53984 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 54992 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 53424 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 54992 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 54992 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 53424 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 52416 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 54992 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 53984 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 53424 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 53984 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 50848 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 52416 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 48048 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 50848 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 50848 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 49280 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 52416 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 52416 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 53984 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 54992 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 53424 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform -1 0 55552 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 48272 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 52752 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 54992 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 52416 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 50064 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 46704 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 52416 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 44800 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 49616 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 51968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 51184 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 51856 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 53424 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 54208 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 2800 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 3248 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 3024 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 3808 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 4592 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 3024 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 2912 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4592 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 4480 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 7056 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 8624 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 6720 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 7728 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 8512 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 10192 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 8288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 9296 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 15792 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 12768 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 16016 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 11760 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 12432 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 14224 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 22960 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 21616 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 23184 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 25312 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 16688 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 17808 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 18256 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 19824 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform 1 0 47040 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  S_term_single_106
timestamp 1486834041
transform -1 0 25760 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 53984 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 57344 0 57456 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 57344 4480 57456 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 57344 4928 57456 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 57344 5376 57456 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 57344 5824 57456 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 57344 6272 57456 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 57344 6720 57456 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 57344 7168 57456 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 57344 7616 57456 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 57344 8064 57456 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 57344 8512 57456 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 57344 448 57456 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 57344 8960 57456 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 57344 9408 57456 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 57344 9856 57456 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 57344 10304 57456 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 57344 10752 57456 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 57344 11200 57456 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 57344 11648 57456 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 57344 12096 57456 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 57344 12544 57456 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 57344 12992 57456 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 57344 896 57456 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 57344 13440 57456 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 57344 13888 57456 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 57344 1344 57456 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 57344 1792 57456 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 57344 2240 57456 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 57344 2688 57456 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 57344 3136 57456 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 57344 3584 57456 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 57344 4032 57456 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 4480 0 4592 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 31360 0 31472 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 34048 0 34160 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 36736 0 36848 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 39424 0 39536 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 42112 0 42224 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 44800 0 44912 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 47488 0 47600 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 50176 0 50288 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 52864 0 52976 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 55552 0 55664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 7168 0 7280 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 9856 0 9968 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 12544 0 12656 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 15232 0 15344 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 17920 0 18032 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 20608 0 20720 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 23296 0 23408 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 25984 0 26096 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 28672 0 28784 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 48160 14112 48272 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 52640 14112 52752 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 53088 14112 53200 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 53536 14112 53648 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 53984 14112 54096 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 54432 14112 54544 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 54880 14112 54992 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 55328 14112 55440 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 55776 14112 55888 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 56224 14112 56336 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 56672 14112 56784 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 48608 14112 48720 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 49056 14112 49168 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 49504 14112 49616 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 49952 14112 50064 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 50400 14112 50512 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 50848 14112 50960 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 51296 14112 51408 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 51744 14112 51856 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 52192 14112 52304 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 672 14112 784 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal2 s 1120 14112 1232 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal2 s 1568 14112 1680 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal2 s 2016 14112 2128 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal2 s 2464 14112 2576 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal2 s 2912 14112 3024 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal2 s 3360 14112 3472 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal2 s 3808 14112 3920 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal2 s 4256 14112 4368 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal2 s 4704 14112 4816 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal2 s 5152 14112 5264 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal2 s 5600 14112 5712 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal2 s 6048 14112 6160 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal2 s 6496 14112 6608 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal2 s 6944 14112 7056 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal2 s 7392 14112 7504 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal2 s 7840 14112 7952 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal2 s 8288 14112 8400 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal2 s 8736 14112 8848 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal2 s 9184 14112 9296 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal2 s 9632 14112 9744 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal2 s 10080 14112 10192 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal2 s 10528 14112 10640 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal2 s 10976 14112 11088 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal2 s 11424 14112 11536 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal2 s 11872 14112 11984 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal2 s 40544 14112 40656 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal2 s 45024 14112 45136 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal2 s 45472 14112 45584 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal2 s 45920 14112 46032 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal2 s 46368 14112 46480 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal2 s 46816 14112 46928 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal2 s 47264 14112 47376 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal2 s 40992 14112 41104 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal2 s 41440 14112 41552 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal2 s 41888 14112 42000 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal2 s 42336 14112 42448 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal2 s 42784 14112 42896 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal2 s 43232 14112 43344 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal2 s 43680 14112 43792 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal2 s 44128 14112 44240 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal2 s 44576 14112 44688 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal2 s 1792 0 1904 112 0 FreeSans 448 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 47712 14112 47824 14224 0 FreeSans 448 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
rlabel metal1 28728 12544 28728 12544 0 VDD
rlabel metal1 28728 13328 28728 13328 0 VSS
rlabel metal3 630 56 630 56 0 FrameData[0]
rlabel metal3 742 4536 742 4536 0 FrameData[10]
rlabel metal4 15176 5400 15176 5400 0 FrameData[11]
rlabel metal3 854 5432 854 5432 0 FrameData[12]
rlabel metal3 1694 5880 1694 5880 0 FrameData[13]
rlabel metal3 742 6328 742 6328 0 FrameData[14]
rlabel metal2 17080 8400 17080 8400 0 FrameData[15]
rlabel metal3 854 7224 854 7224 0 FrameData[16]
rlabel metal3 630 7672 630 7672 0 FrameData[17]
rlabel metal3 1694 8120 1694 8120 0 FrameData[18]
rlabel metal3 686 8568 686 8568 0 FrameData[19]
rlabel metal3 1246 504 1246 504 0 FrameData[1]
rlabel metal2 52360 4760 52360 4760 0 FrameData[20]
rlabel metal3 630 9464 630 9464 0 FrameData[21]
rlabel metal3 126 9912 126 9912 0 FrameData[22]
rlabel metal3 1470 10360 1470 10360 0 FrameData[23]
rlabel metal3 854 10808 854 10808 0 FrameData[24]
rlabel metal2 896 8344 896 8344 0 FrameData[25]
rlabel metal2 20216 12656 20216 12656 0 FrameData[26]
rlabel metal3 350 12152 350 12152 0 FrameData[27]
rlabel metal3 294 12600 294 12600 0 FrameData[28]
rlabel metal3 238 13048 238 13048 0 FrameData[29]
rlabel metal3 518 952 518 952 0 FrameData[2]
rlabel metal3 574 13496 574 13496 0 FrameData[30]
rlabel metal3 40096 3304 40096 3304 0 FrameData[31]
rlabel metal3 1302 1400 1302 1400 0 FrameData[3]
rlabel metal3 574 1848 574 1848 0 FrameData[4]
rlabel metal3 574 2296 574 2296 0 FrameData[5]
rlabel metal3 518 2744 518 2744 0 FrameData[6]
rlabel metal3 854 3192 854 3192 0 FrameData[7]
rlabel metal2 54488 8120 54488 8120 0 FrameData[8]
rlabel metal3 1694 4088 1694 4088 0 FrameData[9]
rlabel metal3 56938 56 56938 56 0 FrameData_O[0]
rlabel metal3 55986 4536 55986 4536 0 FrameData_O[10]
rlabel metal3 55188 5096 55188 5096 0 FrameData_O[11]
rlabel metal2 56168 4984 56168 4984 0 FrameData_O[12]
rlabel metal2 54600 5936 54600 5936 0 FrameData_O[13]
rlabel metal2 55160 6384 55160 6384 0 FrameData_O[14]
rlabel metal2 56168 6440 56168 6440 0 FrameData_O[15]
rlabel metal2 54600 7392 54600 7392 0 FrameData_O[16]
rlabel metal3 56770 7672 56770 7672 0 FrameData_O[17]
rlabel metal3 56658 8120 56658 8120 0 FrameData_O[18]
rlabel metal2 54376 8736 54376 8736 0 FrameData_O[19]
rlabel metal3 57106 504 57106 504 0 FrameData_O[1]
rlabel metal3 56770 9016 56770 9016 0 FrameData_O[20]
rlabel metal2 55160 9520 55160 9520 0 FrameData_O[21]
rlabel metal2 54600 10416 54600 10416 0 FrameData_O[22]
rlabel metal3 55328 8120 55328 8120 0 FrameData_O[23]
rlabel metal3 57050 10808 57050 10808 0 FrameData_O[24]
rlabel metal3 54544 8344 54544 8344 0 FrameData_O[25]
rlabel metal2 49224 11480 49224 11480 0 FrameData_O[26]
rlabel metal2 53032 7784 53032 7784 0 FrameData_O[27]
rlabel metal3 53088 10584 53088 10584 0 FrameData_O[28]
rlabel metal3 57162 13048 57162 13048 0 FrameData_O[29]
rlabel metal2 52024 1120 52024 1120 0 FrameData_O[2]
rlabel metal2 54712 11648 54712 11648 0 FrameData_O[30]
rlabel metal2 51240 9296 51240 9296 0 FrameData_O[31]
rlabel metal3 55482 1400 55482 1400 0 FrameData_O[3]
rlabel metal3 55482 1848 55482 1848 0 FrameData_O[4]
rlabel metal2 54936 2184 54936 2184 0 FrameData_O[5]
rlabel metal2 56168 2072 56168 2072 0 FrameData_O[6]
rlabel metal2 54600 3080 54600 3080 0 FrameData_O[7]
rlabel metal2 54824 3696 54824 3696 0 FrameData_O[8]
rlabel metal2 56168 3528 56168 3528 0 FrameData_O[9]
rlabel metal2 4536 238 4536 238 0 FrameStrobe[0]
rlabel metal2 31416 686 31416 686 0 FrameStrobe[10]
rlabel metal2 34104 1022 34104 1022 0 FrameStrobe[11]
rlabel metal3 34552 4536 34552 4536 0 FrameStrobe[12]
rlabel metal2 39480 686 39480 686 0 FrameStrobe[13]
rlabel metal2 42168 1722 42168 1722 0 FrameStrobe[14]
rlabel metal3 21896 1680 21896 1680 0 FrameStrobe[15]
rlabel metal2 51464 2856 51464 2856 0 FrameStrobe[16]
rlabel metal2 50008 4200 50008 4200 0 FrameStrobe[17]
rlabel metal2 52920 126 52920 126 0 FrameStrobe[18]
rlabel metal2 55608 182 55608 182 0 FrameStrobe[19]
rlabel metal2 7224 854 7224 854 0 FrameStrobe[1]
rlabel metal3 10192 3528 10192 3528 0 FrameStrobe[2]
rlabel metal2 15176 5600 15176 5600 0 FrameStrobe[3]
rlabel metal2 15232 3528 15232 3528 0 FrameStrobe[4]
rlabel metal2 16520 6720 16520 6720 0 FrameStrobe[5]
rlabel metal2 20664 630 20664 630 0 FrameStrobe[6]
rlabel metal2 2016 4536 2016 4536 0 FrameStrobe[7]
rlabel metal2 26040 182 26040 182 0 FrameStrobe[8]
rlabel metal2 20048 6888 20048 6888 0 FrameStrobe[9]
rlabel metal2 48216 13650 48216 13650 0 FrameStrobe_O[0]
rlabel metal2 52696 13538 52696 13538 0 FrameStrobe_O[10]
rlabel metal2 53144 13762 53144 13762 0 FrameStrobe_O[11]
rlabel metal2 53648 9688 53648 9688 0 FrameStrobe_O[12]
rlabel metal3 53536 9240 53536 9240 0 FrameStrobe_O[13]
rlabel metal2 51240 11312 51240 11312 0 FrameStrobe_O[14]
rlabel metal2 54936 13874 54936 13874 0 FrameStrobe_O[15]
rlabel metal2 55384 13034 55384 13034 0 FrameStrobe_O[16]
rlabel metal2 53648 6552 53648 6552 0 FrameStrobe_O[17]
rlabel metal2 56280 13482 56280 13482 0 FrameStrobe_O[18]
rlabel metal3 53480 6104 53480 6104 0 FrameStrobe_O[19]
rlabel metal2 48664 13258 48664 13258 0 FrameStrobe_O[1]
rlabel metal2 51128 13328 51128 13328 0 FrameStrobe_O[2]
rlabel metal3 49952 11592 49952 11592 0 FrameStrobe_O[3]
rlabel metal2 50008 13594 50008 13594 0 FrameStrobe_O[4]
rlabel metal2 50456 13258 50456 13258 0 FrameStrobe_O[5]
rlabel metal2 50904 12866 50904 12866 0 FrameStrobe_O[6]
rlabel metal2 51352 13202 51352 13202 0 FrameStrobe_O[7]
rlabel metal2 51800 13706 51800 13706 0 FrameStrobe_O[8]
rlabel metal2 52248 13650 52248 13650 0 FrameStrobe_O[9]
rlabel metal2 728 12698 728 12698 0 N1BEG[0]
rlabel metal2 1736 10360 1736 10360 0 N1BEG[1]
rlabel metal2 1624 13034 1624 13034 0 N1BEG[2]
rlabel metal2 2184 11256 2184 11256 0 N1BEG[3]
rlabel metal2 2520 13650 2520 13650 0 N2BEG[0]
rlabel metal2 2968 13034 2968 13034 0 N2BEG[1]
rlabel metal2 3416 13258 3416 13258 0 N2BEG[2]
rlabel metal2 3864 13426 3864 13426 0 N2BEG[3]
rlabel metal2 2184 13216 2184 13216 0 N2BEG[4]
rlabel metal2 4760 13818 4760 13818 0 N2BEG[5]
rlabel metal3 4928 11592 4928 11592 0 N2BEG[6]
rlabel metal2 5656 13650 5656 13650 0 N2BEG[7]
rlabel metal2 6104 12418 6104 12418 0 N2BEGb[0]
rlabel metal2 6216 12376 6216 12376 0 N2BEGb[1]
rlabel metal2 7448 11704 7448 11704 0 N2BEGb[2]
rlabel metal2 5992 13216 5992 13216 0 N2BEGb[3]
rlabel metal2 7896 13258 7896 13258 0 N2BEGb[4]
rlabel metal2 7784 11872 7784 11872 0 N2BEGb[5]
rlabel metal2 8904 10808 8904 10808 0 N2BEGb[6]
rlabel metal3 8400 13160 8400 13160 0 N2BEGb[7]
rlabel metal2 9688 13258 9688 13258 0 N4BEG[0]
rlabel metal3 14392 10808 14392 10808 0 N4BEG[10]
rlabel metal3 14280 12824 14280 12824 0 N4BEG[11]
rlabel metal2 15064 13258 15064 13258 0 N4BEG[12]
rlabel metal2 15512 12866 15512 12866 0 N4BEG[13]
rlabel metal2 15960 13202 15960 13202 0 N4BEG[14]
rlabel metal2 16408 13594 16408 13594 0 N4BEG[15]
rlabel metal2 10584 11480 10584 11480 0 N4BEG[1]
rlabel metal2 10584 13258 10584 13258 0 N4BEG[2]
rlabel metal2 10976 11592 10976 11592 0 N4BEG[3]
rlabel metal3 10640 13160 10640 13160 0 N4BEG[4]
rlabel metal2 11928 13762 11928 13762 0 N4BEG[5]
rlabel metal2 12376 12698 12376 12698 0 N4BEG[6]
rlabel metal2 12992 10808 12992 10808 0 N4BEG[7]
rlabel metal2 11368 13272 11368 13272 0 N4BEG[8]
rlabel metal2 13720 12866 13720 12866 0 N4BEG[9]
rlabel metal2 16800 12376 16800 12376 0 NN4BEG[0]
rlabel metal2 21336 12698 21336 12698 0 NN4BEG[10]
rlabel metal3 21504 13160 21504 13160 0 NN4BEG[11]
rlabel metal2 22232 13258 22232 13258 0 NN4BEG[12]
rlabel metal2 22680 13650 22680 13650 0 NN4BEG[13]
rlabel metal2 23128 13258 23128 13258 0 NN4BEG[14]
rlabel metal2 23576 13818 23576 13818 0 NN4BEG[15]
rlabel metal2 17304 13538 17304 13538 0 NN4BEG[1]
rlabel metal2 17752 13258 17752 13258 0 NN4BEG[2]
rlabel metal2 18200 13202 18200 13202 0 NN4BEG[3]
rlabel metal3 18088 13048 18088 13048 0 NN4BEG[4]
rlabel metal2 19096 12698 19096 12698 0 NN4BEG[5]
rlabel metal2 19544 13202 19544 13202 0 NN4BEG[6]
rlabel metal3 19656 12824 19656 12824 0 NN4BEG[7]
rlabel metal2 20440 12866 20440 12866 0 NN4BEG[8]
rlabel metal2 20888 13202 20888 13202 0 NN4BEG[9]
rlabel metal2 24472 13818 24472 13818 0 S1END[0]
rlabel metal2 24920 13762 24920 13762 0 S1END[1]
rlabel metal2 25368 12306 25368 12306 0 S1END[2]
rlabel metal2 53256 4256 53256 4256 0 S1END[3]
rlabel metal2 41608 7168 41608 7168 0 S2END[0]
rlabel metal2 51688 2408 51688 2408 0 S2END[1]
rlabel metal2 52248 5712 52248 5712 0 S2END[2]
rlabel metal2 31192 13034 31192 13034 0 S2END[3]
rlabel metal2 31640 12922 31640 12922 0 S2END[4]
rlabel metal2 24696 2744 24696 2744 0 S2END[5]
rlabel metal2 32536 12978 32536 12978 0 S2END[6]
rlabel metal2 25592 8344 25592 8344 0 S2END[7]
rlabel metal2 26264 12698 26264 12698 0 S2MID[0]
rlabel metal2 26712 13762 26712 13762 0 S2MID[1]
rlabel metal2 37688 11032 37688 11032 0 S2MID[2]
rlabel metal3 34608 3304 34608 3304 0 S2MID[3]
rlabel metal2 28056 12978 28056 12978 0 S2MID[4]
rlabel metal2 50456 10976 50456 10976 0 S2MID[5]
rlabel metal2 39816 7112 39816 7112 0 S2MID[6]
rlabel metal2 51800 7224 51800 7224 0 S2MID[7]
rlabel metal2 25144 5376 25144 5376 0 S4END[0]
rlabel metal2 37912 13034 37912 13034 0 S4END[10]
rlabel metal2 46424 12600 46424 12600 0 S4END[11]
rlabel metal2 33208 9856 33208 9856 0 S4END[12]
rlabel metal2 39256 10906 39256 10906 0 S4END[13]
rlabel metal2 26824 8512 26824 8512 0 S4END[14]
rlabel metal3 26600 10080 26600 10080 0 S4END[15]
rlabel metal2 24248 5824 24248 5824 0 S4END[1]
rlabel metal3 21000 8400 21000 8400 0 S4END[2]
rlabel metal2 17640 11872 17640 11872 0 S4END[3]
rlabel metal2 15512 8904 15512 8904 0 S4END[4]
rlabel metal3 22848 1400 22848 1400 0 S4END[5]
rlabel metal3 18984 3024 18984 3024 0 S4END[6]
rlabel metal2 50904 7616 50904 7616 0 S4END[7]
rlabel metal2 19432 9800 19432 9800 0 S4END[8]
rlabel metal2 42504 10920 42504 10920 0 S4END[9]
rlabel metal2 26152 10752 26152 10752 0 SS4END[0]
rlabel metal4 15288 7952 15288 7952 0 SS4END[10]
rlabel metal2 15736 2436 15736 2436 0 SS4END[11]
rlabel metal2 3304 1680 3304 1680 0 SS4END[12]
rlabel metal4 21000 13776 21000 13776 0 SS4END[13]
rlabel metal3 21000 5600 21000 5600 0 SS4END[14]
rlabel metal3 43176 3024 43176 3024 0 SS4END[15]
rlabel metal2 16072 10808 16072 10808 0 SS4END[1]
rlabel metal3 21952 3192 21952 3192 0 SS4END[2]
rlabel metal3 21000 840 21000 840 0 SS4END[3]
rlabel metal2 42392 11130 42392 11130 0 SS4END[4]
rlabel metal2 42840 13426 42840 13426 0 SS4END[5]
rlabel metal2 21896 6832 21896 6832 0 SS4END[6]
rlabel metal2 25592 2072 25592 2072 0 SS4END[7]
rlabel metal2 24472 11144 24472 11144 0 SS4END[8]
rlabel metal4 15512 5417 15512 5417 0 SS4END[9]
rlabel metal3 1568 9800 1568 9800 0 UserCLK
rlabel metal2 47656 11592 47656 11592 0 UserCLKo
rlabel metal3 50792 2744 50792 2744 0 net1
rlabel metal2 55272 9296 55272 9296 0 net10
rlabel metal2 18648 12040 18648 12040 0 net100
rlabel metal2 18872 12880 18872 12880 0 net101
rlabel metal2 2968 9352 2968 9352 0 net102
rlabel metal2 16856 6664 16856 6664 0 net103
rlabel metal2 21112 10752 21112 10752 0 net104
rlabel metal2 1512 7504 1512 7504 0 net105
rlabel metal3 24752 13160 24752 13160 0 net106
rlabel metal2 53368 6272 53368 6272 0 net11
rlabel metal2 52584 4872 52584 4872 0 net12
rlabel metal3 54152 5208 54152 5208 0 net13
rlabel metal2 54264 6048 54264 6048 0 net14
rlabel metal2 53480 9632 53480 9632 0 net15
rlabel metal2 54152 7784 54152 7784 0 net16
rlabel metal2 51128 5768 51128 5768 0 net17
rlabel metal2 52584 7616 52584 7616 0 net18
rlabel metal3 41944 10080 41944 10080 0 net19
rlabel metal3 47936 4200 47936 4200 0 net2
rlabel metal2 52136 7112 52136 7112 0 net20
rlabel metal3 50008 8232 50008 8232 0 net21
rlabel metal2 22120 3584 22120 3584 0 net22
rlabel metal3 50708 1176 50708 1176 0 net23
rlabel metal2 45528 11424 45528 11424 0 net24
rlabel metal2 49952 4424 49952 4424 0 net25
rlabel metal2 52584 1344 52584 1344 0 net26
rlabel metal3 50120 2072 50120 2072 0 net27
rlabel metal2 54152 2240 54152 2240 0 net28
rlabel metal2 55160 1400 55160 1400 0 net29
rlabel metal3 52920 6440 52920 6440 0 net3
rlabel metal2 53592 2968 53592 2968 0 net30
rlabel metal2 55104 3528 55104 3528 0 net31
rlabel metal2 55160 2912 55160 2912 0 net32
rlabel metal3 19544 6776 19544 6776 0 net33
rlabel metal2 52920 10640 52920 10640 0 net34
rlabel metal2 52360 2408 52360 2408 0 net35
rlabel metal2 52528 9800 52528 9800 0 net36
rlabel metal2 52136 8848 52136 8848 0 net37
rlabel metal3 43624 10472 43624 10472 0 net38
rlabel metal4 41832 1400 41832 1400 0 net39
rlabel metal3 52472 3696 52472 3696 0 net4
rlabel metal2 48664 7616 48664 7616 0 net40
rlabel metal2 52696 7784 52696 7784 0 net41
rlabel metal2 20776 6608 20776 6608 0 net42
rlabel metal2 52136 5600 52136 5600 0 net43
rlabel metal2 18424 1400 18424 1400 0 net44
rlabel metal2 50456 5964 50456 5964 0 net45
rlabel metal2 18816 952 18816 952 0 net46
rlabel metal2 52360 11088 52360 11088 0 net47
rlabel metal2 52248 10808 52248 10808 0 net48
rlabel metal2 51352 11088 51352 11088 0 net49
rlabel metal4 35336 5880 35336 5880 0 net5
rlabel metal2 52136 10360 52136 10360 0 net50
rlabel metal2 53592 11704 53592 11704 0 net51
rlabel metal2 54376 12096 54376 12096 0 net52
rlabel metal4 2296 5544 2296 5544 0 net53
rlabel metal2 15512 1568 15512 1568 0 net54
rlabel metal2 3080 9520 3080 9520 0 net55
rlabel metal4 2856 6888 2856 6888 0 net56
rlabel metal3 44856 2520 44856 2520 0 net57
rlabel metal2 16184 12264 16184 12264 0 net58
rlabel metal2 2744 7840 2744 7840 0 net59
rlabel metal3 52276 6664 52276 6664 0 net6
rlabel metal2 19880 10584 19880 10584 0 net60
rlabel metal2 2576 4760 2576 4760 0 net61
rlabel metal4 15400 1915 15400 1915 0 net62
rlabel metal4 15848 3330 15848 3330 0 net63
rlabel metal2 18424 8848 18424 8848 0 net64
rlabel metal3 12376 8960 12376 8960 0 net65
rlabel metal3 13496 8064 13496 8064 0 net66
rlabel metal3 11424 1624 11424 1624 0 net67
rlabel metal4 20552 14056 20552 14056 0 net68
rlabel metal4 13720 5488 13720 5488 0 net69
rlabel metal3 53816 5824 53816 5824 0 net7
rlabel metal2 52696 4480 52696 4480 0 net70
rlabel metal2 52248 3696 52248 3696 0 net71
rlabel metal2 16520 11144 16520 11144 0 net72
rlabel metal2 19992 8008 19992 8008 0 net73
rlabel metal2 19656 7224 19656 7224 0 net74
rlabel metal2 9464 11424 9464 11424 0 net75
rlabel metal3 16128 9912 16128 9912 0 net76
rlabel metal2 14392 8680 14392 8680 0 net77
rlabel metal2 15512 5432 15512 5432 0 net78
rlabel metal3 20664 8232 20664 8232 0 net79
rlabel metal2 50568 3752 50568 3752 0 net8
rlabel metal2 20328 9520 20328 9520 0 net80
rlabel metal4 25032 2296 25032 2296 0 net81
rlabel metal2 24024 3696 24024 3696 0 net82
rlabel metal2 16632 7392 16632 7392 0 net83
rlabel metal2 23688 4592 23688 4592 0 net84
rlabel metal2 22064 2296 22064 2296 0 net85
rlabel metal2 14112 7560 14112 7560 0 net86
rlabel metal3 16520 11872 16520 11872 0 net87
rlabel metal2 13552 5992 13552 5992 0 net88
rlabel metal2 3976 5432 3976 5432 0 net89
rlabel metal2 55160 7112 55160 7112 0 net9
rlabel metal2 22792 10864 22792 10864 0 net90
rlabel metal2 21784 12880 21784 12880 0 net91
rlabel metal2 2072 6804 2072 6804 0 net92
rlabel metal3 18648 12880 18648 12880 0 net93
rlabel metal4 15288 5843 15288 5843 0 net94
rlabel metal2 25592 11424 25592 11424 0 net95
rlabel metal2 16856 10976 16856 10976 0 net96
rlabel metal2 1960 3136 1960 3136 0 net97
rlabel metal3 16800 12040 16800 12040 0 net98
rlabel metal2 16968 12712 16968 12712 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 14224
<< end >>
