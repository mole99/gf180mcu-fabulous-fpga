magic
tech gf180mcuD
magscale 1 5
timestamp 1764971535
<< metal1 >>
rect 336 6677 15512 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 15512 6677
rect 336 6634 15512 6651
rect 6735 6593 6761 6599
rect 1185 6567 1191 6593
rect 1217 6567 1223 6593
rect 6735 6561 6761 6567
rect 7519 6593 7545 6599
rect 7519 6561 7545 6567
rect 8135 6537 8161 6543
rect 8135 6505 8161 6511
rect 1359 6481 1385 6487
rect 9423 6481 9449 6487
rect 2137 6455 2143 6481
rect 2169 6455 2175 6481
rect 3089 6455 3095 6481
rect 3121 6455 3127 6481
rect 3873 6455 3879 6481
rect 3905 6455 3911 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 5329 6455 5335 6481
rect 5361 6455 5367 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 7233 6455 7239 6481
rect 7265 6455 7271 6481
rect 9193 6455 9199 6481
rect 9225 6455 9231 6481
rect 10593 6455 10599 6481
rect 10625 6455 10631 6481
rect 11321 6455 11327 6481
rect 11353 6455 11359 6481
rect 12553 6455 12559 6481
rect 12585 6455 12591 6481
rect 13393 6455 13399 6481
rect 13425 6455 13431 6481
rect 14513 6455 14519 6481
rect 14545 6455 14551 6481
rect 1359 6449 1385 6455
rect 9423 6449 9449 6455
rect 2591 6425 2617 6431
rect 1801 6399 1807 6425
rect 1833 6399 1839 6425
rect 2591 6393 2617 6399
rect 3375 6425 3401 6431
rect 3375 6393 3401 6399
rect 4663 6425 4689 6431
rect 4663 6393 4689 6399
rect 5839 6425 5865 6431
rect 8751 6425 8777 6431
rect 8353 6399 8359 6425
rect 8385 6399 8391 6425
rect 5839 6393 5865 6399
rect 8751 6393 8777 6399
rect 9703 6425 9729 6431
rect 9703 6393 9729 6399
rect 10151 6425 10177 6431
rect 10151 6393 10177 6399
rect 10935 6425 10961 6431
rect 10935 6393 10961 6399
rect 12111 6425 12137 6431
rect 12111 6393 12137 6399
rect 12895 6425 12921 6431
rect 12895 6393 12921 6399
rect 14127 6425 14153 6431
rect 14127 6393 14153 6399
rect 336 6285 15512 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 15512 6285
rect 336 6242 15512 6259
rect 4047 6201 4073 6207
rect 4047 6169 4073 6175
rect 5559 6201 5585 6207
rect 5559 6169 5585 6175
rect 8079 6201 8105 6207
rect 8079 6169 8105 6175
rect 11439 6201 11465 6207
rect 11439 6169 11465 6175
rect 13455 6201 13481 6207
rect 13455 6169 13481 6175
rect 13063 6145 13089 6151
rect 7513 6119 7519 6145
rect 7545 6119 7551 6145
rect 9473 6119 9479 6145
rect 9505 6119 9511 6145
rect 15129 6119 15135 6145
rect 15161 6119 15167 6145
rect 13063 6113 13089 6119
rect 7295 6089 7321 6095
rect 7295 6057 7321 6063
rect 8751 6089 8777 6095
rect 8751 6057 8777 6063
rect 9031 6089 9057 6095
rect 12609 6063 12615 6089
rect 12641 6063 12647 6089
rect 9031 6057 9057 6063
rect 4545 6007 4551 6033
rect 4577 6007 4583 6033
rect 5273 6007 5279 6033
rect 5305 6007 5311 6033
rect 8577 6007 8583 6033
rect 8609 6007 8615 6033
rect 9921 6007 9927 6033
rect 9953 6007 9959 6033
rect 11937 6007 11943 6033
rect 11969 6007 11975 6033
rect 13953 6007 13959 6033
rect 13985 6007 13991 6033
rect 14681 6007 14687 6033
rect 14713 6007 14719 6033
rect 336 5893 15512 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 15512 5893
rect 336 5850 15512 5867
rect 7071 5753 7097 5759
rect 13337 5727 13343 5753
rect 13369 5727 13375 5753
rect 7071 5721 7097 5727
rect 6791 5697 6817 5703
rect 6791 5665 6817 5671
rect 7239 5697 7265 5703
rect 7239 5665 7265 5671
rect 7687 5697 7713 5703
rect 7687 5665 7713 5671
rect 8471 5697 8497 5703
rect 8471 5665 8497 5671
rect 8751 5697 8777 5703
rect 12329 5671 12335 5697
rect 12361 5671 12367 5697
rect 13729 5671 13735 5697
rect 13761 5671 13767 5697
rect 14009 5671 14015 5697
rect 14041 5671 14047 5697
rect 14681 5671 14687 5697
rect 14713 5671 14719 5697
rect 8751 5665 8777 5671
rect 7519 5641 7545 5647
rect 7519 5609 7545 5615
rect 7967 5641 7993 5647
rect 7967 5609 7993 5615
rect 12839 5641 12865 5647
rect 12839 5609 12865 5615
rect 14407 5585 14433 5591
rect 14407 5553 14433 5559
rect 15191 5585 15217 5591
rect 15191 5553 15217 5559
rect 336 5501 15512 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 15512 5501
rect 336 5458 15512 5475
rect 13847 5417 13873 5423
rect 13847 5385 13873 5391
rect 8135 5305 8161 5311
rect 8135 5273 8161 5279
rect 8415 5305 8441 5311
rect 13337 5279 13343 5305
rect 13369 5279 13375 5305
rect 14737 5279 14743 5305
rect 14769 5279 14775 5305
rect 8415 5273 8441 5279
rect 8695 5249 8721 5255
rect 15073 5223 15079 5249
rect 15105 5223 15111 5249
rect 8695 5217 8721 5223
rect 7855 5193 7881 5199
rect 7855 5161 7881 5167
rect 336 5109 15512 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 15512 5109
rect 336 5066 15512 5083
rect 13505 4943 13511 4969
rect 13537 4943 13543 4969
rect 13897 4943 13903 4969
rect 13929 4943 13935 4969
rect 14289 4943 14295 4969
rect 14321 4943 14327 4969
rect 7351 4913 7377 4919
rect 7351 4881 7377 4887
rect 7631 4913 7657 4919
rect 7631 4881 7657 4887
rect 8471 4913 8497 4919
rect 13113 4887 13119 4913
rect 13145 4887 13151 4913
rect 14681 4887 14687 4913
rect 14713 4887 14719 4913
rect 8471 4881 8497 4887
rect 8751 4857 8777 4863
rect 8751 4825 8777 4831
rect 15191 4801 15217 4807
rect 15191 4769 15217 4775
rect 336 4717 15512 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 15512 4717
rect 336 4674 15512 4691
rect 5217 4551 5223 4577
rect 5249 4551 5255 4577
rect 7569 4551 7575 4577
rect 7601 4551 7607 4577
rect 13785 4551 13791 4577
rect 13817 4551 13823 4577
rect 5447 4521 5473 4527
rect 5447 4489 5473 4495
rect 8863 4521 8889 4527
rect 13337 4495 13343 4521
rect 13369 4495 13375 4521
rect 14681 4495 14687 4521
rect 14713 4495 14719 4521
rect 8863 4489 8889 4495
rect 15073 4439 15079 4465
rect 15105 4439 15111 4465
rect 7351 4409 7377 4415
rect 7351 4377 7377 4383
rect 8583 4409 8609 4415
rect 8583 4377 8609 4383
rect 336 4325 15512 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 15512 4325
rect 336 4282 15512 4299
rect 6567 4185 6593 4191
rect 6567 4153 6593 4159
rect 7743 4185 7769 4191
rect 7743 4153 7769 4159
rect 9535 4185 9561 4191
rect 9535 4153 9561 4159
rect 9983 4185 10009 4191
rect 9983 4153 10009 4159
rect 10431 4185 10457 4191
rect 10431 4153 10457 4159
rect 11439 4185 11465 4191
rect 11439 4153 11465 4159
rect 13623 4185 13649 4191
rect 13897 4159 13903 4185
rect 13929 4159 13935 4185
rect 13623 4153 13649 4159
rect 6847 4129 6873 4135
rect 6847 4097 6873 4103
rect 7183 4129 7209 4135
rect 7183 4097 7209 4103
rect 8023 4129 8049 4135
rect 8023 4097 8049 4103
rect 8471 4129 8497 4135
rect 8471 4097 8497 4103
rect 9815 4129 9841 4135
rect 10711 4129 10737 4135
rect 10201 4103 10207 4129
rect 10233 4103 10239 4129
rect 9815 4097 9841 4103
rect 10711 4097 10737 4103
rect 11719 4129 11745 4135
rect 11719 4097 11745 4103
rect 13343 4129 13369 4135
rect 14681 4103 14687 4129
rect 14713 4103 14719 4129
rect 13343 4097 13369 4103
rect 7463 4073 7489 4079
rect 7463 4041 7489 4047
rect 8751 4073 8777 4079
rect 14345 4047 14351 4073
rect 14377 4047 14383 4073
rect 8751 4041 8777 4047
rect 15191 4017 15217 4023
rect 15191 3985 15217 3991
rect 336 3933 15512 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 15512 3933
rect 336 3890 15512 3907
rect 8975 3793 9001 3799
rect 10711 3793 10737 3799
rect 4993 3767 4999 3793
rect 5025 3767 5031 3793
rect 5889 3767 5895 3793
rect 5921 3767 5927 3793
rect 7513 3767 7519 3793
rect 7545 3767 7551 3793
rect 9697 3767 9703 3793
rect 9729 3767 9735 3793
rect 8975 3761 9001 3767
rect 10711 3761 10737 3767
rect 11383 3793 11409 3799
rect 14457 3767 14463 3793
rect 14489 3767 14495 3793
rect 15129 3767 15135 3793
rect 15161 3767 15167 3793
rect 11383 3761 11409 3767
rect 5223 3737 5249 3743
rect 9193 3711 9199 3737
rect 9225 3711 9231 3737
rect 14289 3711 14295 3737
rect 14321 3711 14327 3737
rect 14793 3711 14799 3737
rect 14825 3711 14831 3737
rect 5223 3705 5249 3711
rect 9479 3681 9505 3687
rect 9479 3649 9505 3655
rect 6119 3625 6145 3631
rect 6119 3593 6145 3599
rect 7295 3625 7321 3631
rect 7295 3593 7321 3599
rect 10991 3625 11017 3631
rect 10991 3593 11017 3599
rect 11663 3625 11689 3631
rect 11663 3593 11689 3599
rect 336 3541 15512 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 15512 3541
rect 336 3498 15512 3515
rect 7743 3457 7769 3463
rect 7743 3425 7769 3431
rect 8919 3457 8945 3463
rect 8919 3425 8945 3431
rect 10151 3457 10177 3463
rect 10705 3431 10711 3457
rect 10737 3431 10743 3457
rect 10151 3425 10177 3431
rect 8415 3401 8441 3407
rect 8415 3369 8441 3375
rect 7015 3345 7041 3351
rect 7015 3313 7041 3319
rect 9703 3345 9729 3351
rect 9703 3313 9729 3319
rect 10879 3345 10905 3351
rect 10879 3313 10905 3319
rect 11159 3345 11185 3351
rect 11159 3313 11185 3319
rect 11439 3345 11465 3351
rect 11439 3313 11465 3319
rect 12335 3345 12361 3351
rect 13455 3345 13481 3351
rect 12553 3319 12559 3345
rect 12585 3319 12591 3345
rect 12335 3313 12361 3319
rect 13455 3313 13481 3319
rect 13735 3345 13761 3351
rect 13897 3319 13903 3345
rect 13929 3319 13935 3345
rect 14681 3319 14687 3345
rect 14713 3319 14719 3345
rect 13735 3313 13761 3319
rect 7295 3289 7321 3295
rect 8695 3289 8721 3295
rect 7961 3263 7967 3289
rect 7993 3263 7999 3289
rect 7295 3257 7321 3263
rect 8695 3257 8721 3263
rect 9199 3289 9225 3295
rect 10431 3289 10457 3295
rect 9921 3263 9927 3289
rect 9953 3263 9959 3289
rect 9199 3257 9225 3263
rect 10431 3257 10457 3263
rect 15191 3289 15217 3295
rect 15191 3257 15217 3263
rect 14407 3233 14433 3239
rect 14407 3201 14433 3207
rect 336 3149 15512 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 15512 3149
rect 336 3106 15512 3123
rect 12055 3009 12081 3015
rect 10593 2983 10599 3009
rect 10625 2983 10631 3009
rect 12055 2977 12081 2983
rect 13959 3009 13985 3015
rect 13959 2977 13985 2983
rect 14519 3009 14545 3015
rect 15129 2983 15135 3009
rect 15161 2983 15167 3009
rect 14519 2977 14545 2983
rect 7519 2953 7545 2959
rect 7519 2921 7545 2927
rect 8191 2953 8217 2959
rect 8191 2921 8217 2927
rect 9143 2953 9169 2959
rect 9143 2921 9169 2927
rect 9311 2953 9337 2959
rect 9311 2921 9337 2927
rect 9759 2953 9785 2959
rect 9759 2921 9785 2927
rect 10823 2953 10849 2959
rect 14289 2927 14295 2953
rect 14321 2927 14327 2953
rect 14681 2927 14687 2953
rect 14713 2927 14719 2953
rect 10823 2921 10849 2927
rect 7351 2897 7377 2903
rect 7351 2865 7377 2871
rect 7799 2897 7825 2903
rect 7799 2865 7825 2871
rect 8471 2897 8497 2903
rect 8471 2865 8497 2871
rect 9591 2897 9617 2903
rect 9591 2865 9617 2871
rect 10039 2897 10065 2903
rect 10039 2865 10065 2871
rect 11103 2897 11129 2903
rect 11103 2865 11129 2871
rect 7071 2841 7097 2847
rect 7071 2809 7097 2815
rect 8863 2841 8889 2847
rect 8863 2809 8889 2815
rect 10375 2841 10401 2847
rect 10375 2809 10401 2815
rect 12335 2841 12361 2847
rect 12335 2809 12361 2815
rect 13679 2841 13705 2847
rect 13679 2809 13705 2815
rect 336 2757 15512 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 15512 2757
rect 336 2714 15512 2731
rect 7351 2673 7377 2679
rect 7351 2641 7377 2647
rect 8471 2673 8497 2679
rect 8471 2641 8497 2647
rect 8919 2673 8945 2679
rect 8919 2641 8945 2647
rect 9367 2673 9393 2679
rect 9367 2641 9393 2647
rect 11439 2673 11465 2679
rect 11439 2641 11465 2647
rect 12279 2673 12305 2679
rect 12279 2641 12305 2647
rect 8751 2617 8777 2623
rect 12559 2617 12585 2623
rect 10481 2591 10487 2617
rect 10513 2591 10519 2617
rect 11265 2591 11271 2617
rect 11297 2591 11303 2617
rect 13897 2591 13903 2617
rect 13929 2591 13935 2617
rect 15073 2591 15079 2617
rect 15105 2591 15111 2617
rect 8751 2585 8777 2591
rect 12559 2585 12585 2591
rect 6847 2561 6873 2567
rect 6847 2529 6873 2535
rect 7799 2561 7825 2567
rect 7799 2529 7825 2535
rect 11719 2561 11745 2567
rect 14737 2535 14743 2561
rect 14769 2535 14775 2561
rect 11719 2529 11745 2535
rect 7127 2505 7153 2511
rect 9199 2505 9225 2511
rect 7569 2479 7575 2505
rect 7601 2479 7607 2505
rect 8017 2479 8023 2505
rect 8049 2479 8055 2505
rect 7127 2473 7153 2479
rect 9199 2473 9225 2479
rect 9647 2505 9673 2511
rect 9647 2473 9673 2479
rect 14407 2505 14433 2511
rect 14407 2473 14433 2479
rect 9983 2449 10009 2455
rect 9983 2417 10009 2423
rect 10767 2449 10793 2455
rect 10767 2417 10793 2423
rect 336 2365 15512 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 15512 2365
rect 336 2322 15512 2339
rect 8359 2225 8385 2231
rect 10481 2199 10487 2225
rect 10513 2199 10519 2225
rect 11377 2199 11383 2225
rect 11409 2199 11415 2225
rect 12553 2199 12559 2225
rect 12585 2199 12591 2225
rect 15129 2199 15135 2225
rect 15161 2199 15167 2225
rect 8359 2193 8385 2199
rect 8079 2169 8105 2175
rect 5889 2143 5895 2169
rect 5921 2143 5927 2169
rect 7289 2143 7295 2169
rect 7321 2143 7327 2169
rect 9305 2143 9311 2169
rect 9337 2143 9343 2169
rect 10873 2143 10879 2169
rect 10905 2143 10911 2169
rect 14681 2143 14687 2169
rect 14713 2143 14719 2169
rect 8079 2137 8105 2143
rect 5503 2113 5529 2119
rect 5503 2081 5529 2087
rect 6119 2113 6145 2119
rect 8863 2113 8889 2119
rect 12167 2113 12193 2119
rect 6505 2087 6511 2113
rect 6537 2087 6543 2113
rect 11713 2087 11719 2113
rect 11745 2087 11751 2113
rect 6119 2081 6145 2087
rect 8863 2081 8889 2087
rect 12167 2081 12193 2087
rect 5223 2057 5249 2063
rect 5223 2025 5249 2031
rect 6791 2057 6817 2063
rect 6791 2025 6817 2031
rect 7575 2057 7601 2063
rect 7575 2025 7601 2031
rect 8583 2057 8609 2063
rect 8583 2025 8609 2031
rect 9479 2057 9505 2063
rect 9479 2025 9505 2031
rect 11887 2057 11913 2063
rect 11887 2025 11913 2031
rect 12335 2057 12361 2063
rect 12335 2025 12361 2031
rect 336 1973 15512 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 15512 1973
rect 336 1930 15512 1947
rect 6231 1889 6257 1895
rect 6231 1857 6257 1863
rect 6511 1833 6537 1839
rect 9641 1807 9647 1833
rect 9673 1807 9679 1833
rect 11209 1807 11215 1833
rect 11241 1807 11247 1833
rect 13113 1807 13119 1833
rect 13145 1807 13151 1833
rect 14289 1807 14295 1833
rect 14321 1807 14327 1833
rect 6511 1801 6537 1807
rect 4775 1777 4801 1783
rect 4775 1745 4801 1751
rect 5783 1777 5809 1783
rect 12279 1777 12305 1783
rect 6729 1751 6735 1777
rect 6761 1751 6767 1777
rect 7457 1751 7463 1777
rect 7489 1751 7495 1777
rect 8409 1751 8415 1777
rect 8441 1751 8447 1777
rect 9473 1751 9479 1777
rect 9505 1751 9511 1777
rect 11041 1751 11047 1777
rect 11073 1751 11079 1777
rect 13897 1751 13903 1777
rect 13929 1751 13935 1777
rect 14737 1751 14743 1777
rect 14769 1751 14775 1777
rect 5783 1745 5809 1751
rect 12279 1745 12305 1751
rect 6063 1721 6089 1727
rect 8639 1721 8665 1727
rect 4993 1695 4999 1721
rect 5025 1695 5031 1721
rect 7065 1695 7071 1721
rect 7097 1695 7103 1721
rect 6063 1689 6089 1695
rect 8639 1689 8665 1695
rect 12559 1721 12585 1727
rect 15191 1721 15217 1727
rect 13561 1695 13567 1721
rect 13593 1695 13599 1721
rect 12559 1689 12585 1695
rect 15191 1689 15217 1695
rect 7743 1665 7769 1671
rect 7743 1633 7769 1639
rect 8975 1665 9001 1671
rect 8975 1633 9001 1639
rect 9927 1665 9953 1671
rect 9927 1633 9953 1639
rect 10543 1665 10569 1671
rect 10543 1633 10569 1639
rect 11719 1665 11745 1671
rect 11719 1633 11745 1639
rect 336 1581 15512 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 15512 1581
rect 336 1538 15512 1555
rect 13847 1441 13873 1447
rect 3369 1415 3375 1441
rect 3401 1415 3407 1441
rect 15129 1415 15135 1441
rect 15161 1415 15167 1441
rect 13847 1409 13873 1415
rect 5889 1359 5895 1385
rect 5921 1359 5927 1385
rect 7401 1359 7407 1385
rect 7433 1359 7439 1385
rect 8185 1359 8191 1385
rect 8217 1359 8223 1385
rect 9585 1359 9591 1385
rect 9617 1359 9623 1385
rect 11881 1359 11887 1385
rect 11913 1359 11919 1385
rect 12721 1359 12727 1385
rect 12753 1359 12759 1385
rect 14681 1359 14687 1385
rect 14713 1359 14719 1385
rect 3767 1329 3793 1335
rect 3767 1297 3793 1303
rect 4775 1329 4801 1335
rect 4775 1297 4801 1303
rect 5223 1329 5249 1335
rect 5223 1297 5249 1303
rect 5391 1329 5417 1335
rect 5391 1297 5417 1303
rect 6119 1329 6145 1335
rect 10039 1329 10065 1335
rect 12951 1329 12977 1335
rect 6617 1303 6623 1329
rect 6649 1303 6655 1329
rect 7009 1303 7015 1329
rect 7041 1303 7047 1329
rect 9193 1303 9199 1329
rect 9225 1303 9231 1329
rect 10313 1303 10319 1329
rect 10345 1303 10351 1329
rect 11713 1303 11719 1329
rect 11745 1303 11751 1329
rect 13337 1303 13343 1329
rect 13369 1303 13375 1329
rect 6119 1297 6145 1303
rect 10039 1297 10065 1303
rect 12951 1297 12977 1303
rect 3599 1273 3625 1279
rect 3599 1241 3625 1247
rect 4047 1273 4073 1279
rect 4047 1241 4073 1247
rect 4495 1273 4521 1279
rect 4495 1241 4521 1247
rect 4943 1273 4969 1279
rect 4943 1241 4969 1247
rect 5671 1273 5697 1279
rect 5671 1241 5697 1247
rect 7687 1273 7713 1279
rect 7687 1241 7713 1247
rect 8471 1273 8497 1279
rect 8471 1241 8497 1247
rect 9759 1273 9785 1279
rect 9759 1241 9785 1247
rect 10599 1273 10625 1279
rect 10599 1241 10625 1247
rect 11439 1273 11465 1279
rect 11439 1241 11465 1247
rect 12167 1273 12193 1279
rect 12167 1241 12193 1247
rect 336 1189 15512 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 15512 1189
rect 336 1146 15512 1163
rect 12615 1105 12641 1111
rect 12615 1073 12641 1079
rect 4831 1049 4857 1055
rect 4831 1017 4857 1023
rect 5447 1049 5473 1055
rect 5889 1023 5895 1049
rect 5921 1023 5927 1049
rect 6673 1023 6679 1049
rect 6705 1023 6711 1049
rect 7457 1023 7463 1049
rect 7489 1023 7495 1049
rect 9977 1023 9983 1049
rect 10009 1023 10015 1049
rect 13113 1023 13119 1049
rect 13145 1023 13151 1049
rect 13897 1023 13903 1049
rect 13929 1023 13935 1049
rect 14681 1023 14687 1049
rect 14713 1023 14719 1049
rect 15073 1023 15079 1049
rect 15105 1023 15111 1049
rect 5447 1017 5473 1023
rect 4551 993 4577 999
rect 5727 993 5753 999
rect 11551 993 11577 999
rect 5217 967 5223 993
rect 5249 967 5255 993
rect 8521 967 8527 993
rect 8553 967 8559 993
rect 9697 967 9703 993
rect 9729 967 9735 993
rect 10761 967 10767 993
rect 10793 967 10799 993
rect 12777 967 12783 993
rect 12809 967 12815 993
rect 4551 961 4577 967
rect 5727 961 5753 967
rect 11551 961 11577 967
rect 14407 937 14433 943
rect 5049 911 5055 937
rect 5081 911 5087 937
rect 7849 911 7855 937
rect 7881 911 7887 937
rect 11097 911 11103 937
rect 11129 911 11135 937
rect 11769 911 11775 937
rect 11801 911 11807 937
rect 14407 905 14433 911
rect 6399 881 6425 887
rect 6399 849 6425 855
rect 7183 881 7209 887
rect 7183 849 7209 855
rect 8695 881 8721 887
rect 8695 849 8721 855
rect 9311 881 9337 887
rect 9311 849 9337 855
rect 10263 881 10289 887
rect 10263 849 10289 855
rect 13623 881 13649 887
rect 13623 849 13649 855
rect 336 797 15512 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 15512 797
rect 336 754 15512 771
rect 15191 713 15217 719
rect 15191 681 15217 687
rect 4047 657 4073 663
rect 2921 631 2927 657
rect 2953 631 2959 657
rect 3369 631 3375 657
rect 3401 631 3407 657
rect 4047 625 4073 631
rect 4887 657 4913 663
rect 4887 625 4913 631
rect 6959 657 6985 663
rect 6959 625 6985 631
rect 12055 657 12081 663
rect 14345 631 14351 657
rect 14377 631 14383 657
rect 12055 625 12081 631
rect 6449 575 6455 601
rect 6481 575 6487 601
rect 7345 575 7351 601
rect 7377 575 7383 601
rect 8297 575 8303 601
rect 8329 575 8335 601
rect 9137 575 9143 601
rect 9169 575 9175 601
rect 10089 575 10095 601
rect 10121 575 10127 601
rect 10817 575 10823 601
rect 10849 575 10855 601
rect 12553 575 12559 601
rect 12585 575 12591 601
rect 13057 575 13063 601
rect 13089 575 13095 601
rect 13897 575 13903 601
rect 13929 575 13935 601
rect 14681 575 14687 601
rect 14713 575 14719 601
rect 4719 545 4745 551
rect 5329 519 5335 545
rect 5361 519 5367 545
rect 5721 519 5727 545
rect 5753 519 5759 545
rect 7625 519 7631 545
rect 7657 519 7663 545
rect 13337 519 13343 545
rect 13369 519 13375 545
rect 4719 513 4745 519
rect 3151 489 3177 495
rect 3151 457 3177 463
rect 3599 489 3625 495
rect 3599 457 3625 463
rect 3767 489 3793 495
rect 3767 457 3793 463
rect 4439 489 4465 495
rect 4439 457 4465 463
rect 5167 489 5193 495
rect 5167 457 5193 463
rect 8583 489 8609 495
rect 8583 457 8609 463
rect 9367 489 9393 495
rect 9367 457 9393 463
rect 10319 489 10345 495
rect 10319 457 10345 463
rect 11103 489 11129 495
rect 11103 457 11129 463
rect 336 405 15512 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 15512 405
rect 336 362 15512 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 1191 6567 1217 6593
rect 6735 6567 6761 6593
rect 7519 6567 7545 6593
rect 8135 6511 8161 6537
rect 1359 6455 1385 6481
rect 2143 6455 2169 6481
rect 3095 6455 3121 6481
rect 3879 6455 3905 6481
rect 5167 6455 5193 6481
rect 5335 6455 5361 6481
rect 6455 6455 6481 6481
rect 7239 6455 7265 6481
rect 9199 6455 9225 6481
rect 9423 6455 9449 6481
rect 10599 6455 10625 6481
rect 11327 6455 11353 6481
rect 12559 6455 12585 6481
rect 13399 6455 13425 6481
rect 14519 6455 14545 6481
rect 1807 6399 1833 6425
rect 2591 6399 2617 6425
rect 3375 6399 3401 6425
rect 4663 6399 4689 6425
rect 5839 6399 5865 6425
rect 8359 6399 8385 6425
rect 8751 6399 8777 6425
rect 9703 6399 9729 6425
rect 10151 6399 10177 6425
rect 10935 6399 10961 6425
rect 12111 6399 12137 6425
rect 12895 6399 12921 6425
rect 14127 6399 14153 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 4047 6175 4073 6201
rect 5559 6175 5585 6201
rect 8079 6175 8105 6201
rect 11439 6175 11465 6201
rect 13455 6175 13481 6201
rect 7519 6119 7545 6145
rect 9479 6119 9505 6145
rect 13063 6119 13089 6145
rect 15135 6119 15161 6145
rect 7295 6063 7321 6089
rect 8751 6063 8777 6089
rect 9031 6063 9057 6089
rect 12615 6063 12641 6089
rect 4551 6007 4577 6033
rect 5279 6007 5305 6033
rect 8583 6007 8609 6033
rect 9927 6007 9953 6033
rect 11943 6007 11969 6033
rect 13959 6007 13985 6033
rect 14687 6007 14713 6033
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 7071 5727 7097 5753
rect 13343 5727 13369 5753
rect 6791 5671 6817 5697
rect 7239 5671 7265 5697
rect 7687 5671 7713 5697
rect 8471 5671 8497 5697
rect 8751 5671 8777 5697
rect 12335 5671 12361 5697
rect 13735 5671 13761 5697
rect 14015 5671 14041 5697
rect 14687 5671 14713 5697
rect 7519 5615 7545 5641
rect 7967 5615 7993 5641
rect 12839 5615 12865 5641
rect 14407 5559 14433 5585
rect 15191 5559 15217 5585
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 13847 5391 13873 5417
rect 8135 5279 8161 5305
rect 8415 5279 8441 5305
rect 13343 5279 13369 5305
rect 14743 5279 14769 5305
rect 8695 5223 8721 5249
rect 15079 5223 15105 5249
rect 7855 5167 7881 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 13511 4943 13537 4969
rect 13903 4943 13929 4969
rect 14295 4943 14321 4969
rect 7351 4887 7377 4913
rect 7631 4887 7657 4913
rect 8471 4887 8497 4913
rect 13119 4887 13145 4913
rect 14687 4887 14713 4913
rect 8751 4831 8777 4857
rect 15191 4775 15217 4801
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 5223 4551 5249 4577
rect 7575 4551 7601 4577
rect 13791 4551 13817 4577
rect 5447 4495 5473 4521
rect 8863 4495 8889 4521
rect 13343 4495 13369 4521
rect 14687 4495 14713 4521
rect 15079 4439 15105 4465
rect 7351 4383 7377 4409
rect 8583 4383 8609 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 6567 4159 6593 4185
rect 7743 4159 7769 4185
rect 9535 4159 9561 4185
rect 9983 4159 10009 4185
rect 10431 4159 10457 4185
rect 11439 4159 11465 4185
rect 13623 4159 13649 4185
rect 13903 4159 13929 4185
rect 6847 4103 6873 4129
rect 7183 4103 7209 4129
rect 8023 4103 8049 4129
rect 8471 4103 8497 4129
rect 9815 4103 9841 4129
rect 10207 4103 10233 4129
rect 10711 4103 10737 4129
rect 11719 4103 11745 4129
rect 13343 4103 13369 4129
rect 14687 4103 14713 4129
rect 7463 4047 7489 4073
rect 8751 4047 8777 4073
rect 14351 4047 14377 4073
rect 15191 3991 15217 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 4999 3767 5025 3793
rect 5895 3767 5921 3793
rect 7519 3767 7545 3793
rect 8975 3767 9001 3793
rect 9703 3767 9729 3793
rect 10711 3767 10737 3793
rect 11383 3767 11409 3793
rect 14463 3767 14489 3793
rect 15135 3767 15161 3793
rect 5223 3711 5249 3737
rect 9199 3711 9225 3737
rect 14295 3711 14321 3737
rect 14799 3711 14825 3737
rect 9479 3655 9505 3681
rect 6119 3599 6145 3625
rect 7295 3599 7321 3625
rect 10991 3599 11017 3625
rect 11663 3599 11689 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 7743 3431 7769 3457
rect 8919 3431 8945 3457
rect 10151 3431 10177 3457
rect 10711 3431 10737 3457
rect 8415 3375 8441 3401
rect 7015 3319 7041 3345
rect 9703 3319 9729 3345
rect 10879 3319 10905 3345
rect 11159 3319 11185 3345
rect 11439 3319 11465 3345
rect 12335 3319 12361 3345
rect 12559 3319 12585 3345
rect 13455 3319 13481 3345
rect 13735 3319 13761 3345
rect 13903 3319 13929 3345
rect 14687 3319 14713 3345
rect 7295 3263 7321 3289
rect 7967 3263 7993 3289
rect 8695 3263 8721 3289
rect 9199 3263 9225 3289
rect 9927 3263 9953 3289
rect 10431 3263 10457 3289
rect 15191 3263 15217 3289
rect 14407 3207 14433 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 10599 2983 10625 3009
rect 12055 2983 12081 3009
rect 13959 2983 13985 3009
rect 14519 2983 14545 3009
rect 15135 2983 15161 3009
rect 7519 2927 7545 2953
rect 8191 2927 8217 2953
rect 9143 2927 9169 2953
rect 9311 2927 9337 2953
rect 9759 2927 9785 2953
rect 10823 2927 10849 2953
rect 14295 2927 14321 2953
rect 14687 2927 14713 2953
rect 7351 2871 7377 2897
rect 7799 2871 7825 2897
rect 8471 2871 8497 2897
rect 9591 2871 9617 2897
rect 10039 2871 10065 2897
rect 11103 2871 11129 2897
rect 7071 2815 7097 2841
rect 8863 2815 8889 2841
rect 10375 2815 10401 2841
rect 12335 2815 12361 2841
rect 13679 2815 13705 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 7351 2647 7377 2673
rect 8471 2647 8497 2673
rect 8919 2647 8945 2673
rect 9367 2647 9393 2673
rect 11439 2647 11465 2673
rect 12279 2647 12305 2673
rect 8751 2591 8777 2617
rect 10487 2591 10513 2617
rect 11271 2591 11297 2617
rect 12559 2591 12585 2617
rect 13903 2591 13929 2617
rect 15079 2591 15105 2617
rect 6847 2535 6873 2561
rect 7799 2535 7825 2561
rect 11719 2535 11745 2561
rect 14743 2535 14769 2561
rect 7127 2479 7153 2505
rect 7575 2479 7601 2505
rect 8023 2479 8049 2505
rect 9199 2479 9225 2505
rect 9647 2479 9673 2505
rect 14407 2479 14433 2505
rect 9983 2423 10009 2449
rect 10767 2423 10793 2449
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 8359 2199 8385 2225
rect 10487 2199 10513 2225
rect 11383 2199 11409 2225
rect 12559 2199 12585 2225
rect 15135 2199 15161 2225
rect 5895 2143 5921 2169
rect 7295 2143 7321 2169
rect 8079 2143 8105 2169
rect 9311 2143 9337 2169
rect 10879 2143 10905 2169
rect 14687 2143 14713 2169
rect 5503 2087 5529 2113
rect 6119 2087 6145 2113
rect 6511 2087 6537 2113
rect 8863 2087 8889 2113
rect 11719 2087 11745 2113
rect 12167 2087 12193 2113
rect 5223 2031 5249 2057
rect 6791 2031 6817 2057
rect 7575 2031 7601 2057
rect 8583 2031 8609 2057
rect 9479 2031 9505 2057
rect 11887 2031 11913 2057
rect 12335 2031 12361 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 6231 1863 6257 1889
rect 6511 1807 6537 1833
rect 9647 1807 9673 1833
rect 11215 1807 11241 1833
rect 13119 1807 13145 1833
rect 14295 1807 14321 1833
rect 4775 1751 4801 1777
rect 5783 1751 5809 1777
rect 6735 1751 6761 1777
rect 7463 1751 7489 1777
rect 8415 1751 8441 1777
rect 9479 1751 9505 1777
rect 11047 1751 11073 1777
rect 12279 1751 12305 1777
rect 13903 1751 13929 1777
rect 14743 1751 14769 1777
rect 4999 1695 5025 1721
rect 6063 1695 6089 1721
rect 7071 1695 7097 1721
rect 8639 1695 8665 1721
rect 12559 1695 12585 1721
rect 13567 1695 13593 1721
rect 15191 1695 15217 1721
rect 7743 1639 7769 1665
rect 8975 1639 9001 1665
rect 9927 1639 9953 1665
rect 10543 1639 10569 1665
rect 11719 1639 11745 1665
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 3375 1415 3401 1441
rect 13847 1415 13873 1441
rect 15135 1415 15161 1441
rect 5895 1359 5921 1385
rect 7407 1359 7433 1385
rect 8191 1359 8217 1385
rect 9591 1359 9617 1385
rect 11887 1359 11913 1385
rect 12727 1359 12753 1385
rect 14687 1359 14713 1385
rect 3767 1303 3793 1329
rect 4775 1303 4801 1329
rect 5223 1303 5249 1329
rect 5391 1303 5417 1329
rect 6119 1303 6145 1329
rect 6623 1303 6649 1329
rect 7015 1303 7041 1329
rect 9199 1303 9225 1329
rect 10039 1303 10065 1329
rect 10319 1303 10345 1329
rect 11719 1303 11745 1329
rect 12951 1303 12977 1329
rect 13343 1303 13369 1329
rect 3599 1247 3625 1273
rect 4047 1247 4073 1273
rect 4495 1247 4521 1273
rect 4943 1247 4969 1273
rect 5671 1247 5697 1273
rect 7687 1247 7713 1273
rect 8471 1247 8497 1273
rect 9759 1247 9785 1273
rect 10599 1247 10625 1273
rect 11439 1247 11465 1273
rect 12167 1247 12193 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 12615 1079 12641 1105
rect 4831 1023 4857 1049
rect 5447 1023 5473 1049
rect 5895 1023 5921 1049
rect 6679 1023 6705 1049
rect 7463 1023 7489 1049
rect 9983 1023 10009 1049
rect 13119 1023 13145 1049
rect 13903 1023 13929 1049
rect 14687 1023 14713 1049
rect 15079 1023 15105 1049
rect 4551 967 4577 993
rect 5223 967 5249 993
rect 5727 967 5753 993
rect 8527 967 8553 993
rect 9703 967 9729 993
rect 10767 967 10793 993
rect 11551 967 11577 993
rect 12783 967 12809 993
rect 5055 911 5081 937
rect 7855 911 7881 937
rect 11103 911 11129 937
rect 11775 911 11801 937
rect 14407 911 14433 937
rect 6399 855 6425 881
rect 7183 855 7209 881
rect 8695 855 8721 881
rect 9311 855 9337 881
rect 10263 855 10289 881
rect 13623 855 13649 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 15191 687 15217 713
rect 2927 631 2953 657
rect 3375 631 3401 657
rect 4047 631 4073 657
rect 4887 631 4913 657
rect 6959 631 6985 657
rect 12055 631 12081 657
rect 14351 631 14377 657
rect 6455 575 6481 601
rect 7351 575 7377 601
rect 8303 575 8329 601
rect 9143 575 9169 601
rect 10095 575 10121 601
rect 10823 575 10849 601
rect 12559 575 12585 601
rect 13063 575 13089 601
rect 13903 575 13929 601
rect 14687 575 14713 601
rect 4719 519 4745 545
rect 5335 519 5361 545
rect 5727 519 5753 545
rect 7631 519 7657 545
rect 13343 519 13369 545
rect 3151 463 3177 489
rect 3599 463 3625 489
rect 3767 463 3793 489
rect 4439 463 4465 489
rect 5167 463 5193 489
rect 8583 463 8609 489
rect 9367 463 9393 489
rect 10319 463 10345 489
rect 11103 463 11129 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
<< metal2 >>
rect 1120 7056 1176 7112
rect 1792 7056 1848 7112
rect 2464 7056 2520 7112
rect 3136 7056 3192 7112
rect 3808 7056 3864 7112
rect 4480 7056 4536 7112
rect 5152 7056 5208 7112
rect 5824 7056 5880 7112
rect 6496 7056 6552 7112
rect 7168 7056 7224 7112
rect 7840 7056 7896 7112
rect 8512 7056 8568 7112
rect 9184 7056 9240 7112
rect 9856 7056 9912 7112
rect 10528 7056 10584 7112
rect 11200 7056 11256 7112
rect 11872 7056 11928 7112
rect 12544 7056 12600 7112
rect 13216 7056 13272 7112
rect 13888 7056 13944 7112
rect 14560 7056 14616 7112
rect 742 6986 770 6991
rect 742 5754 770 6958
rect 1134 6594 1162 7056
rect 1190 6594 1218 6599
rect 1134 6593 1218 6594
rect 1134 6567 1191 6593
rect 1217 6567 1218 6593
rect 1134 6566 1218 6567
rect 1190 6561 1218 6566
rect 1358 6481 1386 6487
rect 1358 6455 1359 6481
rect 1385 6455 1386 6481
rect 742 5721 770 5726
rect 798 6314 826 6319
rect 798 5698 826 6286
rect 798 5665 826 5670
rect 1358 4634 1386 6455
rect 1806 6425 1834 7056
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 1806 6399 1807 6425
rect 1833 6399 1834 6425
rect 1806 6393 1834 6399
rect 2142 6481 2170 6487
rect 2142 6455 2143 6481
rect 2169 6455 2170 6481
rect 2142 6370 2170 6455
rect 2478 6426 2506 7056
rect 3150 7042 3178 7056
rect 3150 7009 3178 7014
rect 3374 7042 3402 7047
rect 3094 6481 3122 6487
rect 3094 6455 3095 6481
rect 3121 6455 3122 6481
rect 2590 6426 2618 6431
rect 2478 6425 2618 6426
rect 2478 6399 2591 6425
rect 2617 6399 2618 6425
rect 2478 6398 2618 6399
rect 2590 6393 2618 6398
rect 2142 6337 2170 6342
rect 3094 6314 3122 6455
rect 3374 6425 3402 7014
rect 3822 6594 3850 7056
rect 4494 7042 4522 7056
rect 4494 7009 4522 7014
rect 4662 7042 4690 7047
rect 3822 6566 4074 6594
rect 3374 6399 3375 6425
rect 3401 6399 3402 6425
rect 3374 6393 3402 6399
rect 3878 6481 3906 6487
rect 3878 6455 3879 6481
rect 3905 6455 3906 6481
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 3094 6281 3122 6286
rect 1902 6253 2034 6258
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 3878 5530 3906 6455
rect 4046 6201 4074 6566
rect 4662 6425 4690 7014
rect 5166 7042 5194 7056
rect 5166 7009 5194 7014
rect 5558 7042 5586 7047
rect 4662 6399 4663 6425
rect 4689 6399 4690 6425
rect 4662 6393 4690 6399
rect 4998 6482 5026 6487
rect 4046 6175 4047 6201
rect 4073 6175 4074 6201
rect 4046 6169 4074 6175
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 3878 5497 3906 5502
rect 4550 6033 4578 6039
rect 4550 6007 4551 6033
rect 4577 6007 4578 6033
rect 1902 5469 2034 5474
rect 4550 5474 4578 6007
rect 4550 5441 4578 5446
rect 4886 5978 4914 5983
rect 4662 5138 4690 5143
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 1358 4601 1386 4606
rect 742 4578 770 4583
rect 182 4186 210 4191
rect 182 2506 210 4158
rect 182 2473 210 2478
rect 742 1162 770 4550
rect 2982 4466 3010 4471
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 1358 3738 1386 3743
rect 798 1778 826 1783
rect 798 1386 826 1750
rect 798 1353 826 1358
rect 742 1129 770 1134
rect 1358 266 1386 3710
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 2926 2226 2954 2231
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 2702 1442 2730 1447
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 1358 233 1386 238
rect 2702 56 2730 1414
rect 2814 714 2842 719
rect 2814 56 2842 686
rect 2926 657 2954 2198
rect 2982 938 3010 4438
rect 4270 3682 4298 3687
rect 3990 3570 4018 3575
rect 2982 905 3010 910
rect 3206 2786 3234 2791
rect 2926 631 2927 657
rect 2953 631 2954 657
rect 2926 625 2954 631
rect 3150 489 3178 495
rect 3150 463 3151 489
rect 3177 463 3178 489
rect 3150 434 3178 463
rect 3150 401 3178 406
rect 2926 322 2954 327
rect 2926 56 2954 294
rect 3038 266 3066 271
rect 3038 56 3066 238
rect 3206 210 3234 2758
rect 3150 182 3234 210
rect 3262 2562 3290 2567
rect 3150 56 3178 182
rect 3262 56 3290 2534
rect 3430 1778 3458 1783
rect 3374 1554 3402 1559
rect 3374 1441 3402 1526
rect 3374 1415 3375 1441
rect 3401 1415 3402 1441
rect 3374 1409 3402 1415
rect 3374 657 3402 663
rect 3374 631 3375 657
rect 3401 631 3402 657
rect 3374 602 3402 631
rect 3374 569 3402 574
rect 3430 490 3458 1750
rect 3766 1329 3794 1335
rect 3766 1303 3767 1329
rect 3793 1303 3794 1329
rect 3374 462 3458 490
rect 3486 1274 3514 1279
rect 3374 56 3402 462
rect 3486 56 3514 1246
rect 3598 1273 3626 1279
rect 3598 1247 3599 1273
rect 3625 1247 3626 1273
rect 3598 658 3626 1247
rect 3598 625 3626 630
rect 3710 994 3738 999
rect 3598 490 3626 495
rect 3598 443 3626 462
rect 3598 378 3626 383
rect 3598 56 3626 350
rect 3710 56 3738 966
rect 3766 770 3794 1303
rect 3766 737 3794 742
rect 3990 546 4018 3542
rect 4158 3346 4186 3351
rect 4046 1274 4074 1279
rect 4046 1273 4130 1274
rect 4046 1247 4047 1273
rect 4073 1247 4130 1273
rect 4046 1246 4130 1247
rect 4046 1241 4074 1246
rect 4046 826 4074 831
rect 4046 657 4074 798
rect 4046 631 4047 657
rect 4073 631 4074 657
rect 4046 625 4074 631
rect 3990 518 4074 546
rect 3766 489 3794 495
rect 3766 463 3767 489
rect 3793 463 3794 489
rect 3766 266 3794 463
rect 3766 233 3794 238
rect 3822 490 3850 495
rect 3822 56 3850 462
rect 3934 434 3962 439
rect 3934 56 3962 406
rect 4046 56 4074 518
rect 4102 434 4130 1246
rect 4102 401 4130 406
rect 4158 56 4186 3318
rect 4270 56 4298 3654
rect 4326 3514 4354 3519
rect 4326 1274 4354 3486
rect 4550 2618 4578 2623
rect 4550 1722 4578 2590
rect 4550 1689 4578 1694
rect 4606 2170 4634 2175
rect 4326 1246 4410 1274
rect 4382 56 4410 1246
rect 4494 1273 4522 1279
rect 4494 1247 4495 1273
rect 4521 1247 4522 1273
rect 4494 714 4522 1247
rect 4550 994 4578 999
rect 4550 947 4578 966
rect 4494 681 4522 686
rect 4438 489 4466 495
rect 4438 463 4439 489
rect 4465 463 4466 489
rect 4438 322 4466 463
rect 4438 289 4466 294
rect 4494 98 4522 103
rect 4494 56 4522 70
rect 4606 56 4634 2142
rect 4662 154 4690 5110
rect 4718 1946 4746 1951
rect 4718 938 4746 1918
rect 4774 1777 4802 1783
rect 4774 1751 4775 1777
rect 4801 1751 4802 1777
rect 4774 1442 4802 1751
rect 4774 1409 4802 1414
rect 4830 1498 4858 1503
rect 4774 1329 4802 1335
rect 4774 1303 4775 1329
rect 4801 1303 4802 1329
rect 4774 1050 4802 1303
rect 4774 1017 4802 1022
rect 4830 1049 4858 1470
rect 4886 1162 4914 5950
rect 4998 3793 5026 6454
rect 5166 6481 5194 6487
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 5166 5922 5194 6455
rect 5334 6482 5362 6487
rect 5334 6435 5362 6454
rect 5558 6201 5586 7014
rect 5838 6425 5866 7056
rect 6510 7042 6538 7056
rect 6510 7009 6538 7014
rect 6734 7042 6762 7047
rect 6734 6593 6762 7014
rect 6734 6567 6735 6593
rect 6761 6567 6762 6593
rect 6734 6561 6762 6567
rect 7182 6594 7210 7056
rect 7182 6561 7210 6566
rect 7294 6762 7322 6767
rect 6454 6482 6482 6487
rect 7238 6482 7266 6487
rect 5838 6399 5839 6425
rect 5865 6399 5866 6425
rect 5838 6393 5866 6399
rect 5894 6481 6482 6482
rect 5894 6455 6455 6481
rect 6481 6455 6482 6481
rect 5894 6454 6482 6455
rect 5558 6175 5559 6201
rect 5585 6175 5586 6201
rect 5558 6169 5586 6175
rect 5166 5889 5194 5894
rect 5278 6033 5306 6039
rect 5278 6007 5279 6033
rect 5305 6007 5306 6033
rect 5222 4578 5250 4583
rect 5278 4578 5306 6007
rect 5222 4577 5306 4578
rect 5222 4551 5223 4577
rect 5249 4551 5306 4577
rect 5222 4550 5306 4551
rect 5446 4858 5474 4863
rect 5222 4545 5250 4550
rect 5446 4521 5474 4830
rect 5446 4495 5447 4521
rect 5473 4495 5474 4521
rect 5446 4489 5474 4495
rect 4998 3767 4999 3793
rect 5025 3767 5026 3793
rect 4998 3761 5026 3767
rect 5222 4354 5250 4359
rect 5222 3737 5250 4326
rect 5222 3711 5223 3737
rect 5249 3711 5250 3737
rect 5222 3705 5250 3711
rect 5334 4298 5362 4303
rect 5054 3458 5082 3463
rect 4942 2730 4970 2735
rect 4942 1666 4970 2702
rect 5054 2674 5082 3430
rect 5054 2641 5082 2646
rect 5222 2057 5250 2063
rect 5222 2031 5223 2057
rect 5249 2031 5250 2057
rect 4998 1722 5026 1741
rect 5222 1694 5250 2031
rect 4998 1689 5026 1694
rect 4942 1633 4970 1638
rect 5110 1666 5250 1694
rect 4942 1274 4970 1279
rect 4942 1227 4970 1246
rect 5054 1162 5082 1167
rect 4886 1134 4970 1162
rect 4830 1023 4831 1049
rect 4857 1023 4858 1049
rect 4830 1017 4858 1023
rect 4718 910 4914 938
rect 4830 658 4858 663
rect 4718 546 4746 551
rect 4718 499 4746 518
rect 4662 121 4690 126
rect 4718 434 4746 439
rect 4718 56 4746 406
rect 4830 56 4858 630
rect 4886 657 4914 910
rect 4886 631 4887 657
rect 4913 631 4914 657
rect 4886 625 4914 631
rect 4942 56 4970 1134
rect 5054 937 5082 1134
rect 5054 911 5055 937
rect 5081 911 5082 937
rect 5054 905 5082 911
rect 5110 378 5138 1666
rect 5222 1330 5250 1335
rect 5222 1283 5250 1302
rect 5222 993 5250 999
rect 5222 967 5223 993
rect 5249 967 5250 993
rect 5166 938 5194 943
rect 5166 770 5194 910
rect 5222 882 5250 967
rect 5334 882 5362 4270
rect 5894 3793 5922 6454
rect 6454 6449 6482 6454
rect 7126 6481 7266 6482
rect 7126 6455 7239 6481
rect 7265 6455 7266 6481
rect 7126 6454 7266 6455
rect 7070 5754 7098 5759
rect 7070 5707 7098 5726
rect 6790 5697 6818 5703
rect 6790 5671 6791 5697
rect 6817 5671 6818 5697
rect 6790 5194 6818 5671
rect 6790 5161 6818 5166
rect 6566 4186 6594 4191
rect 6566 4139 6594 4158
rect 7126 4186 7154 6454
rect 7238 6449 7266 6454
rect 7294 6089 7322 6734
rect 7518 6594 7546 6599
rect 7518 6547 7546 6566
rect 7854 6538 7882 7056
rect 8526 7042 8554 7056
rect 8526 7009 8554 7014
rect 8750 7042 8778 7047
rect 8134 6538 8162 6543
rect 7854 6510 8106 6538
rect 8078 6201 8106 6510
rect 8134 6491 8162 6510
rect 8358 6426 8386 6431
rect 8358 6379 8386 6398
rect 8750 6425 8778 7014
rect 9198 6594 9226 7056
rect 9870 7042 9898 7056
rect 9870 7009 9898 7014
rect 10150 7042 10178 7047
rect 9198 6561 9226 6566
rect 9478 6594 9506 6599
rect 8750 6399 8751 6425
rect 8777 6399 8778 6425
rect 8750 6393 8778 6399
rect 9198 6481 9226 6487
rect 9198 6455 9199 6481
rect 9225 6455 9226 6481
rect 8078 6175 8079 6201
rect 8105 6175 8106 6201
rect 8078 6169 8106 6175
rect 9142 6314 9170 6319
rect 7518 6146 7546 6151
rect 7294 6063 7295 6089
rect 7321 6063 7322 6089
rect 7294 6057 7322 6063
rect 7462 6145 7546 6146
rect 7462 6119 7519 6145
rect 7545 6119 7546 6145
rect 7462 6118 7546 6119
rect 7238 5697 7266 5703
rect 7238 5671 7239 5697
rect 7265 5671 7266 5697
rect 7238 5642 7266 5671
rect 7238 5609 7266 5614
rect 7350 4913 7378 4919
rect 7350 4887 7351 4913
rect 7377 4887 7378 4913
rect 7350 4802 7378 4887
rect 7350 4769 7378 4774
rect 7462 4802 7490 6118
rect 7518 6113 7546 6118
rect 8750 6090 8778 6095
rect 8750 6043 8778 6062
rect 9030 6090 9058 6095
rect 9030 6043 9058 6062
rect 8582 6034 8610 6039
rect 8582 6033 8666 6034
rect 8582 6007 8583 6033
rect 8609 6007 8666 6033
rect 8582 6006 8666 6007
rect 8582 6001 8610 6006
rect 7742 5922 7770 5927
rect 7686 5697 7714 5703
rect 7686 5671 7687 5697
rect 7713 5671 7714 5697
rect 7518 5641 7546 5647
rect 7518 5615 7519 5641
rect 7545 5615 7546 5641
rect 7518 5362 7546 5615
rect 7686 5586 7714 5671
rect 7686 5553 7714 5558
rect 7518 5329 7546 5334
rect 7462 4769 7490 4774
rect 7574 4970 7602 4975
rect 7574 4577 7602 4942
rect 7630 4914 7658 4919
rect 7630 4867 7658 4886
rect 7574 4551 7575 4577
rect 7601 4551 7602 4577
rect 7574 4545 7602 4551
rect 7686 4466 7714 4471
rect 7350 4410 7378 4415
rect 7350 4363 7378 4382
rect 7126 4153 7154 4158
rect 5894 3767 5895 3793
rect 5921 3767 5922 3793
rect 5894 3761 5922 3767
rect 6734 4130 6762 4135
rect 6118 3626 6146 3631
rect 6118 3625 6202 3626
rect 6118 3599 6119 3625
rect 6145 3599 6202 3625
rect 6118 3598 6202 3599
rect 6118 3593 6146 3598
rect 5614 3066 5642 3071
rect 5502 2114 5530 2119
rect 5502 2067 5530 2086
rect 5502 2002 5530 2007
rect 5222 849 5250 854
rect 5278 854 5362 882
rect 5390 1329 5418 1335
rect 5390 1303 5391 1329
rect 5417 1303 5418 1329
rect 5166 742 5250 770
rect 5166 490 5194 495
rect 5166 443 5194 462
rect 5110 345 5138 350
rect 5222 266 5250 742
rect 5054 238 5250 266
rect 5054 56 5082 238
rect 5166 154 5194 159
rect 5166 56 5194 126
rect 5278 56 5306 854
rect 5390 714 5418 1303
rect 5446 1106 5474 1111
rect 5446 1049 5474 1078
rect 5446 1023 5447 1049
rect 5473 1023 5474 1049
rect 5446 1017 5474 1023
rect 5390 681 5418 686
rect 5334 546 5362 551
rect 5446 546 5474 551
rect 5334 499 5362 518
rect 5390 518 5446 546
rect 5390 56 5418 518
rect 5446 513 5474 518
rect 5502 434 5530 1974
rect 5502 401 5530 406
rect 5558 1890 5586 1895
rect 5558 322 5586 1862
rect 5614 546 5642 3038
rect 5838 2842 5866 2847
rect 5782 1778 5810 1783
rect 5782 1731 5810 1750
rect 5670 1273 5698 1279
rect 5670 1247 5671 1273
rect 5697 1247 5698 1273
rect 5670 658 5698 1247
rect 5726 994 5754 999
rect 5726 947 5754 966
rect 5670 625 5698 630
rect 5614 513 5642 518
rect 5726 546 5754 551
rect 5726 499 5754 518
rect 5502 294 5586 322
rect 5614 434 5642 439
rect 5502 56 5530 294
rect 5614 56 5642 406
rect 5726 210 5754 215
rect 5726 56 5754 182
rect 5838 56 5866 2814
rect 5894 2170 5922 2175
rect 5894 2123 5922 2142
rect 6118 2113 6146 2119
rect 6118 2087 6119 2113
rect 6145 2087 6146 2113
rect 6118 1778 6146 2087
rect 6118 1745 6146 1750
rect 6062 1721 6090 1727
rect 6062 1695 6063 1721
rect 6089 1695 6090 1721
rect 5894 1385 5922 1391
rect 5894 1359 5895 1385
rect 5921 1359 5922 1385
rect 5894 1218 5922 1359
rect 6062 1386 6090 1695
rect 6174 1666 6202 3598
rect 6734 2674 6762 4102
rect 6846 4129 6874 4135
rect 6846 4103 6847 4129
rect 6873 4103 6874 4129
rect 6846 3906 6874 4103
rect 6846 3873 6874 3878
rect 7182 4129 7210 4135
rect 7182 4103 7183 4129
rect 7209 4103 7210 4129
rect 7182 3626 7210 4103
rect 7518 4130 7546 4135
rect 7462 4074 7490 4079
rect 7462 4027 7490 4046
rect 7518 3793 7546 4102
rect 7518 3767 7519 3793
rect 7545 3767 7546 3793
rect 7518 3761 7546 3767
rect 7182 3593 7210 3598
rect 7294 3625 7322 3631
rect 7294 3599 7295 3625
rect 7321 3599 7322 3625
rect 7294 3402 7322 3599
rect 7686 3458 7714 4438
rect 7742 4185 7770 5894
rect 8470 5698 8498 5703
rect 8470 5651 8498 5670
rect 7966 5642 7994 5647
rect 7966 5595 7994 5614
rect 8358 5530 8386 5535
rect 8134 5306 8162 5311
rect 8134 5259 8162 5278
rect 7854 5193 7882 5199
rect 7854 5167 7855 5193
rect 7881 5167 7882 5193
rect 7854 5082 7882 5167
rect 7854 5049 7882 5054
rect 7742 4159 7743 4185
rect 7769 4159 7770 4185
rect 7742 4153 7770 4159
rect 8358 4186 8386 5502
rect 8414 5418 8442 5423
rect 8414 5305 8442 5390
rect 8414 5279 8415 5305
rect 8441 5279 8442 5305
rect 8414 5273 8442 5279
rect 8638 4970 8666 6006
rect 8750 5698 8778 5703
rect 8750 5651 8778 5670
rect 8694 5250 8722 5255
rect 8694 5203 8722 5222
rect 9142 5082 9170 6286
rect 9142 5049 9170 5054
rect 8638 4942 9002 4970
rect 8470 4913 8498 4919
rect 8470 4887 8471 4913
rect 8497 4887 8498 4913
rect 8470 4522 8498 4887
rect 8750 4858 8778 4863
rect 8750 4811 8778 4830
rect 8918 4578 8946 4583
rect 8470 4489 8498 4494
rect 8862 4522 8890 4527
rect 8862 4475 8890 4494
rect 8582 4409 8610 4415
rect 8582 4383 8583 4409
rect 8609 4383 8610 4409
rect 8582 4242 8610 4383
rect 8582 4209 8610 4214
rect 8358 4153 8386 4158
rect 8022 4129 8050 4135
rect 8022 4103 8023 4129
rect 8049 4103 8050 4129
rect 8022 3514 8050 4103
rect 8470 4129 8498 4135
rect 8470 4103 8471 4129
rect 8497 4103 8498 4129
rect 8470 3850 8498 4103
rect 8750 4073 8778 4079
rect 8750 4047 8751 4073
rect 8777 4047 8778 4073
rect 8750 4018 8778 4047
rect 8750 3985 8778 3990
rect 8470 3817 8498 3822
rect 8022 3481 8050 3486
rect 8190 3738 8218 3743
rect 7742 3458 7770 3463
rect 7686 3457 7770 3458
rect 7686 3431 7743 3457
rect 7769 3431 7770 3457
rect 7686 3430 7770 3431
rect 7742 3425 7770 3430
rect 7294 3369 7322 3374
rect 7014 3345 7042 3351
rect 7014 3319 7015 3345
rect 7041 3319 7042 3345
rect 7014 3234 7042 3319
rect 7014 3201 7042 3206
rect 7294 3289 7322 3295
rect 7294 3263 7295 3289
rect 7321 3263 7322 3289
rect 7294 3234 7322 3263
rect 7294 3201 7322 3206
rect 7966 3289 7994 3295
rect 7966 3263 7967 3289
rect 7993 3263 7994 3289
rect 7294 2982 7434 3010
rect 7294 2954 7322 2982
rect 7406 2954 7434 2982
rect 7518 2954 7546 2959
rect 7406 2953 7546 2954
rect 7406 2927 7519 2953
rect 7545 2927 7546 2953
rect 7406 2926 7546 2927
rect 7294 2921 7322 2926
rect 7518 2921 7546 2926
rect 7350 2898 7378 2903
rect 7798 2898 7826 2903
rect 7350 2897 7434 2898
rect 7350 2871 7351 2897
rect 7377 2871 7434 2897
rect 7350 2870 7434 2871
rect 7350 2865 7378 2870
rect 7070 2842 7098 2847
rect 6734 2641 6762 2646
rect 6958 2841 7098 2842
rect 6958 2815 7071 2841
rect 7097 2815 7098 2841
rect 6958 2814 7098 2815
rect 6846 2562 6874 2567
rect 6846 2515 6874 2534
rect 6566 2338 6594 2343
rect 6510 2114 6538 2119
rect 6342 2113 6538 2114
rect 6342 2087 6511 2113
rect 6537 2087 6538 2113
rect 6342 2086 6538 2087
rect 6230 2058 6258 2063
rect 6230 1889 6258 2030
rect 6230 1863 6231 1889
rect 6257 1863 6258 1889
rect 6230 1857 6258 1863
rect 6174 1633 6202 1638
rect 6062 1353 6090 1358
rect 6118 1329 6146 1335
rect 6118 1303 6119 1329
rect 6145 1303 6146 1329
rect 5894 1185 5922 1190
rect 6062 1274 6090 1279
rect 5894 1050 5922 1055
rect 5894 1003 5922 1022
rect 5950 322 5978 327
rect 5950 56 5978 294
rect 6062 56 6090 1246
rect 6118 1218 6146 1303
rect 6118 1185 6146 1190
rect 6174 882 6202 887
rect 6174 56 6202 854
rect 6342 826 6370 2086
rect 6510 2081 6538 2086
rect 6510 1834 6538 1839
rect 6566 1834 6594 2310
rect 6510 1833 6594 1834
rect 6510 1807 6511 1833
rect 6537 1807 6594 1833
rect 6510 1806 6594 1807
rect 6678 2114 6706 2119
rect 6510 1801 6538 1806
rect 6454 1330 6482 1335
rect 6622 1330 6650 1335
rect 6398 882 6426 887
rect 6398 835 6426 854
rect 6342 793 6370 798
rect 6398 658 6426 663
rect 6286 490 6314 495
rect 6286 56 6314 462
rect 6398 56 6426 630
rect 6454 601 6482 1302
rect 6566 1329 6650 1330
rect 6566 1303 6623 1329
rect 6649 1303 6650 1329
rect 6566 1302 6650 1303
rect 6454 575 6455 601
rect 6481 575 6482 601
rect 6454 569 6482 575
rect 6510 994 6538 999
rect 6510 56 6538 966
rect 6566 602 6594 1302
rect 6622 1297 6650 1302
rect 6678 1049 6706 2086
rect 6790 2057 6818 2063
rect 6790 2031 6791 2057
rect 6817 2031 6818 2057
rect 6734 1777 6762 1783
rect 6734 1751 6735 1777
rect 6761 1751 6762 1777
rect 6734 1722 6762 1751
rect 6734 1689 6762 1694
rect 6678 1023 6679 1049
rect 6705 1023 6706 1049
rect 6678 1017 6706 1023
rect 6566 569 6594 574
rect 6622 826 6650 831
rect 6622 56 6650 798
rect 6790 378 6818 2031
rect 6902 882 6930 887
rect 6734 350 6818 378
rect 6846 546 6874 551
rect 6734 56 6762 350
rect 6846 56 6874 518
rect 6902 154 6930 854
rect 6958 826 6986 2814
rect 7070 2809 7098 2814
rect 7350 2786 7378 2791
rect 7350 2673 7378 2758
rect 7350 2647 7351 2673
rect 7377 2647 7378 2673
rect 7350 2641 7378 2647
rect 7126 2505 7154 2511
rect 7126 2479 7127 2505
rect 7153 2479 7154 2505
rect 7070 1721 7098 1727
rect 7070 1695 7071 1721
rect 7097 1695 7098 1721
rect 6958 793 6986 798
rect 7014 1329 7042 1335
rect 7014 1303 7015 1329
rect 7041 1303 7042 1329
rect 6958 657 6986 663
rect 6958 631 6959 657
rect 6985 631 6986 657
rect 6958 266 6986 631
rect 7014 658 7042 1303
rect 7014 625 7042 630
rect 6958 233 6986 238
rect 6902 126 6986 154
rect 6958 56 6986 126
rect 7070 56 7098 1695
rect 7126 1050 7154 2479
rect 7294 2226 7322 2231
rect 7294 2169 7322 2198
rect 7294 2143 7295 2169
rect 7321 2143 7322 2169
rect 7294 2137 7322 2143
rect 7406 1610 7434 2870
rect 7798 2851 7826 2870
rect 7798 2562 7826 2567
rect 7798 2515 7826 2534
rect 7574 2506 7602 2511
rect 7518 2505 7602 2506
rect 7518 2479 7575 2505
rect 7601 2479 7602 2505
rect 7518 2478 7602 2479
rect 7406 1577 7434 1582
rect 7462 1777 7490 1783
rect 7462 1751 7463 1777
rect 7489 1751 7490 1777
rect 7462 1498 7490 1751
rect 7462 1465 7490 1470
rect 7406 1386 7434 1391
rect 7406 1339 7434 1358
rect 7462 1050 7490 1055
rect 7126 1049 7490 1050
rect 7126 1023 7463 1049
rect 7489 1023 7490 1049
rect 7126 1022 7490 1023
rect 7462 1017 7490 1022
rect 7238 938 7266 943
rect 7518 938 7546 2478
rect 7574 2473 7602 2478
rect 7182 881 7210 887
rect 7182 855 7183 881
rect 7209 855 7210 881
rect 7182 434 7210 855
rect 7182 401 7210 406
rect 7238 322 7266 910
rect 7350 910 7546 938
rect 7574 2057 7602 2063
rect 7574 2031 7575 2057
rect 7601 2031 7602 2057
rect 7574 938 7602 2031
rect 7742 1665 7770 1671
rect 7742 1639 7743 1665
rect 7769 1639 7770 1665
rect 7182 294 7266 322
rect 7294 658 7322 663
rect 7182 56 7210 294
rect 7294 56 7322 630
rect 7350 601 7378 910
rect 7574 905 7602 910
rect 7686 1273 7714 1279
rect 7686 1247 7687 1273
rect 7713 1247 7714 1273
rect 7350 575 7351 601
rect 7377 575 7378 601
rect 7350 569 7378 575
rect 7406 826 7434 831
rect 7406 56 7434 798
rect 7686 658 7714 1247
rect 7742 882 7770 1639
rect 7742 849 7770 854
rect 7854 937 7882 943
rect 7854 911 7855 937
rect 7881 911 7882 937
rect 7686 630 7770 658
rect 7630 546 7658 551
rect 7630 499 7658 518
rect 7518 434 7546 439
rect 7518 56 7546 406
rect 7630 266 7658 271
rect 7630 56 7658 238
rect 7742 56 7770 630
rect 7854 56 7882 911
rect 7966 826 7994 3263
rect 8190 2953 8218 3710
rect 8918 3457 8946 4550
rect 8974 3793 9002 4942
rect 9198 4242 9226 6455
rect 9422 6481 9450 6487
rect 9422 6455 9423 6481
rect 9449 6455 9450 6481
rect 9422 5810 9450 6455
rect 9478 6145 9506 6566
rect 9478 6119 9479 6145
rect 9505 6119 9506 6145
rect 9478 6113 9506 6119
rect 9702 6425 9730 6431
rect 9702 6399 9703 6425
rect 9729 6399 9730 6425
rect 9422 5777 9450 5782
rect 9534 5474 9562 5479
rect 9198 4209 9226 4214
rect 9310 5138 9338 5143
rect 8974 3767 8975 3793
rect 9001 3767 9002 3793
rect 8974 3761 9002 3767
rect 9198 3738 9226 3743
rect 8918 3431 8919 3457
rect 8945 3431 8946 3457
rect 8918 3425 8946 3431
rect 9030 3737 9226 3738
rect 9030 3711 9199 3737
rect 9225 3711 9226 3737
rect 9030 3710 9226 3711
rect 8414 3402 8442 3407
rect 8414 3355 8442 3374
rect 8190 2927 8191 2953
rect 8217 2927 8218 2953
rect 8190 2921 8218 2927
rect 8694 3289 8722 3295
rect 8694 3263 8695 3289
rect 8721 3263 8722 3289
rect 8470 2898 8498 2903
rect 8470 2897 8554 2898
rect 8470 2871 8471 2897
rect 8497 2871 8554 2897
rect 8470 2870 8554 2871
rect 8470 2865 8498 2870
rect 8470 2674 8498 2679
rect 8470 2627 8498 2646
rect 8022 2505 8050 2511
rect 8022 2479 8023 2505
rect 8049 2479 8050 2505
rect 8022 1386 8050 2479
rect 8526 2506 8554 2870
rect 8526 2473 8554 2478
rect 8358 2394 8386 2399
rect 8078 2282 8106 2287
rect 8078 2169 8106 2254
rect 8358 2225 8386 2366
rect 8358 2199 8359 2225
rect 8385 2199 8386 2225
rect 8358 2193 8386 2199
rect 8694 2226 8722 3263
rect 8750 3010 8778 3015
rect 8750 2617 8778 2982
rect 8750 2591 8751 2617
rect 8777 2591 8778 2617
rect 8750 2585 8778 2591
rect 8862 2841 8890 2847
rect 8862 2815 8863 2841
rect 8889 2815 8890 2841
rect 8862 2618 8890 2815
rect 8918 2786 8946 2791
rect 8918 2673 8946 2758
rect 8918 2647 8919 2673
rect 8945 2647 8946 2673
rect 8918 2641 8946 2647
rect 8862 2585 8890 2590
rect 8694 2193 8722 2198
rect 8078 2143 8079 2169
rect 8105 2143 8106 2169
rect 8078 2137 8106 2143
rect 8862 2113 8890 2119
rect 8862 2087 8863 2113
rect 8889 2087 8890 2113
rect 8582 2057 8610 2063
rect 8582 2031 8583 2057
rect 8609 2031 8610 2057
rect 8582 2002 8610 2031
rect 8582 1969 8610 1974
rect 8414 1834 8442 1839
rect 8414 1777 8442 1806
rect 8414 1751 8415 1777
rect 8441 1751 8442 1777
rect 8414 1745 8442 1751
rect 8526 1778 8554 1783
rect 8022 1353 8050 1358
rect 8190 1554 8218 1559
rect 8190 1385 8218 1526
rect 8190 1359 8191 1385
rect 8217 1359 8218 1385
rect 8190 1353 8218 1359
rect 8470 1273 8498 1279
rect 8470 1247 8471 1273
rect 8497 1247 8498 1273
rect 7966 793 7994 798
rect 8078 938 8106 943
rect 7966 546 7994 551
rect 7966 56 7994 518
rect 8078 56 8106 910
rect 8470 938 8498 1247
rect 8526 993 8554 1750
rect 8638 1722 8666 1741
rect 8638 1689 8666 1694
rect 8862 1666 8890 2087
rect 8974 1666 9002 1671
rect 8862 1633 8890 1638
rect 8918 1665 9002 1666
rect 8918 1639 8975 1665
rect 9001 1639 9002 1665
rect 8918 1638 9002 1639
rect 8526 967 8527 993
rect 8553 967 8554 993
rect 8526 961 8554 967
rect 8638 1330 8666 1335
rect 8470 905 8498 910
rect 8358 882 8386 887
rect 8302 770 8330 775
rect 8302 601 8330 742
rect 8302 575 8303 601
rect 8329 575 8330 601
rect 8302 569 8330 575
rect 8190 490 8218 495
rect 8190 56 8218 462
rect 8358 434 8386 854
rect 8582 490 8610 495
rect 8582 443 8610 462
rect 8302 406 8386 434
rect 8526 434 8554 439
rect 8302 56 8330 406
rect 8414 266 8442 271
rect 8414 56 8442 238
rect 8526 56 8554 406
rect 8638 56 8666 1302
rect 8694 882 8722 887
rect 8918 882 8946 1638
rect 8974 1633 9002 1638
rect 9030 994 9058 3710
rect 9198 3705 9226 3710
rect 9198 3289 9226 3295
rect 9198 3263 9199 3289
rect 9225 3263 9226 3289
rect 9142 2954 9170 2959
rect 9142 2907 9170 2926
rect 9198 2618 9226 3263
rect 9310 2953 9338 5110
rect 9534 4185 9562 5446
rect 9702 4578 9730 6399
rect 10150 6425 10178 7014
rect 10542 7042 10570 7056
rect 10542 7009 10570 7014
rect 10934 7042 10962 7047
rect 10150 6399 10151 6425
rect 10177 6399 10178 6425
rect 10150 6393 10178 6399
rect 10598 6481 10626 6487
rect 10598 6455 10599 6481
rect 10625 6455 10626 6481
rect 9702 4545 9730 4550
rect 9926 6033 9954 6039
rect 9926 6007 9927 6033
rect 9953 6007 9954 6033
rect 9534 4159 9535 4185
rect 9561 4159 9562 4185
rect 9534 4153 9562 4159
rect 9814 4129 9842 4135
rect 9814 4103 9815 4129
rect 9841 4103 9842 4129
rect 9702 3794 9730 3799
rect 9646 3793 9730 3794
rect 9646 3767 9703 3793
rect 9729 3767 9730 3793
rect 9646 3766 9730 3767
rect 9478 3682 9506 3687
rect 9478 3635 9506 3654
rect 9310 2927 9311 2953
rect 9337 2927 9338 2953
rect 9310 2921 9338 2927
rect 9366 3458 9394 3463
rect 9366 2673 9394 3430
rect 9366 2647 9367 2673
rect 9393 2647 9394 2673
rect 9366 2641 9394 2647
rect 9534 3290 9562 3295
rect 9198 2590 9282 2618
rect 9198 2506 9226 2511
rect 9086 2505 9226 2506
rect 9086 2479 9199 2505
rect 9225 2479 9226 2505
rect 9086 2478 9226 2479
rect 9086 1946 9114 2478
rect 9198 2473 9226 2478
rect 9254 2394 9282 2590
rect 9198 2366 9282 2394
rect 9086 1918 9170 1946
rect 9030 961 9058 966
rect 9086 1834 9114 1839
rect 8694 835 8722 854
rect 8750 854 8946 882
rect 8974 882 9002 887
rect 9086 882 9114 1806
rect 8750 56 8778 854
rect 8862 490 8890 495
rect 8862 56 8890 462
rect 8974 56 9002 854
rect 9030 854 9114 882
rect 9030 434 9058 854
rect 9142 601 9170 1918
rect 9198 1442 9226 2366
rect 9198 1409 9226 1414
rect 9310 2169 9338 2175
rect 9310 2143 9311 2169
rect 9337 2143 9338 2169
rect 9198 1330 9226 1335
rect 9198 1283 9226 1302
rect 9310 1106 9338 2143
rect 9478 2057 9506 2063
rect 9478 2031 9479 2057
rect 9505 2031 9506 2057
rect 9478 1890 9506 2031
rect 9478 1857 9506 1862
rect 9478 1778 9506 1783
rect 9534 1778 9562 3262
rect 9590 2897 9618 2903
rect 9590 2871 9591 2897
rect 9617 2871 9618 2897
rect 9590 2786 9618 2871
rect 9590 2753 9618 2758
rect 9646 2674 9674 3766
rect 9702 3761 9730 3766
rect 9758 3570 9786 3575
rect 9702 3346 9730 3351
rect 9702 3299 9730 3318
rect 9758 2953 9786 3542
rect 9758 2927 9759 2953
rect 9785 2927 9786 2953
rect 9758 2921 9786 2927
rect 9478 1777 9562 1778
rect 9478 1751 9479 1777
rect 9505 1751 9562 1777
rect 9478 1750 9562 1751
rect 9590 2646 9674 2674
rect 9478 1745 9506 1750
rect 9590 1385 9618 2646
rect 9814 2562 9842 4103
rect 9926 3794 9954 6007
rect 10150 5978 10178 5983
rect 9982 4242 10010 4247
rect 9982 4185 10010 4214
rect 9982 4159 9983 4185
rect 10009 4159 10010 4185
rect 9982 4153 10010 4159
rect 9926 3761 9954 3766
rect 10150 3457 10178 5950
rect 10542 5082 10570 5087
rect 10486 4634 10514 4639
rect 10430 4186 10458 4191
rect 10430 4139 10458 4158
rect 10150 3431 10151 3457
rect 10177 3431 10178 3457
rect 10150 3425 10178 3431
rect 10206 4129 10234 4135
rect 10206 4103 10207 4129
rect 10233 4103 10234 4129
rect 9926 3290 9954 3295
rect 9926 3243 9954 3262
rect 9758 2534 9842 2562
rect 10038 2897 10066 2903
rect 10038 2871 10039 2897
rect 10065 2871 10066 2897
rect 9646 2506 9674 2511
rect 9646 2505 9730 2506
rect 9646 2479 9647 2505
rect 9673 2479 9730 2505
rect 9646 2478 9730 2479
rect 9646 2473 9674 2478
rect 9646 1946 9674 1951
rect 9646 1833 9674 1918
rect 9646 1807 9647 1833
rect 9673 1807 9674 1833
rect 9646 1801 9674 1807
rect 9590 1359 9591 1385
rect 9617 1359 9618 1385
rect 9590 1353 9618 1359
rect 9310 1073 9338 1078
rect 9534 1050 9562 1055
rect 9142 575 9143 601
rect 9169 575 9170 601
rect 9142 569 9170 575
rect 9198 994 9226 999
rect 9030 406 9114 434
rect 9086 56 9114 406
rect 9198 378 9226 966
rect 9422 938 9450 943
rect 9310 881 9338 887
rect 9310 855 9311 881
rect 9337 855 9338 881
rect 9310 434 9338 855
rect 9310 401 9338 406
rect 9366 489 9394 495
rect 9366 463 9367 489
rect 9393 463 9394 489
rect 9142 350 9226 378
rect 9142 154 9170 350
rect 9310 322 9338 327
rect 9142 121 9170 126
rect 9198 210 9226 215
rect 9198 56 9226 182
rect 9310 56 9338 294
rect 9366 266 9394 463
rect 9366 233 9394 238
rect 9422 56 9450 910
rect 9534 56 9562 1022
rect 9702 993 9730 2478
rect 9758 2170 9786 2534
rect 9982 2450 10010 2455
rect 9758 2137 9786 2142
rect 9814 2449 10010 2450
rect 9814 2423 9983 2449
rect 10009 2423 10010 2449
rect 9814 2422 10010 2423
rect 9758 1274 9786 1279
rect 9758 1227 9786 1246
rect 9702 967 9703 993
rect 9729 967 9730 993
rect 9702 961 9730 967
rect 9814 882 9842 2422
rect 9982 2417 10010 2422
rect 10038 1694 10066 2871
rect 9758 854 9842 882
rect 9926 1665 9954 1671
rect 10038 1666 10122 1694
rect 9926 1639 9927 1665
rect 9953 1639 9954 1665
rect 9646 826 9674 831
rect 9646 56 9674 798
rect 9758 56 9786 854
rect 9870 546 9898 551
rect 9870 56 9898 518
rect 9926 322 9954 1639
rect 9982 1610 10010 1615
rect 9982 1049 10010 1582
rect 9982 1023 9983 1049
rect 10009 1023 10010 1049
rect 9982 1017 10010 1023
rect 10038 1329 10066 1335
rect 10038 1303 10039 1329
rect 10065 1303 10066 1329
rect 10038 994 10066 1303
rect 10038 961 10066 966
rect 10094 601 10122 1666
rect 10206 714 10234 4103
rect 10486 3682 10514 4606
rect 10542 3794 10570 5054
rect 10598 4186 10626 6455
rect 10934 6425 10962 7014
rect 11214 6594 11242 7056
rect 11886 7042 11914 7056
rect 11886 7009 11914 7014
rect 12110 7042 12138 7047
rect 11214 6566 11466 6594
rect 10934 6399 10935 6425
rect 10961 6399 10962 6425
rect 10934 6393 10962 6399
rect 11326 6481 11354 6487
rect 11326 6455 11327 6481
rect 11353 6455 11354 6481
rect 10598 4153 10626 4158
rect 10878 6370 10906 6375
rect 10710 4130 10738 4135
rect 10710 4129 10794 4130
rect 10710 4103 10711 4129
rect 10737 4103 10794 4129
rect 10710 4102 10794 4103
rect 10710 4097 10738 4102
rect 10710 3794 10738 3799
rect 10542 3793 10738 3794
rect 10542 3767 10711 3793
rect 10737 3767 10738 3793
rect 10542 3766 10738 3767
rect 10710 3761 10738 3766
rect 10486 3654 10738 3682
rect 10710 3457 10738 3654
rect 10710 3431 10711 3457
rect 10737 3431 10738 3457
rect 10710 3425 10738 3431
rect 10430 3289 10458 3295
rect 10430 3263 10431 3289
rect 10457 3263 10458 3289
rect 10374 2842 10402 2847
rect 10374 2795 10402 2814
rect 10374 2450 10402 2455
rect 10318 1329 10346 1335
rect 10318 1303 10319 1329
rect 10345 1303 10346 1329
rect 10318 1162 10346 1303
rect 10318 1129 10346 1134
rect 10262 882 10290 887
rect 10262 835 10290 854
rect 10206 686 10290 714
rect 10094 575 10095 601
rect 10121 575 10122 601
rect 10094 569 10122 575
rect 10206 602 10234 607
rect 9926 289 9954 294
rect 9982 434 10010 439
rect 9982 56 10010 406
rect 10094 266 10122 271
rect 10094 56 10122 238
rect 10206 56 10234 574
rect 10262 154 10290 686
rect 10318 490 10346 495
rect 10318 443 10346 462
rect 10374 378 10402 2422
rect 10430 1498 10458 3263
rect 10598 3009 10626 3015
rect 10598 2983 10599 3009
rect 10625 2983 10626 3009
rect 10486 2618 10514 2623
rect 10598 2618 10626 2983
rect 10486 2617 10626 2618
rect 10486 2591 10487 2617
rect 10513 2591 10626 2617
rect 10486 2590 10626 2591
rect 10486 2585 10514 2590
rect 10766 2562 10794 4102
rect 10822 4074 10850 4079
rect 10822 3234 10850 4046
rect 10878 3458 10906 6342
rect 10878 3425 10906 3430
rect 10934 4298 10962 4303
rect 10822 3201 10850 3206
rect 10878 3345 10906 3351
rect 10878 3319 10879 3345
rect 10905 3319 10906 3345
rect 10822 3066 10850 3071
rect 10822 2953 10850 3038
rect 10822 2927 10823 2953
rect 10849 2927 10850 2953
rect 10822 2921 10850 2927
rect 10598 2534 10794 2562
rect 10430 1465 10458 1470
rect 10486 2225 10514 2231
rect 10486 2199 10487 2225
rect 10513 2199 10514 2225
rect 10262 121 10290 126
rect 10318 350 10402 378
rect 10430 1106 10458 1111
rect 10318 56 10346 350
rect 10430 56 10458 1078
rect 10486 546 10514 2199
rect 10542 1665 10570 1671
rect 10542 1639 10543 1665
rect 10569 1639 10570 1665
rect 10542 826 10570 1639
rect 10598 1386 10626 2534
rect 10766 2450 10794 2455
rect 10766 2403 10794 2422
rect 10878 2394 10906 3319
rect 10934 3346 10962 4270
rect 10934 3313 10962 3318
rect 10990 3625 11018 3631
rect 10990 3599 10991 3625
rect 11017 3599 11018 3625
rect 10822 2366 10906 2394
rect 10934 2562 10962 2567
rect 10822 1694 10850 2366
rect 10934 2282 10962 2534
rect 10878 2254 10962 2282
rect 10878 2169 10906 2254
rect 10878 2143 10879 2169
rect 10905 2143 10906 2169
rect 10878 2137 10906 2143
rect 10934 2170 10962 2175
rect 10598 1353 10626 1358
rect 10766 1666 10850 1694
rect 10878 1946 10906 1951
rect 10598 1273 10626 1279
rect 10598 1247 10599 1273
rect 10625 1247 10626 1273
rect 10598 938 10626 1247
rect 10598 905 10626 910
rect 10654 1218 10682 1223
rect 10542 793 10570 798
rect 10486 513 10514 518
rect 10542 658 10570 663
rect 10542 56 10570 630
rect 10654 56 10682 1190
rect 10766 1106 10794 1666
rect 10710 1078 10794 1106
rect 10710 882 10738 1078
rect 10766 994 10794 999
rect 10766 947 10794 966
rect 10710 854 10794 882
rect 10766 56 10794 854
rect 10822 714 10850 719
rect 10822 601 10850 686
rect 10822 575 10823 601
rect 10849 575 10850 601
rect 10822 569 10850 575
rect 10878 56 10906 1918
rect 10934 770 10962 2142
rect 10934 737 10962 742
rect 10990 56 11018 3599
rect 11270 3514 11298 3519
rect 11158 3346 11186 3351
rect 11046 3345 11186 3346
rect 11046 3319 11159 3345
rect 11185 3319 11186 3345
rect 11046 3318 11186 3319
rect 11046 1946 11074 3318
rect 11158 3313 11186 3318
rect 11102 2898 11130 2903
rect 11102 2897 11242 2898
rect 11102 2871 11103 2897
rect 11129 2871 11242 2897
rect 11102 2870 11242 2871
rect 11102 2865 11130 2870
rect 11046 1913 11074 1918
rect 11214 1833 11242 2870
rect 11270 2730 11298 3486
rect 11326 3010 11354 6455
rect 11438 6201 11466 6566
rect 12110 6425 12138 7014
rect 12558 7042 12586 7056
rect 12558 7009 12586 7014
rect 12894 7042 12922 7047
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12110 6399 12111 6425
rect 12137 6399 12138 6425
rect 12110 6393 12138 6399
rect 12558 6481 12586 6487
rect 12558 6455 12559 6481
rect 12585 6455 12586 6481
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11438 6175 11439 6201
rect 11465 6175 11466 6201
rect 11438 6169 11466 6175
rect 11942 6034 11970 6039
rect 11942 6033 12194 6034
rect 11942 6007 11943 6033
rect 11969 6007 12194 6033
rect 11942 6006 12194 6007
rect 11942 6001 11970 6006
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11902 5469 12034 5474
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 11606 4410 11634 4415
rect 11438 4186 11466 4191
rect 11438 4139 11466 4158
rect 11382 3794 11410 3799
rect 11382 3747 11410 3766
rect 11438 3458 11466 3463
rect 11438 3345 11466 3430
rect 11438 3319 11439 3345
rect 11465 3319 11466 3345
rect 11438 3313 11466 3319
rect 11326 2977 11354 2982
rect 11438 2730 11466 2735
rect 11270 2702 11354 2730
rect 11270 2618 11298 2623
rect 11270 2571 11298 2590
rect 11214 1807 11215 1833
rect 11241 1807 11242 1833
rect 11214 1801 11242 1807
rect 11046 1777 11074 1783
rect 11046 1751 11047 1777
rect 11073 1751 11074 1777
rect 11046 994 11074 1751
rect 11326 1694 11354 2702
rect 11438 2673 11466 2702
rect 11438 2647 11439 2673
rect 11465 2647 11466 2673
rect 11438 2641 11466 2647
rect 11214 1666 11354 1694
rect 11382 2225 11410 2231
rect 11382 2199 11383 2225
rect 11409 2199 11410 2225
rect 11158 1386 11186 1391
rect 11046 961 11074 966
rect 11102 1050 11130 1055
rect 11102 937 11130 1022
rect 11102 911 11103 937
rect 11129 911 11130 937
rect 11102 905 11130 911
rect 11102 490 11130 495
rect 11046 489 11130 490
rect 11046 463 11103 489
rect 11129 463 11130 489
rect 11046 462 11130 463
rect 11046 210 11074 462
rect 11102 457 11130 462
rect 11158 378 11186 1358
rect 11214 882 11242 1666
rect 11214 854 11354 882
rect 11046 177 11074 182
rect 11102 350 11186 378
rect 11214 770 11242 775
rect 11102 56 11130 350
rect 11214 56 11242 742
rect 11326 56 11354 854
rect 11382 658 11410 2199
rect 11550 1554 11578 1559
rect 11494 1442 11522 1447
rect 11382 625 11410 630
rect 11438 1273 11466 1279
rect 11438 1247 11439 1273
rect 11465 1247 11466 1273
rect 11438 434 11466 1247
rect 11494 602 11522 1414
rect 11550 1162 11578 1526
rect 11550 1129 11578 1134
rect 11550 993 11578 999
rect 11550 967 11551 993
rect 11577 967 11578 993
rect 11550 938 11578 967
rect 11550 905 11578 910
rect 11606 714 11634 4382
rect 11718 4129 11746 4135
rect 11718 4103 11719 4129
rect 11745 4103 11746 4129
rect 11662 3625 11690 3631
rect 11662 3599 11663 3625
rect 11689 3599 11690 3625
rect 11662 882 11690 3599
rect 11718 2898 11746 4103
rect 11830 4130 11858 4135
rect 11718 2870 11802 2898
rect 11718 2562 11746 2567
rect 11718 2515 11746 2534
rect 11718 2114 11746 2119
rect 11718 2067 11746 2086
rect 11718 1665 11746 1671
rect 11718 1639 11719 1665
rect 11745 1639 11746 1665
rect 11718 1442 11746 1639
rect 11718 1409 11746 1414
rect 11718 1330 11746 1335
rect 11718 1283 11746 1302
rect 11662 849 11690 854
rect 11718 1162 11746 1167
rect 11494 569 11522 574
rect 11550 686 11634 714
rect 11662 714 11690 719
rect 11438 401 11466 406
rect 11438 322 11466 327
rect 11438 56 11466 294
rect 11550 56 11578 686
rect 11662 322 11690 686
rect 11662 289 11690 294
rect 11718 210 11746 1134
rect 11774 1050 11802 2870
rect 11830 1106 11858 4102
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12166 3458 12194 6006
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12334 5698 12362 5703
rect 12334 5651 12362 5670
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 12558 4298 12586 6455
rect 12670 6426 12698 6431
rect 12614 6090 12642 6095
rect 12614 6043 12642 6062
rect 12558 4265 12586 4270
rect 12670 4186 12698 6398
rect 12894 6425 12922 7014
rect 13230 7042 13258 7056
rect 13230 7009 13258 7014
rect 13398 7042 13426 7047
rect 13398 6594 13426 7014
rect 13902 7042 13930 7056
rect 13902 7009 13930 7014
rect 14126 7042 14154 7047
rect 13790 6986 13818 6991
rect 13510 6762 13538 6767
rect 13398 6566 13482 6594
rect 12894 6399 12895 6425
rect 12921 6399 12922 6425
rect 12894 6393 12922 6399
rect 13398 6481 13426 6487
rect 13398 6455 13399 6481
rect 13425 6455 13426 6481
rect 12838 6314 12866 6319
rect 12838 5641 12866 6286
rect 13062 6145 13090 6151
rect 13062 6119 13063 6145
rect 13089 6119 13090 6145
rect 13062 6090 13090 6119
rect 13062 6057 13090 6062
rect 13342 5978 13370 5983
rect 13342 5753 13370 5950
rect 13342 5727 13343 5753
rect 13369 5727 13370 5753
rect 13342 5721 13370 5727
rect 12838 5615 12839 5641
rect 12865 5615 12866 5641
rect 12838 5609 12866 5615
rect 13342 5642 13370 5647
rect 13342 5305 13370 5614
rect 13342 5279 13343 5305
rect 13369 5279 13370 5305
rect 13342 5273 13370 5279
rect 13118 4913 13146 4919
rect 13118 4887 13119 4913
rect 13145 4887 13146 4913
rect 13118 4802 13146 4887
rect 13118 4769 13146 4774
rect 12670 4153 12698 4158
rect 13062 4634 13090 4639
rect 12614 4074 12642 4079
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12166 3430 12362 3458
rect 12166 3346 12194 3351
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 12054 3010 12082 3015
rect 12054 2963 12082 2982
rect 12166 2674 12194 3318
rect 12334 3345 12362 3430
rect 12558 3346 12586 3351
rect 12334 3319 12335 3345
rect 12361 3319 12362 3345
rect 12334 3313 12362 3319
rect 12502 3345 12586 3346
rect 12502 3319 12559 3345
rect 12585 3319 12586 3345
rect 12502 3318 12586 3319
rect 12334 2842 12362 2861
rect 12334 2809 12362 2814
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12278 2674 12306 2679
rect 12166 2673 12306 2674
rect 12166 2647 12279 2673
rect 12305 2647 12306 2673
rect 12166 2646 12306 2647
rect 12278 2641 12306 2646
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 11902 2333 12034 2338
rect 12166 2114 12194 2119
rect 12166 2067 12194 2086
rect 11886 2058 11914 2063
rect 11886 2011 11914 2030
rect 12334 2058 12362 2077
rect 12334 2025 12362 2030
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12278 1778 12306 1783
rect 12278 1731 12306 1750
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 11886 1498 11914 1503
rect 11886 1385 11914 1470
rect 11886 1359 11887 1385
rect 11913 1359 11914 1385
rect 11886 1353 11914 1359
rect 12166 1273 12194 1279
rect 12166 1247 12167 1273
rect 12193 1247 12194 1273
rect 12166 1218 12194 1247
rect 12166 1185 12194 1190
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 11830 1078 12250 1106
rect 11774 1022 12194 1050
rect 11774 938 11802 957
rect 11774 905 11802 910
rect 12110 882 12138 887
rect 11662 182 11746 210
rect 11774 826 11802 831
rect 11662 56 11690 182
rect 11774 56 11802 798
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 12054 657 12082 663
rect 12054 631 12055 657
rect 12081 631 12082 657
rect 12054 266 12082 631
rect 12054 233 12082 238
rect 11998 154 12026 159
rect 11886 98 11914 103
rect 11886 56 11914 70
rect 11998 56 12026 126
rect 12110 56 12138 854
rect 12166 322 12194 1022
rect 12222 490 12250 1078
rect 12502 882 12530 3318
rect 12558 3313 12586 3318
rect 12614 3010 12642 4046
rect 12614 2977 12642 2982
rect 12838 3122 12866 3127
rect 12558 2618 12586 2623
rect 12558 2571 12586 2590
rect 12558 2225 12586 2231
rect 12558 2199 12559 2225
rect 12585 2199 12586 2225
rect 12558 1834 12586 2199
rect 12558 1806 12642 1834
rect 12222 457 12250 462
rect 12446 854 12530 882
rect 12558 1721 12586 1727
rect 12558 1695 12559 1721
rect 12585 1695 12586 1721
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12334 322 12362 327
rect 12166 294 12250 322
rect 12222 56 12250 294
rect 12334 56 12362 294
rect 12446 56 12474 854
rect 12558 601 12586 1695
rect 12614 1694 12642 1806
rect 12614 1666 12810 1694
rect 12726 1385 12754 1391
rect 12726 1359 12727 1385
rect 12753 1359 12754 1385
rect 12614 1106 12642 1111
rect 12614 1059 12642 1078
rect 12558 575 12559 601
rect 12585 575 12586 601
rect 12558 569 12586 575
rect 12670 938 12698 943
rect 12558 490 12586 495
rect 12558 56 12586 462
rect 12670 56 12698 910
rect 12726 546 12754 1359
rect 12782 993 12810 1666
rect 12782 967 12783 993
rect 12809 967 12810 993
rect 12782 961 12810 967
rect 12726 513 12754 518
rect 12782 882 12810 887
rect 12838 882 12866 3094
rect 12894 2954 12922 2959
rect 12894 2562 12922 2926
rect 12894 2529 12922 2534
rect 13006 2954 13034 2959
rect 12950 1330 12978 1335
rect 12950 1283 12978 1302
rect 12838 854 12922 882
rect 12782 56 12810 854
rect 12894 56 12922 854
rect 13006 56 13034 2926
rect 13062 714 13090 4606
rect 13342 4578 13370 4583
rect 13342 4521 13370 4550
rect 13342 4495 13343 4521
rect 13369 4495 13370 4521
rect 13342 4489 13370 4495
rect 13342 4130 13370 4135
rect 13342 4083 13370 4102
rect 13398 3458 13426 6455
rect 13454 6201 13482 6566
rect 13454 6175 13455 6201
rect 13481 6175 13482 6201
rect 13454 6169 13482 6175
rect 13510 4969 13538 6734
rect 13734 5698 13762 5703
rect 13734 5651 13762 5670
rect 13510 4943 13511 4969
rect 13537 4943 13538 4969
rect 13510 4937 13538 4943
rect 13790 4577 13818 6958
rect 14126 6425 14154 7014
rect 14126 6399 14127 6425
rect 14153 6399 14154 6425
rect 14126 6393 14154 6399
rect 14350 6538 14378 6543
rect 13958 6033 13986 6039
rect 13958 6007 13959 6033
rect 13985 6007 13986 6033
rect 13846 5866 13874 5871
rect 13846 5417 13874 5838
rect 13846 5391 13847 5417
rect 13873 5391 13874 5417
rect 13846 5385 13874 5391
rect 13902 5362 13930 5367
rect 13902 4969 13930 5334
rect 13902 4943 13903 4969
rect 13929 4943 13930 4969
rect 13902 4937 13930 4943
rect 13790 4551 13791 4577
rect 13817 4551 13818 4577
rect 13790 4545 13818 4551
rect 13622 4298 13650 4303
rect 13622 4185 13650 4270
rect 13622 4159 13623 4185
rect 13649 4159 13650 4185
rect 13622 4153 13650 4159
rect 13902 4186 13930 4191
rect 13902 4139 13930 4158
rect 13398 3425 13426 3430
rect 13734 3458 13762 3463
rect 13454 3345 13482 3351
rect 13454 3319 13455 3345
rect 13481 3319 13482 3345
rect 13174 2674 13202 2679
rect 13118 2506 13146 2511
rect 13118 1833 13146 2478
rect 13118 1807 13119 1833
rect 13145 1807 13146 1833
rect 13118 1801 13146 1807
rect 13118 1666 13146 1671
rect 13118 1049 13146 1638
rect 13118 1023 13119 1049
rect 13145 1023 13146 1049
rect 13118 1017 13146 1023
rect 13062 681 13090 686
rect 13062 602 13090 607
rect 13174 602 13202 2646
rect 13230 2562 13258 2567
rect 13230 826 13258 2534
rect 13342 1329 13370 1335
rect 13342 1303 13343 1329
rect 13369 1303 13370 1329
rect 13342 1274 13370 1303
rect 13342 1241 13370 1246
rect 13454 938 13482 3319
rect 13734 3345 13762 3430
rect 13734 3319 13735 3345
rect 13761 3319 13762 3345
rect 13734 3313 13762 3319
rect 13902 3345 13930 3351
rect 13902 3319 13903 3345
rect 13929 3319 13930 3345
rect 13902 3290 13930 3319
rect 13902 3257 13930 3262
rect 13902 3066 13930 3071
rect 13678 2841 13706 2847
rect 13678 2815 13679 2841
rect 13705 2815 13706 2841
rect 13510 2282 13538 2287
rect 13510 1386 13538 2254
rect 13510 1353 13538 1358
rect 13566 1721 13594 1727
rect 13566 1695 13567 1721
rect 13593 1695 13594 1721
rect 13454 905 13482 910
rect 13230 793 13258 798
rect 13062 601 13202 602
rect 13062 575 13063 601
rect 13089 575 13202 601
rect 13062 574 13202 575
rect 13062 569 13090 574
rect 13342 545 13370 551
rect 13342 519 13343 545
rect 13369 519 13370 545
rect 13342 490 13370 519
rect 13342 457 13370 462
rect 13566 266 13594 1695
rect 13622 881 13650 887
rect 13622 855 13623 881
rect 13649 855 13650 881
rect 13622 714 13650 855
rect 13678 882 13706 2815
rect 13902 2617 13930 3038
rect 13958 3009 13986 6007
rect 14014 5697 14042 5703
rect 14014 5671 14015 5697
rect 14041 5671 14042 5697
rect 14014 5250 14042 5671
rect 14014 5217 14042 5222
rect 14294 5642 14322 5647
rect 14294 4969 14322 5614
rect 14294 4943 14295 4969
rect 14321 4943 14322 4969
rect 14294 4937 14322 4943
rect 14350 4073 14378 6510
rect 14518 6482 14546 6487
rect 14462 6481 14546 6482
rect 14462 6455 14519 6481
rect 14545 6455 14546 6481
rect 14462 6454 14546 6455
rect 14406 5585 14434 5591
rect 14406 5559 14407 5585
rect 14433 5559 14434 5585
rect 14406 5418 14434 5559
rect 14406 5385 14434 5390
rect 14350 4047 14351 4073
rect 14377 4047 14378 4073
rect 14350 4041 14378 4047
rect 14462 3793 14490 6454
rect 14518 6449 14546 6454
rect 14574 5978 14602 7056
rect 15134 6145 15162 6151
rect 15134 6119 15135 6145
rect 15161 6119 15162 6145
rect 14574 5945 14602 5950
rect 14686 6033 14714 6039
rect 14686 6007 14687 6033
rect 14713 6007 14714 6033
rect 14686 5922 14714 6007
rect 14686 5889 14714 5894
rect 14462 3767 14463 3793
rect 14489 3767 14490 3793
rect 14462 3761 14490 3767
rect 14518 5698 14546 5703
rect 14518 3794 14546 5670
rect 14686 5697 14714 5703
rect 14686 5671 14687 5697
rect 14713 5671 14714 5697
rect 14686 5306 14714 5671
rect 14686 5273 14714 5278
rect 14742 5305 14770 5311
rect 14742 5279 14743 5305
rect 14769 5279 14770 5305
rect 14686 4913 14714 4919
rect 14686 4887 14687 4913
rect 14713 4887 14714 4913
rect 14686 4858 14714 4887
rect 14742 4914 14770 5279
rect 15078 5249 15106 5255
rect 15078 5223 15079 5249
rect 15105 5223 15106 5249
rect 14742 4881 14770 4886
rect 14798 4970 14826 4975
rect 14686 4825 14714 4830
rect 14686 4522 14714 4527
rect 14686 4475 14714 4494
rect 14686 4129 14714 4135
rect 14686 4103 14687 4129
rect 14713 4103 14714 4129
rect 14686 4018 14714 4103
rect 14686 3985 14714 3990
rect 14518 3766 14602 3794
rect 14294 3737 14322 3743
rect 14294 3711 14295 3737
rect 14321 3711 14322 3737
rect 14294 3122 14322 3711
rect 14406 3233 14434 3239
rect 14406 3207 14407 3233
rect 14433 3207 14434 3233
rect 14406 3178 14434 3207
rect 14406 3145 14434 3150
rect 14294 3089 14322 3094
rect 13958 2983 13959 3009
rect 13985 2983 13986 3009
rect 13958 2977 13986 2983
rect 14518 3010 14546 3015
rect 14574 3010 14602 3766
rect 14798 3737 14826 4942
rect 15078 4746 15106 5223
rect 15134 5194 15162 6119
rect 15134 5161 15162 5166
rect 15190 5585 15218 5591
rect 15190 5559 15191 5585
rect 15217 5559 15218 5585
rect 15190 4970 15218 5559
rect 15190 4937 15218 4942
rect 15078 4713 15106 4718
rect 15190 4801 15218 4807
rect 15190 4775 15191 4801
rect 15217 4775 15218 4801
rect 15190 4522 15218 4775
rect 15190 4489 15218 4494
rect 15078 4465 15106 4471
rect 15078 4439 15079 4465
rect 15105 4439 15106 4465
rect 15078 4298 15106 4439
rect 15078 4265 15106 4270
rect 15134 4074 15162 4079
rect 15134 3793 15162 4046
rect 15190 4017 15218 4023
rect 15190 3991 15191 4017
rect 15217 3991 15218 4017
rect 15190 3850 15218 3991
rect 15190 3817 15218 3822
rect 15134 3767 15135 3793
rect 15161 3767 15162 3793
rect 15134 3761 15162 3767
rect 14798 3711 14799 3737
rect 14825 3711 14826 3737
rect 14798 3705 14826 3711
rect 15190 3626 15218 3631
rect 15134 3402 15162 3407
rect 14686 3345 14714 3351
rect 14686 3319 14687 3345
rect 14713 3319 14714 3345
rect 14686 3234 14714 3319
rect 14686 3201 14714 3206
rect 14518 3009 14602 3010
rect 14518 2983 14519 3009
rect 14545 2983 14602 3009
rect 14518 2982 14602 2983
rect 14686 3010 14714 3015
rect 14518 2977 14546 2982
rect 14294 2954 14322 2959
rect 14294 2907 14322 2926
rect 14686 2953 14714 2982
rect 15134 3009 15162 3374
rect 15190 3289 15218 3598
rect 15190 3263 15191 3289
rect 15217 3263 15218 3289
rect 15190 3257 15218 3263
rect 15134 2983 15135 3009
rect 15161 2983 15162 3009
rect 15134 2977 15162 2983
rect 14686 2927 14687 2953
rect 14713 2927 14714 2953
rect 14686 2921 14714 2927
rect 15078 2954 15106 2959
rect 13902 2591 13903 2617
rect 13929 2591 13930 2617
rect 13902 2585 13930 2591
rect 14742 2898 14770 2903
rect 14742 2561 14770 2870
rect 15078 2617 15106 2926
rect 15078 2591 15079 2617
rect 15105 2591 15106 2617
rect 15078 2585 15106 2591
rect 15134 2730 15162 2735
rect 14742 2535 14743 2561
rect 14769 2535 14770 2561
rect 14742 2529 14770 2535
rect 14406 2506 14434 2511
rect 14406 2459 14434 2478
rect 14742 2450 14770 2455
rect 14686 2226 14714 2231
rect 14686 2169 14714 2198
rect 14686 2143 14687 2169
rect 14713 2143 14714 2169
rect 14686 2137 14714 2143
rect 14294 1834 14322 1839
rect 14294 1787 14322 1806
rect 13902 1777 13930 1783
rect 13902 1751 13903 1777
rect 13929 1751 13930 1777
rect 13902 1722 13930 1751
rect 14742 1777 14770 2422
rect 15134 2225 15162 2702
rect 15134 2199 15135 2225
rect 15161 2199 15162 2225
rect 15134 2193 15162 2199
rect 15190 2282 15218 2287
rect 14742 1751 14743 1777
rect 14769 1751 14770 1777
rect 14742 1745 14770 1751
rect 15134 2058 15162 2063
rect 13902 1689 13930 1694
rect 15078 1610 15106 1615
rect 13678 849 13706 854
rect 13846 1441 13874 1447
rect 13846 1415 13847 1441
rect 13873 1415 13874 1441
rect 13622 681 13650 686
rect 13566 233 13594 238
rect 2688 0 2744 56
rect 2800 0 2856 56
rect 2912 0 2968 56
rect 3024 0 3080 56
rect 3136 0 3192 56
rect 3248 0 3304 56
rect 3360 0 3416 56
rect 3472 0 3528 56
rect 3584 0 3640 56
rect 3696 0 3752 56
rect 3808 0 3864 56
rect 3920 0 3976 56
rect 4032 0 4088 56
rect 4144 0 4200 56
rect 4256 0 4312 56
rect 4368 0 4424 56
rect 4480 0 4536 56
rect 4592 0 4648 56
rect 4704 0 4760 56
rect 4816 0 4872 56
rect 4928 0 4984 56
rect 5040 0 5096 56
rect 5152 0 5208 56
rect 5264 0 5320 56
rect 5376 0 5432 56
rect 5488 0 5544 56
rect 5600 0 5656 56
rect 5712 0 5768 56
rect 5824 0 5880 56
rect 5936 0 5992 56
rect 6048 0 6104 56
rect 6160 0 6216 56
rect 6272 0 6328 56
rect 6384 0 6440 56
rect 6496 0 6552 56
rect 6608 0 6664 56
rect 6720 0 6776 56
rect 6832 0 6888 56
rect 6944 0 7000 56
rect 7056 0 7112 56
rect 7168 0 7224 56
rect 7280 0 7336 56
rect 7392 0 7448 56
rect 7504 0 7560 56
rect 7616 0 7672 56
rect 7728 0 7784 56
rect 7840 0 7896 56
rect 7952 0 8008 56
rect 8064 0 8120 56
rect 8176 0 8232 56
rect 8288 0 8344 56
rect 8400 0 8456 56
rect 8512 0 8568 56
rect 8624 0 8680 56
rect 8736 0 8792 56
rect 8848 0 8904 56
rect 8960 0 9016 56
rect 9072 0 9128 56
rect 9184 0 9240 56
rect 9296 0 9352 56
rect 9408 0 9464 56
rect 9520 0 9576 56
rect 9632 0 9688 56
rect 9744 0 9800 56
rect 9856 0 9912 56
rect 9968 0 10024 56
rect 10080 0 10136 56
rect 10192 0 10248 56
rect 10304 0 10360 56
rect 10416 0 10472 56
rect 10528 0 10584 56
rect 10640 0 10696 56
rect 10752 0 10808 56
rect 10864 0 10920 56
rect 10976 0 11032 56
rect 11088 0 11144 56
rect 11200 0 11256 56
rect 11312 0 11368 56
rect 11424 0 11480 56
rect 11536 0 11592 56
rect 11648 0 11704 56
rect 11760 0 11816 56
rect 11872 0 11928 56
rect 11984 0 12040 56
rect 12096 0 12152 56
rect 12208 0 12264 56
rect 12320 0 12376 56
rect 12432 0 12488 56
rect 12544 0 12600 56
rect 12656 0 12712 56
rect 12768 0 12824 56
rect 12880 0 12936 56
rect 12992 0 13048 56
rect 13846 42 13874 1415
rect 13902 1442 13930 1447
rect 13902 1049 13930 1414
rect 14686 1386 14714 1391
rect 14686 1339 14714 1358
rect 13902 1023 13903 1049
rect 13929 1023 13930 1049
rect 13902 1017 13930 1023
rect 14406 1162 14434 1167
rect 14350 938 14378 943
rect 14350 657 14378 910
rect 14406 937 14434 1134
rect 14686 1050 14714 1055
rect 14686 1003 14714 1022
rect 15078 1049 15106 1582
rect 15134 1441 15162 2030
rect 15190 1721 15218 2254
rect 15190 1695 15191 1721
rect 15217 1695 15218 1721
rect 15190 1689 15218 1695
rect 15134 1415 15135 1441
rect 15161 1415 15162 1441
rect 15134 1409 15162 1415
rect 15078 1023 15079 1049
rect 15105 1023 15106 1049
rect 15078 1017 15106 1023
rect 15190 1386 15218 1391
rect 14406 911 14407 937
rect 14433 911 14434 937
rect 14406 905 14434 911
rect 14350 631 14351 657
rect 14377 631 14378 657
rect 14350 625 14378 631
rect 14686 826 14714 831
rect 13902 602 13930 607
rect 13902 555 13930 574
rect 14686 601 14714 798
rect 15190 713 15218 1358
rect 15190 687 15191 713
rect 15217 687 15218 713
rect 15190 681 15218 687
rect 14686 575 14687 601
rect 14713 575 14714 601
rect 14686 569 14714 575
rect 13846 9 13874 14
<< via2 >>
rect 742 6958 770 6986
rect 742 5726 770 5754
rect 798 6286 826 6314
rect 798 5670 826 5698
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 3150 7014 3178 7042
rect 3374 7014 3402 7042
rect 2142 6342 2170 6370
rect 4494 7014 4522 7042
rect 4662 7014 4690 7042
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 3094 6286 3122 6314
rect 2006 6258 2034 6259
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 5166 7014 5194 7042
rect 5558 7014 5586 7042
rect 4998 6454 5026 6482
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 3878 5502 3906 5530
rect 2006 5474 2034 5475
rect 4550 5446 4578 5474
rect 4886 5950 4914 5978
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 4662 5110 4690 5138
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1358 4606 1386 4634
rect 742 4550 770 4578
rect 182 4158 210 4186
rect 182 2478 210 2506
rect 2982 4438 3010 4466
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 1358 3710 1386 3738
rect 798 1750 826 1778
rect 798 1358 826 1386
rect 742 1134 770 1162
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 2926 2198 2954 2226
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 2702 1414 2730 1442
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 1358 238 1386 266
rect 2814 686 2842 714
rect 4270 3654 4298 3682
rect 3990 3542 4018 3570
rect 2982 910 3010 938
rect 3206 2758 3234 2786
rect 3150 406 3178 434
rect 2926 294 2954 322
rect 3038 238 3066 266
rect 3262 2534 3290 2562
rect 3430 1750 3458 1778
rect 3374 1526 3402 1554
rect 3374 574 3402 602
rect 3486 1246 3514 1274
rect 3598 630 3626 658
rect 3710 966 3738 994
rect 3598 489 3626 490
rect 3598 463 3599 489
rect 3599 463 3625 489
rect 3625 463 3626 489
rect 3598 462 3626 463
rect 3598 350 3626 378
rect 3766 742 3794 770
rect 4158 3318 4186 3346
rect 4046 798 4074 826
rect 3766 238 3794 266
rect 3822 462 3850 490
rect 3934 406 3962 434
rect 4102 406 4130 434
rect 4326 3486 4354 3514
rect 4550 2590 4578 2618
rect 4550 1694 4578 1722
rect 4606 2142 4634 2170
rect 4550 993 4578 994
rect 4550 967 4551 993
rect 4551 967 4577 993
rect 4577 967 4578 993
rect 4550 966 4578 967
rect 4494 686 4522 714
rect 4438 294 4466 322
rect 4494 70 4522 98
rect 4718 1918 4746 1946
rect 4774 1414 4802 1442
rect 4830 1470 4858 1498
rect 4774 1022 4802 1050
rect 5334 6481 5362 6482
rect 5334 6455 5335 6481
rect 5335 6455 5361 6481
rect 5361 6455 5362 6481
rect 5334 6454 5362 6455
rect 6510 7014 6538 7042
rect 6734 7014 6762 7042
rect 7182 6566 7210 6594
rect 7294 6734 7322 6762
rect 5166 5894 5194 5922
rect 5446 4830 5474 4858
rect 5222 4326 5250 4354
rect 5334 4270 5362 4298
rect 5054 3430 5082 3458
rect 4942 2702 4970 2730
rect 5054 2646 5082 2674
rect 4998 1721 5026 1722
rect 4998 1695 4999 1721
rect 4999 1695 5025 1721
rect 5025 1695 5026 1721
rect 4998 1694 5026 1695
rect 4942 1638 4970 1666
rect 4942 1273 4970 1274
rect 4942 1247 4943 1273
rect 4943 1247 4969 1273
rect 4969 1247 4970 1273
rect 4942 1246 4970 1247
rect 4830 630 4858 658
rect 4718 545 4746 546
rect 4718 519 4719 545
rect 4719 519 4745 545
rect 4745 519 4746 545
rect 4718 518 4746 519
rect 4662 126 4690 154
rect 4718 406 4746 434
rect 5054 1134 5082 1162
rect 5222 1329 5250 1330
rect 5222 1303 5223 1329
rect 5223 1303 5249 1329
rect 5249 1303 5250 1329
rect 5222 1302 5250 1303
rect 5166 910 5194 938
rect 7070 5753 7098 5754
rect 7070 5727 7071 5753
rect 7071 5727 7097 5753
rect 7097 5727 7098 5753
rect 7070 5726 7098 5727
rect 6790 5166 6818 5194
rect 6566 4185 6594 4186
rect 6566 4159 6567 4185
rect 6567 4159 6593 4185
rect 6593 4159 6594 4185
rect 6566 4158 6594 4159
rect 7518 6593 7546 6594
rect 7518 6567 7519 6593
rect 7519 6567 7545 6593
rect 7545 6567 7546 6593
rect 7518 6566 7546 6567
rect 8526 7014 8554 7042
rect 8750 7014 8778 7042
rect 8134 6537 8162 6538
rect 8134 6511 8135 6537
rect 8135 6511 8161 6537
rect 8161 6511 8162 6537
rect 8134 6510 8162 6511
rect 8358 6425 8386 6426
rect 8358 6399 8359 6425
rect 8359 6399 8385 6425
rect 8385 6399 8386 6425
rect 8358 6398 8386 6399
rect 9870 7014 9898 7042
rect 10150 7014 10178 7042
rect 9198 6566 9226 6594
rect 9478 6566 9506 6594
rect 9142 6286 9170 6314
rect 7238 5614 7266 5642
rect 7350 4774 7378 4802
rect 8750 6089 8778 6090
rect 8750 6063 8751 6089
rect 8751 6063 8777 6089
rect 8777 6063 8778 6089
rect 8750 6062 8778 6063
rect 9030 6089 9058 6090
rect 9030 6063 9031 6089
rect 9031 6063 9057 6089
rect 9057 6063 9058 6089
rect 9030 6062 9058 6063
rect 7742 5894 7770 5922
rect 7686 5558 7714 5586
rect 7518 5334 7546 5362
rect 7462 4774 7490 4802
rect 7574 4942 7602 4970
rect 7630 4913 7658 4914
rect 7630 4887 7631 4913
rect 7631 4887 7657 4913
rect 7657 4887 7658 4913
rect 7630 4886 7658 4887
rect 7686 4438 7714 4466
rect 7350 4409 7378 4410
rect 7350 4383 7351 4409
rect 7351 4383 7377 4409
rect 7377 4383 7378 4409
rect 7350 4382 7378 4383
rect 7126 4158 7154 4186
rect 6734 4102 6762 4130
rect 5614 3038 5642 3066
rect 5502 2113 5530 2114
rect 5502 2087 5503 2113
rect 5503 2087 5529 2113
rect 5529 2087 5530 2113
rect 5502 2086 5530 2087
rect 5502 1974 5530 2002
rect 5222 854 5250 882
rect 5166 489 5194 490
rect 5166 463 5167 489
rect 5167 463 5193 489
rect 5193 463 5194 489
rect 5166 462 5194 463
rect 5110 350 5138 378
rect 5166 126 5194 154
rect 5446 1078 5474 1106
rect 5390 686 5418 714
rect 5334 545 5362 546
rect 5334 519 5335 545
rect 5335 519 5361 545
rect 5361 519 5362 545
rect 5334 518 5362 519
rect 5446 518 5474 546
rect 5502 406 5530 434
rect 5558 1862 5586 1890
rect 5838 2814 5866 2842
rect 5782 1777 5810 1778
rect 5782 1751 5783 1777
rect 5783 1751 5809 1777
rect 5809 1751 5810 1777
rect 5782 1750 5810 1751
rect 5726 993 5754 994
rect 5726 967 5727 993
rect 5727 967 5753 993
rect 5753 967 5754 993
rect 5726 966 5754 967
rect 5670 630 5698 658
rect 5614 518 5642 546
rect 5726 545 5754 546
rect 5726 519 5727 545
rect 5727 519 5753 545
rect 5753 519 5754 545
rect 5726 518 5754 519
rect 5614 406 5642 434
rect 5726 182 5754 210
rect 5894 2169 5922 2170
rect 5894 2143 5895 2169
rect 5895 2143 5921 2169
rect 5921 2143 5922 2169
rect 5894 2142 5922 2143
rect 6118 1750 6146 1778
rect 6846 3878 6874 3906
rect 7518 4102 7546 4130
rect 7462 4073 7490 4074
rect 7462 4047 7463 4073
rect 7463 4047 7489 4073
rect 7489 4047 7490 4073
rect 7462 4046 7490 4047
rect 7182 3598 7210 3626
rect 8470 5697 8498 5698
rect 8470 5671 8471 5697
rect 8471 5671 8497 5697
rect 8497 5671 8498 5697
rect 8470 5670 8498 5671
rect 7966 5641 7994 5642
rect 7966 5615 7967 5641
rect 7967 5615 7993 5641
rect 7993 5615 7994 5641
rect 7966 5614 7994 5615
rect 8358 5502 8386 5530
rect 8134 5305 8162 5306
rect 8134 5279 8135 5305
rect 8135 5279 8161 5305
rect 8161 5279 8162 5305
rect 8134 5278 8162 5279
rect 7854 5054 7882 5082
rect 8414 5390 8442 5418
rect 8750 5697 8778 5698
rect 8750 5671 8751 5697
rect 8751 5671 8777 5697
rect 8777 5671 8778 5697
rect 8750 5670 8778 5671
rect 8694 5249 8722 5250
rect 8694 5223 8695 5249
rect 8695 5223 8721 5249
rect 8721 5223 8722 5249
rect 8694 5222 8722 5223
rect 9142 5054 9170 5082
rect 8750 4857 8778 4858
rect 8750 4831 8751 4857
rect 8751 4831 8777 4857
rect 8777 4831 8778 4857
rect 8750 4830 8778 4831
rect 8918 4550 8946 4578
rect 8470 4494 8498 4522
rect 8862 4521 8890 4522
rect 8862 4495 8863 4521
rect 8863 4495 8889 4521
rect 8889 4495 8890 4521
rect 8862 4494 8890 4495
rect 8582 4214 8610 4242
rect 8358 4158 8386 4186
rect 8750 3990 8778 4018
rect 8470 3822 8498 3850
rect 8022 3486 8050 3514
rect 8190 3710 8218 3738
rect 7294 3374 7322 3402
rect 7014 3206 7042 3234
rect 7294 3206 7322 3234
rect 7294 2926 7322 2954
rect 6734 2646 6762 2674
rect 6846 2561 6874 2562
rect 6846 2535 6847 2561
rect 6847 2535 6873 2561
rect 6873 2535 6874 2561
rect 6846 2534 6874 2535
rect 6566 2310 6594 2338
rect 6230 2030 6258 2058
rect 6174 1638 6202 1666
rect 6062 1358 6090 1386
rect 5894 1190 5922 1218
rect 6062 1246 6090 1274
rect 5894 1049 5922 1050
rect 5894 1023 5895 1049
rect 5895 1023 5921 1049
rect 5921 1023 5922 1049
rect 5894 1022 5922 1023
rect 5950 294 5978 322
rect 6118 1190 6146 1218
rect 6174 854 6202 882
rect 6678 2086 6706 2114
rect 6454 1302 6482 1330
rect 6398 881 6426 882
rect 6398 855 6399 881
rect 6399 855 6425 881
rect 6425 855 6426 881
rect 6398 854 6426 855
rect 6342 798 6370 826
rect 6398 630 6426 658
rect 6286 462 6314 490
rect 6510 966 6538 994
rect 6734 1694 6762 1722
rect 6566 574 6594 602
rect 6622 798 6650 826
rect 6902 854 6930 882
rect 6846 518 6874 546
rect 7350 2758 7378 2786
rect 6958 798 6986 826
rect 7014 630 7042 658
rect 6958 238 6986 266
rect 7294 2198 7322 2226
rect 7798 2897 7826 2898
rect 7798 2871 7799 2897
rect 7799 2871 7825 2897
rect 7825 2871 7826 2897
rect 7798 2870 7826 2871
rect 7798 2561 7826 2562
rect 7798 2535 7799 2561
rect 7799 2535 7825 2561
rect 7825 2535 7826 2561
rect 7798 2534 7826 2535
rect 7406 1582 7434 1610
rect 7462 1470 7490 1498
rect 7406 1385 7434 1386
rect 7406 1359 7407 1385
rect 7407 1359 7433 1385
rect 7433 1359 7434 1385
rect 7406 1358 7434 1359
rect 7238 910 7266 938
rect 7182 406 7210 434
rect 7574 910 7602 938
rect 7294 630 7322 658
rect 7406 798 7434 826
rect 7742 854 7770 882
rect 7630 545 7658 546
rect 7630 519 7631 545
rect 7631 519 7657 545
rect 7657 519 7658 545
rect 7630 518 7658 519
rect 7518 406 7546 434
rect 7630 238 7658 266
rect 9422 5782 9450 5810
rect 9534 5446 9562 5474
rect 9198 4214 9226 4242
rect 9310 5110 9338 5138
rect 8414 3401 8442 3402
rect 8414 3375 8415 3401
rect 8415 3375 8441 3401
rect 8441 3375 8442 3401
rect 8414 3374 8442 3375
rect 8470 2673 8498 2674
rect 8470 2647 8471 2673
rect 8471 2647 8497 2673
rect 8497 2647 8498 2673
rect 8470 2646 8498 2647
rect 8526 2478 8554 2506
rect 8358 2366 8386 2394
rect 8078 2254 8106 2282
rect 8750 2982 8778 3010
rect 8918 2758 8946 2786
rect 8862 2590 8890 2618
rect 8694 2198 8722 2226
rect 8582 1974 8610 2002
rect 8414 1806 8442 1834
rect 8526 1750 8554 1778
rect 8022 1358 8050 1386
rect 8190 1526 8218 1554
rect 7966 798 7994 826
rect 8078 910 8106 938
rect 7966 518 7994 546
rect 8638 1721 8666 1722
rect 8638 1695 8639 1721
rect 8639 1695 8665 1721
rect 8665 1695 8666 1721
rect 8638 1694 8666 1695
rect 8862 1638 8890 1666
rect 8638 1302 8666 1330
rect 8470 910 8498 938
rect 8358 854 8386 882
rect 8302 742 8330 770
rect 8190 462 8218 490
rect 8582 489 8610 490
rect 8582 463 8583 489
rect 8583 463 8609 489
rect 8609 463 8610 489
rect 8582 462 8610 463
rect 8526 406 8554 434
rect 8414 238 8442 266
rect 9142 2953 9170 2954
rect 9142 2927 9143 2953
rect 9143 2927 9169 2953
rect 9169 2927 9170 2953
rect 9142 2926 9170 2927
rect 10542 7014 10570 7042
rect 10934 7014 10962 7042
rect 9702 4550 9730 4578
rect 9478 3681 9506 3682
rect 9478 3655 9479 3681
rect 9479 3655 9505 3681
rect 9505 3655 9506 3681
rect 9478 3654 9506 3655
rect 9366 3430 9394 3458
rect 9534 3262 9562 3290
rect 9030 966 9058 994
rect 9086 1806 9114 1834
rect 8694 881 8722 882
rect 8694 855 8695 881
rect 8695 855 8721 881
rect 8721 855 8722 881
rect 8694 854 8722 855
rect 8974 854 9002 882
rect 8862 462 8890 490
rect 9198 1414 9226 1442
rect 9198 1329 9226 1330
rect 9198 1303 9199 1329
rect 9199 1303 9225 1329
rect 9225 1303 9226 1329
rect 9198 1302 9226 1303
rect 9478 1862 9506 1890
rect 9590 2758 9618 2786
rect 9758 3542 9786 3570
rect 9702 3345 9730 3346
rect 9702 3319 9703 3345
rect 9703 3319 9729 3345
rect 9729 3319 9730 3345
rect 9702 3318 9730 3319
rect 10150 5950 10178 5978
rect 9982 4214 10010 4242
rect 9926 3766 9954 3794
rect 10542 5054 10570 5082
rect 10486 4606 10514 4634
rect 10430 4185 10458 4186
rect 10430 4159 10431 4185
rect 10431 4159 10457 4185
rect 10457 4159 10458 4185
rect 10430 4158 10458 4159
rect 9926 3289 9954 3290
rect 9926 3263 9927 3289
rect 9927 3263 9953 3289
rect 9953 3263 9954 3289
rect 9926 3262 9954 3263
rect 9646 1918 9674 1946
rect 9310 1078 9338 1106
rect 9534 1022 9562 1050
rect 9198 966 9226 994
rect 9422 910 9450 938
rect 9310 406 9338 434
rect 9310 294 9338 322
rect 9142 126 9170 154
rect 9198 182 9226 210
rect 9366 238 9394 266
rect 9758 2142 9786 2170
rect 9758 1273 9786 1274
rect 9758 1247 9759 1273
rect 9759 1247 9785 1273
rect 9785 1247 9786 1273
rect 9758 1246 9786 1247
rect 9646 798 9674 826
rect 9870 518 9898 546
rect 9982 1582 10010 1610
rect 10038 966 10066 994
rect 11886 7014 11914 7042
rect 12110 7014 12138 7042
rect 10598 4158 10626 4186
rect 10878 6342 10906 6370
rect 10374 2841 10402 2842
rect 10374 2815 10375 2841
rect 10375 2815 10401 2841
rect 10401 2815 10402 2841
rect 10374 2814 10402 2815
rect 10374 2422 10402 2450
rect 10318 1134 10346 1162
rect 10262 881 10290 882
rect 10262 855 10263 881
rect 10263 855 10289 881
rect 10289 855 10290 881
rect 10262 854 10290 855
rect 10206 574 10234 602
rect 9926 294 9954 322
rect 9982 406 10010 434
rect 10094 238 10122 266
rect 10318 489 10346 490
rect 10318 463 10319 489
rect 10319 463 10345 489
rect 10345 463 10346 489
rect 10318 462 10346 463
rect 10822 4046 10850 4074
rect 10878 3430 10906 3458
rect 10934 4270 10962 4298
rect 10822 3206 10850 3234
rect 10822 3038 10850 3066
rect 10430 1470 10458 1498
rect 10262 126 10290 154
rect 10430 1078 10458 1106
rect 10766 2449 10794 2450
rect 10766 2423 10767 2449
rect 10767 2423 10793 2449
rect 10793 2423 10794 2449
rect 10766 2422 10794 2423
rect 10934 3318 10962 3346
rect 10934 2534 10962 2562
rect 10934 2142 10962 2170
rect 10598 1358 10626 1386
rect 10878 1918 10906 1946
rect 10598 910 10626 938
rect 10654 1190 10682 1218
rect 10542 798 10570 826
rect 10486 518 10514 546
rect 10542 630 10570 658
rect 10766 993 10794 994
rect 10766 967 10767 993
rect 10767 967 10793 993
rect 10793 967 10794 993
rect 10766 966 10794 967
rect 10822 686 10850 714
rect 10934 742 10962 770
rect 11270 3486 11298 3514
rect 11046 1918 11074 1946
rect 12558 7014 12586 7042
rect 12894 7014 12922 7042
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 11606 4382 11634 4410
rect 11438 4185 11466 4186
rect 11438 4159 11439 4185
rect 11439 4159 11465 4185
rect 11465 4159 11466 4185
rect 11438 4158 11466 4159
rect 11382 3793 11410 3794
rect 11382 3767 11383 3793
rect 11383 3767 11409 3793
rect 11409 3767 11410 3793
rect 11382 3766 11410 3767
rect 11438 3430 11466 3458
rect 11326 2982 11354 3010
rect 11270 2617 11298 2618
rect 11270 2591 11271 2617
rect 11271 2591 11297 2617
rect 11297 2591 11298 2617
rect 11270 2590 11298 2591
rect 11438 2702 11466 2730
rect 11158 1358 11186 1386
rect 11046 966 11074 994
rect 11102 1022 11130 1050
rect 11046 182 11074 210
rect 11214 742 11242 770
rect 11550 1526 11578 1554
rect 11494 1414 11522 1442
rect 11382 630 11410 658
rect 11550 1134 11578 1162
rect 11550 910 11578 938
rect 11830 4102 11858 4130
rect 11718 2561 11746 2562
rect 11718 2535 11719 2561
rect 11719 2535 11745 2561
rect 11745 2535 11746 2561
rect 11718 2534 11746 2535
rect 11718 2113 11746 2114
rect 11718 2087 11719 2113
rect 11719 2087 11745 2113
rect 11745 2087 11746 2113
rect 11718 2086 11746 2087
rect 11718 1414 11746 1442
rect 11718 1329 11746 1330
rect 11718 1303 11719 1329
rect 11719 1303 11745 1329
rect 11745 1303 11746 1329
rect 11718 1302 11746 1303
rect 11662 854 11690 882
rect 11718 1134 11746 1162
rect 11494 574 11522 602
rect 11662 686 11690 714
rect 11438 406 11466 434
rect 11438 294 11466 322
rect 11662 294 11690 322
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12334 5697 12362 5698
rect 12334 5671 12335 5697
rect 12335 5671 12361 5697
rect 12361 5671 12362 5697
rect 12334 5670 12362 5671
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12670 6398 12698 6426
rect 12614 6089 12642 6090
rect 12614 6063 12615 6089
rect 12615 6063 12641 6089
rect 12641 6063 12642 6089
rect 12614 6062 12642 6063
rect 12558 4270 12586 4298
rect 13230 7014 13258 7042
rect 13398 7014 13426 7042
rect 13902 7014 13930 7042
rect 14126 7014 14154 7042
rect 13790 6958 13818 6986
rect 13510 6734 13538 6762
rect 12838 6286 12866 6314
rect 13062 6062 13090 6090
rect 13342 5950 13370 5978
rect 13342 5614 13370 5642
rect 13118 4774 13146 4802
rect 12670 4158 12698 4186
rect 13062 4606 13090 4634
rect 12614 4046 12642 4074
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12166 3318 12194 3346
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 12054 3009 12082 3010
rect 12054 2983 12055 3009
rect 12055 2983 12081 3009
rect 12081 2983 12082 3009
rect 12054 2982 12082 2983
rect 12334 2841 12362 2842
rect 12334 2815 12335 2841
rect 12335 2815 12361 2841
rect 12361 2815 12362 2841
rect 12334 2814 12362 2815
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12006 2338 12034 2339
rect 12166 2113 12194 2114
rect 12166 2087 12167 2113
rect 12167 2087 12193 2113
rect 12193 2087 12194 2113
rect 12166 2086 12194 2087
rect 11886 2057 11914 2058
rect 11886 2031 11887 2057
rect 11887 2031 11913 2057
rect 11913 2031 11914 2057
rect 11886 2030 11914 2031
rect 12334 2057 12362 2058
rect 12334 2031 12335 2057
rect 12335 2031 12361 2057
rect 12361 2031 12362 2057
rect 12334 2030 12362 2031
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 12278 1777 12306 1778
rect 12278 1751 12279 1777
rect 12279 1751 12305 1777
rect 12305 1751 12306 1777
rect 12278 1750 12306 1751
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 11886 1470 11914 1498
rect 12166 1190 12194 1218
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 11774 937 11802 938
rect 11774 911 11775 937
rect 11775 911 11801 937
rect 11801 911 11802 937
rect 11774 910 11802 911
rect 12110 854 12138 882
rect 11774 798 11802 826
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 12054 238 12082 266
rect 11998 126 12026 154
rect 11886 70 11914 98
rect 12614 2982 12642 3010
rect 12838 3094 12866 3122
rect 12558 2617 12586 2618
rect 12558 2591 12559 2617
rect 12559 2591 12585 2617
rect 12585 2591 12586 2617
rect 12558 2590 12586 2591
rect 12222 462 12250 490
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12334 294 12362 322
rect 12614 1105 12642 1106
rect 12614 1079 12615 1105
rect 12615 1079 12641 1105
rect 12641 1079 12642 1105
rect 12614 1078 12642 1079
rect 12670 910 12698 938
rect 12558 462 12586 490
rect 12726 518 12754 546
rect 12782 854 12810 882
rect 12894 2926 12922 2954
rect 12894 2534 12922 2562
rect 13006 2926 13034 2954
rect 12950 1329 12978 1330
rect 12950 1303 12951 1329
rect 12951 1303 12977 1329
rect 12977 1303 12978 1329
rect 12950 1302 12978 1303
rect 13342 4550 13370 4578
rect 13342 4129 13370 4130
rect 13342 4103 13343 4129
rect 13343 4103 13369 4129
rect 13369 4103 13370 4129
rect 13342 4102 13370 4103
rect 13734 5697 13762 5698
rect 13734 5671 13735 5697
rect 13735 5671 13761 5697
rect 13761 5671 13762 5697
rect 13734 5670 13762 5671
rect 14350 6510 14378 6538
rect 13846 5838 13874 5866
rect 13902 5334 13930 5362
rect 13622 4270 13650 4298
rect 13902 4185 13930 4186
rect 13902 4159 13903 4185
rect 13903 4159 13929 4185
rect 13929 4159 13930 4185
rect 13902 4158 13930 4159
rect 13398 3430 13426 3458
rect 13734 3430 13762 3458
rect 13174 2646 13202 2674
rect 13118 2478 13146 2506
rect 13118 1638 13146 1666
rect 13062 686 13090 714
rect 13230 2534 13258 2562
rect 13342 1246 13370 1274
rect 13902 3262 13930 3290
rect 13902 3038 13930 3066
rect 13510 2254 13538 2282
rect 13510 1358 13538 1386
rect 13454 910 13482 938
rect 13230 798 13258 826
rect 13342 462 13370 490
rect 14014 5222 14042 5250
rect 14294 5614 14322 5642
rect 14406 5390 14434 5418
rect 14574 5950 14602 5978
rect 14686 5894 14714 5922
rect 14518 5670 14546 5698
rect 14686 5278 14714 5306
rect 14742 4886 14770 4914
rect 14798 4942 14826 4970
rect 14686 4830 14714 4858
rect 14686 4521 14714 4522
rect 14686 4495 14687 4521
rect 14687 4495 14713 4521
rect 14713 4495 14714 4521
rect 14686 4494 14714 4495
rect 14686 3990 14714 4018
rect 14406 3150 14434 3178
rect 14294 3094 14322 3122
rect 15134 5166 15162 5194
rect 15190 4942 15218 4970
rect 15078 4718 15106 4746
rect 15190 4494 15218 4522
rect 15078 4270 15106 4298
rect 15134 4046 15162 4074
rect 15190 3822 15218 3850
rect 15190 3598 15218 3626
rect 15134 3374 15162 3402
rect 14686 3206 14714 3234
rect 14686 2982 14714 3010
rect 14294 2953 14322 2954
rect 14294 2927 14295 2953
rect 14295 2927 14321 2953
rect 14321 2927 14322 2953
rect 14294 2926 14322 2927
rect 15078 2926 15106 2954
rect 14742 2870 14770 2898
rect 15134 2702 15162 2730
rect 14406 2505 14434 2506
rect 14406 2479 14407 2505
rect 14407 2479 14433 2505
rect 14433 2479 14434 2505
rect 14406 2478 14434 2479
rect 14742 2422 14770 2450
rect 14686 2198 14714 2226
rect 14294 1833 14322 1834
rect 14294 1807 14295 1833
rect 14295 1807 14321 1833
rect 14321 1807 14322 1833
rect 14294 1806 14322 1807
rect 15190 2254 15218 2282
rect 15134 2030 15162 2058
rect 13902 1694 13930 1722
rect 15078 1582 15106 1610
rect 13678 854 13706 882
rect 13622 686 13650 714
rect 13566 238 13594 266
rect 13902 1414 13930 1442
rect 14686 1385 14714 1386
rect 14686 1359 14687 1385
rect 14687 1359 14713 1385
rect 14713 1359 14714 1385
rect 14686 1358 14714 1359
rect 14406 1134 14434 1162
rect 14350 910 14378 938
rect 14686 1049 14714 1050
rect 14686 1023 14687 1049
rect 14687 1023 14713 1049
rect 14713 1023 14714 1049
rect 14686 1022 14714 1023
rect 15190 1358 15218 1386
rect 14686 798 14714 826
rect 13902 601 13930 602
rect 13902 575 13903 601
rect 13903 575 13929 601
rect 13929 575 13930 601
rect 13902 574 13930 575
rect 13846 14 13874 42
<< metal3 >>
rect 3145 7014 3150 7042
rect 3178 7014 3374 7042
rect 3402 7014 3407 7042
rect 4489 7014 4494 7042
rect 4522 7014 4662 7042
rect 4690 7014 4695 7042
rect 5161 7014 5166 7042
rect 5194 7014 5558 7042
rect 5586 7014 5591 7042
rect 6505 7014 6510 7042
rect 6538 7014 6734 7042
rect 6762 7014 6767 7042
rect 8521 7014 8526 7042
rect 8554 7014 8750 7042
rect 8778 7014 8783 7042
rect 9865 7014 9870 7042
rect 9898 7014 10150 7042
rect 10178 7014 10183 7042
rect 10537 7014 10542 7042
rect 10570 7014 10934 7042
rect 10962 7014 10967 7042
rect 11881 7014 11886 7042
rect 11914 7014 12110 7042
rect 12138 7014 12143 7042
rect 12553 7014 12558 7042
rect 12586 7014 12894 7042
rect 12922 7014 12927 7042
rect 13225 7014 13230 7042
rect 13258 7014 13398 7042
rect 13426 7014 13431 7042
rect 13897 7014 13902 7042
rect 13930 7014 14126 7042
rect 14154 7014 14159 7042
rect 0 6986 56 7000
rect 15792 6986 15848 7000
rect 0 6958 742 6986
rect 770 6958 775 6986
rect 13785 6958 13790 6986
rect 13818 6958 15848 6986
rect 0 6944 56 6958
rect 15792 6944 15848 6958
rect 0 6762 56 6776
rect 15792 6762 15848 6776
rect 0 6734 7294 6762
rect 7322 6734 7327 6762
rect 13505 6734 13510 6762
rect 13538 6734 15848 6762
rect 0 6720 56 6734
rect 15792 6720 15848 6734
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 7177 6566 7182 6594
rect 7210 6566 7518 6594
rect 7546 6566 7551 6594
rect 9193 6566 9198 6594
rect 9226 6566 9478 6594
rect 9506 6566 9511 6594
rect 0 6538 56 6552
rect 15792 6538 15848 6552
rect 0 6510 8134 6538
rect 8162 6510 8167 6538
rect 14345 6510 14350 6538
rect 14378 6510 15848 6538
rect 0 6496 56 6510
rect 15792 6496 15848 6510
rect 4993 6454 4998 6482
rect 5026 6454 5334 6482
rect 5362 6454 5367 6482
rect 8353 6398 8358 6426
rect 8386 6398 12670 6426
rect 12698 6398 12703 6426
rect 2137 6342 2142 6370
rect 2170 6342 10878 6370
rect 10906 6342 10911 6370
rect 0 6314 56 6328
rect 15792 6314 15848 6328
rect 0 6286 798 6314
rect 826 6286 831 6314
rect 3089 6286 3094 6314
rect 3122 6286 9142 6314
rect 9170 6286 9175 6314
rect 12833 6286 12838 6314
rect 12866 6286 15848 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 15792 6272 15848 6286
rect 0 6090 56 6104
rect 15792 6090 15848 6104
rect 0 6062 8750 6090
rect 8778 6062 8783 6090
rect 9025 6062 9030 6090
rect 9058 6062 12614 6090
rect 12642 6062 12647 6090
rect 13057 6062 13062 6090
rect 13090 6062 15848 6090
rect 0 6048 56 6062
rect 15792 6048 15848 6062
rect 4881 5950 4886 5978
rect 4914 5950 10150 5978
rect 10178 5950 10183 5978
rect 13337 5950 13342 5978
rect 13370 5950 14574 5978
rect 14602 5950 14607 5978
rect 5161 5894 5166 5922
rect 5194 5894 7742 5922
rect 7770 5894 7775 5922
rect 13426 5894 14686 5922
rect 14714 5894 14719 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 0 5838 2142 5866
rect 2170 5838 2175 5866
rect 0 5824 56 5838
rect 1666 5782 9422 5810
rect 9450 5782 9455 5810
rect 1666 5754 1694 5782
rect 13426 5754 13454 5894
rect 15792 5866 15848 5880
rect 13841 5838 13846 5866
rect 13874 5838 15848 5866
rect 15792 5824 15848 5838
rect 737 5726 742 5754
rect 770 5726 1694 5754
rect 7065 5726 7070 5754
rect 7098 5726 13454 5754
rect 793 5670 798 5698
rect 826 5670 8470 5698
rect 8498 5670 8503 5698
rect 8745 5670 8750 5698
rect 8778 5670 12334 5698
rect 12362 5670 12367 5698
rect 13729 5670 13734 5698
rect 13762 5670 14518 5698
rect 14546 5670 14551 5698
rect 0 5642 56 5656
rect 15792 5642 15848 5656
rect 0 5614 7238 5642
rect 7266 5614 7271 5642
rect 7961 5614 7966 5642
rect 7994 5614 13342 5642
rect 13370 5614 13375 5642
rect 14289 5614 14294 5642
rect 14322 5614 15848 5642
rect 0 5600 56 5614
rect 15792 5600 15848 5614
rect 2137 5558 2142 5586
rect 2170 5558 7686 5586
rect 7714 5558 7719 5586
rect 3873 5502 3878 5530
rect 3906 5502 8358 5530
rect 8386 5502 8391 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 4545 5446 4550 5474
rect 4578 5446 9534 5474
rect 9562 5446 9567 5474
rect 0 5418 56 5432
rect 15792 5418 15848 5432
rect 0 5390 8414 5418
rect 8442 5390 8447 5418
rect 14401 5390 14406 5418
rect 14434 5390 15848 5418
rect 0 5376 56 5390
rect 15792 5376 15848 5390
rect 7513 5334 7518 5362
rect 7546 5334 13902 5362
rect 13930 5334 13935 5362
rect 8129 5278 8134 5306
rect 8162 5278 14686 5306
rect 14714 5278 14719 5306
rect 8689 5222 8694 5250
rect 8722 5222 14014 5250
rect 14042 5222 14047 5250
rect 0 5194 56 5208
rect 15792 5194 15848 5208
rect 0 5166 6790 5194
rect 6818 5166 6823 5194
rect 15129 5166 15134 5194
rect 15162 5166 15848 5194
rect 0 5152 56 5166
rect 15792 5152 15848 5166
rect 4657 5110 4662 5138
rect 4690 5110 9310 5138
rect 9338 5110 9343 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 5054 5054 7854 5082
rect 7882 5054 7887 5082
rect 9137 5054 9142 5082
rect 9170 5054 10542 5082
rect 10570 5054 10575 5082
rect 0 4970 56 4984
rect 5054 4970 5082 5054
rect 15792 4970 15848 4984
rect 0 4942 5082 4970
rect 7569 4942 7574 4970
rect 7602 4942 14798 4970
rect 14826 4942 14831 4970
rect 15185 4942 15190 4970
rect 15218 4942 15848 4970
rect 0 4928 56 4942
rect 15792 4928 15848 4942
rect 7625 4886 7630 4914
rect 7658 4886 14742 4914
rect 14770 4886 14775 4914
rect 5441 4830 5446 4858
rect 5474 4830 8638 4858
rect 8666 4830 8671 4858
rect 8745 4830 8750 4858
rect 8778 4830 14686 4858
rect 14714 4830 14719 4858
rect 1666 4774 7350 4802
rect 7378 4774 7383 4802
rect 7457 4774 7462 4802
rect 7490 4774 13118 4802
rect 13146 4774 13151 4802
rect 0 4746 56 4760
rect 1666 4746 1694 4774
rect 15792 4746 15848 4760
rect 0 4718 1694 4746
rect 15073 4718 15078 4746
rect 15106 4718 15848 4746
rect 0 4704 56 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 15792 4704 15848 4718
rect 8633 4662 8638 4690
rect 8666 4662 10794 4690
rect 10766 4634 10794 4662
rect 1353 4606 1358 4634
rect 1386 4606 10486 4634
rect 10514 4606 10519 4634
rect 10766 4606 13062 4634
rect 13090 4606 13095 4634
rect 737 4550 742 4578
rect 770 4550 8918 4578
rect 8946 4550 8951 4578
rect 9697 4550 9702 4578
rect 9730 4550 13342 4578
rect 13370 4550 13375 4578
rect 0 4522 56 4536
rect 15792 4522 15848 4536
rect 0 4494 8470 4522
rect 8498 4494 8503 4522
rect 8857 4494 8862 4522
rect 8890 4494 14686 4522
rect 14714 4494 14719 4522
rect 15185 4494 15190 4522
rect 15218 4494 15848 4522
rect 0 4480 56 4494
rect 15792 4480 15848 4494
rect 2977 4438 2982 4466
rect 3010 4438 7686 4466
rect 7714 4438 7719 4466
rect 5889 4382 5894 4410
rect 5922 4382 7350 4410
rect 7378 4382 7383 4410
rect 7546 4382 11606 4410
rect 11634 4382 11639 4410
rect 7546 4354 7574 4382
rect 5217 4326 5222 4354
rect 5250 4326 7574 4354
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 15792 4298 15848 4312
rect 0 4270 1694 4298
rect 5329 4270 5334 4298
rect 5362 4270 7462 4298
rect 7490 4270 7495 4298
rect 7569 4270 7574 4298
rect 7602 4270 10934 4298
rect 10962 4270 10967 4298
rect 12553 4270 12558 4298
rect 12586 4270 13622 4298
rect 13650 4270 13655 4298
rect 15073 4270 15078 4298
rect 15106 4270 15848 4298
rect 0 4256 56 4270
rect 1666 4242 1694 4270
rect 15792 4256 15848 4270
rect 1666 4214 8582 4242
rect 8610 4214 8615 4242
rect 9193 4214 9198 4242
rect 9226 4214 9982 4242
rect 10010 4214 10015 4242
rect 177 4158 182 4186
rect 210 4158 1694 4186
rect 6561 4158 6566 4186
rect 6594 4158 7126 4186
rect 7154 4158 7159 4186
rect 8353 4158 8358 4186
rect 8386 4158 10430 4186
rect 10458 4158 10463 4186
rect 10593 4158 10598 4186
rect 10626 4158 11438 4186
rect 11466 4158 11471 4186
rect 12665 4158 12670 4186
rect 12698 4158 13902 4186
rect 13930 4158 13935 4186
rect 1666 4130 1694 4158
rect 1666 4102 6734 4130
rect 6762 4102 6767 4130
rect 7513 4102 7518 4130
rect 7546 4102 10962 4130
rect 11825 4102 11830 4130
rect 11858 4102 13342 4130
rect 13370 4102 13375 4130
rect 0 4074 56 4088
rect 10934 4074 10962 4102
rect 15792 4074 15848 4088
rect 0 4046 5894 4074
rect 5922 4046 5927 4074
rect 7457 4046 7462 4074
rect 7490 4046 10822 4074
rect 10850 4046 10855 4074
rect 10934 4046 12614 4074
rect 12642 4046 12647 4074
rect 15129 4046 15134 4074
rect 15162 4046 15848 4074
rect 0 4032 56 4046
rect 15792 4032 15848 4046
rect 8745 3990 8750 4018
rect 8778 3990 14686 4018
rect 14714 3990 14719 4018
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 6841 3878 6846 3906
rect 6874 3878 11718 3906
rect 11746 3878 11751 3906
rect 0 3850 56 3864
rect 15792 3850 15848 3864
rect 0 3822 8470 3850
rect 8498 3822 8503 3850
rect 15185 3822 15190 3850
rect 15218 3822 15848 3850
rect 0 3808 56 3822
rect 15792 3808 15848 3822
rect 9921 3766 9926 3794
rect 9954 3766 11382 3794
rect 11410 3766 11415 3794
rect 1353 3710 1358 3738
rect 1386 3710 8190 3738
rect 8218 3710 8223 3738
rect 4265 3654 4270 3682
rect 4298 3654 9478 3682
rect 9506 3654 9511 3682
rect 0 3626 56 3640
rect 15792 3626 15848 3640
rect 0 3598 7182 3626
rect 7210 3598 7215 3626
rect 15185 3598 15190 3626
rect 15218 3598 15848 3626
rect 0 3584 56 3598
rect 15792 3584 15848 3598
rect 3985 3542 3990 3570
rect 4018 3542 9758 3570
rect 9786 3542 9791 3570
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 4321 3486 4326 3514
rect 4354 3486 7574 3514
rect 8017 3486 8022 3514
rect 8050 3486 11270 3514
rect 11298 3486 11303 3514
rect 7546 3458 7574 3486
rect 5049 3430 5054 3458
rect 5082 3430 7434 3458
rect 7546 3430 9366 3458
rect 9394 3430 9399 3458
rect 10873 3430 10878 3458
rect 10906 3430 11438 3458
rect 11466 3430 11471 3458
rect 13393 3430 13398 3458
rect 13426 3430 13734 3458
rect 13762 3430 13767 3458
rect 0 3402 56 3416
rect 7406 3402 7434 3430
rect 15792 3402 15848 3416
rect 0 3374 7294 3402
rect 7322 3374 7327 3402
rect 7406 3374 8414 3402
rect 8442 3374 8447 3402
rect 15129 3374 15134 3402
rect 15162 3374 15848 3402
rect 0 3360 56 3374
rect 15792 3360 15848 3374
rect 4153 3318 4158 3346
rect 4186 3318 9702 3346
rect 9730 3318 9735 3346
rect 10929 3318 10934 3346
rect 10962 3318 12166 3346
rect 12194 3318 12199 3346
rect 9529 3262 9534 3290
rect 9562 3262 9926 3290
rect 9954 3262 9959 3290
rect 10542 3262 13902 3290
rect 13930 3262 13935 3290
rect 10542 3234 10570 3262
rect 1666 3206 7014 3234
rect 7042 3206 7047 3234
rect 7289 3206 7294 3234
rect 7322 3206 10570 3234
rect 10817 3206 10822 3234
rect 10850 3206 14686 3234
rect 14714 3206 14719 3234
rect 0 3178 56 3192
rect 1666 3178 1694 3206
rect 15792 3178 15848 3192
rect 0 3150 1694 3178
rect 14401 3150 14406 3178
rect 14434 3150 15848 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 15792 3136 15848 3150
rect 12833 3094 12838 3122
rect 12866 3094 14294 3122
rect 14322 3094 14327 3122
rect 5609 3038 5614 3066
rect 5642 3038 10822 3066
rect 10850 3038 10855 3066
rect 11102 3038 13902 3066
rect 13930 3038 13935 3066
rect 11102 3010 11130 3038
rect 8745 2982 8750 3010
rect 8778 2982 11130 3010
rect 11321 2982 11326 3010
rect 11354 2982 12054 3010
rect 12082 2982 12087 3010
rect 12609 2982 12614 3010
rect 12642 2982 14686 3010
rect 14714 2982 14719 3010
rect 0 2954 56 2968
rect 15792 2954 15848 2968
rect 0 2926 7294 2954
rect 7322 2926 7327 2954
rect 9137 2926 9142 2954
rect 9170 2926 12894 2954
rect 12922 2926 12927 2954
rect 13001 2926 13006 2954
rect 13034 2926 14294 2954
rect 14322 2926 14327 2954
rect 15073 2926 15078 2954
rect 15106 2926 15848 2954
rect 0 2912 56 2926
rect 15792 2912 15848 2926
rect 7793 2870 7798 2898
rect 7826 2870 14742 2898
rect 14770 2870 14775 2898
rect 5833 2814 5838 2842
rect 5866 2814 10374 2842
rect 10402 2814 10407 2842
rect 12329 2814 12334 2842
rect 12362 2814 12446 2842
rect 12474 2814 12479 2842
rect 3201 2758 3206 2786
rect 3234 2758 7350 2786
rect 7378 2758 7383 2786
rect 7457 2758 7462 2786
rect 7490 2758 8918 2786
rect 8946 2758 8951 2786
rect 9585 2758 9590 2786
rect 9618 2758 11578 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 0 2702 1694 2730
rect 4937 2702 4942 2730
rect 4970 2702 6958 2730
rect 6986 2702 6991 2730
rect 7961 2702 7966 2730
rect 7994 2702 11438 2730
rect 11466 2702 11471 2730
rect 0 2688 56 2702
rect 1666 2674 1694 2702
rect 11550 2674 11578 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 15792 2730 15848 2744
rect 15129 2702 15134 2730
rect 15162 2702 15848 2730
rect 15792 2688 15848 2702
rect 1666 2646 5054 2674
rect 5082 2646 5087 2674
rect 6729 2646 6734 2674
rect 6762 2646 8470 2674
rect 8498 2646 8503 2674
rect 11550 2646 13174 2674
rect 13202 2646 13207 2674
rect 4545 2590 4550 2618
rect 4578 2590 8862 2618
rect 8890 2590 8895 2618
rect 11265 2590 11270 2618
rect 11298 2590 12558 2618
rect 12586 2590 12591 2618
rect 3257 2534 3262 2562
rect 3290 2534 6846 2562
rect 6874 2534 6879 2562
rect 6953 2534 6958 2562
rect 6986 2534 7798 2562
rect 7826 2534 7831 2562
rect 10929 2534 10934 2562
rect 10962 2534 11718 2562
rect 11746 2534 11751 2562
rect 12889 2534 12894 2562
rect 12922 2534 13230 2562
rect 13258 2534 13263 2562
rect 0 2506 56 2520
rect 15792 2506 15848 2520
rect 0 2478 182 2506
rect 210 2478 215 2506
rect 8521 2478 8526 2506
rect 8554 2478 13118 2506
rect 13146 2478 13151 2506
rect 14401 2478 14406 2506
rect 14434 2478 15848 2506
rect 0 2464 56 2478
rect 15792 2464 15848 2478
rect 10369 2422 10374 2450
rect 10402 2422 10766 2450
rect 10794 2422 10799 2450
rect 10878 2422 14742 2450
rect 14770 2422 14775 2450
rect 10878 2394 10906 2422
rect 8353 2366 8358 2394
rect 8386 2366 10906 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 6561 2310 6566 2338
rect 6594 2310 9170 2338
rect 0 2282 56 2296
rect 9142 2282 9170 2310
rect 15792 2282 15848 2296
rect 0 2254 8078 2282
rect 8106 2254 8111 2282
rect 9142 2254 13510 2282
rect 13538 2254 13543 2282
rect 15185 2254 15190 2282
rect 15218 2254 15848 2282
rect 0 2240 56 2254
rect 15792 2240 15848 2254
rect 2921 2198 2926 2226
rect 2954 2198 7294 2226
rect 7322 2198 7327 2226
rect 8689 2198 8694 2226
rect 8722 2198 14686 2226
rect 14714 2198 14719 2226
rect 4601 2142 4606 2170
rect 4634 2142 5894 2170
rect 5922 2142 5927 2170
rect 9753 2142 9758 2170
rect 9786 2142 10934 2170
rect 10962 2142 10967 2170
rect 5497 2086 5502 2114
rect 5530 2086 6678 2114
rect 6706 2086 6711 2114
rect 11713 2086 11718 2114
rect 11746 2086 12166 2114
rect 12194 2086 12199 2114
rect 0 2058 56 2072
rect 15792 2058 15848 2072
rect 0 2030 6230 2058
rect 6258 2030 6263 2058
rect 6449 2030 6454 2058
rect 6482 2030 11886 2058
rect 11914 2030 11919 2058
rect 11998 2030 12334 2058
rect 12362 2030 12367 2058
rect 15129 2030 15134 2058
rect 15162 2030 15848 2058
rect 0 2016 56 2030
rect 11998 2002 12026 2030
rect 15792 2016 15848 2030
rect 5497 1974 5502 2002
rect 5530 1974 8582 2002
rect 8610 1974 8615 2002
rect 9249 1974 9254 2002
rect 9282 1974 12026 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 4713 1918 4718 1946
rect 4746 1918 9646 1946
rect 9674 1918 9679 1946
rect 10873 1918 10878 1946
rect 10906 1918 11046 1946
rect 11074 1918 11079 1946
rect 5553 1862 5558 1890
rect 5586 1862 9002 1890
rect 0 1834 56 1848
rect 0 1806 8414 1834
rect 8442 1806 8447 1834
rect 0 1792 56 1806
rect 8974 1778 9002 1862
rect 9086 1862 9478 1890
rect 9506 1862 9511 1890
rect 9086 1834 9114 1862
rect 15792 1834 15848 1848
rect 9081 1806 9086 1834
rect 9114 1806 9119 1834
rect 14289 1806 14294 1834
rect 14322 1806 15848 1834
rect 15792 1792 15848 1806
rect 793 1750 798 1778
rect 826 1750 1694 1778
rect 3425 1750 3430 1778
rect 3458 1750 5782 1778
rect 5810 1750 5815 1778
rect 6113 1750 6118 1778
rect 6146 1750 8526 1778
rect 8554 1750 8559 1778
rect 8974 1750 12278 1778
rect 12306 1750 12311 1778
rect 1666 1722 1694 1750
rect 1666 1694 4550 1722
rect 4578 1694 4583 1722
rect 4993 1694 4998 1722
rect 5026 1694 6734 1722
rect 6762 1694 6767 1722
rect 8633 1694 8638 1722
rect 8666 1694 13902 1722
rect 13930 1694 13935 1722
rect 1806 1638 4942 1666
rect 4970 1638 4975 1666
rect 6169 1638 6174 1666
rect 6202 1638 8750 1666
rect 8778 1638 8783 1666
rect 8857 1638 8862 1666
rect 8890 1638 13118 1666
rect 13146 1638 13151 1666
rect 0 1610 56 1624
rect 1806 1610 1834 1638
rect 15792 1610 15848 1624
rect 0 1582 1834 1610
rect 7401 1582 7406 1610
rect 7434 1582 9982 1610
rect 10010 1582 10015 1610
rect 15073 1582 15078 1610
rect 15106 1582 15848 1610
rect 0 1568 56 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 15792 1568 15848 1582
rect 3369 1526 3374 1554
rect 3402 1526 8190 1554
rect 8218 1526 8223 1554
rect 8745 1526 8750 1554
rect 8778 1526 11550 1554
rect 11578 1526 11583 1554
rect 4825 1470 4830 1498
rect 4858 1470 7462 1498
rect 7490 1470 7495 1498
rect 10425 1470 10430 1498
rect 10458 1470 11886 1498
rect 11914 1470 11919 1498
rect 2697 1414 2702 1442
rect 2730 1414 4774 1442
rect 4802 1414 4807 1442
rect 9193 1414 9198 1442
rect 9226 1414 11298 1442
rect 11489 1414 11494 1442
rect 11522 1414 11718 1442
rect 11746 1414 11751 1442
rect 13426 1414 13902 1442
rect 13930 1414 13935 1442
rect 0 1386 56 1400
rect 11270 1386 11298 1414
rect 13426 1386 13454 1414
rect 15792 1386 15848 1400
rect 0 1358 798 1386
rect 826 1358 831 1386
rect 6057 1358 6062 1386
rect 6090 1358 7406 1386
rect 7434 1358 7439 1386
rect 8017 1358 8022 1386
rect 8050 1358 9338 1386
rect 10593 1358 10598 1386
rect 10626 1358 11158 1386
rect 11186 1358 11191 1386
rect 11270 1358 13454 1386
rect 13505 1358 13510 1386
rect 13538 1358 14686 1386
rect 14714 1358 14719 1386
rect 15185 1358 15190 1386
rect 15218 1358 15848 1386
rect 0 1344 56 1358
rect 9310 1330 9338 1358
rect 15792 1344 15848 1358
rect 5217 1302 5222 1330
rect 5250 1302 6454 1330
rect 6482 1302 6487 1330
rect 8633 1302 8638 1330
rect 8666 1302 9198 1330
rect 9226 1302 9231 1330
rect 9310 1302 11214 1330
rect 11242 1302 11247 1330
rect 11713 1302 11718 1330
rect 11746 1302 12950 1330
rect 12978 1302 12983 1330
rect 3481 1246 3486 1274
rect 3514 1246 4942 1274
rect 4970 1246 4975 1274
rect 6057 1246 6062 1274
rect 6090 1246 9758 1274
rect 9786 1246 9791 1274
rect 10430 1246 13342 1274
rect 13370 1246 13375 1274
rect 10430 1218 10458 1246
rect 2529 1190 2534 1218
rect 2562 1190 5894 1218
rect 5922 1190 5927 1218
rect 6113 1190 6118 1218
rect 6146 1190 10458 1218
rect 10649 1190 10654 1218
rect 10682 1190 12166 1218
rect 12194 1190 12199 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 15792 1162 15848 1176
rect 0 1134 742 1162
rect 770 1134 775 1162
rect 5049 1134 5054 1162
rect 5082 1134 10318 1162
rect 10346 1134 10351 1162
rect 11545 1134 11550 1162
rect 11578 1134 11718 1162
rect 11746 1134 11751 1162
rect 14401 1134 14406 1162
rect 14434 1134 15848 1162
rect 0 1120 56 1134
rect 15792 1120 15848 1134
rect 5441 1078 5446 1106
rect 5474 1078 9310 1106
rect 9338 1078 9343 1106
rect 10425 1078 10430 1106
rect 10458 1078 12614 1106
rect 12642 1078 12647 1106
rect 4769 1022 4774 1050
rect 4802 1022 5894 1050
rect 5922 1022 5927 1050
rect 9529 1022 9534 1050
rect 9562 1022 11102 1050
rect 11130 1022 11135 1050
rect 11209 1022 11214 1050
rect 11242 1022 14686 1050
rect 14714 1022 14719 1050
rect 3705 966 3710 994
rect 3738 966 4550 994
rect 4578 966 4583 994
rect 5721 966 5726 994
rect 5754 966 6510 994
rect 6538 966 6543 994
rect 9025 966 9030 994
rect 9058 966 9198 994
rect 9226 966 9231 994
rect 10033 966 10038 994
rect 10066 966 10766 994
rect 10794 966 10799 994
rect 11041 966 11046 994
rect 11074 966 11802 994
rect 0 938 56 952
rect 11774 938 11802 966
rect 15792 938 15848 952
rect 0 910 2982 938
rect 3010 910 3015 938
rect 5161 910 5166 938
rect 5194 910 6454 938
rect 6482 910 6487 938
rect 7233 910 7238 938
rect 7266 910 7574 938
rect 7602 910 7607 938
rect 8073 910 8078 938
rect 8106 910 8470 938
rect 8498 910 8503 938
rect 9417 910 9422 938
rect 9450 910 10598 938
rect 10626 910 10631 938
rect 11531 910 11550 938
rect 11578 910 11583 938
rect 11769 910 11774 938
rect 11802 910 11807 938
rect 12665 910 12670 938
rect 12698 910 13454 938
rect 13482 910 13487 938
rect 14345 910 14350 938
rect 14378 910 15848 938
rect 0 896 56 910
rect 15792 896 15848 910
rect 5217 854 5222 882
rect 5250 854 6174 882
rect 6202 854 6207 882
rect 6393 854 6398 882
rect 6426 854 6902 882
rect 6930 854 6935 882
rect 7406 854 7742 882
rect 7770 854 7775 882
rect 8353 854 8358 882
rect 8386 854 8694 882
rect 8722 854 8727 882
rect 8969 854 8974 882
rect 9002 854 10262 882
rect 10290 854 10295 882
rect 11657 854 11662 882
rect 11690 854 12110 882
rect 12138 854 12143 882
rect 12777 854 12782 882
rect 12810 854 13678 882
rect 13706 854 13711 882
rect 7406 826 7434 854
rect 4041 798 4046 826
rect 4074 798 6342 826
rect 6370 798 6375 826
rect 6617 798 6622 826
rect 6650 798 6958 826
rect 6986 798 6991 826
rect 7401 798 7406 826
rect 7434 798 7439 826
rect 7961 798 7966 826
rect 7994 798 8442 826
rect 9641 798 9646 826
rect 9674 798 10542 826
rect 10570 798 10575 826
rect 10654 798 11522 826
rect 11713 798 11718 826
rect 11746 798 11774 826
rect 11802 798 11807 826
rect 13225 798 13230 826
rect 13258 798 14686 826
rect 14714 798 14719 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 8414 770 8442 798
rect 10654 770 10682 798
rect 3761 742 3766 770
rect 3794 742 8302 770
rect 8330 742 8335 770
rect 8414 742 10682 770
rect 10929 742 10934 770
rect 10962 742 11214 770
rect 11242 742 11247 770
rect 0 714 56 728
rect 0 686 2114 714
rect 2809 686 2814 714
rect 2842 686 4494 714
rect 4522 686 4527 714
rect 5385 686 5390 714
rect 5418 686 10822 714
rect 10850 686 10855 714
rect 0 672 56 686
rect 2086 546 2114 686
rect 11494 658 11522 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 15792 714 15848 728
rect 11657 686 11662 714
rect 11690 686 13062 714
rect 13090 686 13095 714
rect 13617 686 13622 714
rect 13650 686 15848 714
rect 15792 672 15848 686
rect 3593 630 3598 658
rect 3626 630 4830 658
rect 4858 630 4863 658
rect 5665 630 5670 658
rect 5698 630 6398 658
rect 6426 630 6431 658
rect 7009 630 7014 658
rect 7042 630 7294 658
rect 7322 630 7327 658
rect 7518 630 10430 658
rect 10458 630 10463 658
rect 10537 630 10542 658
rect 10570 630 11382 658
rect 11410 630 11415 658
rect 11494 630 13454 658
rect 3369 574 3374 602
rect 3402 574 6566 602
rect 6594 574 6599 602
rect 2086 518 4214 546
rect 4713 518 4718 546
rect 4746 518 5334 546
rect 5362 518 5367 546
rect 5441 518 5446 546
rect 5474 518 5614 546
rect 5642 518 5647 546
rect 5721 518 5726 546
rect 5754 518 6846 546
rect 6874 518 6879 546
rect 0 490 56 504
rect 4186 490 4214 518
rect 7518 490 7546 630
rect 13426 602 13454 630
rect 10201 574 10206 602
rect 10234 574 11494 602
rect 11522 574 11527 602
rect 13426 574 13902 602
rect 13930 574 13935 602
rect 7625 518 7630 546
rect 7658 518 7966 546
rect 7994 518 7999 546
rect 8078 518 9254 546
rect 9282 518 9287 546
rect 9865 518 9870 546
rect 9898 518 10486 546
rect 10514 518 10519 546
rect 10598 518 12726 546
rect 12754 518 12759 546
rect 0 462 2170 490
rect 3593 462 3598 490
rect 3626 462 3822 490
rect 3850 462 3855 490
rect 4186 462 4858 490
rect 5161 462 5166 490
rect 5194 462 6286 490
rect 6314 462 6319 490
rect 6398 462 7546 490
rect 0 448 56 462
rect 0 266 56 280
rect 0 238 1358 266
rect 1386 238 1391 266
rect 0 224 56 238
rect 2142 154 2170 462
rect 4830 434 4858 462
rect 6398 434 6426 462
rect 8078 434 8106 518
rect 10598 490 10626 518
rect 15792 490 15848 504
rect 8185 462 8190 490
rect 8218 462 8582 490
rect 8610 462 8615 490
rect 8857 462 8862 490
rect 8890 462 10318 490
rect 10346 462 10351 490
rect 10425 462 10430 490
rect 10458 462 10626 490
rect 12217 462 12222 490
rect 12250 462 12558 490
rect 12586 462 12591 490
rect 13337 462 13342 490
rect 13370 462 15848 490
rect 15792 448 15848 462
rect 3145 406 3150 434
rect 3178 406 3934 434
rect 3962 406 3967 434
rect 4097 406 4102 434
rect 4130 406 4718 434
rect 4746 406 4751 434
rect 4830 406 5502 434
rect 5530 406 5535 434
rect 5609 406 5614 434
rect 5642 406 6426 434
rect 7177 406 7182 434
rect 7210 406 7518 434
rect 7546 406 7551 434
rect 7630 406 8106 434
rect 8521 406 8526 434
rect 8554 406 9310 434
rect 9338 406 9343 434
rect 9977 406 9982 434
rect 10010 406 11438 434
rect 11466 406 11471 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 7630 378 7658 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 3593 350 3598 378
rect 3626 350 5110 378
rect 5138 350 5143 378
rect 5222 350 7658 378
rect 9198 350 11550 378
rect 11578 350 11583 378
rect 2921 294 2926 322
rect 2954 294 4438 322
rect 4466 294 4471 322
rect 3033 238 3038 266
rect 3066 238 3766 266
rect 3794 238 3799 266
rect 5222 154 5250 350
rect 9198 322 9226 350
rect 5945 294 5950 322
rect 5978 294 9226 322
rect 9305 294 9310 322
rect 9338 294 9926 322
rect 9954 294 9959 322
rect 11433 294 11438 322
rect 11466 294 11662 322
rect 11690 294 11695 322
rect 12329 294 12334 322
rect 12362 294 12446 322
rect 12474 294 12479 322
rect 15792 266 15848 280
rect 6953 238 6958 266
rect 6986 238 7630 266
rect 7658 238 7663 266
rect 8409 238 8414 266
rect 8442 238 9366 266
rect 9394 238 9399 266
rect 10089 238 10094 266
rect 10122 238 12054 266
rect 12082 238 12087 266
rect 13561 238 13566 266
rect 13594 238 15848 266
rect 15792 224 15848 238
rect 5721 182 5726 210
rect 5754 182 7966 210
rect 7994 182 7999 210
rect 9193 182 9198 210
rect 9226 182 11046 210
rect 11074 182 11079 210
rect 2142 126 4662 154
rect 4690 126 4695 154
rect 5161 126 5166 154
rect 5194 126 5250 154
rect 9137 126 9142 154
rect 9170 126 9175 154
rect 10257 126 10262 154
rect 10290 126 11998 154
rect 12026 126 12031 154
rect 9142 98 9170 126
rect 4489 70 4494 98
rect 4522 70 7462 98
rect 7490 70 7495 98
rect 9142 70 11886 98
rect 11914 70 11919 98
rect 0 42 56 56
rect 15792 42 15848 56
rect 0 14 2534 42
rect 2562 14 2567 42
rect 13841 14 13846 42
rect 13874 14 15848 42
rect 0 0 56 14
rect 15792 0 15848 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 2142 5838 2170 5866
rect 2142 5558 2170 5586
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 8638 4830 8666 4858
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 8638 4662 8666 4690
rect 5894 4382 5922 4410
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 7462 4270 7490 4298
rect 7574 4270 7602 4298
rect 5894 4046 5922 4074
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 11718 3878 11746 3906
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 12446 2814 12474 2842
rect 7462 2758 7490 2786
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 6958 2702 6986 2730
rect 7966 2702 7994 2730
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 6958 2534 6986 2562
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 6454 2030 6482 2058
rect 9254 1974 9282 2002
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 8750 1638 8778 1666
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 8750 1526 8778 1554
rect 11214 1302 11242 1330
rect 2534 1190 2562 1218
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 11214 1022 11242 1050
rect 6454 910 6482 938
rect 11550 910 11578 938
rect 11718 798 11746 826
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 10430 630 10458 658
rect 9254 518 9282 546
rect 10430 462 10458 490
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 11550 350 11578 378
rect 12446 294 12474 322
rect 7966 182 7994 210
rect 7462 70 7490 98
rect 2534 14 2562 42
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 2142 5866 2170 5871
rect 2142 5586 2170 5838
rect 2142 5553 2170 5558
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 5110 2378 5866
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 8638 4858 8666 4863
rect 8638 4690 8666 4830
rect 8638 4657 8666 4662
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 5894 4410 5922 4415
rect 5894 4074 5922 4382
rect 7462 4298 7490 4303
rect 7574 4298 7602 4303
rect 7490 4270 7574 4289
rect 7462 4261 7602 4270
rect 5894 4041 5922 4046
rect 11888 3934 12048 4690
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 11718 3906 11746 3911
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 7462 2786 7490 2791
rect 2218 1974 2378 2730
rect 6958 2730 6986 2735
rect 6958 2562 6986 2702
rect 6958 2529 6986 2534
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 6454 2058 6482 2063
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 2534 1218 2562 1223
rect 2534 42 2562 1190
rect 6454 938 6482 2030
rect 6454 905 6482 910
rect 7462 98 7490 2758
rect 7966 2730 7994 2735
rect 7966 210 7994 2702
rect 9254 2002 9282 2007
rect 8750 1666 8778 1671
rect 8750 1554 8778 1638
rect 8750 1521 8778 1526
rect 9254 546 9282 1974
rect 11214 1330 11242 1335
rect 11214 1050 11242 1302
rect 11214 1017 11242 1022
rect 11550 938 11578 943
rect 9254 513 9282 518
rect 10430 658 10458 663
rect 10430 490 10458 630
rect 10430 457 10458 462
rect 11550 378 11578 910
rect 11718 826 11746 3878
rect 11718 793 11746 798
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 11888 798 12048 1554
rect 11550 345 11578 350
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 7966 177 7994 182
rect 7462 65 7490 70
rect 2534 9 2562 14
rect 11888 0 12048 770
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 12446 2842 12474 2847
rect 12446 322 12474 2814
rect 12446 289 12474 294
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _00_
timestamp 1486834041
transform 1 0 5768 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _01_
timestamp 1486834041
transform 1 0 8120 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _02_
timestamp 1486834041
transform 1 0 9240 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _03_
timestamp 1486834041
transform 1 0 8512 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _04_
timestamp 1486834041
transform 1 0 7672 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _05_
timestamp 1486834041
transform 1 0 8848 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _06_
timestamp 1486834041
transform 1 0 8792 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _07_
timestamp 1486834041
transform 1 0 7728 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _08_
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _09_
timestamp 1486834041
transform 1 0 6160 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _10_
timestamp 1486834041
transform 1 0 8008 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _11_
timestamp 1486834041
transform 1 0 8400 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _12_
timestamp 1486834041
transform 1 0 8344 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _13_
timestamp 1486834041
transform 1 0 7448 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _14_
timestamp 1486834041
transform 1 0 6944 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _15_
timestamp 1486834041
transform 1 0 7224 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _16_
timestamp 1486834041
transform 1 0 7112 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _17_
timestamp 1486834041
transform 1 0 8400 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _18_
timestamp 1486834041
transform 1 0 7280 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _19_
timestamp 1486834041
transform 1 0 8512 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _20_
timestamp 1486834041
transform 1 0 8400 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _21_
timestamp 1486834041
transform 1 0 7280 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _22_
timestamp 1486834041
transform 1 0 7784 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _23_
timestamp 1486834041
transform 1 0 6720 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _24_
timestamp 1486834041
transform 1 0 8344 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _25_
timestamp 1486834041
transform 1 0 7168 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _26_
timestamp 1486834041
transform 1 0 7616 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _27_
timestamp 1486834041
transform 1 0 8680 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _28_
timestamp 1486834041
transform 1 0 8400 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _29_
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _30_
timestamp 1486834041
transform 1 0 7224 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _31_
timestamp 1486834041
transform 1 0 9352 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _32_
timestamp 1486834041
transform 1 0 11088 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _33_
timestamp 1486834041
transform -1 0 11088 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _34_
timestamp 1486834041
transform -1 0 10808 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _35_
timestamp 1486834041
transform -1 0 9912 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _36_
timestamp 1486834041
transform -1 0 8120 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _37_
timestamp 1486834041
transform -1 0 5544 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _38_
timestamp 1486834041
transform -1 0 5320 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _39_
timestamp 1486834041
transform -1 0 6216 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _40_
timestamp 1486834041
transform -1 0 6944 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _41_
timestamp 1486834041
transform -1 0 9352 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _42_
timestamp 1486834041
transform -1 0 10360 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _43_
timestamp 1486834041
transform -1 0 11760 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _44_
timestamp 1486834041
transform -1 0 11816 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _45_
timestamp 1486834041
transform -1 0 12432 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _46_
timestamp 1486834041
transform -1 0 12712 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _47_
timestamp 1486834041
transform 1 0 13272 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _48_
timestamp 1486834041
transform 1 0 13384 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _49_
timestamp 1486834041
transform 1 0 13608 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _50_
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _51_
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _52_
timestamp 1486834041
transform 1 0 3696 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _53_
timestamp 1486834041
transform 1 0 4368 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _54_
timestamp 1486834041
transform 1 0 4424 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _55_
timestamp 1486834041
transform 1 0 4704 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _56_
timestamp 1486834041
transform -1 0 3248 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _57_
timestamp 1486834041
transform -1 0 3696 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _58_
timestamp 1486834041
transform 1 0 4480 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _59_
timestamp 1486834041
transform 1 0 5152 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _60_
timestamp 1486834041
transform 1 0 4872 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _61_
timestamp 1486834041
transform 1 0 5712 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _62_
timestamp 1486834041
transform 1 0 6776 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _63_
timestamp 1486834041
transform 1 0 7280 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _64_
timestamp 1486834041
transform -1 0 3696 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _65_
timestamp 1486834041
transform -1 0 4144 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _66_
timestamp 1486834041
transform 1 0 5768 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _67_
timestamp 1486834041
transform 1 0 8848 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _68_
timestamp 1486834041
transform 1 0 9296 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _69_
timestamp 1486834041
transform 1 0 9408 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _70_
timestamp 1486834041
transform 1 0 9632 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _71_
timestamp 1486834041
transform 1 0 9688 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _72_
timestamp 1486834041
transform 1 0 7000 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _73_
timestamp 1486834041
transform -1 0 5824 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _74_
timestamp 1486834041
transform -1 0 5768 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _75_
timestamp 1486834041
transform -1 0 5264 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _76_
timestamp 1486834041
transform -1 0 5376 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _77_
timestamp 1486834041
transform 1 0 9688 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _78_
timestamp 1486834041
transform 1 0 11480 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _79_
timestamp 1486834041
transform 1 0 10304 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _80_
timestamp 1486834041
transform 1 0 11368 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _81_
timestamp 1486834041
transform 1 0 12600 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _82_
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _83_
timestamp 1486834041
transform 1 0 10752 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _84_
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _85_
timestamp 1486834041
transform 1 0 12264 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _86_
timestamp 1486834041
transform 1 0 11816 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _87_
timestamp 1486834041
transform 1 0 10080 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _88_
timestamp 1486834041
transform -1 0 10976 0 -1 3528
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140
timestamp 1486834041
transform 1 0 8176 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_169
timestamp 1486834041
transform 1 0 9800 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_200
timestamp 1486834041
transform 1 0 11536 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_220
timestamp 1486834041
transform 1 0 12656 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 4032 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_207
timestamp 1486834041
transform 1 0 11928 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 12040 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_226
timestamp 1486834041
transform 1 0 12992 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_45
timestamp 1486834041
transform 1 0 2856 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_49
timestamp 1486834041
transform 1 0 3080 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_51
timestamp 1486834041
transform 1 0 3192 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_68
timestamp 1486834041
transform 1 0 4144 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_72
timestamp 1486834041
transform 1 0 4368 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_227
timestamp 1486834041
transform 1 0 13048 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_247
timestamp 1486834041
transform 1 0 14168 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1486834041
transform 1 0 4592 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_86
timestamp 1486834041
transform 1 0 5152 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_94
timestamp 1486834041
transform 1 0 5600 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_150
timestamp 1486834041
transform 1 0 8736 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_207
timestamp 1486834041
transform 1 0 11928 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 12040 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_220
timestamp 1486834041
transform 1 0 12656 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_224
timestamp 1486834041
transform 1 0 12880 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_226
timestamp 1486834041
transform 1 0 12992 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_69
timestamp 1486834041
transform 1 0 4200 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_85
timestamp 1486834041
transform 1 0 5096 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_94
timestamp 1486834041
transform 1 0 5600 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_96
timestamp 1486834041
transform 1 0 5712 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_145
timestamp 1486834041
transform 1 0 8456 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_154
timestamp 1486834041
transform 1 0 8960 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_156
timestamp 1486834041
transform 1 0 9072 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 9912 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_221
timestamp 1486834041
transform 1 0 12712 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_237
timestamp 1486834041
transform 1 0 13608 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 4032 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_104
timestamp 1486834041
transform 1 0 6160 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_112
timestamp 1486834041
transform 1 0 6608 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_114
timestamp 1486834041
transform 1 0 6720 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_123
timestamp 1486834041
transform 1 0 7224 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_168
timestamp 1486834041
transform 1 0 9744 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_205
timestamp 1486834041
transform 1 0 11816 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_220
timestamp 1486834041
transform 1 0 12656 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 13552 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1486834041
transform 1 0 13776 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 5992 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1486834041
transform 1 0 6776 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_135
timestamp 1486834041
transform 1 0 7896 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_147
timestamp 1486834041
transform 1 0 8568 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_194
timestamp 1486834041
transform 1 0 11200 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_202
timestamp 1486834041
transform 1 0 11648 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_206
timestamp 1486834041
transform 1 0 11872 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_216
timestamp 1486834041
transform 1 0 12432 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_232
timestamp 1486834041
transform 1 0 13328 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_236
timestamp 1486834041
transform 1 0 13552 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 4032 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_104
timestamp 1486834041
transform 1 0 6160 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_112
timestamp 1486834041
transform 1 0 6608 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_116
timestamp 1486834041
transform 1 0 6832 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_126
timestamp 1486834041
transform 1 0 7392 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_130
timestamp 1486834041
transform 1 0 7616 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 8120 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_142
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_151
timestamp 1486834041
transform 1 0 8792 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_160
timestamp 1486834041
transform 1 0 9296 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_164
timestamp 1486834041
transform 1 0 9520 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_182
timestamp 1486834041
transform 1 0 10528 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_190
timestamp 1486834041
transform 1 0 10976 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_200
timestamp 1486834041
transform 1 0 11536 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_208
timestamp 1486834041
transform 1 0 11984 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_221
timestamp 1486834041
transform 1 0 12712 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_229
timestamp 1486834041
transform 1 0 13160 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1486834041
transform 1 0 4200 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1486834041
transform 1 0 4648 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_89
timestamp 1486834041
transform 1 0 5320 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_131
timestamp 1486834041
transform 1 0 7672 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_147
timestamp 1486834041
transform 1 0 8568 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_151
timestamp 1486834041
transform 1 0 8792 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_161
timestamp 1486834041
transform 1 0 9352 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_170
timestamp 1486834041
transform 1 0 9856 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 10080 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_181
timestamp 1486834041
transform 1 0 10472 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_183
timestamp 1486834041
transform 1 0 10584 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_192
timestamp 1486834041
transform 1 0 11088 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_204
timestamp 1486834041
transform 1 0 11760 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_236
timestamp 1486834041
transform 1 0 13552 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_244
timestamp 1486834041
transform 1 0 14000 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 4032 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_104
timestamp 1486834041
transform 1 0 6160 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_108
timestamp 1486834041
transform 1 0 6384 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_118
timestamp 1486834041
transform 1 0 6944 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_120
timestamp 1486834041
transform 1 0 7056 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_129
timestamp 1486834041
transform 1 0 7560 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_139
timestamp 1486834041
transform 1 0 8120 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_152
timestamp 1486834041
transform 1 0 8848 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_160
timestamp 1486834041
transform 1 0 9296 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_162
timestamp 1486834041
transform 1 0 9408 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_187
timestamp 1486834041
transform 1 0 10808 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_195
timestamp 1486834041
transform 1 0 11256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_205
timestamp 1486834041
transform 1 0 11816 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 12040 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_228
timestamp 1486834041
transform 1 0 13104 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_230
timestamp 1486834041
transform 1 0 13216 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_239
timestamp 1486834041
transform 1 0 13720 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 2240 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_69
timestamp 1486834041
transform 1 0 4200 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_93
timestamp 1486834041
transform 1 0 5544 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 5992 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_123
timestamp 1486834041
transform 1 0 7224 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_132
timestamp 1486834041
transform 1 0 7728 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_140
timestamp 1486834041
transform 1 0 8176 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_144
timestamp 1486834041
transform 1 0 8400 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_154
timestamp 1486834041
transform 1 0 8960 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_170
timestamp 1486834041
transform 1 0 9856 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1486834041
transform 1 0 10080 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_209
timestamp 1486834041
transform 1 0 12040 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_225
timestamp 1486834041
transform 1 0 12936 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_229
timestamp 1486834041
transform 1 0 13160 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_247
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 4032 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_104
timestamp 1486834041
transform 1 0 6160 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_120
timestamp 1486834041
transform 1 0 7056 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_132
timestamp 1486834041
transform 1 0 7728 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_152
timestamp 1486834041
transform 1 0 8848 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_184
timestamp 1486834041
transform 1 0 10640 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_200
timestamp 1486834041
transform 1 0 11536 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_208
timestamp 1486834041
transform 1 0 11984 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_220
timestamp 1486834041
transform 1 0 12656 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_224
timestamp 1486834041
transform 1 0 12880 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_226
timestamp 1486834041
transform 1 0 12992 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1486834041
transform 1 0 5992 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_107
timestamp 1486834041
transform 1 0 6328 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_123
timestamp 1486834041
transform 1 0 7224 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_131
timestamp 1486834041
transform 1 0 7672 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_141
timestamp 1486834041
transform 1 0 8232 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_151
timestamp 1486834041
transform 1 0 8792 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_167
timestamp 1486834041
transform 1 0 9688 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_209
timestamp 1486834041
transform 1 0 12040 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_225
timestamp 1486834041
transform 1 0 12936 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_229
timestamp 1486834041
transform 1 0 13160 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1486834041
transform 1 0 4032 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_104
timestamp 1486834041
transform 1 0 6160 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_112
timestamp 1486834041
transform 1 0 6608 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_138
timestamp 1486834041
transform 1 0 8064 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_152
timestamp 1486834041
transform 1 0 8848 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_184
timestamp 1486834041
transform 1 0 10640 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_200
timestamp 1486834041
transform 1 0 11536 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_208
timestamp 1486834041
transform 1 0 11984 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 2240 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_53
timestamp 1486834041
transform 1 0 3304 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_61
timestamp 1486834041
transform 1 0 3752 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_77
timestamp 1486834041
transform 1 0 4648 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_85
timestamp 1486834041
transform 1 0 5096 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1486834041
transform 1 0 5992 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_131
timestamp 1486834041
transform 1 0 7672 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_157
timestamp 1486834041
transform 1 0 9128 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_173
timestamp 1486834041
transform 1 0 10024 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_177
timestamp 1486834041
transform 1 0 10248 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_193
timestamp 1486834041
transform 1 0 11144 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_209
timestamp 1486834041
transform 1 0 12040 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_247
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_10
timestamp 1486834041
transform 1 0 896 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_65
timestamp 1486834041
transform 1 0 3976 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_67
timestamp 1486834041
transform 1 0 4088 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_146
timestamp 1486834041
transform 1 0 8512 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_169
timestamp 1486834041
transform 1 0 9800 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_200
timestamp 1486834041
transform 1 0 11536 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_206
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_235
timestamp 1486834041
transform 1 0 13496 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_237
timestamp 1486834041
transform 1 0 13608 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_240
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_242
timestamp 1486834041
transform 1 0 13888 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_257
timestamp 1486834041
transform 1 0 14728 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_265
timestamp 1486834041
transform 1 0 15176 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 13272 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 14616 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 13832 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 14616 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 14616 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 13832 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 14616 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 14616 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 14616 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 14616 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 13048 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 14616 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 14616 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 14616 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 14616 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 13832 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 13832 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 13272 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 12488 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 12264 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 13832 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 12880 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 13048 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 13272 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 13048 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 13832 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 13832 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 14616 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 14616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 13832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 14616 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 2240 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform -1 0 9352 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform -1 0 10024 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform -1 0 10752 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform -1 0 11536 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 12040 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 12712 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 13496 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 14056 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform -1 0 14728 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform -1 0 13832 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 3192 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 3976 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 4648 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 5208 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 6384 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 7168 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform -1 0 8680 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 6440 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 5264 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 5824 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 6608 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 7224 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 6552 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 7392 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 6608 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 6384 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 7336 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 7392 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 7168 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 8120 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 8232 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 8344 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 9016 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 9912 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 9688 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 9576 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 9912 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 12656 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 11144 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 11368 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 12992 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 11816 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 11816 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 9128 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 10752 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 9576 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 10696 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 11144 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 10584 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 11032 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 11816 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output89
timestamp 1486834041
transform -1 0 1456 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 15512 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 15512 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 15512 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 15512 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 15512 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 15512 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 15512 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 15512 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 15512 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 15512 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 15512 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 15512 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 15512 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 15512 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 15512 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 15512 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_40
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_41
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_42
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_43
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_44
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_45
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_46
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_47
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_48
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_49
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_50
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_51
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_52
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_53
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_54
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_55
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_56
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_57
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_58
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_59
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_60
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_61
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_62
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_63
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_64
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_65
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_66
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_67
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_68
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_69
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_70
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_71
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_72
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_73
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_74
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_75
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_76
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_77
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_78
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_79
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_80
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_81
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_82
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_83
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_84
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_85
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_86
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_87
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_88
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_89
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_90
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_91
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_92
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_93
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_94
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 15792 0 15848 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 15792 2240 15848 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 15792 2464 15848 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 15792 2688 15848 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 15792 2912 15848 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 15792 3136 15848 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 15792 3360 15848 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 15792 3584 15848 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 15792 3808 15848 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 15792 4032 15848 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 15792 4256 15848 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 15792 224 15848 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 15792 4480 15848 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 15792 4704 15848 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 15792 4928 15848 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 15792 5152 15848 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 15792 5376 15848 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 15792 5600 15848 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 15792 5824 15848 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 15792 6048 15848 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 15792 6272 15848 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 15792 6496 15848 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 15792 448 15848 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 15792 6720 15848 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 15792 6944 15848 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 15792 672 15848 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 15792 896 15848 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 15792 1120 15848 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 15792 1344 15848 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 15792 1568 15848 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 15792 1792 15848 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 15792 2016 15848 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 10864 0 10920 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 11984 0 12040 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 12096 0 12152 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 12208 0 12264 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 12320 0 12376 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 12432 0 12488 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 12544 0 12600 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 12656 0 12712 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 12768 0 12824 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 12880 0 12936 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 12992 0 13048 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 10976 0 11032 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 11088 0 11144 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 11200 0 11256 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 11312 0 11368 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 11424 0 11480 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 11536 0 11592 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 11648 0 11704 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 11760 0 11816 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 11872 0 11928 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 1792 7056 1848 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 8512 7056 8568 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 9184 7056 9240 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 9856 7056 9912 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 10528 7056 10584 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 11200 7056 11256 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 11872 7056 11928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 12544 7056 12600 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 13216 7056 13272 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 13888 7056 13944 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 14560 7056 14616 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 2464 7056 2520 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 3136 7056 3192 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 3808 7056 3864 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 4480 7056 4536 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 5152 7056 5208 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 5824 7056 5880 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 6496 7056 6552 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 7168 7056 7224 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 7840 7056 7896 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2688 0 2744 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 2800 0 2856 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 2912 0 2968 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 3024 0 3080 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 4032 0 4088 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 4144 0 4200 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 4256 0 4312 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 4368 0 4424 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 4480 0 4536 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 4592 0 4648 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 4704 0 4760 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 4816 0 4872 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 3136 0 3192 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 3248 0 3304 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 3360 0 3416 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 3472 0 3528 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 3584 0 3640 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 3696 0 3752 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 3808 0 3864 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 3920 0 3976 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 4928 0 4984 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 6048 0 6104 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 6160 0 6216 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 6272 0 6328 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 6384 0 6440 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 6496 0 6552 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 6608 0 6664 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 5040 0 5096 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 5152 0 5208 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 5264 0 5320 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 5376 0 5432 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 5488 0 5544 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 5600 0 5656 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 5712 0 5768 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 5824 0 5880 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 5936 0 5992 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 6720 0 6776 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 140 nsew signal output
flabel metal2 s 6832 0 6888 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 141 nsew signal output
flabel metal2 s 6944 0 7000 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 142 nsew signal output
flabel metal2 s 7056 0 7112 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 143 nsew signal output
flabel metal2 s 7168 0 7224 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 144 nsew signal output
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 145 nsew signal output
flabel metal2 s 7392 0 7448 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 146 nsew signal output
flabel metal2 s 7504 0 7560 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 147 nsew signal output
flabel metal2 s 7616 0 7672 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 148 nsew signal output
flabel metal2 s 7728 0 7784 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 149 nsew signal output
flabel metal2 s 7840 0 7896 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 150 nsew signal output
flabel metal2 s 7952 0 8008 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 151 nsew signal output
flabel metal2 s 8064 0 8120 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 152 nsew signal output
flabel metal2 s 8176 0 8232 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 153 nsew signal output
flabel metal2 s 8288 0 8344 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 154 nsew signal output
flabel metal2 s 8400 0 8456 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 155 nsew signal output
flabel metal2 s 8512 0 8568 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 156 nsew signal output
flabel metal2 s 8624 0 8680 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 157 nsew signal output
flabel metal2 s 8736 0 8792 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 158 nsew signal output
flabel metal2 s 8848 0 8904 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 159 nsew signal output
flabel metal2 s 8960 0 9016 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 160 nsew signal output
flabel metal2 s 10080 0 10136 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 161 nsew signal output
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 162 nsew signal output
flabel metal2 s 10304 0 10360 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 163 nsew signal output
flabel metal2 s 10416 0 10472 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 164 nsew signal output
flabel metal2 s 10528 0 10584 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 165 nsew signal output
flabel metal2 s 10640 0 10696 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 166 nsew signal output
flabel metal2 s 9072 0 9128 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 167 nsew signal output
flabel metal2 s 9184 0 9240 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 168 nsew signal output
flabel metal2 s 9296 0 9352 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 169 nsew signal output
flabel metal2 s 9408 0 9464 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 170 nsew signal output
flabel metal2 s 9520 0 9576 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 171 nsew signal output
flabel metal2 s 9632 0 9688 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 172 nsew signal output
flabel metal2 s 9744 0 9800 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 173 nsew signal output
flabel metal2 s 9856 0 9912 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 174 nsew signal output
flabel metal2 s 9968 0 10024 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 175 nsew signal output
flabel metal2 s 10752 0 10808 56 0 FreeSans 224 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 1120 7056 1176 7112 0 FreeSans 224 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 178 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 179 nsew ground bidirectional
rlabel metal1 7924 6272 7924 6272 0 VDD
rlabel metal1 7924 6664 7924 6664 0 VSS
rlabel metal3 1295 28 1295 28 0 FrameData[0]
rlabel metal2 8092 2212 8092 2212 0 FrameData[10]
rlabel metal3 119 2492 119 2492 0 FrameData[11]
rlabel metal3 861 2716 861 2716 0 FrameData[12]
rlabel metal2 7308 2968 7308 2968 0 FrameData[13]
rlabel metal3 861 3164 861 3164 0 FrameData[14]
rlabel metal2 7308 3500 7308 3500 0 FrameData[15]
rlabel metal2 7196 3864 7196 3864 0 FrameData[16]
rlabel metal2 8484 3976 8484 3976 0 FrameData[17]
rlabel metal4 5908 4228 5908 4228 0 FrameData[18]
rlabel metal2 8596 4312 8596 4312 0 FrameData[19]
rlabel metal3 707 252 707 252 0 FrameData[1]
rlabel metal2 8484 4704 8484 4704 0 FrameData[20]
rlabel metal3 861 4732 861 4732 0 FrameData[21]
rlabel metal2 7868 5124 7868 5124 0 FrameData[22]
rlabel metal2 6804 5432 6804 5432 0 FrameData[23]
rlabel metal2 8428 5348 8428 5348 0 FrameData[24]
rlabel metal2 7252 5656 7252 5656 0 FrameData[25]
rlabel metal2 7700 5628 7700 5628 0 FrameData[26]
rlabel metal3 4403 6076 4403 6076 0 FrameData[27]
rlabel metal3 427 6300 427 6300 0 FrameData[28]
rlabel metal3 4095 6524 4095 6524 0 FrameData[29]
rlabel metal3 1099 476 1099 476 0 FrameData[2]
rlabel metal2 7308 6412 7308 6412 0 FrameData[30]
rlabel metal3 399 6972 399 6972 0 FrameData[31]
rlabel metal3 1071 700 1071 700 0 FrameData[3]
rlabel metal3 1519 924 1519 924 0 FrameData[4]
rlabel metal3 399 1148 399 1148 0 FrameData[5]
rlabel metal3 427 1372 427 1372 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal2 8428 1792 8428 1792 0 FrameData[8]
rlabel metal2 6244 1960 6244 1960 0 FrameData[9]
rlabel metal3 14833 28 14833 28 0 FrameData_O[0]
rlabel metal2 15204 1988 15204 1988 0 FrameData_O[10]
rlabel metal3 15113 2492 15113 2492 0 FrameData_O[11]
rlabel metal2 15148 2464 15148 2464 0 FrameData_O[12]
rlabel metal2 15092 2772 15092 2772 0 FrameData_O[13]
rlabel metal3 15113 3164 15113 3164 0 FrameData_O[14]
rlabel metal2 15148 3192 15148 3192 0 FrameData_O[15]
rlabel metal2 15204 3444 15204 3444 0 FrameData_O[16]
rlabel metal3 15505 3836 15505 3836 0 FrameData_O[17]
rlabel metal2 15148 3920 15148 3920 0 FrameData_O[18]
rlabel metal3 15449 4284 15449 4284 0 FrameData_O[19]
rlabel metal3 14693 252 14693 252 0 FrameData_O[1]
rlabel metal3 15505 4508 15505 4508 0 FrameData_O[20]
rlabel metal3 15449 4732 15449 4732 0 FrameData_O[21]
rlabel metal3 15505 4956 15505 4956 0 FrameData_O[22]
rlabel metal3 15477 5180 15477 5180 0 FrameData_O[23]
rlabel metal3 15113 5404 15113 5404 0 FrameData_O[24]
rlabel metal2 14308 5292 14308 5292 0 FrameData_O[25]
rlabel metal2 13860 5628 13860 5628 0 FrameData_O[26]
rlabel metal2 13076 6104 13076 6104 0 FrameData_O[27]
rlabel metal2 12852 5964 12852 5964 0 FrameData_O[28]
rlabel metal3 15085 6524 15085 6524 0 FrameData_O[29]
rlabel metal2 13356 504 13356 504 0 FrameData_O[2]
rlabel metal2 13524 5852 13524 5852 0 FrameData_O[30]
rlabel metal2 13804 5768 13804 5768 0 FrameData_O[31]
rlabel metal3 14721 700 14721 700 0 FrameData_O[3]
rlabel metal2 14364 784 14364 784 0 FrameData_O[4]
rlabel metal2 14420 1036 14420 1036 0 FrameData_O[5]
rlabel metal2 15204 1036 15204 1036 0 FrameData_O[6]
rlabel metal2 15092 1316 15092 1316 0 FrameData_O[7]
rlabel metal3 15057 1820 15057 1820 0 FrameData_O[8]
rlabel metal2 15148 1736 15148 1736 0 FrameData_O[9]
rlabel metal3 10976 1932 10976 1932 0 FrameStrobe[0]
rlabel metal2 12012 91 12012 91 0 FrameStrobe[10]
rlabel metal2 12124 455 12124 455 0 FrameStrobe[11]
rlabel metal2 12236 175 12236 175 0 FrameStrobe[12]
rlabel metal2 12348 175 12348 175 0 FrameStrobe[13]
rlabel metal2 12460 455 12460 455 0 FrameStrobe[14]
rlabel metal2 12572 259 12572 259 0 FrameStrobe[15]
rlabel metal2 13468 2128 13468 2128 0 FrameStrobe[16]
rlabel metal2 13692 1848 13692 1848 0 FrameStrobe[17]
rlabel metal2 14308 3416 14308 3416 0 FrameStrobe[18]
rlabel metal2 13020 1491 13020 1491 0 FrameStrobe[19]
rlabel metal2 11004 1827 11004 1827 0 FrameStrobe[1]
rlabel metal2 11116 203 11116 203 0 FrameStrobe[2]
rlabel metal2 11228 399 11228 399 0 FrameStrobe[3]
rlabel metal2 11340 455 11340 455 0 FrameStrobe[4]
rlabel metal2 11452 175 11452 175 0 FrameStrobe[5]
rlabel metal2 11564 371 11564 371 0 FrameStrobe[6]
rlabel metal2 11676 119 11676 119 0 FrameStrobe[7]
rlabel metal2 11788 427 11788 427 0 FrameStrobe[8]
rlabel metal2 11900 63 11900 63 0 FrameStrobe[9]
rlabel metal2 1820 6741 1820 6741 0 FrameStrobe_O[0]
rlabel metal2 8540 7049 8540 7049 0 FrameStrobe_O[10]
rlabel metal2 9492 6356 9492 6356 0 FrameStrobe_O[11]
rlabel metal2 9884 7049 9884 7049 0 FrameStrobe_O[12]
rlabel metal2 10556 7049 10556 7049 0 FrameStrobe_O[13]
rlabel metal2 11452 6384 11452 6384 0 FrameStrobe_O[14]
rlabel metal2 11900 7049 11900 7049 0 FrameStrobe_O[15]
rlabel metal2 12572 7049 12572 7049 0 FrameStrobe_O[16]
rlabel metal2 13468 6384 13468 6384 0 FrameStrobe_O[17]
rlabel metal2 13916 7049 13916 7049 0 FrameStrobe_O[18]
rlabel metal2 14588 6517 14588 6517 0 FrameStrobe_O[19]
rlabel metal2 2492 6741 2492 6741 0 FrameStrobe_O[1]
rlabel metal2 3164 7049 3164 7049 0 FrameStrobe_O[2]
rlabel metal2 4060 6384 4060 6384 0 FrameStrobe_O[3]
rlabel metal2 4508 7049 4508 7049 0 FrameStrobe_O[4]
rlabel metal2 5180 7049 5180 7049 0 FrameStrobe_O[5]
rlabel metal2 5852 6741 5852 6741 0 FrameStrobe_O[6]
rlabel metal2 6524 7049 6524 7049 0 FrameStrobe_O[7]
rlabel metal3 7364 6580 7364 6580 0 FrameStrobe_O[8]
rlabel metal2 8092 6356 8092 6356 0 FrameStrobe_O[9]
rlabel metal2 2716 735 2716 735 0 N1END[0]
rlabel metal2 2828 371 2828 371 0 N1END[1]
rlabel metal2 2940 175 2940 175 0 N1END[2]
rlabel metal2 3052 147 3052 147 0 N1END[3]
rlabel metal2 4060 287 4060 287 0 N2END[0]
rlabel metal2 4172 1687 4172 1687 0 N2END[1]
rlabel metal2 4284 1855 4284 1855 0 N2END[2]
rlabel metal2 4396 651 4396 651 0 N2END[3]
rlabel metal2 8932 2716 8932 2716 0 N2END[4]
rlabel metal3 5264 2156 5264 2156 0 N2END[5]
rlabel metal2 4116 840 4116 840 0 N2END[6]
rlabel metal2 3612 952 3612 952 0 N2END[7]
rlabel metal2 3164 119 3164 119 0 N2MID[0]
rlabel metal3 5068 2548 5068 2548 0 N2MID[1]
rlabel metal2 3388 259 3388 259 0 N2MID[2]
rlabel metal2 3500 651 3500 651 0 N2MID[3]
rlabel metal2 3612 203 3612 203 0 N2MID[4]
rlabel metal2 3724 511 3724 511 0 N2MID[5]
rlabel metal2 3836 259 3836 259 0 N2MID[6]
rlabel metal2 3948 231 3948 231 0 N2MID[7]
rlabel metal2 4956 595 4956 595 0 N4END[0]
rlabel metal2 6076 651 6076 651 0 N4END[10]
rlabel metal2 6188 455 6188 455 0 N4END[11]
rlabel metal2 6300 259 6300 259 0 N4END[12]
rlabel metal2 6412 343 6412 343 0 N4END[13]
rlabel metal2 6524 511 6524 511 0 N4END[14]
rlabel metal2 6636 427 6636 427 0 N4END[15]
rlabel metal2 5068 147 5068 147 0 N4END[1]
rlabel metal2 5180 91 5180 91 0 N4END[2]
rlabel metal2 5292 455 5292 455 0 N4END[3]
rlabel metal2 5404 287 5404 287 0 N4END[4]
rlabel metal2 5516 175 5516 175 0 N4END[5]
rlabel metal2 5628 231 5628 231 0 N4END[6]
rlabel metal2 5740 119 5740 119 0 N4END[7]
rlabel metal2 5852 1435 5852 1435 0 N4END[8]
rlabel metal2 5964 175 5964 175 0 N4END[9]
rlabel metal2 6748 203 6748 203 0 S1BEG[0]
rlabel metal2 6860 287 6860 287 0 S1BEG[1]
rlabel metal2 6972 91 6972 91 0 S1BEG[2]
rlabel metal2 7084 875 7084 875 0 S1BEG[3]
rlabel metal2 7196 175 7196 175 0 S2BEG[0]
rlabel metal2 7308 343 7308 343 0 S2BEG[1]
rlabel metal2 7420 427 7420 427 0 S2BEG[2]
rlabel metal2 7532 231 7532 231 0 S2BEG[3]
rlabel metal2 6972 448 6972 448 0 S2BEG[4]
rlabel metal2 7756 343 7756 343 0 S2BEG[5]
rlabel metal2 7868 483 7868 483 0 S2BEG[6]
rlabel metal2 7980 287 7980 287 0 S2BEG[7]
rlabel metal2 8092 483 8092 483 0 S2BEGb[0]
rlabel metal2 8204 259 8204 259 0 S2BEGb[1]
rlabel metal2 8316 231 8316 231 0 S2BEGb[2]
rlabel metal2 8428 147 8428 147 0 S2BEGb[3]
rlabel metal2 8540 231 8540 231 0 S2BEGb[4]
rlabel metal2 8652 679 8652 679 0 S2BEGb[5]
rlabel metal2 8764 455 8764 455 0 S2BEGb[6]
rlabel metal2 8876 259 8876 259 0 S2BEGb[7]
rlabel metal2 8988 455 8988 455 0 S4BEG[0]
rlabel metal2 10108 147 10108 147 0 S4BEG[10]
rlabel metal2 10220 315 10220 315 0 S4BEG[11]
rlabel metal2 10332 203 10332 203 0 S4BEG[12]
rlabel metal2 10444 567 10444 567 0 S4BEG[13]
rlabel metal2 10556 343 10556 343 0 S4BEG[14]
rlabel metal2 10668 623 10668 623 0 S4BEG[15]
rlabel metal2 9100 231 9100 231 0 S4BEG[1]
rlabel metal2 9212 119 9212 119 0 S4BEG[2]
rlabel metal2 9324 175 9324 175 0 S4BEG[3]
rlabel metal2 9436 483 9436 483 0 S4BEG[4]
rlabel metal2 9548 539 9548 539 0 S4BEG[5]
rlabel metal2 9660 427 9660 427 0 S4BEG[6]
rlabel metal2 9772 455 9772 455 0 S4BEG[7]
rlabel metal2 9884 287 9884 287 0 S4BEG[8]
rlabel metal2 9996 231 9996 231 0 S4BEG[9]
rlabel metal2 10780 455 10780 455 0 UserCLK
rlabel metal2 1176 6580 1176 6580 0 UserCLKo
rlabel metal2 6132 1260 6132 1260 0 net1
rlabel metal2 14812 4340 14812 4340 0 net10
rlabel metal3 11788 4508 11788 4508 0 net11
rlabel metal2 13132 2156 13132 2156 0 net12
rlabel metal2 14700 4872 14700 4872 0 net13
rlabel metal2 14756 5096 14756 5096 0 net14
rlabel metal2 14700 5488 14700 5488 0 net15
rlabel metal2 14700 5964 14700 5964 0 net16
rlabel metal2 14028 5460 14028 5460 0 net17
rlabel metal2 13916 5152 13916 5152 0 net18
rlabel metal2 13356 5460 13356 5460 0 net19
rlabel metal2 14756 2100 14756 2100 0 net2
rlabel metal3 10836 6076 10836 6076 0 net20
rlabel metal3 10556 5684 10556 5684 0 net21
rlabel metal2 12684 5292 12684 5292 0 net22
rlabel metal2 13132 588 13132 588 0 net23
rlabel metal2 13132 4844 13132 4844 0 net24
rlabel metal2 13356 4536 13356 4536 0 net25
rlabel metal3 11004 1652 11004 1652 0 net26
rlabel metal3 13678 588 13678 588 0 net27
rlabel metal2 13916 1232 13916 1232 0 net28
rlabel metal2 14700 700 14700 700 0 net29
rlabel metal2 13916 2828 13916 2828 0 net3
rlabel metal3 8680 1372 8680 1372 0 net30
rlabel metal2 13916 1736 13916 1736 0 net31
rlabel metal2 13524 1820 13524 1820 0 net32
rlabel metal2 11452 3388 11452 3388 0 net33
rlabel metal2 9996 4200 9996 4200 0 net34
rlabel metal3 10668 3780 10668 3780 0 net35
rlabel metal3 11032 4172 11032 4172 0 net36
rlabel metal3 11704 2996 11704 2996 0 net37
rlabel metal2 12348 3388 12348 3388 0 net38
rlabel metal2 13636 4228 13636 4228 0 net39
rlabel metal2 14700 2184 14700 2184 0 net4
rlabel metal2 13748 3388 13748 3388 0 net40
rlabel metal2 13972 4508 13972 4508 0 net41
rlabel metal2 14504 6468 14504 6468 0 net42
rlabel metal2 14560 2996 14560 2996 0 net43
rlabel metal2 10640 3780 10640 3780 0 net44
rlabel metal2 8372 4844 8372 4844 0 net45
rlabel metal2 9548 4816 9548 4816 0 net46
rlabel metal2 7756 5040 7756 5040 0 net47
rlabel metal2 5264 4564 5264 4564 0 net48
rlabel metal2 5012 5124 5012 5124 0 net49
rlabel metal2 14756 2716 14756 2716 0 net5
rlabel metal2 5908 5124 5908 5124 0 net50
rlabel metal3 6860 4172 6860 4172 0 net51
rlabel metal2 8988 4368 8988 4368 0 net52
rlabel metal2 4060 728 4060 728 0 net53
rlabel metal3 5040 532 5040 532 0 net54
rlabel metal3 5348 1036 5348 1036 0 net55
rlabel metal3 5880 1708 5880 1708 0 net56
rlabel metal3 5124 2212 5124 2212 0 net57
rlabel metal2 3388 616 3388 616 0 net58
rlabel metal2 4844 1260 4844 1260 0 net59
rlabel metal2 13916 3304 13916 3304 0 net6
rlabel metal3 6104 2100 6104 2100 0 net60
rlabel metal2 6468 952 6468 952 0 net61
rlabel metal3 6748 1372 6748 1372 0 net62
rlabel metal2 7308 1036 7308 1036 0 net63
rlabel metal2 7364 756 7364 756 0 net64
rlabel metal2 3388 1484 3388 1484 0 net65
rlabel metal2 3780 1036 3780 1036 0 net66
rlabel metal2 8540 1372 8540 1372 0 net67
rlabel metal2 9128 1932 9128 1932 0 net68
rlabel metal2 9688 2492 9688 2492 0 net69
rlabel metal2 14700 2968 14700 2968 0 net7
rlabel metal2 9632 2660 9632 2660 0 net70
rlabel metal3 9744 3276 9744 3276 0 net71
rlabel metal2 10108 1134 10108 1134 0 net72
rlabel metal2 9996 1316 9996 1316 0 net73
rlabel metal2 12572 1148 12572 1148 0 net74
rlabel metal2 11228 2352 11228 2352 0 net75
rlabel metal3 11928 2604 11928 2604 0 net76
rlabel metal2 12796 1330 12796 1330 0 net77
rlabel metal3 11956 2100 11956 2100 0 net78
rlabel metal3 11172 1484 11172 1484 0 net79
rlabel metal2 14700 3276 14700 3276 0 net8
rlabel metal2 5460 1064 5460 1064 0 net80
rlabel metal2 5404 1008 5404 1008 0 net81
rlabel metal2 4900 784 4900 784 0 net82
rlabel metal2 5068 1036 5068 1036 0 net83
rlabel metal3 10416 980 10416 980 0 net84
rlabel metal3 11788 952 11788 952 0 net85
rlabel metal2 10612 2800 10612 2800 0 net86
rlabel metal2 10892 2212 10892 2212 0 net87
rlabel metal3 12348 1316 12348 1316 0 net88
rlabel metal2 1372 5544 1372 5544 0 net89
rlabel metal2 14700 4060 14700 4060 0 net9
<< properties >>
string FIXED_BBOX 0 0 15848 7112
<< end >>
