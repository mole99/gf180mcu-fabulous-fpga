magic
tech gf180mcuD
magscale 1 10
timestamp 1765465586
<< metal2 >>
rect 1820 719124 1876 719134
rect 1820 717444 1876 719068
rect 1820 717378 1876 717388
rect 812 196 868 15372
rect 812 112 868 140
rect 2156 112 2212 15372
rect 3500 112 3556 15372
rect 4844 112 4900 15372
rect 6188 112 6244 15372
rect 7532 112 7588 15372
rect 8876 112 8932 15372
rect 10220 112 10276 15372
rect 11564 112 11620 15372
rect 12908 112 12964 15372
rect 14252 112 14308 15372
rect 15596 112 15652 15372
rect 16940 112 16996 15372
rect 18284 112 18340 15372
rect 19628 112 19684 15372
rect 20972 112 21028 15372
rect 22316 112 22372 15372
rect 23660 112 23716 15372
rect 25004 112 25060 15372
rect 26348 112 26404 15372
rect 27692 112 27748 15372
rect 30044 112 30100 1148
rect 32060 112 32116 1148
rect 34076 112 34132 1148
rect 36092 112 36148 1148
rect 38108 112 38164 1148
rect 40124 112 40180 1148
rect 42140 112 42196 1148
rect 44184 980 44240 1148
rect 44156 924 44184 980
rect 44156 914 44240 924
rect 784 0 896 112
rect 2128 0 2240 112
rect 3472 0 3584 112
rect 4816 0 4928 112
rect 6160 0 6272 112
rect 7504 0 7616 112
rect 8848 0 8960 112
rect 10192 0 10304 112
rect 11536 0 11648 112
rect 12880 0 12992 112
rect 14224 0 14336 112
rect 15568 0 15680 112
rect 16912 0 17024 112
rect 18256 0 18368 112
rect 19600 0 19712 112
rect 20944 0 21056 112
rect 22288 0 22400 112
rect 23632 0 23744 112
rect 24976 0 25088 112
rect 26320 0 26432 112
rect 27664 0 27776 112
rect 30016 0 30128 112
rect 32032 0 32144 112
rect 34048 0 34160 112
rect 36064 0 36176 112
rect 38080 0 38192 112
rect 40096 0 40208 112
rect 42112 0 42224 112
rect 44156 84 44212 914
rect 46172 112 46228 1148
rect 48188 112 48244 1148
rect 50204 112 50260 1148
rect 52220 112 52276 1148
rect 54236 112 54292 1148
rect 56252 112 56308 1148
rect 58268 112 58324 1148
rect 60284 112 60340 1148
rect 62300 112 62356 1148
rect 64316 112 64372 1148
rect 66332 112 66388 1148
rect 68348 112 68404 1148
rect 70364 112 70420 1148
rect 72380 112 72436 1148
rect 74396 112 74452 1148
rect 76412 112 76468 1148
rect 78428 112 78484 1148
rect 80444 112 80500 1148
rect 82460 112 82516 1148
rect 84476 112 84532 1148
rect 87920 980 87976 1148
rect 87920 914 87976 924
rect 90636 112 90692 1148
rect 93324 112 93380 1148
rect 96012 112 96068 1148
rect 98700 112 98756 1148
rect 101388 112 101444 1148
rect 104076 112 104132 1148
rect 106764 112 106820 1148
rect 109452 112 109508 1148
rect 112140 112 112196 1148
rect 114828 112 114884 1148
rect 117516 112 117572 1148
rect 120204 112 120260 1148
rect 122892 112 122948 1148
rect 125580 112 125636 1148
rect 128268 112 128324 1148
rect 130956 112 131012 1148
rect 133644 112 133700 1148
rect 136332 112 136388 1148
rect 139020 112 139076 1148
rect 141708 112 141764 1148
rect 145376 980 145432 1148
rect 145376 914 145432 924
rect 148092 112 148148 1148
rect 150780 112 150836 1148
rect 153468 112 153524 1148
rect 156156 112 156212 1148
rect 158844 112 158900 1148
rect 161532 112 161588 1148
rect 164220 112 164276 1148
rect 166908 112 166964 1148
rect 169596 112 169652 1148
rect 172284 112 172340 1148
rect 174972 112 175028 1148
rect 177660 112 177716 1148
rect 180348 112 180404 1148
rect 183036 112 183092 1148
rect 185724 112 185780 1148
rect 188412 112 188468 1148
rect 191100 112 191156 1148
rect 193788 112 193844 1148
rect 196476 112 196532 1148
rect 199164 112 199220 1148
rect 203952 980 204008 1148
rect 203952 914 204008 924
rect 206892 112 206948 1148
rect 209804 112 209860 1148
rect 212716 112 212772 1148
rect 215628 112 215684 1148
rect 218540 112 218596 1148
rect 221452 112 221508 1148
rect 224364 112 224420 1148
rect 227276 112 227332 1148
rect 230188 112 230244 1148
rect 233100 112 233156 1148
rect 236012 112 236068 1148
rect 238924 112 238980 1148
rect 241836 112 241892 1148
rect 244748 112 244804 1148
rect 247660 112 247716 1148
rect 250572 112 250628 1148
rect 253484 112 253540 1148
rect 256396 112 256452 1148
rect 259308 112 259364 1148
rect 262220 112 262276 1148
rect 267288 980 267344 1148
rect 267288 914 267344 924
rect 269948 112 270004 1148
rect 272636 112 272692 1148
rect 275324 112 275380 1148
rect 278012 112 278068 1148
rect 280700 112 280756 1148
rect 283388 112 283444 1148
rect 286076 112 286132 1148
rect 288764 112 288820 1148
rect 291452 112 291508 1148
rect 294140 112 294196 1148
rect 296828 112 296884 1148
rect 299516 112 299572 1148
rect 302204 112 302260 1148
rect 304892 112 304948 1148
rect 307580 112 307636 1148
rect 310268 112 310324 1148
rect 312956 112 313012 1148
rect 315644 112 315700 1148
rect 318332 112 318388 1148
rect 321020 112 321076 1148
rect 324464 980 324520 1148
rect 324464 914 324520 924
rect 326956 112 327012 1148
rect 329420 112 329476 1148
rect 331884 112 331940 1148
rect 334348 112 334404 1148
rect 336812 112 336868 1148
rect 339276 112 339332 1148
rect 341740 112 341796 1148
rect 344204 112 344260 1148
rect 346668 112 346724 1148
rect 349132 112 349188 1148
rect 351596 112 351652 1148
rect 354060 112 354116 1148
rect 356524 112 356580 1148
rect 358988 112 359044 1148
rect 361452 112 361508 1148
rect 363916 112 363972 1148
rect 366380 112 366436 1148
rect 368844 112 368900 1148
rect 371308 112 371364 1148
rect 373772 112 373828 1148
rect 377496 980 377552 1148
rect 377496 914 377552 924
rect 380156 112 380212 1148
rect 382844 112 382900 1148
rect 385532 112 385588 1148
rect 388220 112 388276 1148
rect 390908 112 390964 1148
rect 393596 112 393652 1148
rect 396284 112 396340 1148
rect 398972 112 399028 1148
rect 401660 112 401716 1148
rect 404348 112 404404 1148
rect 407036 112 407092 1148
rect 409724 112 409780 1148
rect 412412 112 412468 1148
rect 415100 112 415156 1148
rect 417788 112 417844 1148
rect 420476 112 420532 1148
rect 423164 112 423220 1148
rect 425852 112 425908 1148
rect 428540 112 428596 1148
rect 431228 112 431284 1148
rect 435344 980 435400 1148
rect 435344 914 435400 924
rect 436716 112 436772 1148
rect 438060 112 438116 1148
rect 439404 112 439460 1148
rect 440748 112 440804 1148
rect 442092 112 442148 1148
rect 443436 112 443492 1148
rect 444780 112 444836 1148
rect 446124 112 446180 1148
rect 447468 196 447524 1148
rect 447468 130 447524 140
rect 448252 196 448308 206
rect 448252 112 448308 140
rect 448812 112 448868 1148
rect 450156 112 450212 1148
rect 451500 112 451556 1148
rect 452844 112 452900 1148
rect 454188 112 454244 1148
rect 455532 112 455588 1148
rect 456876 112 456932 1148
rect 458220 112 458276 1148
rect 459564 112 459620 1148
rect 460908 112 460964 1148
rect 462252 112 462308 1148
rect 44156 18 44212 28
rect 46144 0 46256 112
rect 48160 0 48272 112
rect 50176 0 50288 112
rect 52192 0 52304 112
rect 54208 0 54320 112
rect 56224 0 56336 112
rect 58240 0 58352 112
rect 60256 0 60368 112
rect 62272 0 62384 112
rect 64288 0 64400 112
rect 66304 0 66416 112
rect 68320 0 68432 112
rect 70336 0 70448 112
rect 72352 0 72464 112
rect 74368 0 74480 112
rect 76384 0 76496 112
rect 78400 0 78512 112
rect 80416 0 80528 112
rect 82432 0 82544 112
rect 84448 0 84560 112
rect 90608 0 90720 112
rect 93296 0 93408 112
rect 95984 0 96096 112
rect 98672 0 98784 112
rect 101360 0 101472 112
rect 104048 0 104160 112
rect 106736 0 106848 112
rect 109424 0 109536 112
rect 112112 0 112224 112
rect 114800 0 114912 112
rect 117488 0 117600 112
rect 120176 0 120288 112
rect 122864 0 122976 112
rect 125552 0 125664 112
rect 128240 0 128352 112
rect 130928 0 131040 112
rect 133616 0 133728 112
rect 136304 0 136416 112
rect 138992 0 139104 112
rect 141680 0 141792 112
rect 148064 0 148176 112
rect 150752 0 150864 112
rect 153440 0 153552 112
rect 156128 0 156240 112
rect 158816 0 158928 112
rect 161504 0 161616 112
rect 164192 0 164304 112
rect 166880 0 166992 112
rect 169568 0 169680 112
rect 172256 0 172368 112
rect 174944 0 175056 112
rect 177632 0 177744 112
rect 180320 0 180432 112
rect 183008 0 183120 112
rect 185696 0 185808 112
rect 188384 0 188496 112
rect 191072 0 191184 112
rect 193760 0 193872 112
rect 196448 0 196560 112
rect 199136 0 199248 112
rect 206864 0 206976 112
rect 209776 0 209888 112
rect 212688 0 212800 112
rect 215600 0 215712 112
rect 218512 0 218624 112
rect 221424 0 221536 112
rect 224336 0 224448 112
rect 227248 0 227360 112
rect 230160 0 230272 112
rect 233072 0 233184 112
rect 235984 0 236096 112
rect 238896 0 239008 112
rect 241808 0 241920 112
rect 244720 0 244832 112
rect 247632 0 247744 112
rect 250544 0 250656 112
rect 253456 0 253568 112
rect 256368 0 256480 112
rect 259280 0 259392 112
rect 262192 0 262304 112
rect 269920 0 270032 112
rect 272608 0 272720 112
rect 275296 0 275408 112
rect 277984 0 278096 112
rect 280672 0 280784 112
rect 283360 0 283472 112
rect 286048 0 286160 112
rect 288736 0 288848 112
rect 291424 0 291536 112
rect 294112 0 294224 112
rect 296800 0 296912 112
rect 299488 0 299600 112
rect 302176 0 302288 112
rect 304864 0 304976 112
rect 307552 0 307664 112
rect 310240 0 310352 112
rect 312928 0 313040 112
rect 315616 0 315728 112
rect 318304 0 318416 112
rect 320992 0 321104 112
rect 326928 0 327040 112
rect 329392 0 329504 112
rect 331856 0 331968 112
rect 334320 0 334432 112
rect 336784 0 336896 112
rect 339248 0 339360 112
rect 341712 0 341824 112
rect 344176 0 344288 112
rect 346640 0 346752 112
rect 349104 0 349216 112
rect 351568 0 351680 112
rect 354032 0 354144 112
rect 356496 0 356608 112
rect 358960 0 359072 112
rect 361424 0 361536 112
rect 363888 0 364000 112
rect 366352 0 366464 112
rect 368816 0 368928 112
rect 371280 0 371392 112
rect 373744 0 373856 112
rect 380128 0 380240 112
rect 382816 0 382928 112
rect 385504 0 385616 112
rect 388192 0 388304 112
rect 390880 0 390992 112
rect 393568 0 393680 112
rect 396256 0 396368 112
rect 398944 0 399056 112
rect 401632 0 401744 112
rect 404320 0 404432 112
rect 407008 0 407120 112
rect 409696 0 409808 112
rect 412384 0 412496 112
rect 415072 0 415184 112
rect 417760 0 417872 112
rect 420448 0 420560 112
rect 423136 0 423248 112
rect 425824 0 425936 112
rect 428512 0 428624 112
rect 431200 0 431312 112
rect 436688 0 436800 112
rect 438032 0 438144 112
rect 439376 0 439488 112
rect 440720 0 440832 112
rect 442064 0 442176 112
rect 443408 0 443520 112
rect 444752 0 444864 112
rect 446096 0 446208 112
rect 448224 0 448336 112
rect 448784 0 448896 112
rect 450128 0 450240 112
rect 451472 0 451584 112
rect 452816 0 452928 112
rect 454160 0 454272 112
rect 455504 0 455616 112
rect 456848 0 456960 112
rect 458192 0 458304 112
rect 459536 0 459648 112
rect 460880 0 460992 112
rect 462224 0 462336 112
<< via2 >>
rect 1820 719068 1876 719124
rect 1820 717388 1876 717444
rect 812 140 868 196
rect 44184 924 44240 980
rect 87920 924 87976 980
rect 145376 924 145432 980
rect 203952 924 204008 980
rect 267288 924 267344 980
rect 324464 924 324520 980
rect 377496 924 377552 980
rect 435344 924 435400 980
rect 447468 140 447524 196
rect 448252 140 448308 196
rect 44156 28 44212 84
<< metal3 >>
rect 1810 719068 1820 719124
rect 1876 719068 28140 719124
rect 28196 719068 28206 719124
rect 0 718788 112 718816
rect 0 718732 28728 718788
rect 0 718704 112 718732
rect 0 718340 112 718368
rect 0 718284 28728 718340
rect 0 718256 112 718284
rect 0 717892 112 717920
rect 0 717836 28728 717892
rect 0 717808 112 717836
rect 0 717444 112 717472
rect 28130 717444 28140 717500
rect 28196 717444 28728 717500
rect 0 717388 1820 717444
rect 1876 717388 1886 717444
rect 0 717360 112 717388
rect 0 716996 112 717024
rect 0 716940 28728 716996
rect 0 716912 112 716940
rect 0 716548 112 716576
rect 0 716492 28728 716548
rect 0 716464 112 716492
rect 0 716100 112 716128
rect 0 716044 28728 716100
rect 0 716016 112 716044
rect 0 715652 112 715680
rect 0 715596 28728 715652
rect 0 715568 112 715596
rect 0 715204 112 715232
rect 0 715148 28728 715204
rect 0 715120 112 715148
rect 0 714756 112 714784
rect 0 714700 28728 714756
rect 0 714672 112 714700
rect 0 714308 112 714336
rect 0 714252 28728 714308
rect 0 714224 112 714252
rect 0 713860 112 713888
rect 0 713804 28728 713860
rect 0 713776 112 713804
rect 0 713412 112 713440
rect 0 713356 28728 713412
rect 0 713328 112 713356
rect 0 712964 112 712992
rect 0 712908 28728 712964
rect 0 712880 112 712908
rect 0 712516 112 712544
rect 0 712460 28728 712516
rect 0 712432 112 712460
rect 0 712068 112 712096
rect 0 712012 28728 712068
rect 0 711984 112 712012
rect 0 711620 112 711648
rect 0 711564 28728 711620
rect 0 711536 112 711564
rect 0 711172 112 711200
rect 0 711116 28728 711172
rect 0 711088 112 711116
rect 0 710724 112 710752
rect 0 710668 28728 710724
rect 0 710640 112 710668
rect 0 710276 112 710304
rect 0 710220 28728 710276
rect 0 710192 112 710220
rect 0 709828 112 709856
rect 0 709772 28728 709828
rect 0 709744 112 709772
rect 0 709380 112 709408
rect 0 709324 28728 709380
rect 0 709296 112 709324
rect 0 708932 112 708960
rect 0 708876 28728 708932
rect 0 708848 112 708876
rect 0 708484 112 708512
rect 0 708428 28728 708484
rect 0 708400 112 708428
rect 0 708036 112 708064
rect 0 707980 28728 708036
rect 0 707952 112 707980
rect 0 707588 112 707616
rect 0 707532 28728 707588
rect 0 707504 112 707532
rect 0 707140 112 707168
rect 0 707084 28728 707140
rect 0 707056 112 707084
rect 0 706692 112 706720
rect 0 706636 28728 706692
rect 0 706608 112 706636
rect 0 706244 112 706272
rect 0 706188 28728 706244
rect 0 706160 112 706188
rect 0 705796 112 705824
rect 0 705740 28728 705796
rect 0 705712 112 705740
rect 0 705348 112 705376
rect 0 705292 28728 705348
rect 0 705264 112 705292
rect 0 704900 112 704928
rect 0 704844 8428 704900
rect 0 704816 112 704844
rect 8372 704788 8428 704844
rect 28028 704788 28728 704844
rect 8372 704732 28084 704788
rect 0 702548 112 702576
rect 0 702492 168 702548
rect 0 702464 112 702492
rect 0 701652 112 701680
rect 0 701596 168 701652
rect 0 701568 112 701596
rect 0 700756 112 700784
rect 0 700700 168 700756
rect 0 700672 112 700700
rect 0 699860 112 699888
rect 0 699804 168 699860
rect 0 699776 112 699804
rect 0 698964 112 698992
rect 0 698908 168 698964
rect 0 698880 112 698908
rect 0 698068 112 698096
rect 0 698012 168 698068
rect 0 697984 112 698012
rect 0 697172 112 697200
rect 0 697116 168 697172
rect 0 697088 112 697116
rect 0 696276 112 696304
rect 0 696220 168 696276
rect 0 696192 112 696220
rect 0 695380 112 695408
rect 0 695324 168 695380
rect 0 695296 112 695324
rect 0 694484 112 694512
rect 0 694428 168 694484
rect 0 694400 112 694428
rect 0 693588 112 693616
rect 0 693532 168 693588
rect 0 693504 112 693532
rect 0 692692 112 692720
rect 0 692636 168 692692
rect 0 692608 112 692636
rect 0 691796 112 691824
rect 0 691740 168 691796
rect 0 691712 112 691740
rect 0 690900 112 690928
rect 0 690844 168 690900
rect 0 690816 112 690844
rect 0 690004 112 690032
rect 0 689948 168 690004
rect 0 689920 112 689948
rect 0 689108 112 689136
rect 0 689052 168 689108
rect 0 689024 112 689052
rect 0 688212 112 688240
rect 0 688156 168 688212
rect 0 688128 112 688156
rect 0 687316 112 687344
rect 0 687260 168 687316
rect 0 687232 112 687260
rect 0 686420 112 686448
rect 0 686364 168 686420
rect 0 686336 112 686364
rect 0 685524 112 685552
rect 0 685468 168 685524
rect 0 685440 112 685468
rect 0 684628 112 684656
rect 0 684572 168 684628
rect 0 684544 112 684572
rect 0 683732 112 683760
rect 0 683676 168 683732
rect 0 683648 112 683676
rect 0 682836 112 682864
rect 0 682780 168 682836
rect 0 682752 112 682780
rect 0 681940 112 681968
rect 0 681884 168 681940
rect 0 681856 112 681884
rect 0 681044 112 681072
rect 0 680988 168 681044
rect 0 680960 112 680988
rect 0 680148 112 680176
rect 0 680092 168 680148
rect 0 680064 112 680092
rect 0 679252 112 679280
rect 0 679196 168 679252
rect 0 679168 112 679196
rect 0 678356 112 678384
rect 0 678300 168 678356
rect 0 678272 112 678300
rect 0 677460 112 677488
rect 0 677404 168 677460
rect 0 677376 112 677404
rect 0 676564 112 676592
rect 0 676508 168 676564
rect 0 676480 112 676508
rect 0 675668 112 675696
rect 0 675612 168 675668
rect 0 675584 112 675612
rect 0 674772 112 674800
rect 0 674716 168 674772
rect 0 674688 112 674716
rect 0 673876 112 673904
rect 0 673820 168 673876
rect 0 673792 112 673820
rect 0 672980 112 673008
rect 0 672924 168 672980
rect 0 672896 112 672924
rect 0 672084 112 672112
rect 0 672028 168 672084
rect 0 672000 112 672028
rect 0 671188 112 671216
rect 0 671132 168 671188
rect 0 671104 112 671132
rect 0 670292 112 670320
rect 0 670236 168 670292
rect 0 670208 112 670236
rect 0 669396 112 669424
rect 0 669340 168 669396
rect 0 669312 112 669340
rect 0 668500 112 668528
rect 0 668444 168 668500
rect 0 668416 112 668444
rect 0 667604 112 667632
rect 0 667548 168 667604
rect 0 667520 112 667548
rect 0 666708 112 666736
rect 0 666652 168 666708
rect 0 666624 112 666652
rect 0 665812 112 665840
rect 0 665756 168 665812
rect 0 665728 112 665756
rect 0 664916 112 664944
rect 0 664860 168 664916
rect 0 664832 112 664860
rect 0 664020 112 664048
rect 0 663964 168 664020
rect 0 663936 112 663964
rect 0 663124 112 663152
rect 0 663068 168 663124
rect 0 663040 112 663068
rect 0 662228 112 662256
rect 0 662172 168 662228
rect 0 662144 112 662172
rect 0 661332 112 661360
rect 0 661276 168 661332
rect 0 661248 112 661276
rect 0 660436 112 660464
rect 0 660380 168 660436
rect 0 660352 112 660380
rect 0 659540 112 659568
rect 0 659484 168 659540
rect 0 659456 112 659484
rect 0 658644 112 658672
rect 0 658588 168 658644
rect 0 658560 112 658588
rect 0 657748 112 657776
rect 0 657692 168 657748
rect 0 657664 112 657692
rect 0 656852 112 656880
rect 0 656796 168 656852
rect 0 656768 112 656796
rect 0 655956 112 655984
rect 0 655900 168 655956
rect 0 655872 112 655900
rect 0 655060 112 655088
rect 0 655004 168 655060
rect 0 654976 112 655004
rect 0 654164 112 654192
rect 0 654108 168 654164
rect 0 654080 112 654108
rect 0 653268 112 653296
rect 0 653212 168 653268
rect 0 653184 112 653212
rect 0 652372 112 652400
rect 0 652316 168 652372
rect 0 652288 112 652316
rect 0 651476 112 651504
rect 0 651420 168 651476
rect 0 651392 112 651420
rect 0 650580 112 650608
rect 0 650524 168 650580
rect 0 650496 112 650524
rect 0 649684 112 649712
rect 0 649628 168 649684
rect 0 649600 112 649628
rect 0 645092 112 645120
rect 0 645036 168 645092
rect 0 645008 112 645036
rect 0 644196 112 644224
rect 0 644140 168 644196
rect 0 644112 112 644140
rect 0 643300 112 643328
rect 0 643244 168 643300
rect 0 643216 112 643244
rect 0 642404 112 642432
rect 0 642348 168 642404
rect 0 642320 112 642348
rect 0 641508 112 641536
rect 0 641452 168 641508
rect 0 641424 112 641452
rect 0 640612 112 640640
rect 0 640556 168 640612
rect 0 640528 112 640556
rect 0 639716 112 639744
rect 0 639660 168 639716
rect 0 639632 112 639660
rect 0 638820 112 638848
rect 0 638764 168 638820
rect 0 638736 112 638764
rect 0 637924 112 637952
rect 0 637868 168 637924
rect 0 637840 112 637868
rect 0 637028 112 637056
rect 0 636972 168 637028
rect 0 636944 112 636972
rect 0 636132 112 636160
rect 0 636076 168 636132
rect 0 636048 112 636076
rect 0 635236 112 635264
rect 0 635180 168 635236
rect 0 635152 112 635180
rect 0 634340 112 634368
rect 0 634284 168 634340
rect 0 634256 112 634284
rect 0 633444 112 633472
rect 0 633388 168 633444
rect 0 633360 112 633388
rect 0 632548 112 632576
rect 0 632492 168 632548
rect 0 632464 112 632492
rect 0 631652 112 631680
rect 0 631596 168 631652
rect 0 631568 112 631596
rect 0 630756 112 630784
rect 0 630700 168 630756
rect 0 630672 112 630700
rect 0 629860 112 629888
rect 0 629804 168 629860
rect 0 629776 112 629804
rect 0 628964 112 628992
rect 0 628908 168 628964
rect 0 628880 112 628908
rect 0 628068 112 628096
rect 0 628012 168 628068
rect 0 627984 112 628012
rect 0 627172 112 627200
rect 0 627116 168 627172
rect 0 627088 112 627116
rect 0 626276 112 626304
rect 0 626220 168 626276
rect 0 626192 112 626220
rect 0 625380 112 625408
rect 0 625324 168 625380
rect 0 625296 112 625324
rect 464800 625156 464912 625184
rect 464772 625100 464912 625156
rect 464800 625072 464912 625100
rect 0 624484 112 624512
rect 0 624428 168 624484
rect 0 624400 112 624428
rect 464800 624260 464912 624288
rect 464772 624204 464912 624260
rect 464800 624176 464912 624204
rect 0 623588 112 623616
rect 0 623532 168 623588
rect 0 623504 112 623532
rect 464800 623364 464912 623392
rect 464772 623308 464912 623364
rect 464800 623280 464912 623308
rect 0 622692 112 622720
rect 0 622636 168 622692
rect 0 622608 112 622636
rect 464800 622468 464912 622496
rect 464772 622412 464912 622468
rect 464800 622384 464912 622412
rect 0 621796 112 621824
rect 0 621740 168 621796
rect 0 621712 112 621740
rect 464800 621572 464912 621600
rect 464772 621516 464912 621572
rect 464800 621488 464912 621516
rect 0 620900 112 620928
rect 0 620844 168 620900
rect 0 620816 112 620844
rect 464800 620676 464912 620704
rect 464772 620620 464912 620676
rect 464800 620592 464912 620620
rect 0 620004 112 620032
rect 0 619948 168 620004
rect 0 619920 112 619948
rect 464800 619780 464912 619808
rect 464772 619724 464912 619780
rect 464800 619696 464912 619724
rect 0 619108 112 619136
rect 0 619052 168 619108
rect 0 619024 112 619052
rect 464800 618884 464912 618912
rect 464772 618828 464912 618884
rect 464800 618800 464912 618828
rect 0 618212 112 618240
rect 0 618156 168 618212
rect 0 618128 112 618156
rect 464800 617988 464912 618016
rect 464772 617932 464912 617988
rect 464800 617904 464912 617932
rect 0 617316 112 617344
rect 0 617260 168 617316
rect 0 617232 112 617260
rect 464800 617092 464912 617120
rect 464772 617036 464912 617092
rect 464800 617008 464912 617036
rect 0 616420 112 616448
rect 0 616364 168 616420
rect 0 616336 112 616364
rect 464800 616196 464912 616224
rect 464772 616140 464912 616196
rect 464800 616112 464912 616140
rect 0 615524 112 615552
rect 0 615468 168 615524
rect 0 615440 112 615468
rect 464800 615300 464912 615328
rect 464772 615244 464912 615300
rect 464800 615216 464912 615244
rect 0 614628 112 614656
rect 0 614572 168 614628
rect 0 614544 112 614572
rect 464800 614404 464912 614432
rect 464772 614348 464912 614404
rect 464800 614320 464912 614348
rect 0 613732 112 613760
rect 0 613676 168 613732
rect 0 613648 112 613676
rect 464800 613508 464912 613536
rect 464772 613452 464912 613508
rect 464800 613424 464912 613452
rect 0 612836 112 612864
rect 0 612780 168 612836
rect 0 612752 112 612780
rect 464800 612612 464912 612640
rect 464772 612556 464912 612612
rect 464800 612528 464912 612556
rect 0 611940 112 611968
rect 0 611884 168 611940
rect 0 611856 112 611884
rect 464800 611716 464912 611744
rect 464772 611660 464912 611716
rect 464800 611632 464912 611660
rect 0 611044 112 611072
rect 0 610988 168 611044
rect 0 610960 112 610988
rect 464800 610820 464912 610848
rect 464772 610764 464912 610820
rect 464800 610736 464912 610764
rect 0 610148 112 610176
rect 0 610092 168 610148
rect 0 610064 112 610092
rect 464800 609924 464912 609952
rect 464772 609868 464912 609924
rect 464800 609840 464912 609868
rect 0 609252 112 609280
rect 0 609196 168 609252
rect 0 609168 112 609196
rect 464800 609028 464912 609056
rect 464772 608972 464912 609028
rect 464800 608944 464912 608972
rect 0 608356 112 608384
rect 0 608300 168 608356
rect 0 608272 112 608300
rect 464800 608132 464912 608160
rect 464772 608076 464912 608132
rect 464800 608048 464912 608076
rect 0 607460 112 607488
rect 0 607404 168 607460
rect 0 607376 112 607404
rect 464800 607236 464912 607264
rect 464772 607180 464912 607236
rect 464800 607152 464912 607180
rect 0 606564 112 606592
rect 0 606508 168 606564
rect 0 606480 112 606508
rect 464800 606340 464912 606368
rect 464772 606284 464912 606340
rect 464800 606256 464912 606284
rect 0 605668 112 605696
rect 0 605612 168 605668
rect 0 605584 112 605612
rect 464800 605444 464912 605472
rect 464772 605388 464912 605444
rect 464800 605360 464912 605388
rect 0 604772 112 604800
rect 0 604716 168 604772
rect 0 604688 112 604716
rect 464800 604548 464912 604576
rect 464772 604492 464912 604548
rect 464800 604464 464912 604492
rect 0 603876 112 603904
rect 0 603820 168 603876
rect 0 603792 112 603820
rect 464800 603652 464912 603680
rect 464772 603596 464912 603652
rect 464800 603568 464912 603596
rect 0 602980 112 603008
rect 0 602924 168 602980
rect 0 602896 112 602924
rect 464800 602756 464912 602784
rect 464772 602700 464912 602756
rect 464800 602672 464912 602700
rect 0 602084 112 602112
rect 0 602028 168 602084
rect 0 602000 112 602028
rect 464800 601860 464912 601888
rect 464772 601804 464912 601860
rect 464800 601776 464912 601804
rect 0 601188 112 601216
rect 0 601132 168 601188
rect 0 601104 112 601132
rect 464800 600964 464912 600992
rect 464772 600908 464912 600964
rect 464800 600880 464912 600908
rect 0 600292 112 600320
rect 0 600236 168 600292
rect 0 600208 112 600236
rect 464800 600068 464912 600096
rect 464772 600012 464912 600068
rect 464800 599984 464912 600012
rect 0 599396 112 599424
rect 0 599340 168 599396
rect 0 599312 112 599340
rect 464800 599172 464912 599200
rect 464772 599116 464912 599172
rect 464800 599088 464912 599116
rect 0 598500 112 598528
rect 0 598444 168 598500
rect 0 598416 112 598444
rect 464800 598276 464912 598304
rect 464772 598220 464912 598276
rect 464800 598192 464912 598220
rect 0 597604 112 597632
rect 0 597548 168 597604
rect 0 597520 112 597548
rect 464800 597380 464912 597408
rect 464772 597324 464912 597380
rect 464800 597296 464912 597324
rect 0 596708 112 596736
rect 0 596652 168 596708
rect 0 596624 112 596652
rect 464800 596484 464912 596512
rect 464772 596428 464912 596484
rect 464800 596400 464912 596428
rect 0 595812 112 595840
rect 0 595756 168 595812
rect 0 595728 112 595756
rect 464800 595588 464912 595616
rect 464772 595532 464912 595588
rect 464800 595504 464912 595532
rect 0 594916 112 594944
rect 0 594860 168 594916
rect 0 594832 112 594860
rect 464800 594692 464912 594720
rect 464772 594636 464912 594692
rect 464800 594608 464912 594636
rect 0 594020 112 594048
rect 0 593964 168 594020
rect 0 593936 112 593964
rect 464800 593796 464912 593824
rect 464772 593740 464912 593796
rect 464800 593712 464912 593740
rect 0 593124 112 593152
rect 0 593068 168 593124
rect 0 593040 112 593068
rect 464800 592900 464912 592928
rect 464772 592844 464912 592900
rect 464800 592816 464912 592844
rect 0 592228 112 592256
rect 0 592172 168 592228
rect 0 592144 112 592172
rect 0 587636 112 587664
rect 0 587580 168 587636
rect 0 587552 112 587580
rect 0 586740 112 586768
rect 0 586684 168 586740
rect 0 586656 112 586684
rect 0 585844 112 585872
rect 0 585788 168 585844
rect 0 585760 112 585788
rect 0 584948 112 584976
rect 0 584892 168 584948
rect 0 584864 112 584892
rect 0 584052 112 584080
rect 0 583996 168 584052
rect 0 583968 112 583996
rect 0 583156 112 583184
rect 0 583100 168 583156
rect 0 583072 112 583100
rect 0 582260 112 582288
rect 0 582204 168 582260
rect 0 582176 112 582204
rect 0 581364 112 581392
rect 0 581308 168 581364
rect 0 581280 112 581308
rect 0 580468 112 580496
rect 0 580412 168 580468
rect 0 580384 112 580412
rect 0 579572 112 579600
rect 0 579516 168 579572
rect 0 579488 112 579516
rect 0 578676 112 578704
rect 0 578620 168 578676
rect 0 578592 112 578620
rect 0 577780 112 577808
rect 0 577724 168 577780
rect 0 577696 112 577724
rect 0 576884 112 576912
rect 0 576828 168 576884
rect 0 576800 112 576828
rect 0 575988 112 576016
rect 0 575932 168 575988
rect 0 575904 112 575932
rect 0 575092 112 575120
rect 0 575036 168 575092
rect 0 575008 112 575036
rect 0 574196 112 574224
rect 0 574140 168 574196
rect 0 574112 112 574140
rect 0 573300 112 573328
rect 0 573244 168 573300
rect 0 573216 112 573244
rect 0 572404 112 572432
rect 0 572348 168 572404
rect 0 572320 112 572348
rect 0 571508 112 571536
rect 0 571452 168 571508
rect 0 571424 112 571452
rect 0 570612 112 570640
rect 0 570556 168 570612
rect 0 570528 112 570556
rect 0 569716 112 569744
rect 0 569660 168 569716
rect 0 569632 112 569660
rect 0 568820 112 568848
rect 0 568764 168 568820
rect 0 568736 112 568764
rect 0 567924 112 567952
rect 0 567868 168 567924
rect 0 567840 112 567868
rect 0 567028 112 567056
rect 0 566972 168 567028
rect 0 566944 112 566972
rect 0 566132 112 566160
rect 0 566076 168 566132
rect 0 566048 112 566076
rect 0 565236 112 565264
rect 0 565180 168 565236
rect 0 565152 112 565180
rect 0 564340 112 564368
rect 0 564284 168 564340
rect 0 564256 112 564284
rect 0 563444 112 563472
rect 0 563388 168 563444
rect 0 563360 112 563388
rect 0 562548 112 562576
rect 0 562492 168 562548
rect 0 562464 112 562492
rect 0 561652 112 561680
rect 0 561596 168 561652
rect 0 561568 112 561596
rect 0 560756 112 560784
rect 0 560700 168 560756
rect 0 560672 112 560700
rect 0 559860 112 559888
rect 0 559804 168 559860
rect 0 559776 112 559804
rect 0 558964 112 558992
rect 0 558908 168 558964
rect 0 558880 112 558908
rect 0 558068 112 558096
rect 0 558012 168 558068
rect 0 557984 112 558012
rect 0 557172 112 557200
rect 0 557116 168 557172
rect 0 557088 112 557116
rect 0 556276 112 556304
rect 0 556220 168 556276
rect 0 556192 112 556220
rect 0 555380 112 555408
rect 0 555324 168 555380
rect 0 555296 112 555324
rect 0 554484 112 554512
rect 0 554428 168 554484
rect 0 554400 112 554428
rect 0 553588 112 553616
rect 0 553532 168 553588
rect 0 553504 112 553532
rect 0 552692 112 552720
rect 0 552636 168 552692
rect 0 552608 112 552636
rect 0 551796 112 551824
rect 0 551740 168 551796
rect 0 551712 112 551740
rect 0 550900 112 550928
rect 0 550844 168 550900
rect 0 550816 112 550844
rect 0 550004 112 550032
rect 0 549948 168 550004
rect 0 549920 112 549948
rect 0 549108 112 549136
rect 0 549052 168 549108
rect 0 549024 112 549052
rect 0 548212 112 548240
rect 0 548156 168 548212
rect 0 548128 112 548156
rect 0 547316 112 547344
rect 0 547260 168 547316
rect 0 547232 112 547260
rect 0 546420 112 546448
rect 0 546364 168 546420
rect 0 546336 112 546364
rect 0 545524 112 545552
rect 0 545468 168 545524
rect 0 545440 112 545468
rect 0 544628 112 544656
rect 0 544572 168 544628
rect 0 544544 112 544572
rect 0 543732 112 543760
rect 0 543676 168 543732
rect 0 543648 112 543676
rect 0 542836 112 542864
rect 0 542780 168 542836
rect 0 542752 112 542780
rect 0 541940 112 541968
rect 0 541884 168 541940
rect 0 541856 112 541884
rect 0 541044 112 541072
rect 0 540988 168 541044
rect 0 540960 112 540988
rect 0 540148 112 540176
rect 0 540092 168 540148
rect 0 540064 112 540092
rect 0 539252 112 539280
rect 0 539196 168 539252
rect 0 539168 112 539196
rect 0 538356 112 538384
rect 0 538300 168 538356
rect 0 538272 112 538300
rect 0 537460 112 537488
rect 0 537404 168 537460
rect 0 537376 112 537404
rect 0 536564 112 536592
rect 0 536508 168 536564
rect 0 536480 112 536508
rect 0 535668 112 535696
rect 0 535612 168 535668
rect 0 535584 112 535612
rect 0 534772 112 534800
rect 0 534716 168 534772
rect 0 534688 112 534716
rect 0 530180 112 530208
rect 0 530124 168 530180
rect 0 530096 112 530124
rect 0 529284 112 529312
rect 0 529228 168 529284
rect 0 529200 112 529228
rect 0 528388 112 528416
rect 0 528332 168 528388
rect 0 528304 112 528332
rect 0 527492 112 527520
rect 0 527436 168 527492
rect 0 527408 112 527436
rect 0 526596 112 526624
rect 0 526540 168 526596
rect 0 526512 112 526540
rect 0 525700 112 525728
rect 0 525644 168 525700
rect 0 525616 112 525644
rect 0 524804 112 524832
rect 0 524748 168 524804
rect 0 524720 112 524748
rect 0 523908 112 523936
rect 0 523852 168 523908
rect 0 523824 112 523852
rect 0 523012 112 523040
rect 0 522956 168 523012
rect 0 522928 112 522956
rect 0 522116 112 522144
rect 0 522060 168 522116
rect 0 522032 112 522060
rect 0 521220 112 521248
rect 0 521164 168 521220
rect 0 521136 112 521164
rect 0 520324 112 520352
rect 0 520268 168 520324
rect 0 520240 112 520268
rect 0 519428 112 519456
rect 0 519372 168 519428
rect 0 519344 112 519372
rect 0 518532 112 518560
rect 0 518476 168 518532
rect 0 518448 112 518476
rect 0 517636 112 517664
rect 0 517580 168 517636
rect 0 517552 112 517580
rect 0 516740 112 516768
rect 0 516684 168 516740
rect 0 516656 112 516684
rect 0 515844 112 515872
rect 0 515788 168 515844
rect 0 515760 112 515788
rect 0 514948 112 514976
rect 0 514892 168 514948
rect 0 514864 112 514892
rect 0 514052 112 514080
rect 0 513996 168 514052
rect 0 513968 112 513996
rect 0 513156 112 513184
rect 0 513100 168 513156
rect 0 513072 112 513100
rect 0 512260 112 512288
rect 0 512204 168 512260
rect 0 512176 112 512204
rect 0 511364 112 511392
rect 0 511308 168 511364
rect 0 511280 112 511308
rect 0 510468 112 510496
rect 0 510412 168 510468
rect 0 510384 112 510412
rect 464800 510244 464912 510272
rect 464772 510188 464912 510244
rect 464800 510160 464912 510188
rect 0 509572 112 509600
rect 0 509516 168 509572
rect 0 509488 112 509516
rect 464800 509348 464912 509376
rect 464772 509292 464912 509348
rect 464800 509264 464912 509292
rect 0 508676 112 508704
rect 0 508620 168 508676
rect 0 508592 112 508620
rect 464800 508452 464912 508480
rect 464772 508396 464912 508452
rect 464800 508368 464912 508396
rect 0 507780 112 507808
rect 0 507724 168 507780
rect 0 507696 112 507724
rect 464800 507556 464912 507584
rect 464772 507500 464912 507556
rect 464800 507472 464912 507500
rect 0 506884 112 506912
rect 0 506828 168 506884
rect 0 506800 112 506828
rect 464800 506660 464912 506688
rect 464772 506604 464912 506660
rect 464800 506576 464912 506604
rect 0 505988 112 506016
rect 0 505932 168 505988
rect 0 505904 112 505932
rect 464800 505764 464912 505792
rect 464772 505708 464912 505764
rect 464800 505680 464912 505708
rect 0 505092 112 505120
rect 0 505036 168 505092
rect 0 505008 112 505036
rect 464800 504868 464912 504896
rect 464772 504812 464912 504868
rect 464800 504784 464912 504812
rect 0 504196 112 504224
rect 0 504140 168 504196
rect 0 504112 112 504140
rect 464800 503972 464912 504000
rect 464772 503916 464912 503972
rect 464800 503888 464912 503916
rect 0 503300 112 503328
rect 0 503244 168 503300
rect 0 503216 112 503244
rect 464800 503076 464912 503104
rect 464772 503020 464912 503076
rect 464800 502992 464912 503020
rect 0 502404 112 502432
rect 0 502348 168 502404
rect 0 502320 112 502348
rect 464800 502180 464912 502208
rect 464772 502124 464912 502180
rect 464800 502096 464912 502124
rect 0 501508 112 501536
rect 0 501452 168 501508
rect 0 501424 112 501452
rect 464800 501284 464912 501312
rect 464772 501228 464912 501284
rect 464800 501200 464912 501228
rect 0 500612 112 500640
rect 0 500556 168 500612
rect 0 500528 112 500556
rect 464800 500388 464912 500416
rect 464772 500332 464912 500388
rect 464800 500304 464912 500332
rect 0 499716 112 499744
rect 0 499660 168 499716
rect 0 499632 112 499660
rect 464800 499492 464912 499520
rect 464772 499436 464912 499492
rect 464800 499408 464912 499436
rect 0 498820 112 498848
rect 0 498764 168 498820
rect 0 498736 112 498764
rect 464800 498596 464912 498624
rect 464772 498540 464912 498596
rect 464800 498512 464912 498540
rect 0 497924 112 497952
rect 0 497868 168 497924
rect 0 497840 112 497868
rect 464800 497700 464912 497728
rect 464772 497644 464912 497700
rect 464800 497616 464912 497644
rect 0 497028 112 497056
rect 0 496972 168 497028
rect 0 496944 112 496972
rect 464800 496804 464912 496832
rect 464772 496748 464912 496804
rect 464800 496720 464912 496748
rect 0 496132 112 496160
rect 0 496076 168 496132
rect 0 496048 112 496076
rect 464800 495908 464912 495936
rect 464772 495852 464912 495908
rect 464800 495824 464912 495852
rect 0 495236 112 495264
rect 0 495180 168 495236
rect 0 495152 112 495180
rect 464800 495012 464912 495040
rect 464772 494956 464912 495012
rect 464800 494928 464912 494956
rect 0 494340 112 494368
rect 0 494284 168 494340
rect 0 494256 112 494284
rect 464800 494116 464912 494144
rect 464772 494060 464912 494116
rect 464800 494032 464912 494060
rect 0 493444 112 493472
rect 0 493388 168 493444
rect 0 493360 112 493388
rect 464800 493220 464912 493248
rect 464772 493164 464912 493220
rect 464800 493136 464912 493164
rect 0 492548 112 492576
rect 0 492492 168 492548
rect 0 492464 112 492492
rect 464800 492324 464912 492352
rect 464772 492268 464912 492324
rect 464800 492240 464912 492268
rect 0 491652 112 491680
rect 0 491596 168 491652
rect 0 491568 112 491596
rect 464800 491428 464912 491456
rect 464772 491372 464912 491428
rect 464800 491344 464912 491372
rect 0 490756 112 490784
rect 0 490700 168 490756
rect 0 490672 112 490700
rect 464800 490532 464912 490560
rect 464772 490476 464912 490532
rect 464800 490448 464912 490476
rect 0 489860 112 489888
rect 0 489804 168 489860
rect 0 489776 112 489804
rect 464800 489636 464912 489664
rect 464772 489580 464912 489636
rect 464800 489552 464912 489580
rect 0 488964 112 488992
rect 0 488908 168 488964
rect 0 488880 112 488908
rect 464800 488740 464912 488768
rect 464772 488684 464912 488740
rect 464800 488656 464912 488684
rect 0 488068 112 488096
rect 0 488012 168 488068
rect 0 487984 112 488012
rect 464800 487844 464912 487872
rect 464772 487788 464912 487844
rect 464800 487760 464912 487788
rect 0 487172 112 487200
rect 0 487116 168 487172
rect 0 487088 112 487116
rect 464800 486948 464912 486976
rect 464772 486892 464912 486948
rect 464800 486864 464912 486892
rect 0 486276 112 486304
rect 0 486220 168 486276
rect 0 486192 112 486220
rect 464800 486052 464912 486080
rect 464772 485996 464912 486052
rect 464800 485968 464912 485996
rect 0 485380 112 485408
rect 0 485324 168 485380
rect 0 485296 112 485324
rect 464800 485156 464912 485184
rect 464772 485100 464912 485156
rect 464800 485072 464912 485100
rect 0 484484 112 484512
rect 0 484428 168 484484
rect 0 484400 112 484428
rect 464800 484260 464912 484288
rect 464772 484204 464912 484260
rect 464800 484176 464912 484204
rect 0 483588 112 483616
rect 0 483532 168 483588
rect 0 483504 112 483532
rect 464800 483364 464912 483392
rect 464772 483308 464912 483364
rect 464800 483280 464912 483308
rect 0 482692 112 482720
rect 0 482636 168 482692
rect 0 482608 112 482636
rect 464800 482468 464912 482496
rect 464772 482412 464912 482468
rect 464800 482384 464912 482412
rect 0 481796 112 481824
rect 0 481740 168 481796
rect 0 481712 112 481740
rect 464800 481572 464912 481600
rect 464772 481516 464912 481572
rect 464800 481488 464912 481516
rect 0 480900 112 480928
rect 0 480844 168 480900
rect 0 480816 112 480844
rect 464800 480676 464912 480704
rect 464772 480620 464912 480676
rect 464800 480592 464912 480620
rect 0 480004 112 480032
rect 0 479948 168 480004
rect 0 479920 112 479948
rect 464800 479780 464912 479808
rect 464772 479724 464912 479780
rect 464800 479696 464912 479724
rect 0 479108 112 479136
rect 0 479052 168 479108
rect 0 479024 112 479052
rect 464800 478884 464912 478912
rect 464772 478828 464912 478884
rect 464800 478800 464912 478828
rect 0 478212 112 478240
rect 0 478156 168 478212
rect 0 478128 112 478156
rect 464800 477988 464912 478016
rect 464772 477932 464912 477988
rect 464800 477904 464912 477932
rect 0 477316 112 477344
rect 0 477260 168 477316
rect 0 477232 112 477260
rect 0 472724 112 472752
rect 0 472668 168 472724
rect 0 472640 112 472668
rect 0 471828 112 471856
rect 0 471772 168 471828
rect 0 471744 112 471772
rect 0 470932 112 470960
rect 0 470876 168 470932
rect 0 470848 112 470876
rect 0 470036 112 470064
rect 0 469980 168 470036
rect 0 469952 112 469980
rect 0 469140 112 469168
rect 0 469084 168 469140
rect 0 469056 112 469084
rect 0 468244 112 468272
rect 0 468188 168 468244
rect 0 468160 112 468188
rect 0 467348 112 467376
rect 0 467292 168 467348
rect 0 467264 112 467292
rect 0 466452 112 466480
rect 0 466396 168 466452
rect 0 466368 112 466396
rect 0 465556 112 465584
rect 0 465500 168 465556
rect 0 465472 112 465500
rect 0 464660 112 464688
rect 0 464604 168 464660
rect 0 464576 112 464604
rect 0 463764 112 463792
rect 0 463708 168 463764
rect 0 463680 112 463708
rect 0 462868 112 462896
rect 0 462812 168 462868
rect 0 462784 112 462812
rect 0 461972 112 462000
rect 0 461916 168 461972
rect 0 461888 112 461916
rect 0 461076 112 461104
rect 0 461020 168 461076
rect 0 460992 112 461020
rect 0 460180 112 460208
rect 0 460124 168 460180
rect 0 460096 112 460124
rect 0 459284 112 459312
rect 0 459228 168 459284
rect 0 459200 112 459228
rect 0 458388 112 458416
rect 0 458332 168 458388
rect 0 458304 112 458332
rect 0 457492 112 457520
rect 0 457436 168 457492
rect 0 457408 112 457436
rect 0 456596 112 456624
rect 0 456540 168 456596
rect 0 456512 112 456540
rect 0 455700 112 455728
rect 0 455644 168 455700
rect 0 455616 112 455644
rect 0 454804 112 454832
rect 0 454748 168 454804
rect 0 454720 112 454748
rect 0 453908 112 453936
rect 0 453852 168 453908
rect 0 453824 112 453852
rect 0 453012 112 453040
rect 0 452956 168 453012
rect 0 452928 112 452956
rect 0 452116 112 452144
rect 0 452060 168 452116
rect 0 452032 112 452060
rect 0 451220 112 451248
rect 0 451164 168 451220
rect 0 451136 112 451164
rect 0 450324 112 450352
rect 0 450268 168 450324
rect 0 450240 112 450268
rect 0 449428 112 449456
rect 0 449372 168 449428
rect 0 449344 112 449372
rect 0 448532 112 448560
rect 0 448476 168 448532
rect 0 448448 112 448476
rect 0 447636 112 447664
rect 0 447580 168 447636
rect 0 447552 112 447580
rect 0 446740 112 446768
rect 0 446684 168 446740
rect 0 446656 112 446684
rect 0 445844 112 445872
rect 0 445788 168 445844
rect 0 445760 112 445788
rect 0 444948 112 444976
rect 0 444892 168 444948
rect 0 444864 112 444892
rect 0 444052 112 444080
rect 0 443996 168 444052
rect 0 443968 112 443996
rect 0 443156 112 443184
rect 0 443100 168 443156
rect 0 443072 112 443100
rect 0 442260 112 442288
rect 0 442204 168 442260
rect 0 442176 112 442204
rect 0 441364 112 441392
rect 0 441308 168 441364
rect 0 441280 112 441308
rect 0 440468 112 440496
rect 0 440412 168 440468
rect 0 440384 112 440412
rect 0 439572 112 439600
rect 0 439516 168 439572
rect 0 439488 112 439516
rect 0 438676 112 438704
rect 0 438620 168 438676
rect 0 438592 112 438620
rect 0 437780 112 437808
rect 0 437724 168 437780
rect 0 437696 112 437724
rect 0 436884 112 436912
rect 0 436828 168 436884
rect 0 436800 112 436828
rect 0 435988 112 436016
rect 0 435932 168 435988
rect 0 435904 112 435932
rect 0 435092 112 435120
rect 0 435036 168 435092
rect 0 435008 112 435036
rect 0 434196 112 434224
rect 0 434140 168 434196
rect 0 434112 112 434140
rect 0 433300 112 433328
rect 0 433244 168 433300
rect 0 433216 112 433244
rect 0 432404 112 432432
rect 0 432348 168 432404
rect 0 432320 112 432348
rect 0 431508 112 431536
rect 0 431452 168 431508
rect 0 431424 112 431452
rect 0 430612 112 430640
rect 0 430556 168 430612
rect 0 430528 112 430556
rect 0 429716 112 429744
rect 0 429660 168 429716
rect 0 429632 112 429660
rect 0 428820 112 428848
rect 0 428764 168 428820
rect 0 428736 112 428764
rect 0 427924 112 427952
rect 0 427868 168 427924
rect 0 427840 112 427868
rect 0 427028 112 427056
rect 0 426972 168 427028
rect 0 426944 112 426972
rect 0 426132 112 426160
rect 0 426076 168 426132
rect 0 426048 112 426076
rect 0 425236 112 425264
rect 0 425180 168 425236
rect 0 425152 112 425180
rect 0 424340 112 424368
rect 0 424284 168 424340
rect 0 424256 112 424284
rect 0 423444 112 423472
rect 0 423388 168 423444
rect 0 423360 112 423388
rect 0 422548 112 422576
rect 0 422492 168 422548
rect 0 422464 112 422492
rect 0 421652 112 421680
rect 0 421596 168 421652
rect 0 421568 112 421596
rect 0 420756 112 420784
rect 0 420700 168 420756
rect 0 420672 112 420700
rect 0 419860 112 419888
rect 0 419804 168 419860
rect 0 419776 112 419804
rect 0 415268 112 415296
rect 0 415212 168 415268
rect 0 415184 112 415212
rect 0 414372 112 414400
rect 0 414316 168 414372
rect 0 414288 112 414316
rect 0 413476 112 413504
rect 0 413420 168 413476
rect 0 413392 112 413420
rect 0 412580 112 412608
rect 0 412524 168 412580
rect 0 412496 112 412524
rect 0 411684 112 411712
rect 0 411628 168 411684
rect 0 411600 112 411628
rect 0 410788 112 410816
rect 0 410732 168 410788
rect 0 410704 112 410732
rect 0 409892 112 409920
rect 0 409836 168 409892
rect 0 409808 112 409836
rect 0 408996 112 409024
rect 0 408940 168 408996
rect 0 408912 112 408940
rect 0 408100 112 408128
rect 0 408044 168 408100
rect 0 408016 112 408044
rect 0 407204 112 407232
rect 0 407148 168 407204
rect 0 407120 112 407148
rect 0 406308 112 406336
rect 0 406252 168 406308
rect 0 406224 112 406252
rect 0 405412 112 405440
rect 0 405356 168 405412
rect 0 405328 112 405356
rect 0 404516 112 404544
rect 0 404460 168 404516
rect 0 404432 112 404460
rect 0 403620 112 403648
rect 0 403564 168 403620
rect 0 403536 112 403564
rect 0 402724 112 402752
rect 0 402668 168 402724
rect 0 402640 112 402668
rect 0 401828 112 401856
rect 0 401772 168 401828
rect 0 401744 112 401772
rect 0 400932 112 400960
rect 0 400876 168 400932
rect 0 400848 112 400876
rect 0 400036 112 400064
rect 0 399980 168 400036
rect 0 399952 112 399980
rect 0 399140 112 399168
rect 0 399084 168 399140
rect 0 399056 112 399084
rect 0 398244 112 398272
rect 0 398188 168 398244
rect 0 398160 112 398188
rect 0 397348 112 397376
rect 0 397292 168 397348
rect 0 397264 112 397292
rect 0 396452 112 396480
rect 0 396396 168 396452
rect 0 396368 112 396396
rect 0 395556 112 395584
rect 0 395500 168 395556
rect 0 395472 112 395500
rect 464800 395332 464912 395360
rect 464772 395276 464912 395332
rect 464800 395248 464912 395276
rect 0 394660 112 394688
rect 0 394604 168 394660
rect 0 394576 112 394604
rect 464800 394436 464912 394464
rect 464772 394380 464912 394436
rect 464800 394352 464912 394380
rect 0 393764 112 393792
rect 0 393708 168 393764
rect 0 393680 112 393708
rect 464800 393540 464912 393568
rect 464772 393484 464912 393540
rect 464800 393456 464912 393484
rect 0 392868 112 392896
rect 0 392812 168 392868
rect 0 392784 112 392812
rect 464800 392644 464912 392672
rect 464772 392588 464912 392644
rect 464800 392560 464912 392588
rect 0 391972 112 392000
rect 0 391916 168 391972
rect 0 391888 112 391916
rect 464800 391748 464912 391776
rect 464772 391692 464912 391748
rect 464800 391664 464912 391692
rect 0 391076 112 391104
rect 0 391020 168 391076
rect 0 390992 112 391020
rect 464800 390852 464912 390880
rect 464772 390796 464912 390852
rect 464800 390768 464912 390796
rect 0 390180 112 390208
rect 0 390124 168 390180
rect 0 390096 112 390124
rect 464800 389956 464912 389984
rect 464772 389900 464912 389956
rect 464800 389872 464912 389900
rect 0 389284 112 389312
rect 0 389228 168 389284
rect 0 389200 112 389228
rect 464800 389060 464912 389088
rect 464772 389004 464912 389060
rect 464800 388976 464912 389004
rect 0 388388 112 388416
rect 0 388332 168 388388
rect 0 388304 112 388332
rect 464800 388164 464912 388192
rect 464772 388108 464912 388164
rect 464800 388080 464912 388108
rect 0 387492 112 387520
rect 0 387436 168 387492
rect 0 387408 112 387436
rect 464800 387268 464912 387296
rect 464772 387212 464912 387268
rect 464800 387184 464912 387212
rect 0 386596 112 386624
rect 0 386540 168 386596
rect 0 386512 112 386540
rect 464800 386372 464912 386400
rect 464772 386316 464912 386372
rect 464800 386288 464912 386316
rect 0 385700 112 385728
rect 0 385644 168 385700
rect 0 385616 112 385644
rect 464800 385476 464912 385504
rect 464772 385420 464912 385476
rect 464800 385392 464912 385420
rect 0 384804 112 384832
rect 0 384748 168 384804
rect 0 384720 112 384748
rect 464800 384580 464912 384608
rect 464772 384524 464912 384580
rect 464800 384496 464912 384524
rect 0 383908 112 383936
rect 0 383852 168 383908
rect 0 383824 112 383852
rect 464800 383684 464912 383712
rect 464772 383628 464912 383684
rect 464800 383600 464912 383628
rect 0 383012 112 383040
rect 0 382956 168 383012
rect 0 382928 112 382956
rect 464800 382788 464912 382816
rect 464772 382732 464912 382788
rect 464800 382704 464912 382732
rect 0 382116 112 382144
rect 0 382060 168 382116
rect 0 382032 112 382060
rect 464800 381892 464912 381920
rect 464772 381836 464912 381892
rect 464800 381808 464912 381836
rect 0 381220 112 381248
rect 0 381164 168 381220
rect 0 381136 112 381164
rect 464800 380996 464912 381024
rect 464772 380940 464912 380996
rect 464800 380912 464912 380940
rect 0 380324 112 380352
rect 0 380268 168 380324
rect 0 380240 112 380268
rect 464800 380100 464912 380128
rect 464772 380044 464912 380100
rect 464800 380016 464912 380044
rect 0 379428 112 379456
rect 0 379372 168 379428
rect 0 379344 112 379372
rect 464800 379204 464912 379232
rect 464772 379148 464912 379204
rect 464800 379120 464912 379148
rect 0 378532 112 378560
rect 0 378476 168 378532
rect 0 378448 112 378476
rect 464800 378308 464912 378336
rect 464772 378252 464912 378308
rect 464800 378224 464912 378252
rect 0 377636 112 377664
rect 0 377580 168 377636
rect 0 377552 112 377580
rect 464800 377412 464912 377440
rect 464772 377356 464912 377412
rect 464800 377328 464912 377356
rect 0 376740 112 376768
rect 0 376684 168 376740
rect 0 376656 112 376684
rect 464800 376516 464912 376544
rect 464772 376460 464912 376516
rect 464800 376432 464912 376460
rect 0 375844 112 375872
rect 0 375788 168 375844
rect 0 375760 112 375788
rect 464800 375620 464912 375648
rect 464772 375564 464912 375620
rect 464800 375536 464912 375564
rect 0 374948 112 374976
rect 0 374892 168 374948
rect 0 374864 112 374892
rect 464800 374724 464912 374752
rect 464772 374668 464912 374724
rect 464800 374640 464912 374668
rect 0 374052 112 374080
rect 0 373996 168 374052
rect 0 373968 112 373996
rect 464800 373828 464912 373856
rect 464772 373772 464912 373828
rect 464800 373744 464912 373772
rect 0 373156 112 373184
rect 0 373100 168 373156
rect 0 373072 112 373100
rect 464800 372932 464912 372960
rect 464772 372876 464912 372932
rect 464800 372848 464912 372876
rect 0 372260 112 372288
rect 0 372204 168 372260
rect 0 372176 112 372204
rect 464800 372036 464912 372064
rect 464772 371980 464912 372036
rect 464800 371952 464912 371980
rect 0 371364 112 371392
rect 0 371308 168 371364
rect 0 371280 112 371308
rect 464800 371140 464912 371168
rect 464772 371084 464912 371140
rect 464800 371056 464912 371084
rect 0 370468 112 370496
rect 0 370412 168 370468
rect 0 370384 112 370412
rect 464800 370244 464912 370272
rect 464772 370188 464912 370244
rect 464800 370160 464912 370188
rect 0 369572 112 369600
rect 0 369516 168 369572
rect 0 369488 112 369516
rect 464800 369348 464912 369376
rect 464772 369292 464912 369348
rect 464800 369264 464912 369292
rect 0 368676 112 368704
rect 0 368620 168 368676
rect 0 368592 112 368620
rect 464800 368452 464912 368480
rect 464772 368396 464912 368452
rect 464800 368368 464912 368396
rect 0 367780 112 367808
rect 0 367724 168 367780
rect 0 367696 112 367724
rect 464800 367556 464912 367584
rect 464772 367500 464912 367556
rect 464800 367472 464912 367500
rect 0 366884 112 366912
rect 0 366828 168 366884
rect 0 366800 112 366828
rect 464800 366660 464912 366688
rect 464772 366604 464912 366660
rect 464800 366576 464912 366604
rect 0 365988 112 366016
rect 0 365932 168 365988
rect 0 365904 112 365932
rect 464800 365764 464912 365792
rect 464772 365708 464912 365764
rect 464800 365680 464912 365708
rect 0 365092 112 365120
rect 0 365036 168 365092
rect 0 365008 112 365036
rect 464800 364868 464912 364896
rect 464772 364812 464912 364868
rect 464800 364784 464912 364812
rect 0 364196 112 364224
rect 0 364140 168 364196
rect 0 364112 112 364140
rect 464800 363972 464912 364000
rect 464772 363916 464912 363972
rect 464800 363888 464912 363916
rect 0 363300 112 363328
rect 0 363244 168 363300
rect 0 363216 112 363244
rect 464800 363076 464912 363104
rect 464772 363020 464912 363076
rect 464800 362992 464912 363020
rect 0 362404 112 362432
rect 0 362348 168 362404
rect 0 362320 112 362348
rect 0 357812 112 357840
rect 0 357756 168 357812
rect 0 357728 112 357756
rect 0 356916 112 356944
rect 0 356860 168 356916
rect 0 356832 112 356860
rect 0 356020 112 356048
rect 0 355964 168 356020
rect 0 355936 112 355964
rect 0 355124 112 355152
rect 0 355068 168 355124
rect 0 355040 112 355068
rect 0 354228 112 354256
rect 0 354172 168 354228
rect 0 354144 112 354172
rect 0 353332 112 353360
rect 0 353276 168 353332
rect 0 353248 112 353276
rect 0 352436 112 352464
rect 0 352380 168 352436
rect 0 352352 112 352380
rect 0 351540 112 351568
rect 0 351484 168 351540
rect 0 351456 112 351484
rect 0 350644 112 350672
rect 0 350588 168 350644
rect 0 350560 112 350588
rect 0 349748 112 349776
rect 0 349692 168 349748
rect 0 349664 112 349692
rect 0 348852 112 348880
rect 0 348796 168 348852
rect 0 348768 112 348796
rect 0 347956 112 347984
rect 0 347900 168 347956
rect 0 347872 112 347900
rect 0 347060 112 347088
rect 0 347004 168 347060
rect 0 346976 112 347004
rect 0 346164 112 346192
rect 0 346108 168 346164
rect 0 346080 112 346108
rect 0 345268 112 345296
rect 0 345212 168 345268
rect 0 345184 112 345212
rect 0 344372 112 344400
rect 0 344316 168 344372
rect 0 344288 112 344316
rect 0 343476 112 343504
rect 0 343420 168 343476
rect 0 343392 112 343420
rect 0 342580 112 342608
rect 0 342524 168 342580
rect 0 342496 112 342524
rect 0 341684 112 341712
rect 0 341628 168 341684
rect 0 341600 112 341628
rect 0 340788 112 340816
rect 0 340732 168 340788
rect 0 340704 112 340732
rect 0 339892 112 339920
rect 0 339836 168 339892
rect 0 339808 112 339836
rect 0 338996 112 339024
rect 0 338940 168 338996
rect 0 338912 112 338940
rect 0 338100 112 338128
rect 0 338044 168 338100
rect 0 338016 112 338044
rect 0 337204 112 337232
rect 0 337148 168 337204
rect 0 337120 112 337148
rect 0 336308 112 336336
rect 0 336252 168 336308
rect 0 336224 112 336252
rect 0 335412 112 335440
rect 0 335356 168 335412
rect 0 335328 112 335356
rect 0 334516 112 334544
rect 0 334460 168 334516
rect 0 334432 112 334460
rect 0 333620 112 333648
rect 0 333564 168 333620
rect 0 333536 112 333564
rect 0 332724 112 332752
rect 0 332668 168 332724
rect 0 332640 112 332668
rect 0 331828 112 331856
rect 0 331772 168 331828
rect 0 331744 112 331772
rect 0 330932 112 330960
rect 0 330876 168 330932
rect 0 330848 112 330876
rect 0 330036 112 330064
rect 0 329980 168 330036
rect 0 329952 112 329980
rect 0 329140 112 329168
rect 0 329084 168 329140
rect 0 329056 112 329084
rect 0 328244 112 328272
rect 0 328188 168 328244
rect 0 328160 112 328188
rect 0 327348 112 327376
rect 0 327292 168 327348
rect 0 327264 112 327292
rect 0 326452 112 326480
rect 0 326396 168 326452
rect 0 326368 112 326396
rect 0 325556 112 325584
rect 0 325500 168 325556
rect 0 325472 112 325500
rect 0 324660 112 324688
rect 0 324604 168 324660
rect 0 324576 112 324604
rect 0 323764 112 323792
rect 0 323708 168 323764
rect 0 323680 112 323708
rect 0 322868 112 322896
rect 0 322812 168 322868
rect 0 322784 112 322812
rect 0 321972 112 322000
rect 0 321916 168 321972
rect 0 321888 112 321916
rect 0 321076 112 321104
rect 0 321020 168 321076
rect 0 320992 112 321020
rect 0 320180 112 320208
rect 0 320124 168 320180
rect 0 320096 112 320124
rect 0 319284 112 319312
rect 0 319228 168 319284
rect 0 319200 112 319228
rect 0 318388 112 318416
rect 0 318332 168 318388
rect 0 318304 112 318332
rect 0 317492 112 317520
rect 0 317436 168 317492
rect 0 317408 112 317436
rect 0 316596 112 316624
rect 0 316540 168 316596
rect 0 316512 112 316540
rect 0 315700 112 315728
rect 0 315644 168 315700
rect 0 315616 112 315644
rect 0 314804 112 314832
rect 0 314748 168 314804
rect 0 314720 112 314748
rect 0 313908 112 313936
rect 0 313852 168 313908
rect 0 313824 112 313852
rect 0 313012 112 313040
rect 0 312956 168 313012
rect 0 312928 112 312956
rect 0 312116 112 312144
rect 0 312060 168 312116
rect 0 312032 112 312060
rect 0 311220 112 311248
rect 0 311164 168 311220
rect 0 311136 112 311164
rect 0 310324 112 310352
rect 0 310268 168 310324
rect 0 310240 112 310268
rect 0 309428 112 309456
rect 0 309372 168 309428
rect 0 309344 112 309372
rect 0 308532 112 308560
rect 0 308476 168 308532
rect 0 308448 112 308476
rect 0 307636 112 307664
rect 0 307580 168 307636
rect 0 307552 112 307580
rect 0 306740 112 306768
rect 0 306684 168 306740
rect 0 306656 112 306684
rect 0 305844 112 305872
rect 0 305788 168 305844
rect 0 305760 112 305788
rect 0 304948 112 304976
rect 0 304892 168 304948
rect 0 304864 112 304892
rect 0 300356 112 300384
rect 0 300300 168 300356
rect 0 300272 112 300300
rect 0 299460 112 299488
rect 0 299404 168 299460
rect 0 299376 112 299404
rect 0 298564 112 298592
rect 0 298508 168 298564
rect 0 298480 112 298508
rect 0 297668 112 297696
rect 0 297612 168 297668
rect 0 297584 112 297612
rect 0 296772 112 296800
rect 0 296716 168 296772
rect 0 296688 112 296716
rect 0 295876 112 295904
rect 0 295820 168 295876
rect 0 295792 112 295820
rect 0 294980 112 295008
rect 0 294924 168 294980
rect 0 294896 112 294924
rect 0 294084 112 294112
rect 0 294028 168 294084
rect 0 294000 112 294028
rect 0 293188 112 293216
rect 0 293132 168 293188
rect 0 293104 112 293132
rect 0 292292 112 292320
rect 0 292236 168 292292
rect 0 292208 112 292236
rect 0 291396 112 291424
rect 0 291340 168 291396
rect 0 291312 112 291340
rect 0 290500 112 290528
rect 0 290444 168 290500
rect 0 290416 112 290444
rect 0 289604 112 289632
rect 0 289548 168 289604
rect 0 289520 112 289548
rect 0 288708 112 288736
rect 0 288652 168 288708
rect 0 288624 112 288652
rect 0 287812 112 287840
rect 0 287756 168 287812
rect 0 287728 112 287756
rect 0 286916 112 286944
rect 0 286860 168 286916
rect 0 286832 112 286860
rect 0 286020 112 286048
rect 0 285964 168 286020
rect 0 285936 112 285964
rect 0 285124 112 285152
rect 0 285068 168 285124
rect 0 285040 112 285068
rect 0 284228 112 284256
rect 0 284172 168 284228
rect 0 284144 112 284172
rect 0 283332 112 283360
rect 0 283276 168 283332
rect 0 283248 112 283276
rect 0 282436 112 282464
rect 0 282380 168 282436
rect 0 282352 112 282380
rect 0 281540 112 281568
rect 0 281484 168 281540
rect 0 281456 112 281484
rect 0 280644 112 280672
rect 0 280588 168 280644
rect 0 280560 112 280588
rect 464800 280420 464912 280448
rect 464772 280364 464912 280420
rect 464800 280336 464912 280364
rect 0 279748 112 279776
rect 0 279692 168 279748
rect 0 279664 112 279692
rect 464800 279524 464912 279552
rect 464772 279468 464912 279524
rect 464800 279440 464912 279468
rect 0 278852 112 278880
rect 0 278796 168 278852
rect 0 278768 112 278796
rect 464800 278628 464912 278656
rect 464772 278572 464912 278628
rect 464800 278544 464912 278572
rect 0 277956 112 277984
rect 0 277900 168 277956
rect 0 277872 112 277900
rect 464800 277732 464912 277760
rect 464772 277676 464912 277732
rect 464800 277648 464912 277676
rect 0 277060 112 277088
rect 0 277004 168 277060
rect 0 276976 112 277004
rect 464800 276836 464912 276864
rect 464772 276780 464912 276836
rect 464800 276752 464912 276780
rect 0 276164 112 276192
rect 0 276108 168 276164
rect 0 276080 112 276108
rect 464800 275940 464912 275968
rect 464772 275884 464912 275940
rect 464800 275856 464912 275884
rect 0 275268 112 275296
rect 0 275212 168 275268
rect 0 275184 112 275212
rect 464800 275044 464912 275072
rect 464772 274988 464912 275044
rect 464800 274960 464912 274988
rect 0 274372 112 274400
rect 0 274316 168 274372
rect 0 274288 112 274316
rect 464800 274148 464912 274176
rect 464772 274092 464912 274148
rect 464800 274064 464912 274092
rect 0 273476 112 273504
rect 0 273420 168 273476
rect 0 273392 112 273420
rect 464800 273252 464912 273280
rect 464772 273196 464912 273252
rect 464800 273168 464912 273196
rect 0 272580 112 272608
rect 0 272524 168 272580
rect 0 272496 112 272524
rect 464800 272356 464912 272384
rect 464772 272300 464912 272356
rect 464800 272272 464912 272300
rect 0 271684 112 271712
rect 0 271628 168 271684
rect 0 271600 112 271628
rect 464800 271460 464912 271488
rect 464772 271404 464912 271460
rect 464800 271376 464912 271404
rect 0 270788 112 270816
rect 0 270732 168 270788
rect 0 270704 112 270732
rect 464800 270564 464912 270592
rect 464772 270508 464912 270564
rect 464800 270480 464912 270508
rect 0 269892 112 269920
rect 0 269836 168 269892
rect 0 269808 112 269836
rect 464800 269668 464912 269696
rect 464772 269612 464912 269668
rect 464800 269584 464912 269612
rect 0 268996 112 269024
rect 0 268940 168 268996
rect 0 268912 112 268940
rect 464800 268772 464912 268800
rect 464772 268716 464912 268772
rect 464800 268688 464912 268716
rect 0 268100 112 268128
rect 0 268044 168 268100
rect 0 268016 112 268044
rect 464800 267876 464912 267904
rect 464772 267820 464912 267876
rect 464800 267792 464912 267820
rect 0 267204 112 267232
rect 0 267148 168 267204
rect 0 267120 112 267148
rect 464800 266980 464912 267008
rect 464772 266924 464912 266980
rect 464800 266896 464912 266924
rect 0 266308 112 266336
rect 0 266252 168 266308
rect 0 266224 112 266252
rect 464800 266084 464912 266112
rect 464772 266028 464912 266084
rect 464800 266000 464912 266028
rect 0 265412 112 265440
rect 0 265356 168 265412
rect 0 265328 112 265356
rect 464800 265188 464912 265216
rect 464772 265132 464912 265188
rect 464800 265104 464912 265132
rect 0 264516 112 264544
rect 0 264460 168 264516
rect 0 264432 112 264460
rect 464800 264292 464912 264320
rect 464772 264236 464912 264292
rect 464800 264208 464912 264236
rect 0 263620 112 263648
rect 0 263564 168 263620
rect 0 263536 112 263564
rect 464800 263396 464912 263424
rect 464772 263340 464912 263396
rect 464800 263312 464912 263340
rect 0 262724 112 262752
rect 0 262668 168 262724
rect 0 262640 112 262668
rect 464800 262500 464912 262528
rect 464772 262444 464912 262500
rect 464800 262416 464912 262444
rect 0 261828 112 261856
rect 0 261772 168 261828
rect 0 261744 112 261772
rect 464800 261604 464912 261632
rect 464772 261548 464912 261604
rect 464800 261520 464912 261548
rect 0 260932 112 260960
rect 0 260876 168 260932
rect 0 260848 112 260876
rect 464800 260708 464912 260736
rect 464772 260652 464912 260708
rect 464800 260624 464912 260652
rect 0 260036 112 260064
rect 0 259980 168 260036
rect 0 259952 112 259980
rect 464800 259812 464912 259840
rect 464772 259756 464912 259812
rect 464800 259728 464912 259756
rect 0 259140 112 259168
rect 0 259084 168 259140
rect 0 259056 112 259084
rect 464800 258916 464912 258944
rect 464772 258860 464912 258916
rect 464800 258832 464912 258860
rect 0 258244 112 258272
rect 0 258188 168 258244
rect 0 258160 112 258188
rect 464800 258020 464912 258048
rect 464772 257964 464912 258020
rect 464800 257936 464912 257964
rect 0 257348 112 257376
rect 0 257292 168 257348
rect 0 257264 112 257292
rect 464800 257124 464912 257152
rect 464772 257068 464912 257124
rect 464800 257040 464912 257068
rect 0 256452 112 256480
rect 0 256396 168 256452
rect 0 256368 112 256396
rect 464800 256228 464912 256256
rect 464772 256172 464912 256228
rect 464800 256144 464912 256172
rect 0 255556 112 255584
rect 0 255500 168 255556
rect 0 255472 112 255500
rect 464800 255332 464912 255360
rect 464772 255276 464912 255332
rect 464800 255248 464912 255276
rect 0 254660 112 254688
rect 0 254604 168 254660
rect 0 254576 112 254604
rect 464800 254436 464912 254464
rect 464772 254380 464912 254436
rect 464800 254352 464912 254380
rect 0 253764 112 253792
rect 0 253708 168 253764
rect 0 253680 112 253708
rect 464800 253540 464912 253568
rect 464772 253484 464912 253540
rect 464800 253456 464912 253484
rect 0 252868 112 252896
rect 0 252812 168 252868
rect 0 252784 112 252812
rect 464800 252644 464912 252672
rect 464772 252588 464912 252644
rect 464800 252560 464912 252588
rect 0 251972 112 252000
rect 0 251916 168 251972
rect 0 251888 112 251916
rect 464800 251748 464912 251776
rect 464772 251692 464912 251748
rect 464800 251664 464912 251692
rect 0 251076 112 251104
rect 0 251020 168 251076
rect 0 250992 112 251020
rect 464800 250852 464912 250880
rect 464772 250796 464912 250852
rect 464800 250768 464912 250796
rect 0 250180 112 250208
rect 0 250124 168 250180
rect 0 250096 112 250124
rect 464800 249956 464912 249984
rect 464772 249900 464912 249956
rect 464800 249872 464912 249900
rect 0 249284 112 249312
rect 0 249228 168 249284
rect 0 249200 112 249228
rect 464800 249060 464912 249088
rect 464772 249004 464912 249060
rect 464800 248976 464912 249004
rect 0 248388 112 248416
rect 0 248332 168 248388
rect 0 248304 112 248332
rect 464800 248164 464912 248192
rect 464772 248108 464912 248164
rect 464800 248080 464912 248108
rect 0 247492 112 247520
rect 0 247436 168 247492
rect 0 247408 112 247436
rect 0 242900 112 242928
rect 0 242844 168 242900
rect 0 242816 112 242844
rect 0 242004 112 242032
rect 0 241948 168 242004
rect 0 241920 112 241948
rect 0 241108 112 241136
rect 0 241052 168 241108
rect 0 241024 112 241052
rect 0 240212 112 240240
rect 0 240156 168 240212
rect 0 240128 112 240156
rect 0 239316 112 239344
rect 0 239260 168 239316
rect 0 239232 112 239260
rect 0 238420 112 238448
rect 0 238364 168 238420
rect 0 238336 112 238364
rect 0 237524 112 237552
rect 0 237468 168 237524
rect 0 237440 112 237468
rect 0 236628 112 236656
rect 0 236572 168 236628
rect 0 236544 112 236572
rect 0 235732 112 235760
rect 0 235676 168 235732
rect 0 235648 112 235676
rect 0 234836 112 234864
rect 0 234780 168 234836
rect 0 234752 112 234780
rect 0 233940 112 233968
rect 0 233884 168 233940
rect 0 233856 112 233884
rect 0 233044 112 233072
rect 0 232988 168 233044
rect 0 232960 112 232988
rect 0 232148 112 232176
rect 0 232092 168 232148
rect 0 232064 112 232092
rect 0 231252 112 231280
rect 0 231196 168 231252
rect 0 231168 112 231196
rect 0 230356 112 230384
rect 0 230300 168 230356
rect 0 230272 112 230300
rect 0 229460 112 229488
rect 0 229404 168 229460
rect 0 229376 112 229404
rect 0 228564 112 228592
rect 0 228508 168 228564
rect 0 228480 112 228508
rect 0 227668 112 227696
rect 0 227612 168 227668
rect 0 227584 112 227612
rect 0 226772 112 226800
rect 0 226716 168 226772
rect 0 226688 112 226716
rect 0 225876 112 225904
rect 0 225820 168 225876
rect 0 225792 112 225820
rect 0 224980 112 225008
rect 0 224924 168 224980
rect 0 224896 112 224924
rect 0 224084 112 224112
rect 0 224028 168 224084
rect 0 224000 112 224028
rect 0 223188 112 223216
rect 0 223132 168 223188
rect 0 223104 112 223132
rect 0 222292 112 222320
rect 0 222236 168 222292
rect 0 222208 112 222236
rect 0 221396 112 221424
rect 0 221340 168 221396
rect 0 221312 112 221340
rect 0 220500 112 220528
rect 0 220444 168 220500
rect 0 220416 112 220444
rect 0 219604 112 219632
rect 0 219548 168 219604
rect 0 219520 112 219548
rect 0 218708 112 218736
rect 0 218652 168 218708
rect 0 218624 112 218652
rect 0 217812 112 217840
rect 0 217756 168 217812
rect 0 217728 112 217756
rect 0 216916 112 216944
rect 0 216860 168 216916
rect 0 216832 112 216860
rect 0 216020 112 216048
rect 0 215964 168 216020
rect 0 215936 112 215964
rect 0 215124 112 215152
rect 0 215068 168 215124
rect 0 215040 112 215068
rect 0 214228 112 214256
rect 0 214172 168 214228
rect 0 214144 112 214172
rect 0 213332 112 213360
rect 0 213276 168 213332
rect 0 213248 112 213276
rect 0 212436 112 212464
rect 0 212380 168 212436
rect 0 212352 112 212380
rect 0 211540 112 211568
rect 0 211484 168 211540
rect 0 211456 112 211484
rect 0 210644 112 210672
rect 0 210588 168 210644
rect 0 210560 112 210588
rect 0 209748 112 209776
rect 0 209692 168 209748
rect 0 209664 112 209692
rect 0 208852 112 208880
rect 0 208796 168 208852
rect 0 208768 112 208796
rect 0 207956 112 207984
rect 0 207900 168 207956
rect 0 207872 112 207900
rect 0 207060 112 207088
rect 0 207004 168 207060
rect 0 206976 112 207004
rect 0 206164 112 206192
rect 0 206108 168 206164
rect 0 206080 112 206108
rect 0 205268 112 205296
rect 0 205212 168 205268
rect 0 205184 112 205212
rect 0 204372 112 204400
rect 0 204316 168 204372
rect 0 204288 112 204316
rect 0 203476 112 203504
rect 0 203420 168 203476
rect 0 203392 112 203420
rect 0 202580 112 202608
rect 0 202524 168 202580
rect 0 202496 112 202524
rect 0 201684 112 201712
rect 0 201628 168 201684
rect 0 201600 112 201628
rect 0 200788 112 200816
rect 0 200732 168 200788
rect 0 200704 112 200732
rect 0 199892 112 199920
rect 0 199836 168 199892
rect 0 199808 112 199836
rect 0 198996 112 199024
rect 0 198940 168 198996
rect 0 198912 112 198940
rect 0 198100 112 198128
rect 0 198044 168 198100
rect 0 198016 112 198044
rect 0 197204 112 197232
rect 0 197148 168 197204
rect 0 197120 112 197148
rect 0 196308 112 196336
rect 0 196252 168 196308
rect 0 196224 112 196252
rect 0 195412 112 195440
rect 0 195356 168 195412
rect 0 195328 112 195356
rect 0 194516 112 194544
rect 0 194460 168 194516
rect 0 194432 112 194460
rect 0 193620 112 193648
rect 0 193564 168 193620
rect 0 193536 112 193564
rect 0 192724 112 192752
rect 0 192668 168 192724
rect 0 192640 112 192668
rect 0 191828 112 191856
rect 0 191772 168 191828
rect 0 191744 112 191772
rect 0 190932 112 190960
rect 0 190876 168 190932
rect 0 190848 112 190876
rect 0 190036 112 190064
rect 0 189980 168 190036
rect 0 189952 112 189980
rect 0 185444 112 185472
rect 0 185388 168 185444
rect 0 185360 112 185388
rect 0 184548 112 184576
rect 0 184492 168 184548
rect 0 184464 112 184492
rect 0 183652 112 183680
rect 0 183596 168 183652
rect 0 183568 112 183596
rect 0 182756 112 182784
rect 0 182700 168 182756
rect 0 182672 112 182700
rect 0 181860 112 181888
rect 0 181804 168 181860
rect 0 181776 112 181804
rect 0 180964 112 180992
rect 0 180908 168 180964
rect 0 180880 112 180908
rect 0 180068 112 180096
rect 0 180012 168 180068
rect 0 179984 112 180012
rect 0 179172 112 179200
rect 0 179116 168 179172
rect 0 179088 112 179116
rect 0 178276 112 178304
rect 0 178220 168 178276
rect 0 178192 112 178220
rect 0 177380 112 177408
rect 0 177324 168 177380
rect 0 177296 112 177324
rect 0 176484 112 176512
rect 0 176428 168 176484
rect 0 176400 112 176428
rect 0 175588 112 175616
rect 0 175532 168 175588
rect 0 175504 112 175532
rect 0 174692 112 174720
rect 0 174636 168 174692
rect 0 174608 112 174636
rect 0 173796 112 173824
rect 0 173740 168 173796
rect 0 173712 112 173740
rect 0 172900 112 172928
rect 0 172844 168 172900
rect 0 172816 112 172844
rect 0 172004 112 172032
rect 0 171948 168 172004
rect 0 171920 112 171948
rect 0 171108 112 171136
rect 0 171052 168 171108
rect 0 171024 112 171052
rect 0 170212 112 170240
rect 0 170156 168 170212
rect 0 170128 112 170156
rect 0 169316 112 169344
rect 0 169260 168 169316
rect 0 169232 112 169260
rect 0 168420 112 168448
rect 0 168364 168 168420
rect 0 168336 112 168364
rect 0 167524 112 167552
rect 0 167468 168 167524
rect 0 167440 112 167468
rect 0 166628 112 166656
rect 0 166572 168 166628
rect 0 166544 112 166572
rect 0 165732 112 165760
rect 0 165676 168 165732
rect 0 165648 112 165676
rect 464800 165508 464912 165536
rect 464772 165452 464912 165508
rect 464800 165424 464912 165452
rect 0 164836 112 164864
rect 0 164780 168 164836
rect 0 164752 112 164780
rect 464800 164612 464912 164640
rect 464772 164556 464912 164612
rect 464800 164528 464912 164556
rect 0 163940 112 163968
rect 0 163884 168 163940
rect 0 163856 112 163884
rect 464800 163716 464912 163744
rect 464772 163660 464912 163716
rect 464800 163632 464912 163660
rect 0 163044 112 163072
rect 0 162988 168 163044
rect 0 162960 112 162988
rect 464800 162820 464912 162848
rect 464772 162764 464912 162820
rect 464800 162736 464912 162764
rect 0 162148 112 162176
rect 0 162092 168 162148
rect 0 162064 112 162092
rect 464800 161924 464912 161952
rect 464772 161868 464912 161924
rect 464800 161840 464912 161868
rect 0 161252 112 161280
rect 0 161196 168 161252
rect 0 161168 112 161196
rect 464800 161028 464912 161056
rect 464772 160972 464912 161028
rect 464800 160944 464912 160972
rect 0 160356 112 160384
rect 0 160300 168 160356
rect 0 160272 112 160300
rect 464800 160132 464912 160160
rect 464772 160076 464912 160132
rect 464800 160048 464912 160076
rect 0 159460 112 159488
rect 0 159404 168 159460
rect 0 159376 112 159404
rect 464800 159236 464912 159264
rect 464772 159180 464912 159236
rect 464800 159152 464912 159180
rect 0 158564 112 158592
rect 0 158508 168 158564
rect 0 158480 112 158508
rect 464800 158340 464912 158368
rect 464772 158284 464912 158340
rect 464800 158256 464912 158284
rect 0 157668 112 157696
rect 0 157612 168 157668
rect 0 157584 112 157612
rect 464800 157444 464912 157472
rect 464772 157388 464912 157444
rect 464800 157360 464912 157388
rect 0 156772 112 156800
rect 0 156716 168 156772
rect 0 156688 112 156716
rect 464800 156548 464912 156576
rect 464772 156492 464912 156548
rect 464800 156464 464912 156492
rect 0 155876 112 155904
rect 0 155820 168 155876
rect 0 155792 112 155820
rect 464800 155652 464912 155680
rect 464772 155596 464912 155652
rect 464800 155568 464912 155596
rect 0 154980 112 155008
rect 0 154924 168 154980
rect 0 154896 112 154924
rect 464800 154756 464912 154784
rect 464772 154700 464912 154756
rect 464800 154672 464912 154700
rect 0 154084 112 154112
rect 0 154028 168 154084
rect 0 154000 112 154028
rect 464800 153860 464912 153888
rect 464772 153804 464912 153860
rect 464800 153776 464912 153804
rect 0 153188 112 153216
rect 0 153132 168 153188
rect 0 153104 112 153132
rect 464800 152964 464912 152992
rect 464772 152908 464912 152964
rect 464800 152880 464912 152908
rect 0 152292 112 152320
rect 0 152236 168 152292
rect 0 152208 112 152236
rect 464800 152068 464912 152096
rect 464772 152012 464912 152068
rect 464800 151984 464912 152012
rect 0 151396 112 151424
rect 0 151340 168 151396
rect 0 151312 112 151340
rect 464800 151172 464912 151200
rect 464772 151116 464912 151172
rect 464800 151088 464912 151116
rect 0 150500 112 150528
rect 0 150444 168 150500
rect 0 150416 112 150444
rect 464800 150276 464912 150304
rect 464772 150220 464912 150276
rect 464800 150192 464912 150220
rect 0 149604 112 149632
rect 0 149548 168 149604
rect 0 149520 112 149548
rect 464800 149380 464912 149408
rect 464772 149324 464912 149380
rect 464800 149296 464912 149324
rect 0 148708 112 148736
rect 0 148652 168 148708
rect 0 148624 112 148652
rect 464800 148484 464912 148512
rect 464772 148428 464912 148484
rect 464800 148400 464912 148428
rect 0 147812 112 147840
rect 0 147756 168 147812
rect 0 147728 112 147756
rect 464800 147588 464912 147616
rect 464772 147532 464912 147588
rect 464800 147504 464912 147532
rect 0 146916 112 146944
rect 0 146860 168 146916
rect 0 146832 112 146860
rect 464800 146692 464912 146720
rect 464772 146636 464912 146692
rect 464800 146608 464912 146636
rect 0 146020 112 146048
rect 0 145964 168 146020
rect 0 145936 112 145964
rect 464800 145796 464912 145824
rect 464772 145740 464912 145796
rect 464800 145712 464912 145740
rect 0 145124 112 145152
rect 0 145068 168 145124
rect 0 145040 112 145068
rect 464800 144900 464912 144928
rect 464772 144844 464912 144900
rect 464800 144816 464912 144844
rect 0 144228 112 144256
rect 0 144172 168 144228
rect 0 144144 112 144172
rect 464800 144004 464912 144032
rect 464772 143948 464912 144004
rect 464800 143920 464912 143948
rect 0 143332 112 143360
rect 0 143276 168 143332
rect 0 143248 112 143276
rect 464800 143108 464912 143136
rect 464772 143052 464912 143108
rect 464800 143024 464912 143052
rect 0 142436 112 142464
rect 0 142380 168 142436
rect 0 142352 112 142380
rect 464800 142212 464912 142240
rect 464772 142156 464912 142212
rect 464800 142128 464912 142156
rect 0 141540 112 141568
rect 0 141484 168 141540
rect 0 141456 112 141484
rect 464800 141316 464912 141344
rect 464772 141260 464912 141316
rect 464800 141232 464912 141260
rect 0 140644 112 140672
rect 0 140588 168 140644
rect 0 140560 112 140588
rect 464800 140420 464912 140448
rect 464772 140364 464912 140420
rect 464800 140336 464912 140364
rect 0 139748 112 139776
rect 0 139692 168 139748
rect 0 139664 112 139692
rect 464800 139524 464912 139552
rect 464772 139468 464912 139524
rect 464800 139440 464912 139468
rect 0 138852 112 138880
rect 0 138796 168 138852
rect 0 138768 112 138796
rect 464800 138628 464912 138656
rect 464772 138572 464912 138628
rect 464800 138544 464912 138572
rect 0 137956 112 137984
rect 0 137900 168 137956
rect 0 137872 112 137900
rect 464800 137732 464912 137760
rect 464772 137676 464912 137732
rect 464800 137648 464912 137676
rect 0 137060 112 137088
rect 0 137004 168 137060
rect 0 136976 112 137004
rect 464800 136836 464912 136864
rect 464772 136780 464912 136836
rect 464800 136752 464912 136780
rect 0 136164 112 136192
rect 0 136108 168 136164
rect 0 136080 112 136108
rect 464800 135940 464912 135968
rect 464772 135884 464912 135940
rect 464800 135856 464912 135884
rect 0 135268 112 135296
rect 0 135212 168 135268
rect 0 135184 112 135212
rect 464800 135044 464912 135072
rect 464772 134988 464912 135044
rect 464800 134960 464912 134988
rect 0 134372 112 134400
rect 0 134316 168 134372
rect 0 134288 112 134316
rect 464800 134148 464912 134176
rect 464772 134092 464912 134148
rect 464800 134064 464912 134092
rect 0 133476 112 133504
rect 0 133420 168 133476
rect 0 133392 112 133420
rect 464800 133252 464912 133280
rect 464772 133196 464912 133252
rect 464800 133168 464912 133196
rect 0 132580 112 132608
rect 0 132524 168 132580
rect 0 132496 112 132524
rect 0 127988 112 128016
rect 0 127932 168 127988
rect 0 127904 112 127932
rect 0 127092 112 127120
rect 0 127036 168 127092
rect 0 127008 112 127036
rect 0 126196 112 126224
rect 0 126140 168 126196
rect 0 126112 112 126140
rect 0 125300 112 125328
rect 0 125244 168 125300
rect 0 125216 112 125244
rect 0 124404 112 124432
rect 0 124348 168 124404
rect 0 124320 112 124348
rect 0 123508 112 123536
rect 0 123452 168 123508
rect 0 123424 112 123452
rect 0 122612 112 122640
rect 0 122556 168 122612
rect 0 122528 112 122556
rect 0 121716 112 121744
rect 0 121660 168 121716
rect 0 121632 112 121660
rect 0 120820 112 120848
rect 0 120764 168 120820
rect 0 120736 112 120764
rect 0 119924 112 119952
rect 0 119868 168 119924
rect 0 119840 112 119868
rect 0 119028 112 119056
rect 0 118972 168 119028
rect 0 118944 112 118972
rect 0 118132 112 118160
rect 0 118076 168 118132
rect 0 118048 112 118076
rect 0 117236 112 117264
rect 0 117180 168 117236
rect 0 117152 112 117180
rect 0 116340 112 116368
rect 0 116284 168 116340
rect 0 116256 112 116284
rect 0 115444 112 115472
rect 0 115388 168 115444
rect 0 115360 112 115388
rect 0 114548 112 114576
rect 0 114492 168 114548
rect 0 114464 112 114492
rect 0 113652 112 113680
rect 0 113596 168 113652
rect 0 113568 112 113596
rect 0 112756 112 112784
rect 0 112700 168 112756
rect 0 112672 112 112700
rect 0 111860 112 111888
rect 0 111804 168 111860
rect 0 111776 112 111804
rect 0 110964 112 110992
rect 0 110908 168 110964
rect 0 110880 112 110908
rect 0 110068 112 110096
rect 0 110012 168 110068
rect 0 109984 112 110012
rect 0 109172 112 109200
rect 0 109116 168 109172
rect 0 109088 112 109116
rect 0 108276 112 108304
rect 0 108220 168 108276
rect 0 108192 112 108220
rect 0 107380 112 107408
rect 0 107324 168 107380
rect 0 107296 112 107324
rect 0 106484 112 106512
rect 0 106428 168 106484
rect 0 106400 112 106428
rect 0 105588 112 105616
rect 0 105532 168 105588
rect 0 105504 112 105532
rect 0 104692 112 104720
rect 0 104636 168 104692
rect 0 104608 112 104636
rect 0 103796 112 103824
rect 0 103740 168 103796
rect 0 103712 112 103740
rect 0 102900 112 102928
rect 0 102844 168 102900
rect 0 102816 112 102844
rect 0 102004 112 102032
rect 0 101948 168 102004
rect 0 101920 112 101948
rect 0 101108 112 101136
rect 0 101052 168 101108
rect 0 101024 112 101052
rect 0 100212 112 100240
rect 0 100156 168 100212
rect 0 100128 112 100156
rect 0 99316 112 99344
rect 0 99260 168 99316
rect 0 99232 112 99260
rect 0 98420 112 98448
rect 0 98364 168 98420
rect 0 98336 112 98364
rect 0 97524 112 97552
rect 0 97468 168 97524
rect 0 97440 112 97468
rect 0 96628 112 96656
rect 0 96572 168 96628
rect 0 96544 112 96572
rect 0 95732 112 95760
rect 0 95676 168 95732
rect 0 95648 112 95676
rect 0 94836 112 94864
rect 0 94780 168 94836
rect 0 94752 112 94780
rect 0 93940 112 93968
rect 0 93884 168 93940
rect 0 93856 112 93884
rect 0 93044 112 93072
rect 0 92988 168 93044
rect 0 92960 112 92988
rect 0 92148 112 92176
rect 0 92092 168 92148
rect 0 92064 112 92092
rect 0 91252 112 91280
rect 0 91196 168 91252
rect 0 91168 112 91196
rect 0 90356 112 90384
rect 0 90300 168 90356
rect 0 90272 112 90300
rect 0 89460 112 89488
rect 0 89404 168 89460
rect 0 89376 112 89404
rect 0 88564 112 88592
rect 0 88508 168 88564
rect 0 88480 112 88508
rect 0 87668 112 87696
rect 0 87612 168 87668
rect 0 87584 112 87612
rect 0 86772 112 86800
rect 0 86716 168 86772
rect 0 86688 112 86716
rect 0 85876 112 85904
rect 0 85820 168 85876
rect 0 85792 112 85820
rect 0 84980 112 85008
rect 0 84924 168 84980
rect 0 84896 112 84924
rect 0 84084 112 84112
rect 0 84028 168 84084
rect 0 84000 112 84028
rect 0 83188 112 83216
rect 0 83132 168 83188
rect 0 83104 112 83132
rect 0 82292 112 82320
rect 0 82236 168 82292
rect 0 82208 112 82236
rect 0 81396 112 81424
rect 0 81340 168 81396
rect 0 81312 112 81340
rect 0 80500 112 80528
rect 0 80444 168 80500
rect 0 80416 112 80444
rect 0 79604 112 79632
rect 0 79548 168 79604
rect 0 79520 112 79548
rect 0 78708 112 78736
rect 0 78652 168 78708
rect 0 78624 112 78652
rect 0 77812 112 77840
rect 0 77756 168 77812
rect 0 77728 112 77756
rect 0 76916 112 76944
rect 0 76860 168 76916
rect 0 76832 112 76860
rect 0 76020 112 76048
rect 0 75964 168 76020
rect 0 75936 112 75964
rect 0 75124 112 75152
rect 0 75068 168 75124
rect 0 75040 112 75068
rect 0 70532 112 70560
rect 0 70476 168 70532
rect 0 70448 112 70476
rect 0 69636 112 69664
rect 0 69580 168 69636
rect 0 69552 112 69580
rect 0 68740 112 68768
rect 0 68684 168 68740
rect 0 68656 112 68684
rect 0 67844 112 67872
rect 0 67788 168 67844
rect 0 67760 112 67788
rect 0 66948 112 66976
rect 0 66892 168 66948
rect 0 66864 112 66892
rect 0 66052 112 66080
rect 0 65996 168 66052
rect 0 65968 112 65996
rect 0 65156 112 65184
rect 0 65100 168 65156
rect 0 65072 112 65100
rect 0 64260 112 64288
rect 0 64204 168 64260
rect 0 64176 112 64204
rect 0 63364 112 63392
rect 0 63308 168 63364
rect 0 63280 112 63308
rect 0 62468 112 62496
rect 0 62412 168 62468
rect 0 62384 112 62412
rect 0 61572 112 61600
rect 0 61516 168 61572
rect 0 61488 112 61516
rect 0 60676 112 60704
rect 0 60620 168 60676
rect 0 60592 112 60620
rect 0 59780 112 59808
rect 0 59724 168 59780
rect 0 59696 112 59724
rect 0 58884 112 58912
rect 0 58828 168 58884
rect 0 58800 112 58828
rect 0 57988 112 58016
rect 0 57932 168 57988
rect 0 57904 112 57932
rect 0 57092 112 57120
rect 0 57036 168 57092
rect 0 57008 112 57036
rect 0 56196 112 56224
rect 0 56140 168 56196
rect 0 56112 112 56140
rect 0 55300 112 55328
rect 0 55244 168 55300
rect 0 55216 112 55244
rect 0 54404 112 54432
rect 0 54348 168 54404
rect 0 54320 112 54348
rect 0 53508 112 53536
rect 0 53452 168 53508
rect 0 53424 112 53452
rect 0 52612 112 52640
rect 0 52556 168 52612
rect 0 52528 112 52556
rect 0 51716 112 51744
rect 0 51660 168 51716
rect 0 51632 112 51660
rect 0 50820 112 50848
rect 0 50764 168 50820
rect 0 50736 112 50764
rect 464800 50596 464912 50624
rect 464772 50540 464912 50596
rect 464800 50512 464912 50540
rect 0 49924 112 49952
rect 0 49868 168 49924
rect 0 49840 112 49868
rect 464800 49700 464912 49728
rect 464772 49644 464912 49700
rect 464800 49616 464912 49644
rect 0 49028 112 49056
rect 0 48972 168 49028
rect 0 48944 112 48972
rect 464800 48804 464912 48832
rect 464772 48748 464912 48804
rect 464800 48720 464912 48748
rect 0 48132 112 48160
rect 0 48076 168 48132
rect 0 48048 112 48076
rect 464800 47908 464912 47936
rect 464772 47852 464912 47908
rect 464800 47824 464912 47852
rect 0 47236 112 47264
rect 0 47180 168 47236
rect 0 47152 112 47180
rect 464800 47012 464912 47040
rect 464772 46956 464912 47012
rect 464800 46928 464912 46956
rect 0 46340 112 46368
rect 0 46284 168 46340
rect 0 46256 112 46284
rect 464800 46116 464912 46144
rect 464772 46060 464912 46116
rect 464800 46032 464912 46060
rect 0 45444 112 45472
rect 0 45388 168 45444
rect 0 45360 112 45388
rect 464800 45220 464912 45248
rect 464772 45164 464912 45220
rect 464800 45136 464912 45164
rect 0 44548 112 44576
rect 0 44492 168 44548
rect 0 44464 112 44492
rect 464800 44324 464912 44352
rect 464772 44268 464912 44324
rect 464800 44240 464912 44268
rect 0 43652 112 43680
rect 0 43596 168 43652
rect 0 43568 112 43596
rect 464800 43428 464912 43456
rect 464772 43372 464912 43428
rect 464800 43344 464912 43372
rect 0 42756 112 42784
rect 0 42700 168 42756
rect 0 42672 112 42700
rect 464800 42532 464912 42560
rect 464772 42476 464912 42532
rect 464800 42448 464912 42476
rect 0 41860 112 41888
rect 0 41804 168 41860
rect 0 41776 112 41804
rect 464800 41636 464912 41664
rect 464772 41580 464912 41636
rect 464800 41552 464912 41580
rect 0 40964 112 40992
rect 0 40908 168 40964
rect 0 40880 112 40908
rect 464800 40740 464912 40768
rect 464772 40684 464912 40740
rect 464800 40656 464912 40684
rect 0 40068 112 40096
rect 0 40012 168 40068
rect 0 39984 112 40012
rect 464800 39844 464912 39872
rect 464772 39788 464912 39844
rect 464800 39760 464912 39788
rect 0 39172 112 39200
rect 0 39116 168 39172
rect 0 39088 112 39116
rect 464800 38948 464912 38976
rect 464772 38892 464912 38948
rect 464800 38864 464912 38892
rect 0 38276 112 38304
rect 0 38220 168 38276
rect 0 38192 112 38220
rect 464800 38052 464912 38080
rect 464772 37996 464912 38052
rect 464800 37968 464912 37996
rect 0 37380 112 37408
rect 0 37324 168 37380
rect 0 37296 112 37324
rect 464800 37156 464912 37184
rect 464772 37100 464912 37156
rect 464800 37072 464912 37100
rect 0 36484 112 36512
rect 0 36428 168 36484
rect 0 36400 112 36428
rect 464800 36260 464912 36288
rect 464772 36204 464912 36260
rect 464800 36176 464912 36204
rect 0 35588 112 35616
rect 0 35532 168 35588
rect 0 35504 112 35532
rect 464800 35364 464912 35392
rect 464772 35308 464912 35364
rect 464800 35280 464912 35308
rect 0 34692 112 34720
rect 0 34636 168 34692
rect 0 34608 112 34636
rect 464800 34468 464912 34496
rect 464772 34412 464912 34468
rect 464800 34384 464912 34412
rect 0 33796 112 33824
rect 0 33740 168 33796
rect 0 33712 112 33740
rect 464800 33572 464912 33600
rect 464772 33516 464912 33572
rect 464800 33488 464912 33516
rect 0 32900 112 32928
rect 0 32844 168 32900
rect 0 32816 112 32844
rect 464800 32676 464912 32704
rect 464772 32620 464912 32676
rect 464800 32592 464912 32620
rect 0 32004 112 32032
rect 0 31948 168 32004
rect 0 31920 112 31948
rect 464800 31780 464912 31808
rect 464772 31724 464912 31780
rect 464800 31696 464912 31724
rect 0 31108 112 31136
rect 0 31052 168 31108
rect 0 31024 112 31052
rect 464800 30884 464912 30912
rect 464772 30828 464912 30884
rect 464800 30800 464912 30828
rect 0 30212 112 30240
rect 0 30156 168 30212
rect 0 30128 112 30156
rect 464800 29988 464912 30016
rect 464772 29932 464912 29988
rect 464800 29904 464912 29932
rect 0 29316 112 29344
rect 0 29260 168 29316
rect 0 29232 112 29260
rect 464800 29092 464912 29120
rect 464772 29036 464912 29092
rect 464800 29008 464912 29036
rect 0 28420 112 28448
rect 0 28364 168 28420
rect 0 28336 112 28364
rect 464800 28196 464912 28224
rect 464772 28140 464912 28196
rect 464800 28112 464912 28140
rect 0 27524 112 27552
rect 0 27468 168 27524
rect 0 27440 112 27468
rect 464800 27300 464912 27328
rect 464772 27244 464912 27300
rect 464800 27216 464912 27244
rect 0 26628 112 26656
rect 0 26572 168 26628
rect 0 26544 112 26572
rect 464800 26404 464912 26432
rect 464772 26348 464912 26404
rect 464800 26320 464912 26348
rect 0 25732 112 25760
rect 0 25676 168 25732
rect 0 25648 112 25676
rect 464800 25508 464912 25536
rect 464772 25452 464912 25508
rect 464800 25424 464912 25452
rect 0 24836 112 24864
rect 0 24780 168 24836
rect 0 24752 112 24780
rect 464800 24612 464912 24640
rect 464772 24556 464912 24612
rect 464800 24528 464912 24556
rect 0 23940 112 23968
rect 0 23884 168 23940
rect 0 23856 112 23884
rect 464800 23716 464912 23744
rect 464772 23660 464912 23716
rect 464800 23632 464912 23660
rect 0 23044 112 23072
rect 0 22988 168 23044
rect 0 22960 112 22988
rect 464800 22820 464912 22848
rect 464772 22764 464912 22820
rect 464800 22736 464912 22764
rect 0 22148 112 22176
rect 0 22092 168 22148
rect 0 22064 112 22092
rect 464800 21924 464912 21952
rect 464772 21868 464912 21924
rect 464800 21840 464912 21868
rect 0 21252 112 21280
rect 0 21196 168 21252
rect 0 21168 112 21196
rect 464800 21028 464912 21056
rect 464772 20972 464912 21028
rect 464800 20944 464912 20972
rect 0 20356 112 20384
rect 0 20300 168 20356
rect 0 20272 112 20300
rect 464800 20132 464912 20160
rect 464772 20076 464912 20132
rect 464800 20048 464912 20076
rect 0 19460 112 19488
rect 0 19404 168 19460
rect 0 19376 112 19404
rect 464800 19236 464912 19264
rect 464772 19180 464912 19236
rect 464800 19152 464912 19180
rect 0 18564 112 18592
rect 0 18508 168 18564
rect 0 18480 112 18508
rect 464800 18340 464912 18368
rect 464772 18284 464912 18340
rect 464800 18256 464912 18284
rect 0 17668 112 17696
rect 0 17612 168 17668
rect 0 17584 112 17612
rect 0 15092 112 15120
rect 0 15036 28728 15092
rect 0 15008 112 15036
rect 0 14644 112 14672
rect 0 14588 28728 14644
rect 0 14560 112 14588
rect 0 14196 112 14224
rect 0 14140 28728 14196
rect 0 14112 112 14140
rect 0 13748 112 13776
rect 0 13692 28728 13748
rect 0 13664 112 13692
rect 0 13300 112 13328
rect 0 13244 28728 13300
rect 0 13216 112 13244
rect 0 12852 112 12880
rect 0 12796 28728 12852
rect 0 12768 112 12796
rect 0 12404 112 12432
rect 0 12348 28728 12404
rect 0 12320 112 12348
rect 0 11956 112 11984
rect 0 11900 28728 11956
rect 0 11872 112 11900
rect 0 11508 112 11536
rect 0 11452 28728 11508
rect 0 11424 112 11452
rect 0 11060 112 11088
rect 0 11004 28728 11060
rect 0 10976 112 11004
rect 0 10612 112 10640
rect 0 10556 28728 10612
rect 0 10528 112 10556
rect 0 10164 112 10192
rect 0 10108 28728 10164
rect 0 10080 112 10108
rect 0 9716 112 9744
rect 0 9660 28728 9716
rect 0 9632 112 9660
rect 0 9268 112 9296
rect 0 9212 28728 9268
rect 0 9184 112 9212
rect 0 8820 112 8848
rect 0 8764 28728 8820
rect 0 8736 112 8764
rect 0 8372 112 8400
rect 0 8316 28728 8372
rect 0 8288 112 8316
rect 0 7924 112 7952
rect 0 7868 28728 7924
rect 0 7840 112 7868
rect 0 7476 112 7504
rect 0 7420 28728 7476
rect 0 7392 112 7420
rect 0 7028 112 7056
rect 0 6972 28728 7028
rect 0 6944 112 6972
rect 0 6580 112 6608
rect 0 6524 28728 6580
rect 0 6496 112 6524
rect 0 6132 112 6160
rect 0 6076 28728 6132
rect 0 6048 112 6076
rect 0 5684 112 5712
rect 0 5628 28728 5684
rect 0 5600 112 5628
rect 0 5236 112 5264
rect 0 5180 28728 5236
rect 0 5152 112 5180
rect 0 4788 112 4816
rect 0 4732 28728 4788
rect 0 4704 112 4732
rect 0 4340 112 4368
rect 0 4284 28728 4340
rect 0 4256 112 4284
rect 0 3892 112 3920
rect 0 3836 28728 3892
rect 0 3808 112 3836
rect 0 3444 112 3472
rect 0 3388 28728 3444
rect 0 3360 112 3388
rect 0 2996 112 3024
rect 0 2940 28728 2996
rect 0 2912 112 2940
rect 0 2548 112 2576
rect 0 2492 28728 2548
rect 0 2464 112 2492
rect 0 2100 112 2128
rect 0 2044 28728 2100
rect 0 2016 112 2044
rect 0 1652 112 1680
rect 0 1596 20188 1652
rect 0 1568 112 1596
rect 0 1204 112 1232
rect 0 1148 8428 1204
rect 0 1120 112 1148
rect 8372 868 8428 1148
rect 20132 980 20188 1596
rect 28028 1540 28728 1596
rect 28028 980 28084 1540
rect 20132 924 28084 980
rect 28700 868 28756 1120
rect 44174 924 44184 980
rect 44240 924 87920 980
rect 87976 924 145376 980
rect 145432 924 203952 980
rect 204008 924 267288 980
rect 267344 924 324464 980
rect 324520 924 377496 980
rect 377552 924 435344 980
rect 435400 924 435410 980
rect 8372 812 28756 868
rect 802 140 812 196
rect 868 140 8428 196
rect 447458 140 447468 196
rect 447524 140 448252 196
rect 448308 140 448318 196
rect 8372 84 8428 140
rect 8372 28 44156 84
rect 44212 28 44222 84
<< via3 >>
rect 28140 719068 28196 719124
rect 28140 717444 28196 717500
<< metal4 >>
rect 28140 719124 28196 719134
rect 28140 717500 28196 719068
rect 28140 717434 28196 717444
rect 3888 15344 4208 704816
rect 4548 15344 4868 704816
rect 23888 15344 24208 704816
rect 24548 15344 24868 704816
rect 32448 1120 32768 719040
rect 33108 1120 33428 719040
rect 52448 1120 52768 719040
rect 53108 1120 53428 719040
rect 72448 1120 72768 719040
rect 73108 1120 73428 719040
rect 89904 1120 90224 719040
rect 90564 1120 90884 719040
rect 109904 1120 110224 719040
rect 110564 1120 110884 719040
rect 129904 1120 130224 719040
rect 130564 1120 130884 719040
rect 147360 1120 147680 719040
rect 148020 1120 148340 719040
rect 167360 1120 167680 719040
rect 168020 1120 168340 719040
rect 187360 1120 187680 719040
rect 188020 1120 188340 719040
rect 204816 1120 205136 719040
rect 205476 1120 205796 719040
rect 224816 1120 225136 719040
rect 225476 1120 225796 719040
rect 244816 1120 245136 719040
rect 245476 1120 245796 719040
rect 269216 1120 269536 719040
rect 269876 1120 270196 719040
rect 289216 1120 289536 719040
rect 289876 1120 290196 719040
rect 309216 1120 309536 719040
rect 309876 1120 310196 719040
rect 326672 1120 326992 719040
rect 327332 1120 327652 719040
rect 346672 1120 346992 719040
rect 347332 1120 347652 719040
rect 366672 1120 366992 719040
rect 367332 1120 367652 719040
rect 379424 1120 379744 719040
rect 380084 1120 380404 719040
rect 399424 1120 399744 719040
rect 400084 1120 400404 719040
rect 419424 1120 419744 719040
rect 420084 1120 420404 719040
rect 436880 1120 437200 719040
rect 437540 1120 437860 719040
rect 456880 1120 457200 719040
rect 457540 1120 457860 719040
use W_IO4  Tile_X0Y1_W_IO4
timestamp 0
transform 1 0 112 0 1 647360
box 0 0 1 1
use W_IO4  Tile_X0Y2_W_IO4
timestamp 0
transform 1 0 112 0 1 589904
box 0 0 1 1
use W_IO4  Tile_X0Y3_W_IO4
timestamp 0
transform 1 0 112 0 1 532448
box 0 0 1 1
use W_IO4  Tile_X0Y4_W_IO4
timestamp 0
transform 1 0 112 0 1 474992
box 0 0 1 1
use W_IO4  Tile_X0Y5_W_IO4
timestamp 0
transform 1 0 112 0 1 417536
box 0 0 1 1
use W_IO4  Tile_X0Y6_W_IO4
timestamp 0
transform 1 0 112 0 1 360080
box 0 0 1 1
use W_IO4  Tile_X0Y7_W_IO4
timestamp 0
transform 1 0 112 0 1 302624
box 0 0 1 1
use W_IO4  Tile_X0Y8_W_IO4
timestamp 0
transform 1 0 112 0 1 245168
box 0 0 1 1
use W_IO4  Tile_X0Y9_W_IO4
timestamp 0
transform 1 0 112 0 1 187712
box 0 0 1 1
use W_IO4  Tile_X0Y10_W_IO4
timestamp 0
transform 1 0 112 0 1 130256
box 0 0 1 1
use W_IO4  Tile_X0Y11_W_IO4
timestamp 0
transform 1 0 112 0 1 72800
box 0 0 1 1
use W_IO4  Tile_X0Y12_W_IO4
timestamp 0
transform 1 0 112 0 1 15344
box 0 0 1 1
use N_term_single  Tile_X1Y0_N_term_single
timestamp 0
transform 1 0 28672 0 1 704816
box 0 0 1 1
use LUT4AB  Tile_X1Y1_LUT4AB
timestamp 0
transform 1 0 28672 0 1 647360
box 0 0 1 1
use LUT4AB  Tile_X1Y2_LUT4AB
timestamp 0
transform 1 0 28672 0 1 589904
box 0 0 1 1
use LUT4AB  Tile_X1Y3_LUT4AB
timestamp 0
transform 1 0 28672 0 1 532448
box 0 0 1 1
use LUT4AB  Tile_X1Y4_LUT4AB
timestamp 0
transform 1 0 28672 0 1 474992
box 0 0 1 1
use LUT4AB  Tile_X1Y5_LUT4AB
timestamp 0
transform 1 0 28672 0 1 417536
box 0 0 1 1
use LUT4AB  Tile_X1Y6_LUT4AB
timestamp 0
transform 1 0 28672 0 1 360080
box 0 0 1 1
use LUT4AB  Tile_X1Y7_LUT4AB
timestamp 0
transform 1 0 28672 0 1 302624
box 0 0 1 1
use LUT4AB  Tile_X1Y8_LUT4AB
timestamp 0
transform 1 0 28672 0 1 245168
box 0 0 1 1
use LUT4AB  Tile_X1Y9_LUT4AB
timestamp 0
transform 1 0 28672 0 1 187712
box 0 0 1 1
use LUT4AB  Tile_X1Y10_LUT4AB
timestamp 0
transform 1 0 28672 0 1 130256
box 0 0 1 1
use LUT4AB  Tile_X1Y11_LUT4AB
timestamp 0
transform 1 0 28672 0 1 72800
box 0 0 1 1
use LUT4AB  Tile_X1Y12_LUT4AB
timestamp 0
transform 1 0 28672 0 1 15344
box 0 0 1 1
use S_WARMBOOT  Tile_X1Y13_S_WARMBOOT
timestamp 0
transform 1 0 28672 0 1 1120
box 0 0 1 1
use N_term_single  Tile_X2Y0_N_term_single
timestamp 0
transform 1 0 86128 0 1 704816
box 0 0 1 1
use LUT4AB  Tile_X2Y1_LUT4AB
timestamp 0
transform 1 0 86128 0 1 647360
box 0 0 1 1
use LUT4AB  Tile_X2Y2_LUT4AB
timestamp 0
transform 1 0 86128 0 1 589904
box 0 0 1 1
use LUT4AB  Tile_X2Y3_LUT4AB
timestamp 0
transform 1 0 86128 0 1 532448
box 0 0 1 1
use LUT4AB  Tile_X2Y4_LUT4AB
timestamp 0
transform 1 0 86128 0 1 474992
box 0 0 1 1
use LUT4AB  Tile_X2Y5_LUT4AB
timestamp 0
transform 1 0 86128 0 1 417536
box 0 0 1 1
use LUT4AB  Tile_X2Y6_LUT4AB
timestamp 0
transform 1 0 86128 0 1 360080
box 0 0 1 1
use LUT4AB  Tile_X2Y7_LUT4AB
timestamp 0
transform 1 0 86128 0 1 302624
box 0 0 1 1
use LUT4AB  Tile_X2Y8_LUT4AB
timestamp 0
transform 1 0 86128 0 1 245168
box 0 0 1 1
use LUT4AB  Tile_X2Y9_LUT4AB
timestamp 0
transform 1 0 86128 0 1 187712
box 0 0 1 1
use LUT4AB  Tile_X2Y10_LUT4AB
timestamp 0
transform 1 0 86128 0 1 130256
box 0 0 1 1
use LUT4AB  Tile_X2Y11_LUT4AB
timestamp 0
transform 1 0 86128 0 1 72800
box 0 0 1 1
use LUT4AB  Tile_X2Y12_LUT4AB
timestamp 0
transform 1 0 86128 0 1 15344
box 0 0 1 1
use S_term_single  Tile_X2Y13_S_term_single
timestamp 0
transform 1 0 86128 0 1 1120
box 0 0 1 1
use N_term_single  Tile_X3Y0_N_term_single
timestamp 0
transform 1 0 143584 0 1 704816
box 0 0 1 1
use LUT4AB  Tile_X3Y1_LUT4AB
timestamp 0
transform 1 0 143584 0 1 647360
box 0 0 1 1
use LUT4AB  Tile_X3Y2_LUT4AB
timestamp 0
transform 1 0 143584 0 1 589904
box 0 0 1 1
use LUT4AB  Tile_X3Y3_LUT4AB
timestamp 0
transform 1 0 143584 0 1 532448
box 0 0 1 1
use LUT4AB  Tile_X3Y4_LUT4AB
timestamp 0
transform 1 0 143584 0 1 474992
box 0 0 1 1
use LUT4AB  Tile_X3Y5_LUT4AB
timestamp 0
transform 1 0 143584 0 1 417536
box 0 0 1 1
use LUT4AB  Tile_X3Y6_LUT4AB
timestamp 0
transform 1 0 143584 0 1 360080
box 0 0 1 1
use LUT4AB  Tile_X3Y7_LUT4AB
timestamp 0
transform 1 0 143584 0 1 302624
box 0 0 1 1
use LUT4AB  Tile_X3Y8_LUT4AB
timestamp 0
transform 1 0 143584 0 1 245168
box 0 0 1 1
use LUT4AB  Tile_X3Y9_LUT4AB
timestamp 0
transform 1 0 143584 0 1 187712
box 0 0 1 1
use LUT4AB  Tile_X3Y10_LUT4AB
timestamp 0
transform 1 0 143584 0 1 130256
box 0 0 1 1
use LUT4AB  Tile_X3Y11_LUT4AB
timestamp 0
transform 1 0 143584 0 1 72800
box 0 0 1 1
use LUT4AB  Tile_X3Y12_LUT4AB
timestamp 0
transform 1 0 143584 0 1 15344
box 0 0 1 1
use S_term_single  Tile_X3Y13_S_term_single
timestamp 0
transform 1 0 143584 0 1 1120
box 0 0 1 1
use N_term_single2  Tile_X4Y0_N_term_single2
timestamp 0
transform 1 0 201040 0 1 704816
box 0 0 1 1
use RegFile  Tile_X4Y1_RegFile
timestamp 0
transform 1 0 201040 0 1 647360
box 0 0 1 1
use RegFile  Tile_X4Y2_RegFile
timestamp 0
transform 1 0 201040 0 1 589904
box 0 0 1 1
use RegFile  Tile_X4Y3_RegFile
timestamp 0
transform 1 0 201040 0 1 532448
box 0 0 1 1
use RegFile  Tile_X4Y4_RegFile
timestamp 0
transform 1 0 201040 0 1 474992
box 0 0 1 1
use RegFile  Tile_X4Y5_RegFile
timestamp 0
transform 1 0 201040 0 1 417536
box 0 0 1 1
use RegFile  Tile_X4Y6_RegFile
timestamp 0
transform 1 0 201040 0 1 360080
box 0 0 1 1
use RegFile  Tile_X4Y7_RegFile
timestamp 0
transform 1 0 201040 0 1 302624
box 0 0 1 1
use RegFile  Tile_X4Y8_RegFile
timestamp 0
transform 1 0 201040 0 1 245168
box 0 0 1 1
use RegFile  Tile_X4Y9_RegFile
timestamp 0
transform 1 0 201040 0 1 187712
box 0 0 1 1
use RegFile  Tile_X4Y10_RegFile
timestamp 0
transform 1 0 201040 0 1 130256
box 0 0 1 1
use RegFile  Tile_X4Y11_RegFile
timestamp 0
transform 1 0 201040 0 1 72800
box 0 0 1 1
use RegFile  Tile_X4Y12_RegFile
timestamp 0
transform 1 0 201040 0 1 15344
box 0 0 1 1
use S_term_single2  Tile_X4Y13_S_term_single2
timestamp 0
transform 1 0 201040 0 1 1120
box 0 0 1 1
use N_term_single  Tile_X5Y0_N_term_single
timestamp 0
transform 1 0 265440 0 1 704816
box 0 0 1 1
use LUT4AB  Tile_X5Y1_LUT4AB
timestamp 0
transform 1 0 265440 0 1 647360
box 0 0 1 1
use LUT4AB  Tile_X5Y2_LUT4AB
timestamp 0
transform 1 0 265440 0 1 589904
box 0 0 1 1
use LUT4AB  Tile_X5Y3_LUT4AB
timestamp 0
transform 1 0 265440 0 1 532448
box 0 0 1 1
use LUT4AB  Tile_X5Y4_LUT4AB
timestamp 0
transform 1 0 265440 0 1 474992
box 0 0 1 1
use LUT4AB  Tile_X5Y5_LUT4AB
timestamp 0
transform 1 0 265440 0 1 417536
box 0 0 1 1
use LUT4AB  Tile_X5Y6_LUT4AB
timestamp 0
transform 1 0 265440 0 1 360080
box 0 0 1 1
use LUT4AB  Tile_X5Y7_LUT4AB
timestamp 0
transform 1 0 265440 0 1 302624
box 0 0 1 1
use LUT4AB  Tile_X5Y8_LUT4AB
timestamp 0
transform 1 0 265440 0 1 245168
box 0 0 1 1
use LUT4AB  Tile_X5Y9_LUT4AB
timestamp 0
transform 1 0 265440 0 1 187712
box 0 0 1 1
use LUT4AB  Tile_X5Y10_LUT4AB
timestamp 0
transform 1 0 265440 0 1 130256
box 0 0 1 1
use LUT4AB  Tile_X5Y11_LUT4AB
timestamp 0
transform 1 0 265440 0 1 72800
box 0 0 1 1
use LUT4AB  Tile_X5Y12_LUT4AB
timestamp 0
transform 1 0 265440 0 1 15344
box 0 0 1 1
use S_term_single  Tile_X5Y13_S_term_single
timestamp 0
transform 1 0 265440 0 1 1120
box 0 0 1 1
use N_term_DSP  Tile_X6Y0_N_term_DSP
timestamp 0
transform 1 0 322896 0 1 704816
box 0 0 1 1
use DSP  Tile_X6Y1_DSP
timestamp 0
transform 1 0 322896 0 1 589904
box 0 0 1 1
use DSP  Tile_X6Y3_DSP
timestamp 0
transform 1 0 322896 0 1 474992
box 0 0 1 1
use DSP  Tile_X6Y5_DSP
timestamp 0
transform 1 0 322896 0 1 360080
box 0 0 1 1
use DSP  Tile_X6Y7_DSP
timestamp 0
transform 1 0 322896 0 1 245168
box 0 0 1 1
use DSP  Tile_X6Y9_DSP
timestamp 0
transform 1 0 322896 0 1 130256
box 0 0 1 1
use DSP  Tile_X6Y11_DSP
timestamp 0
transform 1 0 322896 0 1 15344
box 0 0 1 1
use S_term_DSP  Tile_X6Y13_S_term_DSP
timestamp 0
transform 1 0 322896 0 1 1120
box 0 0 1 1
use N_term_single  Tile_X7Y0_N_term_single
timestamp 0
transform 1 0 375648 0 1 704816
box 0 0 1 1
use LUT4AB  Tile_X7Y1_LUT4AB
timestamp 0
transform 1 0 375648 0 1 647360
box 0 0 1 1
use LUT4AB  Tile_X7Y2_LUT4AB
timestamp 0
transform 1 0 375648 0 1 589904
box 0 0 1 1
use LUT4AB  Tile_X7Y3_LUT4AB
timestamp 0
transform 1 0 375648 0 1 532448
box 0 0 1 1
use LUT4AB  Tile_X7Y4_LUT4AB
timestamp 0
transform 1 0 375648 0 1 474992
box 0 0 1 1
use LUT4AB  Tile_X7Y5_LUT4AB
timestamp 0
transform 1 0 375648 0 1 417536
box 0 0 1 1
use LUT4AB  Tile_X7Y6_LUT4AB
timestamp 0
transform 1 0 375648 0 1 360080
box 0 0 1 1
use LUT4AB  Tile_X7Y7_LUT4AB
timestamp 0
transform 1 0 375648 0 1 302624
box 0 0 1 1
use LUT4AB  Tile_X7Y8_LUT4AB
timestamp 0
transform 1 0 375648 0 1 245168
box 0 0 1 1
use LUT4AB  Tile_X7Y9_LUT4AB
timestamp 0
transform 1 0 375648 0 1 187712
box 0 0 1 1
use LUT4AB  Tile_X7Y10_LUT4AB
timestamp 0
transform 1 0 375648 0 1 130256
box 0 0 1 1
use LUT4AB  Tile_X7Y11_LUT4AB
timestamp 0
transform 1 0 375648 0 1 72800
box 0 0 1 1
use LUT4AB  Tile_X7Y12_LUT4AB
timestamp 0
transform 1 0 375648 0 1 15344
box 0 0 1 1
use S_term_single  Tile_X7Y13_S_term_single
timestamp 0
transform 1 0 375648 0 1 1120
box 0 0 1 1
use N_term_SRAM  Tile_X8Y0_N_term_SRAM
timestamp 0
transform 1 0 433104 0 1 704816
box 0 0 1 1
use GF_SRAM  Tile_X8Y1_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 589904
box 0 0 1 1
use GF_SRAM  Tile_X8Y3_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 474992
box 0 0 1 1
use GF_SRAM  Tile_X8Y5_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 360080
box 0 0 1 1
use GF_SRAM  Tile_X8Y7_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 245168
box 0 0 1 1
use GF_SRAM  Tile_X8Y9_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 130256
box 0 0 1 1
use GF_SRAM  Tile_X8Y11_GF_SRAM
timestamp 0
transform 1 0 433104 0 1 15344
box 0 0 1 1
use S_term_SRAM  Tile_X8Y13_S_term_SRAM
timestamp 0
transform 1 0 433104 0 1 1120
box 0 0 1 1
<< labels >>
flabel metal3 s 0 704816 112 704928 0 FreeSans 448 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 563360 112 563472 0 FreeSans 448 0 0 0 FrameData[100]
port 1 nsew signal input
flabel metal3 s 0 564256 112 564368 0 FreeSans 448 0 0 0 FrameData[101]
port 2 nsew signal input
flabel metal3 s 0 565152 112 565264 0 FreeSans 448 0 0 0 FrameData[102]
port 3 nsew signal input
flabel metal3 s 0 566048 112 566160 0 FreeSans 448 0 0 0 FrameData[103]
port 4 nsew signal input
flabel metal3 s 0 566944 112 567056 0 FreeSans 448 0 0 0 FrameData[104]
port 5 nsew signal input
flabel metal3 s 0 567840 112 567952 0 FreeSans 448 0 0 0 FrameData[105]
port 6 nsew signal input
flabel metal3 s 0 568736 112 568848 0 FreeSans 448 0 0 0 FrameData[106]
port 7 nsew signal input
flabel metal3 s 0 569632 112 569744 0 FreeSans 448 0 0 0 FrameData[107]
port 8 nsew signal input
flabel metal3 s 0 570528 112 570640 0 FreeSans 448 0 0 0 FrameData[108]
port 9 nsew signal input
flabel metal3 s 0 571424 112 571536 0 FreeSans 448 0 0 0 FrameData[109]
port 10 nsew signal input
flabel metal3 s 0 709296 112 709408 0 FreeSans 448 0 0 0 FrameData[10]
port 11 nsew signal input
flabel metal3 s 0 572320 112 572432 0 FreeSans 448 0 0 0 FrameData[110]
port 12 nsew signal input
flabel metal3 s 0 573216 112 573328 0 FreeSans 448 0 0 0 FrameData[111]
port 13 nsew signal input
flabel metal3 s 0 574112 112 574224 0 FreeSans 448 0 0 0 FrameData[112]
port 14 nsew signal input
flabel metal3 s 0 575008 112 575120 0 FreeSans 448 0 0 0 FrameData[113]
port 15 nsew signal input
flabel metal3 s 0 575904 112 576016 0 FreeSans 448 0 0 0 FrameData[114]
port 16 nsew signal input
flabel metal3 s 0 576800 112 576912 0 FreeSans 448 0 0 0 FrameData[115]
port 17 nsew signal input
flabel metal3 s 0 577696 112 577808 0 FreeSans 448 0 0 0 FrameData[116]
port 18 nsew signal input
flabel metal3 s 0 578592 112 578704 0 FreeSans 448 0 0 0 FrameData[117]
port 19 nsew signal input
flabel metal3 s 0 579488 112 579600 0 FreeSans 448 0 0 0 FrameData[118]
port 20 nsew signal input
flabel metal3 s 0 580384 112 580496 0 FreeSans 448 0 0 0 FrameData[119]
port 21 nsew signal input
flabel metal3 s 0 709744 112 709856 0 FreeSans 448 0 0 0 FrameData[11]
port 22 nsew signal input
flabel metal3 s 0 581280 112 581392 0 FreeSans 448 0 0 0 FrameData[120]
port 23 nsew signal input
flabel metal3 s 0 582176 112 582288 0 FreeSans 448 0 0 0 FrameData[121]
port 24 nsew signal input
flabel metal3 s 0 583072 112 583184 0 FreeSans 448 0 0 0 FrameData[122]
port 25 nsew signal input
flabel metal3 s 0 583968 112 584080 0 FreeSans 448 0 0 0 FrameData[123]
port 26 nsew signal input
flabel metal3 s 0 584864 112 584976 0 FreeSans 448 0 0 0 FrameData[124]
port 27 nsew signal input
flabel metal3 s 0 585760 112 585872 0 FreeSans 448 0 0 0 FrameData[125]
port 28 nsew signal input
flabel metal3 s 0 586656 112 586768 0 FreeSans 448 0 0 0 FrameData[126]
port 29 nsew signal input
flabel metal3 s 0 587552 112 587664 0 FreeSans 448 0 0 0 FrameData[127]
port 30 nsew signal input
flabel metal3 s 0 502320 112 502432 0 FreeSans 448 0 0 0 FrameData[128]
port 31 nsew signal input
flabel metal3 s 0 503216 112 503328 0 FreeSans 448 0 0 0 FrameData[129]
port 32 nsew signal input
flabel metal3 s 0 710192 112 710304 0 FreeSans 448 0 0 0 FrameData[12]
port 33 nsew signal input
flabel metal3 s 0 504112 112 504224 0 FreeSans 448 0 0 0 FrameData[130]
port 34 nsew signal input
flabel metal3 s 0 505008 112 505120 0 FreeSans 448 0 0 0 FrameData[131]
port 35 nsew signal input
flabel metal3 s 0 505904 112 506016 0 FreeSans 448 0 0 0 FrameData[132]
port 36 nsew signal input
flabel metal3 s 0 506800 112 506912 0 FreeSans 448 0 0 0 FrameData[133]
port 37 nsew signal input
flabel metal3 s 0 507696 112 507808 0 FreeSans 448 0 0 0 FrameData[134]
port 38 nsew signal input
flabel metal3 s 0 508592 112 508704 0 FreeSans 448 0 0 0 FrameData[135]
port 39 nsew signal input
flabel metal3 s 0 509488 112 509600 0 FreeSans 448 0 0 0 FrameData[136]
port 40 nsew signal input
flabel metal3 s 0 510384 112 510496 0 FreeSans 448 0 0 0 FrameData[137]
port 41 nsew signal input
flabel metal3 s 0 511280 112 511392 0 FreeSans 448 0 0 0 FrameData[138]
port 42 nsew signal input
flabel metal3 s 0 512176 112 512288 0 FreeSans 448 0 0 0 FrameData[139]
port 43 nsew signal input
flabel metal3 s 0 710640 112 710752 0 FreeSans 448 0 0 0 FrameData[13]
port 44 nsew signal input
flabel metal3 s 0 513072 112 513184 0 FreeSans 448 0 0 0 FrameData[140]
port 45 nsew signal input
flabel metal3 s 0 513968 112 514080 0 FreeSans 448 0 0 0 FrameData[141]
port 46 nsew signal input
flabel metal3 s 0 514864 112 514976 0 FreeSans 448 0 0 0 FrameData[142]
port 47 nsew signal input
flabel metal3 s 0 515760 112 515872 0 FreeSans 448 0 0 0 FrameData[143]
port 48 nsew signal input
flabel metal3 s 0 516656 112 516768 0 FreeSans 448 0 0 0 FrameData[144]
port 49 nsew signal input
flabel metal3 s 0 517552 112 517664 0 FreeSans 448 0 0 0 FrameData[145]
port 50 nsew signal input
flabel metal3 s 0 518448 112 518560 0 FreeSans 448 0 0 0 FrameData[146]
port 51 nsew signal input
flabel metal3 s 0 519344 112 519456 0 FreeSans 448 0 0 0 FrameData[147]
port 52 nsew signal input
flabel metal3 s 0 520240 112 520352 0 FreeSans 448 0 0 0 FrameData[148]
port 53 nsew signal input
flabel metal3 s 0 521136 112 521248 0 FreeSans 448 0 0 0 FrameData[149]
port 54 nsew signal input
flabel metal3 s 0 711088 112 711200 0 FreeSans 448 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 522032 112 522144 0 FreeSans 448 0 0 0 FrameData[150]
port 56 nsew signal input
flabel metal3 s 0 522928 112 523040 0 FreeSans 448 0 0 0 FrameData[151]
port 57 nsew signal input
flabel metal3 s 0 523824 112 523936 0 FreeSans 448 0 0 0 FrameData[152]
port 58 nsew signal input
flabel metal3 s 0 524720 112 524832 0 FreeSans 448 0 0 0 FrameData[153]
port 59 nsew signal input
flabel metal3 s 0 525616 112 525728 0 FreeSans 448 0 0 0 FrameData[154]
port 60 nsew signal input
flabel metal3 s 0 526512 112 526624 0 FreeSans 448 0 0 0 FrameData[155]
port 61 nsew signal input
flabel metal3 s 0 527408 112 527520 0 FreeSans 448 0 0 0 FrameData[156]
port 62 nsew signal input
flabel metal3 s 0 528304 112 528416 0 FreeSans 448 0 0 0 FrameData[157]
port 63 nsew signal input
flabel metal3 s 0 529200 112 529312 0 FreeSans 448 0 0 0 FrameData[158]
port 64 nsew signal input
flabel metal3 s 0 530096 112 530208 0 FreeSans 448 0 0 0 FrameData[159]
port 65 nsew signal input
flabel metal3 s 0 711536 112 711648 0 FreeSans 448 0 0 0 FrameData[15]
port 66 nsew signal input
flabel metal3 s 0 444864 112 444976 0 FreeSans 448 0 0 0 FrameData[160]
port 67 nsew signal input
flabel metal3 s 0 445760 112 445872 0 FreeSans 448 0 0 0 FrameData[161]
port 68 nsew signal input
flabel metal3 s 0 446656 112 446768 0 FreeSans 448 0 0 0 FrameData[162]
port 69 nsew signal input
flabel metal3 s 0 447552 112 447664 0 FreeSans 448 0 0 0 FrameData[163]
port 70 nsew signal input
flabel metal3 s 0 448448 112 448560 0 FreeSans 448 0 0 0 FrameData[164]
port 71 nsew signal input
flabel metal3 s 0 449344 112 449456 0 FreeSans 448 0 0 0 FrameData[165]
port 72 nsew signal input
flabel metal3 s 0 450240 112 450352 0 FreeSans 448 0 0 0 FrameData[166]
port 73 nsew signal input
flabel metal3 s 0 451136 112 451248 0 FreeSans 448 0 0 0 FrameData[167]
port 74 nsew signal input
flabel metal3 s 0 452032 112 452144 0 FreeSans 448 0 0 0 FrameData[168]
port 75 nsew signal input
flabel metal3 s 0 452928 112 453040 0 FreeSans 448 0 0 0 FrameData[169]
port 76 nsew signal input
flabel metal3 s 0 711984 112 712096 0 FreeSans 448 0 0 0 FrameData[16]
port 77 nsew signal input
flabel metal3 s 0 453824 112 453936 0 FreeSans 448 0 0 0 FrameData[170]
port 78 nsew signal input
flabel metal3 s 0 454720 112 454832 0 FreeSans 448 0 0 0 FrameData[171]
port 79 nsew signal input
flabel metal3 s 0 455616 112 455728 0 FreeSans 448 0 0 0 FrameData[172]
port 80 nsew signal input
flabel metal3 s 0 456512 112 456624 0 FreeSans 448 0 0 0 FrameData[173]
port 81 nsew signal input
flabel metal3 s 0 457408 112 457520 0 FreeSans 448 0 0 0 FrameData[174]
port 82 nsew signal input
flabel metal3 s 0 458304 112 458416 0 FreeSans 448 0 0 0 FrameData[175]
port 83 nsew signal input
flabel metal3 s 0 459200 112 459312 0 FreeSans 448 0 0 0 FrameData[176]
port 84 nsew signal input
flabel metal3 s 0 460096 112 460208 0 FreeSans 448 0 0 0 FrameData[177]
port 85 nsew signal input
flabel metal3 s 0 460992 112 461104 0 FreeSans 448 0 0 0 FrameData[178]
port 86 nsew signal input
flabel metal3 s 0 461888 112 462000 0 FreeSans 448 0 0 0 FrameData[179]
port 87 nsew signal input
flabel metal3 s 0 712432 112 712544 0 FreeSans 448 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 462784 112 462896 0 FreeSans 448 0 0 0 FrameData[180]
port 89 nsew signal input
flabel metal3 s 0 463680 112 463792 0 FreeSans 448 0 0 0 FrameData[181]
port 90 nsew signal input
flabel metal3 s 0 464576 112 464688 0 FreeSans 448 0 0 0 FrameData[182]
port 91 nsew signal input
flabel metal3 s 0 465472 112 465584 0 FreeSans 448 0 0 0 FrameData[183]
port 92 nsew signal input
flabel metal3 s 0 466368 112 466480 0 FreeSans 448 0 0 0 FrameData[184]
port 93 nsew signal input
flabel metal3 s 0 467264 112 467376 0 FreeSans 448 0 0 0 FrameData[185]
port 94 nsew signal input
flabel metal3 s 0 468160 112 468272 0 FreeSans 448 0 0 0 FrameData[186]
port 95 nsew signal input
flabel metal3 s 0 469056 112 469168 0 FreeSans 448 0 0 0 FrameData[187]
port 96 nsew signal input
flabel metal3 s 0 469952 112 470064 0 FreeSans 448 0 0 0 FrameData[188]
port 97 nsew signal input
flabel metal3 s 0 470848 112 470960 0 FreeSans 448 0 0 0 FrameData[189]
port 98 nsew signal input
flabel metal3 s 0 712880 112 712992 0 FreeSans 448 0 0 0 FrameData[18]
port 99 nsew signal input
flabel metal3 s 0 471744 112 471856 0 FreeSans 448 0 0 0 FrameData[190]
port 100 nsew signal input
flabel metal3 s 0 472640 112 472752 0 FreeSans 448 0 0 0 FrameData[191]
port 101 nsew signal input
flabel metal3 s 0 387408 112 387520 0 FreeSans 448 0 0 0 FrameData[192]
port 102 nsew signal input
flabel metal3 s 0 388304 112 388416 0 FreeSans 448 0 0 0 FrameData[193]
port 103 nsew signal input
flabel metal3 s 0 389200 112 389312 0 FreeSans 448 0 0 0 FrameData[194]
port 104 nsew signal input
flabel metal3 s 0 390096 112 390208 0 FreeSans 448 0 0 0 FrameData[195]
port 105 nsew signal input
flabel metal3 s 0 390992 112 391104 0 FreeSans 448 0 0 0 FrameData[196]
port 106 nsew signal input
flabel metal3 s 0 391888 112 392000 0 FreeSans 448 0 0 0 FrameData[197]
port 107 nsew signal input
flabel metal3 s 0 392784 112 392896 0 FreeSans 448 0 0 0 FrameData[198]
port 108 nsew signal input
flabel metal3 s 0 393680 112 393792 0 FreeSans 448 0 0 0 FrameData[199]
port 109 nsew signal input
flabel metal3 s 0 713328 112 713440 0 FreeSans 448 0 0 0 FrameData[19]
port 110 nsew signal input
flabel metal3 s 0 705264 112 705376 0 FreeSans 448 0 0 0 FrameData[1]
port 111 nsew signal input
flabel metal3 s 0 394576 112 394688 0 FreeSans 448 0 0 0 FrameData[200]
port 112 nsew signal input
flabel metal3 s 0 395472 112 395584 0 FreeSans 448 0 0 0 FrameData[201]
port 113 nsew signal input
flabel metal3 s 0 396368 112 396480 0 FreeSans 448 0 0 0 FrameData[202]
port 114 nsew signal input
flabel metal3 s 0 397264 112 397376 0 FreeSans 448 0 0 0 FrameData[203]
port 115 nsew signal input
flabel metal3 s 0 398160 112 398272 0 FreeSans 448 0 0 0 FrameData[204]
port 116 nsew signal input
flabel metal3 s 0 399056 112 399168 0 FreeSans 448 0 0 0 FrameData[205]
port 117 nsew signal input
flabel metal3 s 0 399952 112 400064 0 FreeSans 448 0 0 0 FrameData[206]
port 118 nsew signal input
flabel metal3 s 0 400848 112 400960 0 FreeSans 448 0 0 0 FrameData[207]
port 119 nsew signal input
flabel metal3 s 0 401744 112 401856 0 FreeSans 448 0 0 0 FrameData[208]
port 120 nsew signal input
flabel metal3 s 0 402640 112 402752 0 FreeSans 448 0 0 0 FrameData[209]
port 121 nsew signal input
flabel metal3 s 0 713776 112 713888 0 FreeSans 448 0 0 0 FrameData[20]
port 122 nsew signal input
flabel metal3 s 0 403536 112 403648 0 FreeSans 448 0 0 0 FrameData[210]
port 123 nsew signal input
flabel metal3 s 0 404432 112 404544 0 FreeSans 448 0 0 0 FrameData[211]
port 124 nsew signal input
flabel metal3 s 0 405328 112 405440 0 FreeSans 448 0 0 0 FrameData[212]
port 125 nsew signal input
flabel metal3 s 0 406224 112 406336 0 FreeSans 448 0 0 0 FrameData[213]
port 126 nsew signal input
flabel metal3 s 0 407120 112 407232 0 FreeSans 448 0 0 0 FrameData[214]
port 127 nsew signal input
flabel metal3 s 0 408016 112 408128 0 FreeSans 448 0 0 0 FrameData[215]
port 128 nsew signal input
flabel metal3 s 0 408912 112 409024 0 FreeSans 448 0 0 0 FrameData[216]
port 129 nsew signal input
flabel metal3 s 0 409808 112 409920 0 FreeSans 448 0 0 0 FrameData[217]
port 130 nsew signal input
flabel metal3 s 0 410704 112 410816 0 FreeSans 448 0 0 0 FrameData[218]
port 131 nsew signal input
flabel metal3 s 0 411600 112 411712 0 FreeSans 448 0 0 0 FrameData[219]
port 132 nsew signal input
flabel metal3 s 0 714224 112 714336 0 FreeSans 448 0 0 0 FrameData[21]
port 133 nsew signal input
flabel metal3 s 0 412496 112 412608 0 FreeSans 448 0 0 0 FrameData[220]
port 134 nsew signal input
flabel metal3 s 0 413392 112 413504 0 FreeSans 448 0 0 0 FrameData[221]
port 135 nsew signal input
flabel metal3 s 0 414288 112 414400 0 FreeSans 448 0 0 0 FrameData[222]
port 136 nsew signal input
flabel metal3 s 0 415184 112 415296 0 FreeSans 448 0 0 0 FrameData[223]
port 137 nsew signal input
flabel metal3 s 0 329952 112 330064 0 FreeSans 448 0 0 0 FrameData[224]
port 138 nsew signal input
flabel metal3 s 0 330848 112 330960 0 FreeSans 448 0 0 0 FrameData[225]
port 139 nsew signal input
flabel metal3 s 0 331744 112 331856 0 FreeSans 448 0 0 0 FrameData[226]
port 140 nsew signal input
flabel metal3 s 0 332640 112 332752 0 FreeSans 448 0 0 0 FrameData[227]
port 141 nsew signal input
flabel metal3 s 0 333536 112 333648 0 FreeSans 448 0 0 0 FrameData[228]
port 142 nsew signal input
flabel metal3 s 0 334432 112 334544 0 FreeSans 448 0 0 0 FrameData[229]
port 143 nsew signal input
flabel metal3 s 0 714672 112 714784 0 FreeSans 448 0 0 0 FrameData[22]
port 144 nsew signal input
flabel metal3 s 0 335328 112 335440 0 FreeSans 448 0 0 0 FrameData[230]
port 145 nsew signal input
flabel metal3 s 0 336224 112 336336 0 FreeSans 448 0 0 0 FrameData[231]
port 146 nsew signal input
flabel metal3 s 0 337120 112 337232 0 FreeSans 448 0 0 0 FrameData[232]
port 147 nsew signal input
flabel metal3 s 0 338016 112 338128 0 FreeSans 448 0 0 0 FrameData[233]
port 148 nsew signal input
flabel metal3 s 0 338912 112 339024 0 FreeSans 448 0 0 0 FrameData[234]
port 149 nsew signal input
flabel metal3 s 0 339808 112 339920 0 FreeSans 448 0 0 0 FrameData[235]
port 150 nsew signal input
flabel metal3 s 0 340704 112 340816 0 FreeSans 448 0 0 0 FrameData[236]
port 151 nsew signal input
flabel metal3 s 0 341600 112 341712 0 FreeSans 448 0 0 0 FrameData[237]
port 152 nsew signal input
flabel metal3 s 0 342496 112 342608 0 FreeSans 448 0 0 0 FrameData[238]
port 153 nsew signal input
flabel metal3 s 0 343392 112 343504 0 FreeSans 448 0 0 0 FrameData[239]
port 154 nsew signal input
flabel metal3 s 0 715120 112 715232 0 FreeSans 448 0 0 0 FrameData[23]
port 155 nsew signal input
flabel metal3 s 0 344288 112 344400 0 FreeSans 448 0 0 0 FrameData[240]
port 156 nsew signal input
flabel metal3 s 0 345184 112 345296 0 FreeSans 448 0 0 0 FrameData[241]
port 157 nsew signal input
flabel metal3 s 0 346080 112 346192 0 FreeSans 448 0 0 0 FrameData[242]
port 158 nsew signal input
flabel metal3 s 0 346976 112 347088 0 FreeSans 448 0 0 0 FrameData[243]
port 159 nsew signal input
flabel metal3 s 0 347872 112 347984 0 FreeSans 448 0 0 0 FrameData[244]
port 160 nsew signal input
flabel metal3 s 0 348768 112 348880 0 FreeSans 448 0 0 0 FrameData[245]
port 161 nsew signal input
flabel metal3 s 0 349664 112 349776 0 FreeSans 448 0 0 0 FrameData[246]
port 162 nsew signal input
flabel metal3 s 0 350560 112 350672 0 FreeSans 448 0 0 0 FrameData[247]
port 163 nsew signal input
flabel metal3 s 0 351456 112 351568 0 FreeSans 448 0 0 0 FrameData[248]
port 164 nsew signal input
flabel metal3 s 0 352352 112 352464 0 FreeSans 448 0 0 0 FrameData[249]
port 165 nsew signal input
flabel metal3 s 0 715568 112 715680 0 FreeSans 448 0 0 0 FrameData[24]
port 166 nsew signal input
flabel metal3 s 0 353248 112 353360 0 FreeSans 448 0 0 0 FrameData[250]
port 167 nsew signal input
flabel metal3 s 0 354144 112 354256 0 FreeSans 448 0 0 0 FrameData[251]
port 168 nsew signal input
flabel metal3 s 0 355040 112 355152 0 FreeSans 448 0 0 0 FrameData[252]
port 169 nsew signal input
flabel metal3 s 0 355936 112 356048 0 FreeSans 448 0 0 0 FrameData[253]
port 170 nsew signal input
flabel metal3 s 0 356832 112 356944 0 FreeSans 448 0 0 0 FrameData[254]
port 171 nsew signal input
flabel metal3 s 0 357728 112 357840 0 FreeSans 448 0 0 0 FrameData[255]
port 172 nsew signal input
flabel metal3 s 0 272496 112 272608 0 FreeSans 448 0 0 0 FrameData[256]
port 173 nsew signal input
flabel metal3 s 0 273392 112 273504 0 FreeSans 448 0 0 0 FrameData[257]
port 174 nsew signal input
flabel metal3 s 0 274288 112 274400 0 FreeSans 448 0 0 0 FrameData[258]
port 175 nsew signal input
flabel metal3 s 0 275184 112 275296 0 FreeSans 448 0 0 0 FrameData[259]
port 176 nsew signal input
flabel metal3 s 0 716016 112 716128 0 FreeSans 448 0 0 0 FrameData[25]
port 177 nsew signal input
flabel metal3 s 0 276080 112 276192 0 FreeSans 448 0 0 0 FrameData[260]
port 178 nsew signal input
flabel metal3 s 0 276976 112 277088 0 FreeSans 448 0 0 0 FrameData[261]
port 179 nsew signal input
flabel metal3 s 0 277872 112 277984 0 FreeSans 448 0 0 0 FrameData[262]
port 180 nsew signal input
flabel metal3 s 0 278768 112 278880 0 FreeSans 448 0 0 0 FrameData[263]
port 181 nsew signal input
flabel metal3 s 0 279664 112 279776 0 FreeSans 448 0 0 0 FrameData[264]
port 182 nsew signal input
flabel metal3 s 0 280560 112 280672 0 FreeSans 448 0 0 0 FrameData[265]
port 183 nsew signal input
flabel metal3 s 0 281456 112 281568 0 FreeSans 448 0 0 0 FrameData[266]
port 184 nsew signal input
flabel metal3 s 0 282352 112 282464 0 FreeSans 448 0 0 0 FrameData[267]
port 185 nsew signal input
flabel metal3 s 0 283248 112 283360 0 FreeSans 448 0 0 0 FrameData[268]
port 186 nsew signal input
flabel metal3 s 0 284144 112 284256 0 FreeSans 448 0 0 0 FrameData[269]
port 187 nsew signal input
flabel metal3 s 0 716464 112 716576 0 FreeSans 448 0 0 0 FrameData[26]
port 188 nsew signal input
flabel metal3 s 0 285040 112 285152 0 FreeSans 448 0 0 0 FrameData[270]
port 189 nsew signal input
flabel metal3 s 0 285936 112 286048 0 FreeSans 448 0 0 0 FrameData[271]
port 190 nsew signal input
flabel metal3 s 0 286832 112 286944 0 FreeSans 448 0 0 0 FrameData[272]
port 191 nsew signal input
flabel metal3 s 0 287728 112 287840 0 FreeSans 448 0 0 0 FrameData[273]
port 192 nsew signal input
flabel metal3 s 0 288624 112 288736 0 FreeSans 448 0 0 0 FrameData[274]
port 193 nsew signal input
flabel metal3 s 0 289520 112 289632 0 FreeSans 448 0 0 0 FrameData[275]
port 194 nsew signal input
flabel metal3 s 0 290416 112 290528 0 FreeSans 448 0 0 0 FrameData[276]
port 195 nsew signal input
flabel metal3 s 0 291312 112 291424 0 FreeSans 448 0 0 0 FrameData[277]
port 196 nsew signal input
flabel metal3 s 0 292208 112 292320 0 FreeSans 448 0 0 0 FrameData[278]
port 197 nsew signal input
flabel metal3 s 0 293104 112 293216 0 FreeSans 448 0 0 0 FrameData[279]
port 198 nsew signal input
flabel metal3 s 0 716912 112 717024 0 FreeSans 448 0 0 0 FrameData[27]
port 199 nsew signal input
flabel metal3 s 0 294000 112 294112 0 FreeSans 448 0 0 0 FrameData[280]
port 200 nsew signal input
flabel metal3 s 0 294896 112 295008 0 FreeSans 448 0 0 0 FrameData[281]
port 201 nsew signal input
flabel metal3 s 0 295792 112 295904 0 FreeSans 448 0 0 0 FrameData[282]
port 202 nsew signal input
flabel metal3 s 0 296688 112 296800 0 FreeSans 448 0 0 0 FrameData[283]
port 203 nsew signal input
flabel metal3 s 0 297584 112 297696 0 FreeSans 448 0 0 0 FrameData[284]
port 204 nsew signal input
flabel metal3 s 0 298480 112 298592 0 FreeSans 448 0 0 0 FrameData[285]
port 205 nsew signal input
flabel metal3 s 0 299376 112 299488 0 FreeSans 448 0 0 0 FrameData[286]
port 206 nsew signal input
flabel metal3 s 0 300272 112 300384 0 FreeSans 448 0 0 0 FrameData[287]
port 207 nsew signal input
flabel metal3 s 0 215040 112 215152 0 FreeSans 448 0 0 0 FrameData[288]
port 208 nsew signal input
flabel metal3 s 0 215936 112 216048 0 FreeSans 448 0 0 0 FrameData[289]
port 209 nsew signal input
flabel metal3 s 0 717360 112 717472 0 FreeSans 448 0 0 0 FrameData[28]
port 210 nsew signal input
flabel metal3 s 0 216832 112 216944 0 FreeSans 448 0 0 0 FrameData[290]
port 211 nsew signal input
flabel metal3 s 0 217728 112 217840 0 FreeSans 448 0 0 0 FrameData[291]
port 212 nsew signal input
flabel metal3 s 0 218624 112 218736 0 FreeSans 448 0 0 0 FrameData[292]
port 213 nsew signal input
flabel metal3 s 0 219520 112 219632 0 FreeSans 448 0 0 0 FrameData[293]
port 214 nsew signal input
flabel metal3 s 0 220416 112 220528 0 FreeSans 448 0 0 0 FrameData[294]
port 215 nsew signal input
flabel metal3 s 0 221312 112 221424 0 FreeSans 448 0 0 0 FrameData[295]
port 216 nsew signal input
flabel metal3 s 0 222208 112 222320 0 FreeSans 448 0 0 0 FrameData[296]
port 217 nsew signal input
flabel metal3 s 0 223104 112 223216 0 FreeSans 448 0 0 0 FrameData[297]
port 218 nsew signal input
flabel metal3 s 0 224000 112 224112 0 FreeSans 448 0 0 0 FrameData[298]
port 219 nsew signal input
flabel metal3 s 0 224896 112 225008 0 FreeSans 448 0 0 0 FrameData[299]
port 220 nsew signal input
flabel metal3 s 0 717808 112 717920 0 FreeSans 448 0 0 0 FrameData[29]
port 221 nsew signal input
flabel metal3 s 0 705712 112 705824 0 FreeSans 448 0 0 0 FrameData[2]
port 222 nsew signal input
flabel metal3 s 0 225792 112 225904 0 FreeSans 448 0 0 0 FrameData[300]
port 223 nsew signal input
flabel metal3 s 0 226688 112 226800 0 FreeSans 448 0 0 0 FrameData[301]
port 224 nsew signal input
flabel metal3 s 0 227584 112 227696 0 FreeSans 448 0 0 0 FrameData[302]
port 225 nsew signal input
flabel metal3 s 0 228480 112 228592 0 FreeSans 448 0 0 0 FrameData[303]
port 226 nsew signal input
flabel metal3 s 0 229376 112 229488 0 FreeSans 448 0 0 0 FrameData[304]
port 227 nsew signal input
flabel metal3 s 0 230272 112 230384 0 FreeSans 448 0 0 0 FrameData[305]
port 228 nsew signal input
flabel metal3 s 0 231168 112 231280 0 FreeSans 448 0 0 0 FrameData[306]
port 229 nsew signal input
flabel metal3 s 0 232064 112 232176 0 FreeSans 448 0 0 0 FrameData[307]
port 230 nsew signal input
flabel metal3 s 0 232960 112 233072 0 FreeSans 448 0 0 0 FrameData[308]
port 231 nsew signal input
flabel metal3 s 0 233856 112 233968 0 FreeSans 448 0 0 0 FrameData[309]
port 232 nsew signal input
flabel metal3 s 0 718256 112 718368 0 FreeSans 448 0 0 0 FrameData[30]
port 233 nsew signal input
flabel metal3 s 0 234752 112 234864 0 FreeSans 448 0 0 0 FrameData[310]
port 234 nsew signal input
flabel metal3 s 0 235648 112 235760 0 FreeSans 448 0 0 0 FrameData[311]
port 235 nsew signal input
flabel metal3 s 0 236544 112 236656 0 FreeSans 448 0 0 0 FrameData[312]
port 236 nsew signal input
flabel metal3 s 0 237440 112 237552 0 FreeSans 448 0 0 0 FrameData[313]
port 237 nsew signal input
flabel metal3 s 0 238336 112 238448 0 FreeSans 448 0 0 0 FrameData[314]
port 238 nsew signal input
flabel metal3 s 0 239232 112 239344 0 FreeSans 448 0 0 0 FrameData[315]
port 239 nsew signal input
flabel metal3 s 0 240128 112 240240 0 FreeSans 448 0 0 0 FrameData[316]
port 240 nsew signal input
flabel metal3 s 0 241024 112 241136 0 FreeSans 448 0 0 0 FrameData[317]
port 241 nsew signal input
flabel metal3 s 0 241920 112 242032 0 FreeSans 448 0 0 0 FrameData[318]
port 242 nsew signal input
flabel metal3 s 0 242816 112 242928 0 FreeSans 448 0 0 0 FrameData[319]
port 243 nsew signal input
flabel metal3 s 0 718704 112 718816 0 FreeSans 448 0 0 0 FrameData[31]
port 244 nsew signal input
flabel metal3 s 0 157584 112 157696 0 FreeSans 448 0 0 0 FrameData[320]
port 245 nsew signal input
flabel metal3 s 0 158480 112 158592 0 FreeSans 448 0 0 0 FrameData[321]
port 246 nsew signal input
flabel metal3 s 0 159376 112 159488 0 FreeSans 448 0 0 0 FrameData[322]
port 247 nsew signal input
flabel metal3 s 0 160272 112 160384 0 FreeSans 448 0 0 0 FrameData[323]
port 248 nsew signal input
flabel metal3 s 0 161168 112 161280 0 FreeSans 448 0 0 0 FrameData[324]
port 249 nsew signal input
flabel metal3 s 0 162064 112 162176 0 FreeSans 448 0 0 0 FrameData[325]
port 250 nsew signal input
flabel metal3 s 0 162960 112 163072 0 FreeSans 448 0 0 0 FrameData[326]
port 251 nsew signal input
flabel metal3 s 0 163856 112 163968 0 FreeSans 448 0 0 0 FrameData[327]
port 252 nsew signal input
flabel metal3 s 0 164752 112 164864 0 FreeSans 448 0 0 0 FrameData[328]
port 253 nsew signal input
flabel metal3 s 0 165648 112 165760 0 FreeSans 448 0 0 0 FrameData[329]
port 254 nsew signal input
flabel metal3 s 0 674688 112 674800 0 FreeSans 448 0 0 0 FrameData[32]
port 255 nsew signal input
flabel metal3 s 0 166544 112 166656 0 FreeSans 448 0 0 0 FrameData[330]
port 256 nsew signal input
flabel metal3 s 0 167440 112 167552 0 FreeSans 448 0 0 0 FrameData[331]
port 257 nsew signal input
flabel metal3 s 0 168336 112 168448 0 FreeSans 448 0 0 0 FrameData[332]
port 258 nsew signal input
flabel metal3 s 0 169232 112 169344 0 FreeSans 448 0 0 0 FrameData[333]
port 259 nsew signal input
flabel metal3 s 0 170128 112 170240 0 FreeSans 448 0 0 0 FrameData[334]
port 260 nsew signal input
flabel metal3 s 0 171024 112 171136 0 FreeSans 448 0 0 0 FrameData[335]
port 261 nsew signal input
flabel metal3 s 0 171920 112 172032 0 FreeSans 448 0 0 0 FrameData[336]
port 262 nsew signal input
flabel metal3 s 0 172816 112 172928 0 FreeSans 448 0 0 0 FrameData[337]
port 263 nsew signal input
flabel metal3 s 0 173712 112 173824 0 FreeSans 448 0 0 0 FrameData[338]
port 264 nsew signal input
flabel metal3 s 0 174608 112 174720 0 FreeSans 448 0 0 0 FrameData[339]
port 265 nsew signal input
flabel metal3 s 0 675584 112 675696 0 FreeSans 448 0 0 0 FrameData[33]
port 266 nsew signal input
flabel metal3 s 0 175504 112 175616 0 FreeSans 448 0 0 0 FrameData[340]
port 267 nsew signal input
flabel metal3 s 0 176400 112 176512 0 FreeSans 448 0 0 0 FrameData[341]
port 268 nsew signal input
flabel metal3 s 0 177296 112 177408 0 FreeSans 448 0 0 0 FrameData[342]
port 269 nsew signal input
flabel metal3 s 0 178192 112 178304 0 FreeSans 448 0 0 0 FrameData[343]
port 270 nsew signal input
flabel metal3 s 0 179088 112 179200 0 FreeSans 448 0 0 0 FrameData[344]
port 271 nsew signal input
flabel metal3 s 0 179984 112 180096 0 FreeSans 448 0 0 0 FrameData[345]
port 272 nsew signal input
flabel metal3 s 0 180880 112 180992 0 FreeSans 448 0 0 0 FrameData[346]
port 273 nsew signal input
flabel metal3 s 0 181776 112 181888 0 FreeSans 448 0 0 0 FrameData[347]
port 274 nsew signal input
flabel metal3 s 0 182672 112 182784 0 FreeSans 448 0 0 0 FrameData[348]
port 275 nsew signal input
flabel metal3 s 0 183568 112 183680 0 FreeSans 448 0 0 0 FrameData[349]
port 276 nsew signal input
flabel metal3 s 0 676480 112 676592 0 FreeSans 448 0 0 0 FrameData[34]
port 277 nsew signal input
flabel metal3 s 0 184464 112 184576 0 FreeSans 448 0 0 0 FrameData[350]
port 278 nsew signal input
flabel metal3 s 0 185360 112 185472 0 FreeSans 448 0 0 0 FrameData[351]
port 279 nsew signal input
flabel metal3 s 0 100128 112 100240 0 FreeSans 448 0 0 0 FrameData[352]
port 280 nsew signal input
flabel metal3 s 0 101024 112 101136 0 FreeSans 448 0 0 0 FrameData[353]
port 281 nsew signal input
flabel metal3 s 0 101920 112 102032 0 FreeSans 448 0 0 0 FrameData[354]
port 282 nsew signal input
flabel metal3 s 0 102816 112 102928 0 FreeSans 448 0 0 0 FrameData[355]
port 283 nsew signal input
flabel metal3 s 0 103712 112 103824 0 FreeSans 448 0 0 0 FrameData[356]
port 284 nsew signal input
flabel metal3 s 0 104608 112 104720 0 FreeSans 448 0 0 0 FrameData[357]
port 285 nsew signal input
flabel metal3 s 0 105504 112 105616 0 FreeSans 448 0 0 0 FrameData[358]
port 286 nsew signal input
flabel metal3 s 0 106400 112 106512 0 FreeSans 448 0 0 0 FrameData[359]
port 287 nsew signal input
flabel metal3 s 0 677376 112 677488 0 FreeSans 448 0 0 0 FrameData[35]
port 288 nsew signal input
flabel metal3 s 0 107296 112 107408 0 FreeSans 448 0 0 0 FrameData[360]
port 289 nsew signal input
flabel metal3 s 0 108192 112 108304 0 FreeSans 448 0 0 0 FrameData[361]
port 290 nsew signal input
flabel metal3 s 0 109088 112 109200 0 FreeSans 448 0 0 0 FrameData[362]
port 291 nsew signal input
flabel metal3 s 0 109984 112 110096 0 FreeSans 448 0 0 0 FrameData[363]
port 292 nsew signal input
flabel metal3 s 0 110880 112 110992 0 FreeSans 448 0 0 0 FrameData[364]
port 293 nsew signal input
flabel metal3 s 0 111776 112 111888 0 FreeSans 448 0 0 0 FrameData[365]
port 294 nsew signal input
flabel metal3 s 0 112672 112 112784 0 FreeSans 448 0 0 0 FrameData[366]
port 295 nsew signal input
flabel metal3 s 0 113568 112 113680 0 FreeSans 448 0 0 0 FrameData[367]
port 296 nsew signal input
flabel metal3 s 0 114464 112 114576 0 FreeSans 448 0 0 0 FrameData[368]
port 297 nsew signal input
flabel metal3 s 0 115360 112 115472 0 FreeSans 448 0 0 0 FrameData[369]
port 298 nsew signal input
flabel metal3 s 0 678272 112 678384 0 FreeSans 448 0 0 0 FrameData[36]
port 299 nsew signal input
flabel metal3 s 0 116256 112 116368 0 FreeSans 448 0 0 0 FrameData[370]
port 300 nsew signal input
flabel metal3 s 0 117152 112 117264 0 FreeSans 448 0 0 0 FrameData[371]
port 301 nsew signal input
flabel metal3 s 0 118048 112 118160 0 FreeSans 448 0 0 0 FrameData[372]
port 302 nsew signal input
flabel metal3 s 0 118944 112 119056 0 FreeSans 448 0 0 0 FrameData[373]
port 303 nsew signal input
flabel metal3 s 0 119840 112 119952 0 FreeSans 448 0 0 0 FrameData[374]
port 304 nsew signal input
flabel metal3 s 0 120736 112 120848 0 FreeSans 448 0 0 0 FrameData[375]
port 305 nsew signal input
flabel metal3 s 0 121632 112 121744 0 FreeSans 448 0 0 0 FrameData[376]
port 306 nsew signal input
flabel metal3 s 0 122528 112 122640 0 FreeSans 448 0 0 0 FrameData[377]
port 307 nsew signal input
flabel metal3 s 0 123424 112 123536 0 FreeSans 448 0 0 0 FrameData[378]
port 308 nsew signal input
flabel metal3 s 0 124320 112 124432 0 FreeSans 448 0 0 0 FrameData[379]
port 309 nsew signal input
flabel metal3 s 0 679168 112 679280 0 FreeSans 448 0 0 0 FrameData[37]
port 310 nsew signal input
flabel metal3 s 0 125216 112 125328 0 FreeSans 448 0 0 0 FrameData[380]
port 311 nsew signal input
flabel metal3 s 0 126112 112 126224 0 FreeSans 448 0 0 0 FrameData[381]
port 312 nsew signal input
flabel metal3 s 0 127008 112 127120 0 FreeSans 448 0 0 0 FrameData[382]
port 313 nsew signal input
flabel metal3 s 0 127904 112 128016 0 FreeSans 448 0 0 0 FrameData[383]
port 314 nsew signal input
flabel metal3 s 0 42672 112 42784 0 FreeSans 448 0 0 0 FrameData[384]
port 315 nsew signal input
flabel metal3 s 0 43568 112 43680 0 FreeSans 448 0 0 0 FrameData[385]
port 316 nsew signal input
flabel metal3 s 0 44464 112 44576 0 FreeSans 448 0 0 0 FrameData[386]
port 317 nsew signal input
flabel metal3 s 0 45360 112 45472 0 FreeSans 448 0 0 0 FrameData[387]
port 318 nsew signal input
flabel metal3 s 0 46256 112 46368 0 FreeSans 448 0 0 0 FrameData[388]
port 319 nsew signal input
flabel metal3 s 0 47152 112 47264 0 FreeSans 448 0 0 0 FrameData[389]
port 320 nsew signal input
flabel metal3 s 0 680064 112 680176 0 FreeSans 448 0 0 0 FrameData[38]
port 321 nsew signal input
flabel metal3 s 0 48048 112 48160 0 FreeSans 448 0 0 0 FrameData[390]
port 322 nsew signal input
flabel metal3 s 0 48944 112 49056 0 FreeSans 448 0 0 0 FrameData[391]
port 323 nsew signal input
flabel metal3 s 0 49840 112 49952 0 FreeSans 448 0 0 0 FrameData[392]
port 324 nsew signal input
flabel metal3 s 0 50736 112 50848 0 FreeSans 448 0 0 0 FrameData[393]
port 325 nsew signal input
flabel metal3 s 0 51632 112 51744 0 FreeSans 448 0 0 0 FrameData[394]
port 326 nsew signal input
flabel metal3 s 0 52528 112 52640 0 FreeSans 448 0 0 0 FrameData[395]
port 327 nsew signal input
flabel metal3 s 0 53424 112 53536 0 FreeSans 448 0 0 0 FrameData[396]
port 328 nsew signal input
flabel metal3 s 0 54320 112 54432 0 FreeSans 448 0 0 0 FrameData[397]
port 329 nsew signal input
flabel metal3 s 0 55216 112 55328 0 FreeSans 448 0 0 0 FrameData[398]
port 330 nsew signal input
flabel metal3 s 0 56112 112 56224 0 FreeSans 448 0 0 0 FrameData[399]
port 331 nsew signal input
flabel metal3 s 0 680960 112 681072 0 FreeSans 448 0 0 0 FrameData[39]
port 332 nsew signal input
flabel metal3 s 0 706160 112 706272 0 FreeSans 448 0 0 0 FrameData[3]
port 333 nsew signal input
flabel metal3 s 0 57008 112 57120 0 FreeSans 448 0 0 0 FrameData[400]
port 334 nsew signal input
flabel metal3 s 0 57904 112 58016 0 FreeSans 448 0 0 0 FrameData[401]
port 335 nsew signal input
flabel metal3 s 0 58800 112 58912 0 FreeSans 448 0 0 0 FrameData[402]
port 336 nsew signal input
flabel metal3 s 0 59696 112 59808 0 FreeSans 448 0 0 0 FrameData[403]
port 337 nsew signal input
flabel metal3 s 0 60592 112 60704 0 FreeSans 448 0 0 0 FrameData[404]
port 338 nsew signal input
flabel metal3 s 0 61488 112 61600 0 FreeSans 448 0 0 0 FrameData[405]
port 339 nsew signal input
flabel metal3 s 0 62384 112 62496 0 FreeSans 448 0 0 0 FrameData[406]
port 340 nsew signal input
flabel metal3 s 0 63280 112 63392 0 FreeSans 448 0 0 0 FrameData[407]
port 341 nsew signal input
flabel metal3 s 0 64176 112 64288 0 FreeSans 448 0 0 0 FrameData[408]
port 342 nsew signal input
flabel metal3 s 0 65072 112 65184 0 FreeSans 448 0 0 0 FrameData[409]
port 343 nsew signal input
flabel metal3 s 0 681856 112 681968 0 FreeSans 448 0 0 0 FrameData[40]
port 344 nsew signal input
flabel metal3 s 0 65968 112 66080 0 FreeSans 448 0 0 0 FrameData[410]
port 345 nsew signal input
flabel metal3 s 0 66864 112 66976 0 FreeSans 448 0 0 0 FrameData[411]
port 346 nsew signal input
flabel metal3 s 0 67760 112 67872 0 FreeSans 448 0 0 0 FrameData[412]
port 347 nsew signal input
flabel metal3 s 0 68656 112 68768 0 FreeSans 448 0 0 0 FrameData[413]
port 348 nsew signal input
flabel metal3 s 0 69552 112 69664 0 FreeSans 448 0 0 0 FrameData[414]
port 349 nsew signal input
flabel metal3 s 0 70448 112 70560 0 FreeSans 448 0 0 0 FrameData[415]
port 350 nsew signal input
flabel metal3 s 0 1120 112 1232 0 FreeSans 448 0 0 0 FrameData[416]
port 351 nsew signal input
flabel metal3 s 0 1568 112 1680 0 FreeSans 448 0 0 0 FrameData[417]
port 352 nsew signal input
flabel metal3 s 0 2016 112 2128 0 FreeSans 448 0 0 0 FrameData[418]
port 353 nsew signal input
flabel metal3 s 0 2464 112 2576 0 FreeSans 448 0 0 0 FrameData[419]
port 354 nsew signal input
flabel metal3 s 0 682752 112 682864 0 FreeSans 448 0 0 0 FrameData[41]
port 355 nsew signal input
flabel metal3 s 0 2912 112 3024 0 FreeSans 448 0 0 0 FrameData[420]
port 356 nsew signal input
flabel metal3 s 0 3360 112 3472 0 FreeSans 448 0 0 0 FrameData[421]
port 357 nsew signal input
flabel metal3 s 0 3808 112 3920 0 FreeSans 448 0 0 0 FrameData[422]
port 358 nsew signal input
flabel metal3 s 0 4256 112 4368 0 FreeSans 448 0 0 0 FrameData[423]
port 359 nsew signal input
flabel metal3 s 0 4704 112 4816 0 FreeSans 448 0 0 0 FrameData[424]
port 360 nsew signal input
flabel metal3 s 0 5152 112 5264 0 FreeSans 448 0 0 0 FrameData[425]
port 361 nsew signal input
flabel metal3 s 0 5600 112 5712 0 FreeSans 448 0 0 0 FrameData[426]
port 362 nsew signal input
flabel metal3 s 0 6048 112 6160 0 FreeSans 448 0 0 0 FrameData[427]
port 363 nsew signal input
flabel metal3 s 0 6496 112 6608 0 FreeSans 448 0 0 0 FrameData[428]
port 364 nsew signal input
flabel metal3 s 0 6944 112 7056 0 FreeSans 448 0 0 0 FrameData[429]
port 365 nsew signal input
flabel metal3 s 0 683648 112 683760 0 FreeSans 448 0 0 0 FrameData[42]
port 366 nsew signal input
flabel metal3 s 0 7392 112 7504 0 FreeSans 448 0 0 0 FrameData[430]
port 367 nsew signal input
flabel metal3 s 0 7840 112 7952 0 FreeSans 448 0 0 0 FrameData[431]
port 368 nsew signal input
flabel metal3 s 0 8288 112 8400 0 FreeSans 448 0 0 0 FrameData[432]
port 369 nsew signal input
flabel metal3 s 0 8736 112 8848 0 FreeSans 448 0 0 0 FrameData[433]
port 370 nsew signal input
flabel metal3 s 0 9184 112 9296 0 FreeSans 448 0 0 0 FrameData[434]
port 371 nsew signal input
flabel metal3 s 0 9632 112 9744 0 FreeSans 448 0 0 0 FrameData[435]
port 372 nsew signal input
flabel metal3 s 0 10080 112 10192 0 FreeSans 448 0 0 0 FrameData[436]
port 373 nsew signal input
flabel metal3 s 0 10528 112 10640 0 FreeSans 448 0 0 0 FrameData[437]
port 374 nsew signal input
flabel metal3 s 0 10976 112 11088 0 FreeSans 448 0 0 0 FrameData[438]
port 375 nsew signal input
flabel metal3 s 0 11424 112 11536 0 FreeSans 448 0 0 0 FrameData[439]
port 376 nsew signal input
flabel metal3 s 0 684544 112 684656 0 FreeSans 448 0 0 0 FrameData[43]
port 377 nsew signal input
flabel metal3 s 0 11872 112 11984 0 FreeSans 448 0 0 0 FrameData[440]
port 378 nsew signal input
flabel metal3 s 0 12320 112 12432 0 FreeSans 448 0 0 0 FrameData[441]
port 379 nsew signal input
flabel metal3 s 0 12768 112 12880 0 FreeSans 448 0 0 0 FrameData[442]
port 380 nsew signal input
flabel metal3 s 0 13216 112 13328 0 FreeSans 448 0 0 0 FrameData[443]
port 381 nsew signal input
flabel metal3 s 0 13664 112 13776 0 FreeSans 448 0 0 0 FrameData[444]
port 382 nsew signal input
flabel metal3 s 0 14112 112 14224 0 FreeSans 448 0 0 0 FrameData[445]
port 383 nsew signal input
flabel metal3 s 0 14560 112 14672 0 FreeSans 448 0 0 0 FrameData[446]
port 384 nsew signal input
flabel metal3 s 0 15008 112 15120 0 FreeSans 448 0 0 0 FrameData[447]
port 385 nsew signal input
flabel metal3 s 0 685440 112 685552 0 FreeSans 448 0 0 0 FrameData[44]
port 386 nsew signal input
flabel metal3 s 0 686336 112 686448 0 FreeSans 448 0 0 0 FrameData[45]
port 387 nsew signal input
flabel metal3 s 0 687232 112 687344 0 FreeSans 448 0 0 0 FrameData[46]
port 388 nsew signal input
flabel metal3 s 0 688128 112 688240 0 FreeSans 448 0 0 0 FrameData[47]
port 389 nsew signal input
flabel metal3 s 0 689024 112 689136 0 FreeSans 448 0 0 0 FrameData[48]
port 390 nsew signal input
flabel metal3 s 0 689920 112 690032 0 FreeSans 448 0 0 0 FrameData[49]
port 391 nsew signal input
flabel metal3 s 0 706608 112 706720 0 FreeSans 448 0 0 0 FrameData[4]
port 392 nsew signal input
flabel metal3 s 0 690816 112 690928 0 FreeSans 448 0 0 0 FrameData[50]
port 393 nsew signal input
flabel metal3 s 0 691712 112 691824 0 FreeSans 448 0 0 0 FrameData[51]
port 394 nsew signal input
flabel metal3 s 0 692608 112 692720 0 FreeSans 448 0 0 0 FrameData[52]
port 395 nsew signal input
flabel metal3 s 0 693504 112 693616 0 FreeSans 448 0 0 0 FrameData[53]
port 396 nsew signal input
flabel metal3 s 0 694400 112 694512 0 FreeSans 448 0 0 0 FrameData[54]
port 397 nsew signal input
flabel metal3 s 0 695296 112 695408 0 FreeSans 448 0 0 0 FrameData[55]
port 398 nsew signal input
flabel metal3 s 0 696192 112 696304 0 FreeSans 448 0 0 0 FrameData[56]
port 399 nsew signal input
flabel metal3 s 0 697088 112 697200 0 FreeSans 448 0 0 0 FrameData[57]
port 400 nsew signal input
flabel metal3 s 0 697984 112 698096 0 FreeSans 448 0 0 0 FrameData[58]
port 401 nsew signal input
flabel metal3 s 0 698880 112 698992 0 FreeSans 448 0 0 0 FrameData[59]
port 402 nsew signal input
flabel metal3 s 0 707056 112 707168 0 FreeSans 448 0 0 0 FrameData[5]
port 403 nsew signal input
flabel metal3 s 0 699776 112 699888 0 FreeSans 448 0 0 0 FrameData[60]
port 404 nsew signal input
flabel metal3 s 0 700672 112 700784 0 FreeSans 448 0 0 0 FrameData[61]
port 405 nsew signal input
flabel metal3 s 0 701568 112 701680 0 FreeSans 448 0 0 0 FrameData[62]
port 406 nsew signal input
flabel metal3 s 0 702464 112 702576 0 FreeSans 448 0 0 0 FrameData[63]
port 407 nsew signal input
flabel metal3 s 0 617232 112 617344 0 FreeSans 448 0 0 0 FrameData[64]
port 408 nsew signal input
flabel metal3 s 0 618128 112 618240 0 FreeSans 448 0 0 0 FrameData[65]
port 409 nsew signal input
flabel metal3 s 0 619024 112 619136 0 FreeSans 448 0 0 0 FrameData[66]
port 410 nsew signal input
flabel metal3 s 0 619920 112 620032 0 FreeSans 448 0 0 0 FrameData[67]
port 411 nsew signal input
flabel metal3 s 0 620816 112 620928 0 FreeSans 448 0 0 0 FrameData[68]
port 412 nsew signal input
flabel metal3 s 0 621712 112 621824 0 FreeSans 448 0 0 0 FrameData[69]
port 413 nsew signal input
flabel metal3 s 0 707504 112 707616 0 FreeSans 448 0 0 0 FrameData[6]
port 414 nsew signal input
flabel metal3 s 0 622608 112 622720 0 FreeSans 448 0 0 0 FrameData[70]
port 415 nsew signal input
flabel metal3 s 0 623504 112 623616 0 FreeSans 448 0 0 0 FrameData[71]
port 416 nsew signal input
flabel metal3 s 0 624400 112 624512 0 FreeSans 448 0 0 0 FrameData[72]
port 417 nsew signal input
flabel metal3 s 0 625296 112 625408 0 FreeSans 448 0 0 0 FrameData[73]
port 418 nsew signal input
flabel metal3 s 0 626192 112 626304 0 FreeSans 448 0 0 0 FrameData[74]
port 419 nsew signal input
flabel metal3 s 0 627088 112 627200 0 FreeSans 448 0 0 0 FrameData[75]
port 420 nsew signal input
flabel metal3 s 0 627984 112 628096 0 FreeSans 448 0 0 0 FrameData[76]
port 421 nsew signal input
flabel metal3 s 0 628880 112 628992 0 FreeSans 448 0 0 0 FrameData[77]
port 422 nsew signal input
flabel metal3 s 0 629776 112 629888 0 FreeSans 448 0 0 0 FrameData[78]
port 423 nsew signal input
flabel metal3 s 0 630672 112 630784 0 FreeSans 448 0 0 0 FrameData[79]
port 424 nsew signal input
flabel metal3 s 0 707952 112 708064 0 FreeSans 448 0 0 0 FrameData[7]
port 425 nsew signal input
flabel metal3 s 0 631568 112 631680 0 FreeSans 448 0 0 0 FrameData[80]
port 426 nsew signal input
flabel metal3 s 0 632464 112 632576 0 FreeSans 448 0 0 0 FrameData[81]
port 427 nsew signal input
flabel metal3 s 0 633360 112 633472 0 FreeSans 448 0 0 0 FrameData[82]
port 428 nsew signal input
flabel metal3 s 0 634256 112 634368 0 FreeSans 448 0 0 0 FrameData[83]
port 429 nsew signal input
flabel metal3 s 0 635152 112 635264 0 FreeSans 448 0 0 0 FrameData[84]
port 430 nsew signal input
flabel metal3 s 0 636048 112 636160 0 FreeSans 448 0 0 0 FrameData[85]
port 431 nsew signal input
flabel metal3 s 0 636944 112 637056 0 FreeSans 448 0 0 0 FrameData[86]
port 432 nsew signal input
flabel metal3 s 0 637840 112 637952 0 FreeSans 448 0 0 0 FrameData[87]
port 433 nsew signal input
flabel metal3 s 0 638736 112 638848 0 FreeSans 448 0 0 0 FrameData[88]
port 434 nsew signal input
flabel metal3 s 0 639632 112 639744 0 FreeSans 448 0 0 0 FrameData[89]
port 435 nsew signal input
flabel metal3 s 0 708400 112 708512 0 FreeSans 448 0 0 0 FrameData[8]
port 436 nsew signal input
flabel metal3 s 0 640528 112 640640 0 FreeSans 448 0 0 0 FrameData[90]
port 437 nsew signal input
flabel metal3 s 0 641424 112 641536 0 FreeSans 448 0 0 0 FrameData[91]
port 438 nsew signal input
flabel metal3 s 0 642320 112 642432 0 FreeSans 448 0 0 0 FrameData[92]
port 439 nsew signal input
flabel metal3 s 0 643216 112 643328 0 FreeSans 448 0 0 0 FrameData[93]
port 440 nsew signal input
flabel metal3 s 0 644112 112 644224 0 FreeSans 448 0 0 0 FrameData[94]
port 441 nsew signal input
flabel metal3 s 0 645008 112 645120 0 FreeSans 448 0 0 0 FrameData[95]
port 442 nsew signal input
flabel metal3 s 0 559776 112 559888 0 FreeSans 448 0 0 0 FrameData[96]
port 443 nsew signal input
flabel metal3 s 0 560672 112 560784 0 FreeSans 448 0 0 0 FrameData[97]
port 444 nsew signal input
flabel metal3 s 0 561568 112 561680 0 FreeSans 448 0 0 0 FrameData[98]
port 445 nsew signal input
flabel metal3 s 0 562464 112 562576 0 FreeSans 448 0 0 0 FrameData[99]
port 446 nsew signal input
flabel metal3 s 0 708848 112 708960 0 FreeSans 448 0 0 0 FrameData[9]
port 447 nsew signal input
flabel metal2 s 2128 0 2240 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 448 nsew signal input
flabel metal2 s 269920 0 270032 112 0 FreeSans 448 0 0 0 FrameStrobe[100]
port 449 nsew signal input
flabel metal2 s 272608 0 272720 112 0 FreeSans 448 0 0 0 FrameStrobe[101]
port 450 nsew signal input
flabel metal2 s 275296 0 275408 112 0 FreeSans 448 0 0 0 FrameStrobe[102]
port 451 nsew signal input
flabel metal2 s 277984 0 278096 112 0 FreeSans 448 0 0 0 FrameStrobe[103]
port 452 nsew signal input
flabel metal2 s 280672 0 280784 112 0 FreeSans 448 0 0 0 FrameStrobe[104]
port 453 nsew signal input
flabel metal2 s 283360 0 283472 112 0 FreeSans 448 0 0 0 FrameStrobe[105]
port 454 nsew signal input
flabel metal2 s 286048 0 286160 112 0 FreeSans 448 0 0 0 FrameStrobe[106]
port 455 nsew signal input
flabel metal2 s 288736 0 288848 112 0 FreeSans 448 0 0 0 FrameStrobe[107]
port 456 nsew signal input
flabel metal2 s 291424 0 291536 112 0 FreeSans 448 0 0 0 FrameStrobe[108]
port 457 nsew signal input
flabel metal2 s 294112 0 294224 112 0 FreeSans 448 0 0 0 FrameStrobe[109]
port 458 nsew signal input
flabel metal2 s 15568 0 15680 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 459 nsew signal input
flabel metal2 s 296800 0 296912 112 0 FreeSans 448 0 0 0 FrameStrobe[110]
port 460 nsew signal input
flabel metal2 s 299488 0 299600 112 0 FreeSans 448 0 0 0 FrameStrobe[111]
port 461 nsew signal input
flabel metal2 s 302176 0 302288 112 0 FreeSans 448 0 0 0 FrameStrobe[112]
port 462 nsew signal input
flabel metal2 s 304864 0 304976 112 0 FreeSans 448 0 0 0 FrameStrobe[113]
port 463 nsew signal input
flabel metal2 s 307552 0 307664 112 0 FreeSans 448 0 0 0 FrameStrobe[114]
port 464 nsew signal input
flabel metal2 s 310240 0 310352 112 0 FreeSans 448 0 0 0 FrameStrobe[115]
port 465 nsew signal input
flabel metal2 s 312928 0 313040 112 0 FreeSans 448 0 0 0 FrameStrobe[116]
port 466 nsew signal input
flabel metal2 s 315616 0 315728 112 0 FreeSans 448 0 0 0 FrameStrobe[117]
port 467 nsew signal input
flabel metal2 s 318304 0 318416 112 0 FreeSans 448 0 0 0 FrameStrobe[118]
port 468 nsew signal input
flabel metal2 s 320992 0 321104 112 0 FreeSans 448 0 0 0 FrameStrobe[119]
port 469 nsew signal input
flabel metal2 s 16912 0 17024 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 470 nsew signal input
flabel metal2 s 326928 0 327040 112 0 FreeSans 448 0 0 0 FrameStrobe[120]
port 471 nsew signal input
flabel metal2 s 329392 0 329504 112 0 FreeSans 448 0 0 0 FrameStrobe[121]
port 472 nsew signal input
flabel metal2 s 331856 0 331968 112 0 FreeSans 448 0 0 0 FrameStrobe[122]
port 473 nsew signal input
flabel metal2 s 334320 0 334432 112 0 FreeSans 448 0 0 0 FrameStrobe[123]
port 474 nsew signal input
flabel metal2 s 336784 0 336896 112 0 FreeSans 448 0 0 0 FrameStrobe[124]
port 475 nsew signal input
flabel metal2 s 339248 0 339360 112 0 FreeSans 448 0 0 0 FrameStrobe[125]
port 476 nsew signal input
flabel metal2 s 341712 0 341824 112 0 FreeSans 448 0 0 0 FrameStrobe[126]
port 477 nsew signal input
flabel metal2 s 344176 0 344288 112 0 FreeSans 448 0 0 0 FrameStrobe[127]
port 478 nsew signal input
flabel metal2 s 346640 0 346752 112 0 FreeSans 448 0 0 0 FrameStrobe[128]
port 479 nsew signal input
flabel metal2 s 349104 0 349216 112 0 FreeSans 448 0 0 0 FrameStrobe[129]
port 480 nsew signal input
flabel metal2 s 18256 0 18368 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 481 nsew signal input
flabel metal2 s 351568 0 351680 112 0 FreeSans 448 0 0 0 FrameStrobe[130]
port 482 nsew signal input
flabel metal2 s 354032 0 354144 112 0 FreeSans 448 0 0 0 FrameStrobe[131]
port 483 nsew signal input
flabel metal2 s 356496 0 356608 112 0 FreeSans 448 0 0 0 FrameStrobe[132]
port 484 nsew signal input
flabel metal2 s 358960 0 359072 112 0 FreeSans 448 0 0 0 FrameStrobe[133]
port 485 nsew signal input
flabel metal2 s 361424 0 361536 112 0 FreeSans 448 0 0 0 FrameStrobe[134]
port 486 nsew signal input
flabel metal2 s 363888 0 364000 112 0 FreeSans 448 0 0 0 FrameStrobe[135]
port 487 nsew signal input
flabel metal2 s 366352 0 366464 112 0 FreeSans 448 0 0 0 FrameStrobe[136]
port 488 nsew signal input
flabel metal2 s 368816 0 368928 112 0 FreeSans 448 0 0 0 FrameStrobe[137]
port 489 nsew signal input
flabel metal2 s 371280 0 371392 112 0 FreeSans 448 0 0 0 FrameStrobe[138]
port 490 nsew signal input
flabel metal2 s 373744 0 373856 112 0 FreeSans 448 0 0 0 FrameStrobe[139]
port 491 nsew signal input
flabel metal2 s 19600 0 19712 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 492 nsew signal input
flabel metal2 s 380128 0 380240 112 0 FreeSans 448 0 0 0 FrameStrobe[140]
port 493 nsew signal input
flabel metal2 s 382816 0 382928 112 0 FreeSans 448 0 0 0 FrameStrobe[141]
port 494 nsew signal input
flabel metal2 s 385504 0 385616 112 0 FreeSans 448 0 0 0 FrameStrobe[142]
port 495 nsew signal input
flabel metal2 s 388192 0 388304 112 0 FreeSans 448 0 0 0 FrameStrobe[143]
port 496 nsew signal input
flabel metal2 s 390880 0 390992 112 0 FreeSans 448 0 0 0 FrameStrobe[144]
port 497 nsew signal input
flabel metal2 s 393568 0 393680 112 0 FreeSans 448 0 0 0 FrameStrobe[145]
port 498 nsew signal input
flabel metal2 s 396256 0 396368 112 0 FreeSans 448 0 0 0 FrameStrobe[146]
port 499 nsew signal input
flabel metal2 s 398944 0 399056 112 0 FreeSans 448 0 0 0 FrameStrobe[147]
port 500 nsew signal input
flabel metal2 s 401632 0 401744 112 0 FreeSans 448 0 0 0 FrameStrobe[148]
port 501 nsew signal input
flabel metal2 s 404320 0 404432 112 0 FreeSans 448 0 0 0 FrameStrobe[149]
port 502 nsew signal input
flabel metal2 s 20944 0 21056 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 503 nsew signal input
flabel metal2 s 407008 0 407120 112 0 FreeSans 448 0 0 0 FrameStrobe[150]
port 504 nsew signal input
flabel metal2 s 409696 0 409808 112 0 FreeSans 448 0 0 0 FrameStrobe[151]
port 505 nsew signal input
flabel metal2 s 412384 0 412496 112 0 FreeSans 448 0 0 0 FrameStrobe[152]
port 506 nsew signal input
flabel metal2 s 415072 0 415184 112 0 FreeSans 448 0 0 0 FrameStrobe[153]
port 507 nsew signal input
flabel metal2 s 417760 0 417872 112 0 FreeSans 448 0 0 0 FrameStrobe[154]
port 508 nsew signal input
flabel metal2 s 420448 0 420560 112 0 FreeSans 448 0 0 0 FrameStrobe[155]
port 509 nsew signal input
flabel metal2 s 423136 0 423248 112 0 FreeSans 448 0 0 0 FrameStrobe[156]
port 510 nsew signal input
flabel metal2 s 425824 0 425936 112 0 FreeSans 448 0 0 0 FrameStrobe[157]
port 511 nsew signal input
flabel metal2 s 428512 0 428624 112 0 FreeSans 448 0 0 0 FrameStrobe[158]
port 512 nsew signal input
flabel metal2 s 431200 0 431312 112 0 FreeSans 448 0 0 0 FrameStrobe[159]
port 513 nsew signal input
flabel metal2 s 22288 0 22400 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 514 nsew signal input
flabel metal2 s 436688 0 436800 112 0 FreeSans 448 0 0 0 FrameStrobe[160]
port 515 nsew signal input
flabel metal2 s 438032 0 438144 112 0 FreeSans 448 0 0 0 FrameStrobe[161]
port 516 nsew signal input
flabel metal2 s 439376 0 439488 112 0 FreeSans 448 0 0 0 FrameStrobe[162]
port 517 nsew signal input
flabel metal2 s 440720 0 440832 112 0 FreeSans 448 0 0 0 FrameStrobe[163]
port 518 nsew signal input
flabel metal2 s 442064 0 442176 112 0 FreeSans 448 0 0 0 FrameStrobe[164]
port 519 nsew signal input
flabel metal2 s 443408 0 443520 112 0 FreeSans 448 0 0 0 FrameStrobe[165]
port 520 nsew signal input
flabel metal2 s 444752 0 444864 112 0 FreeSans 448 0 0 0 FrameStrobe[166]
port 521 nsew signal input
flabel metal2 s 446096 0 446208 112 0 FreeSans 448 0 0 0 FrameStrobe[167]
port 522 nsew signal input
flabel metal2 s 448224 0 448336 112 0 FreeSans 448 0 0 0 FrameStrobe[168]
port 523 nsew signal input
flabel metal2 s 448784 0 448896 112 0 FreeSans 448 0 0 0 FrameStrobe[169]
port 524 nsew signal input
flabel metal2 s 23632 0 23744 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 525 nsew signal input
flabel metal2 s 450128 0 450240 112 0 FreeSans 448 0 0 0 FrameStrobe[170]
port 526 nsew signal input
flabel metal2 s 451472 0 451584 112 0 FreeSans 448 0 0 0 FrameStrobe[171]
port 527 nsew signal input
flabel metal2 s 452816 0 452928 112 0 FreeSans 448 0 0 0 FrameStrobe[172]
port 528 nsew signal input
flabel metal2 s 454160 0 454272 112 0 FreeSans 448 0 0 0 FrameStrobe[173]
port 529 nsew signal input
flabel metal2 s 455504 0 455616 112 0 FreeSans 448 0 0 0 FrameStrobe[174]
port 530 nsew signal input
flabel metal2 s 456848 0 456960 112 0 FreeSans 448 0 0 0 FrameStrobe[175]
port 531 nsew signal input
flabel metal2 s 458192 0 458304 112 0 FreeSans 448 0 0 0 FrameStrobe[176]
port 532 nsew signal input
flabel metal2 s 459536 0 459648 112 0 FreeSans 448 0 0 0 FrameStrobe[177]
port 533 nsew signal input
flabel metal2 s 460880 0 460992 112 0 FreeSans 448 0 0 0 FrameStrobe[178]
port 534 nsew signal input
flabel metal2 s 462224 0 462336 112 0 FreeSans 448 0 0 0 FrameStrobe[179]
port 535 nsew signal input
flabel metal2 s 24976 0 25088 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 536 nsew signal input
flabel metal2 s 26320 0 26432 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 537 nsew signal input
flabel metal2 s 27664 0 27776 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 538 nsew signal input
flabel metal2 s 3472 0 3584 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 539 nsew signal input
flabel metal2 s 46144 0 46256 112 0 FreeSans 448 0 0 0 FrameStrobe[20]
port 540 nsew signal input
flabel metal2 s 48160 0 48272 112 0 FreeSans 448 0 0 0 FrameStrobe[21]
port 541 nsew signal input
flabel metal2 s 50176 0 50288 112 0 FreeSans 448 0 0 0 FrameStrobe[22]
port 542 nsew signal input
flabel metal2 s 52192 0 52304 112 0 FreeSans 448 0 0 0 FrameStrobe[23]
port 543 nsew signal input
flabel metal2 s 54208 0 54320 112 0 FreeSans 448 0 0 0 FrameStrobe[24]
port 544 nsew signal input
flabel metal2 s 56224 0 56336 112 0 FreeSans 448 0 0 0 FrameStrobe[25]
port 545 nsew signal input
flabel metal2 s 58240 0 58352 112 0 FreeSans 448 0 0 0 FrameStrobe[26]
port 546 nsew signal input
flabel metal2 s 60256 0 60368 112 0 FreeSans 448 0 0 0 FrameStrobe[27]
port 547 nsew signal input
flabel metal2 s 62272 0 62384 112 0 FreeSans 448 0 0 0 FrameStrobe[28]
port 548 nsew signal input
flabel metal2 s 64288 0 64400 112 0 FreeSans 448 0 0 0 FrameStrobe[29]
port 549 nsew signal input
flabel metal2 s 4816 0 4928 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 550 nsew signal input
flabel metal2 s 66304 0 66416 112 0 FreeSans 448 0 0 0 FrameStrobe[30]
port 551 nsew signal input
flabel metal2 s 68320 0 68432 112 0 FreeSans 448 0 0 0 FrameStrobe[31]
port 552 nsew signal input
flabel metal2 s 70336 0 70448 112 0 FreeSans 448 0 0 0 FrameStrobe[32]
port 553 nsew signal input
flabel metal2 s 72352 0 72464 112 0 FreeSans 448 0 0 0 FrameStrobe[33]
port 554 nsew signal input
flabel metal2 s 74368 0 74480 112 0 FreeSans 448 0 0 0 FrameStrobe[34]
port 555 nsew signal input
flabel metal2 s 76384 0 76496 112 0 FreeSans 448 0 0 0 FrameStrobe[35]
port 556 nsew signal input
flabel metal2 s 78400 0 78512 112 0 FreeSans 448 0 0 0 FrameStrobe[36]
port 557 nsew signal input
flabel metal2 s 80416 0 80528 112 0 FreeSans 448 0 0 0 FrameStrobe[37]
port 558 nsew signal input
flabel metal2 s 82432 0 82544 112 0 FreeSans 448 0 0 0 FrameStrobe[38]
port 559 nsew signal input
flabel metal2 s 84448 0 84560 112 0 FreeSans 448 0 0 0 FrameStrobe[39]
port 560 nsew signal input
flabel metal2 s 6160 0 6272 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 561 nsew signal input
flabel metal2 s 90608 0 90720 112 0 FreeSans 448 0 0 0 FrameStrobe[40]
port 562 nsew signal input
flabel metal2 s 93296 0 93408 112 0 FreeSans 448 0 0 0 FrameStrobe[41]
port 563 nsew signal input
flabel metal2 s 95984 0 96096 112 0 FreeSans 448 0 0 0 FrameStrobe[42]
port 564 nsew signal input
flabel metal2 s 98672 0 98784 112 0 FreeSans 448 0 0 0 FrameStrobe[43]
port 565 nsew signal input
flabel metal2 s 101360 0 101472 112 0 FreeSans 448 0 0 0 FrameStrobe[44]
port 566 nsew signal input
flabel metal2 s 104048 0 104160 112 0 FreeSans 448 0 0 0 FrameStrobe[45]
port 567 nsew signal input
flabel metal2 s 106736 0 106848 112 0 FreeSans 448 0 0 0 FrameStrobe[46]
port 568 nsew signal input
flabel metal2 s 109424 0 109536 112 0 FreeSans 448 0 0 0 FrameStrobe[47]
port 569 nsew signal input
flabel metal2 s 112112 0 112224 112 0 FreeSans 448 0 0 0 FrameStrobe[48]
port 570 nsew signal input
flabel metal2 s 114800 0 114912 112 0 FreeSans 448 0 0 0 FrameStrobe[49]
port 571 nsew signal input
flabel metal2 s 7504 0 7616 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 572 nsew signal input
flabel metal2 s 117488 0 117600 112 0 FreeSans 448 0 0 0 FrameStrobe[50]
port 573 nsew signal input
flabel metal2 s 120176 0 120288 112 0 FreeSans 448 0 0 0 FrameStrobe[51]
port 574 nsew signal input
flabel metal2 s 122864 0 122976 112 0 FreeSans 448 0 0 0 FrameStrobe[52]
port 575 nsew signal input
flabel metal2 s 125552 0 125664 112 0 FreeSans 448 0 0 0 FrameStrobe[53]
port 576 nsew signal input
flabel metal2 s 128240 0 128352 112 0 FreeSans 448 0 0 0 FrameStrobe[54]
port 577 nsew signal input
flabel metal2 s 130928 0 131040 112 0 FreeSans 448 0 0 0 FrameStrobe[55]
port 578 nsew signal input
flabel metal2 s 133616 0 133728 112 0 FreeSans 448 0 0 0 FrameStrobe[56]
port 579 nsew signal input
flabel metal2 s 136304 0 136416 112 0 FreeSans 448 0 0 0 FrameStrobe[57]
port 580 nsew signal input
flabel metal2 s 138992 0 139104 112 0 FreeSans 448 0 0 0 FrameStrobe[58]
port 581 nsew signal input
flabel metal2 s 141680 0 141792 112 0 FreeSans 448 0 0 0 FrameStrobe[59]
port 582 nsew signal input
flabel metal2 s 8848 0 8960 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 583 nsew signal input
flabel metal2 s 148064 0 148176 112 0 FreeSans 448 0 0 0 FrameStrobe[60]
port 584 nsew signal input
flabel metal2 s 150752 0 150864 112 0 FreeSans 448 0 0 0 FrameStrobe[61]
port 585 nsew signal input
flabel metal2 s 153440 0 153552 112 0 FreeSans 448 0 0 0 FrameStrobe[62]
port 586 nsew signal input
flabel metal2 s 156128 0 156240 112 0 FreeSans 448 0 0 0 FrameStrobe[63]
port 587 nsew signal input
flabel metal2 s 158816 0 158928 112 0 FreeSans 448 0 0 0 FrameStrobe[64]
port 588 nsew signal input
flabel metal2 s 161504 0 161616 112 0 FreeSans 448 0 0 0 FrameStrobe[65]
port 589 nsew signal input
flabel metal2 s 164192 0 164304 112 0 FreeSans 448 0 0 0 FrameStrobe[66]
port 590 nsew signal input
flabel metal2 s 166880 0 166992 112 0 FreeSans 448 0 0 0 FrameStrobe[67]
port 591 nsew signal input
flabel metal2 s 169568 0 169680 112 0 FreeSans 448 0 0 0 FrameStrobe[68]
port 592 nsew signal input
flabel metal2 s 172256 0 172368 112 0 FreeSans 448 0 0 0 FrameStrobe[69]
port 593 nsew signal input
flabel metal2 s 10192 0 10304 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 594 nsew signal input
flabel metal2 s 174944 0 175056 112 0 FreeSans 448 0 0 0 FrameStrobe[70]
port 595 nsew signal input
flabel metal2 s 177632 0 177744 112 0 FreeSans 448 0 0 0 FrameStrobe[71]
port 596 nsew signal input
flabel metal2 s 180320 0 180432 112 0 FreeSans 448 0 0 0 FrameStrobe[72]
port 597 nsew signal input
flabel metal2 s 183008 0 183120 112 0 FreeSans 448 0 0 0 FrameStrobe[73]
port 598 nsew signal input
flabel metal2 s 185696 0 185808 112 0 FreeSans 448 0 0 0 FrameStrobe[74]
port 599 nsew signal input
flabel metal2 s 188384 0 188496 112 0 FreeSans 448 0 0 0 FrameStrobe[75]
port 600 nsew signal input
flabel metal2 s 191072 0 191184 112 0 FreeSans 448 0 0 0 FrameStrobe[76]
port 601 nsew signal input
flabel metal2 s 193760 0 193872 112 0 FreeSans 448 0 0 0 FrameStrobe[77]
port 602 nsew signal input
flabel metal2 s 196448 0 196560 112 0 FreeSans 448 0 0 0 FrameStrobe[78]
port 603 nsew signal input
flabel metal2 s 199136 0 199248 112 0 FreeSans 448 0 0 0 FrameStrobe[79]
port 604 nsew signal input
flabel metal2 s 11536 0 11648 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 605 nsew signal input
flabel metal2 s 206864 0 206976 112 0 FreeSans 448 0 0 0 FrameStrobe[80]
port 606 nsew signal input
flabel metal2 s 209776 0 209888 112 0 FreeSans 448 0 0 0 FrameStrobe[81]
port 607 nsew signal input
flabel metal2 s 212688 0 212800 112 0 FreeSans 448 0 0 0 FrameStrobe[82]
port 608 nsew signal input
flabel metal2 s 215600 0 215712 112 0 FreeSans 448 0 0 0 FrameStrobe[83]
port 609 nsew signal input
flabel metal2 s 218512 0 218624 112 0 FreeSans 448 0 0 0 FrameStrobe[84]
port 610 nsew signal input
flabel metal2 s 221424 0 221536 112 0 FreeSans 448 0 0 0 FrameStrobe[85]
port 611 nsew signal input
flabel metal2 s 224336 0 224448 112 0 FreeSans 448 0 0 0 FrameStrobe[86]
port 612 nsew signal input
flabel metal2 s 227248 0 227360 112 0 FreeSans 448 0 0 0 FrameStrobe[87]
port 613 nsew signal input
flabel metal2 s 230160 0 230272 112 0 FreeSans 448 0 0 0 FrameStrobe[88]
port 614 nsew signal input
flabel metal2 s 233072 0 233184 112 0 FreeSans 448 0 0 0 FrameStrobe[89]
port 615 nsew signal input
flabel metal2 s 12880 0 12992 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 616 nsew signal input
flabel metal2 s 235984 0 236096 112 0 FreeSans 448 0 0 0 FrameStrobe[90]
port 617 nsew signal input
flabel metal2 s 238896 0 239008 112 0 FreeSans 448 0 0 0 FrameStrobe[91]
port 618 nsew signal input
flabel metal2 s 241808 0 241920 112 0 FreeSans 448 0 0 0 FrameStrobe[92]
port 619 nsew signal input
flabel metal2 s 244720 0 244832 112 0 FreeSans 448 0 0 0 FrameStrobe[93]
port 620 nsew signal input
flabel metal2 s 247632 0 247744 112 0 FreeSans 448 0 0 0 FrameStrobe[94]
port 621 nsew signal input
flabel metal2 s 250544 0 250656 112 0 FreeSans 448 0 0 0 FrameStrobe[95]
port 622 nsew signal input
flabel metal2 s 253456 0 253568 112 0 FreeSans 448 0 0 0 FrameStrobe[96]
port 623 nsew signal input
flabel metal2 s 256368 0 256480 112 0 FreeSans 448 0 0 0 FrameStrobe[97]
port 624 nsew signal input
flabel metal2 s 259280 0 259392 112 0 FreeSans 448 0 0 0 FrameStrobe[98]
port 625 nsew signal input
flabel metal2 s 262192 0 262304 112 0 FreeSans 448 0 0 0 FrameStrobe[99]
port 626 nsew signal input
flabel metal2 s 14224 0 14336 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 627 nsew signal input
flabel metal3 s 0 133392 112 133504 0 FreeSans 448 0 0 0 Tile_X0Y10_A_I_top
port 628 nsew signal output
flabel metal3 s 0 132496 112 132608 0 FreeSans 448 0 0 0 Tile_X0Y10_A_O_top
port 629 nsew signal input
flabel metal3 s 0 134288 112 134400 0 FreeSans 448 0 0 0 Tile_X0Y10_A_T_top
port 630 nsew signal output
flabel metal3 s 0 143248 112 143360 0 FreeSans 448 0 0 0 Tile_X0Y10_A_config_C_bit0
port 631 nsew signal output
flabel metal3 s 0 144144 112 144256 0 FreeSans 448 0 0 0 Tile_X0Y10_A_config_C_bit1
port 632 nsew signal output
flabel metal3 s 0 145040 112 145152 0 FreeSans 448 0 0 0 Tile_X0Y10_A_config_C_bit2
port 633 nsew signal output
flabel metal3 s 0 145936 112 146048 0 FreeSans 448 0 0 0 Tile_X0Y10_A_config_C_bit3
port 634 nsew signal output
flabel metal3 s 0 136080 112 136192 0 FreeSans 448 0 0 0 Tile_X0Y10_B_I_top
port 635 nsew signal output
flabel metal3 s 0 135184 112 135296 0 FreeSans 448 0 0 0 Tile_X0Y10_B_O_top
port 636 nsew signal input
flabel metal3 s 0 136976 112 137088 0 FreeSans 448 0 0 0 Tile_X0Y10_B_T_top
port 637 nsew signal output
flabel metal3 s 0 146832 112 146944 0 FreeSans 448 0 0 0 Tile_X0Y10_B_config_C_bit0
port 638 nsew signal output
flabel metal3 s 0 147728 112 147840 0 FreeSans 448 0 0 0 Tile_X0Y10_B_config_C_bit1
port 639 nsew signal output
flabel metal3 s 0 148624 112 148736 0 FreeSans 448 0 0 0 Tile_X0Y10_B_config_C_bit2
port 640 nsew signal output
flabel metal3 s 0 149520 112 149632 0 FreeSans 448 0 0 0 Tile_X0Y10_B_config_C_bit3
port 641 nsew signal output
flabel metal3 s 0 138768 112 138880 0 FreeSans 448 0 0 0 Tile_X0Y10_C_I_top
port 642 nsew signal output
flabel metal3 s 0 137872 112 137984 0 FreeSans 448 0 0 0 Tile_X0Y10_C_O_top
port 643 nsew signal input
flabel metal3 s 0 139664 112 139776 0 FreeSans 448 0 0 0 Tile_X0Y10_C_T_top
port 644 nsew signal output
flabel metal3 s 0 150416 112 150528 0 FreeSans 448 0 0 0 Tile_X0Y10_C_config_C_bit0
port 645 nsew signal output
flabel metal3 s 0 151312 112 151424 0 FreeSans 448 0 0 0 Tile_X0Y10_C_config_C_bit1
port 646 nsew signal output
flabel metal3 s 0 152208 112 152320 0 FreeSans 448 0 0 0 Tile_X0Y10_C_config_C_bit2
port 647 nsew signal output
flabel metal3 s 0 153104 112 153216 0 FreeSans 448 0 0 0 Tile_X0Y10_C_config_C_bit3
port 648 nsew signal output
flabel metal3 s 0 141456 112 141568 0 FreeSans 448 0 0 0 Tile_X0Y10_D_I_top
port 649 nsew signal output
flabel metal3 s 0 140560 112 140672 0 FreeSans 448 0 0 0 Tile_X0Y10_D_O_top
port 650 nsew signal input
flabel metal3 s 0 142352 112 142464 0 FreeSans 448 0 0 0 Tile_X0Y10_D_T_top
port 651 nsew signal output
flabel metal3 s 0 154000 112 154112 0 FreeSans 448 0 0 0 Tile_X0Y10_D_config_C_bit0
port 652 nsew signal output
flabel metal3 s 0 154896 112 155008 0 FreeSans 448 0 0 0 Tile_X0Y10_D_config_C_bit1
port 653 nsew signal output
flabel metal3 s 0 155792 112 155904 0 FreeSans 448 0 0 0 Tile_X0Y10_D_config_C_bit2
port 654 nsew signal output
flabel metal3 s 0 156688 112 156800 0 FreeSans 448 0 0 0 Tile_X0Y10_D_config_C_bit3
port 655 nsew signal output
flabel metal3 s 0 75936 112 76048 0 FreeSans 448 0 0 0 Tile_X0Y11_A_I_top
port 656 nsew signal output
flabel metal3 s 0 75040 112 75152 0 FreeSans 448 0 0 0 Tile_X0Y11_A_O_top
port 657 nsew signal input
flabel metal3 s 0 76832 112 76944 0 FreeSans 448 0 0 0 Tile_X0Y11_A_T_top
port 658 nsew signal output
flabel metal3 s 0 85792 112 85904 0 FreeSans 448 0 0 0 Tile_X0Y11_A_config_C_bit0
port 659 nsew signal output
flabel metal3 s 0 86688 112 86800 0 FreeSans 448 0 0 0 Tile_X0Y11_A_config_C_bit1
port 660 nsew signal output
flabel metal3 s 0 87584 112 87696 0 FreeSans 448 0 0 0 Tile_X0Y11_A_config_C_bit2
port 661 nsew signal output
flabel metal3 s 0 88480 112 88592 0 FreeSans 448 0 0 0 Tile_X0Y11_A_config_C_bit3
port 662 nsew signal output
flabel metal3 s 0 78624 112 78736 0 FreeSans 448 0 0 0 Tile_X0Y11_B_I_top
port 663 nsew signal output
flabel metal3 s 0 77728 112 77840 0 FreeSans 448 0 0 0 Tile_X0Y11_B_O_top
port 664 nsew signal input
flabel metal3 s 0 79520 112 79632 0 FreeSans 448 0 0 0 Tile_X0Y11_B_T_top
port 665 nsew signal output
flabel metal3 s 0 89376 112 89488 0 FreeSans 448 0 0 0 Tile_X0Y11_B_config_C_bit0
port 666 nsew signal output
flabel metal3 s 0 90272 112 90384 0 FreeSans 448 0 0 0 Tile_X0Y11_B_config_C_bit1
port 667 nsew signal output
flabel metal3 s 0 91168 112 91280 0 FreeSans 448 0 0 0 Tile_X0Y11_B_config_C_bit2
port 668 nsew signal output
flabel metal3 s 0 92064 112 92176 0 FreeSans 448 0 0 0 Tile_X0Y11_B_config_C_bit3
port 669 nsew signal output
flabel metal3 s 0 81312 112 81424 0 FreeSans 448 0 0 0 Tile_X0Y11_C_I_top
port 670 nsew signal output
flabel metal3 s 0 80416 112 80528 0 FreeSans 448 0 0 0 Tile_X0Y11_C_O_top
port 671 nsew signal input
flabel metal3 s 0 82208 112 82320 0 FreeSans 448 0 0 0 Tile_X0Y11_C_T_top
port 672 nsew signal output
flabel metal3 s 0 92960 112 93072 0 FreeSans 448 0 0 0 Tile_X0Y11_C_config_C_bit0
port 673 nsew signal output
flabel metal3 s 0 93856 112 93968 0 FreeSans 448 0 0 0 Tile_X0Y11_C_config_C_bit1
port 674 nsew signal output
flabel metal3 s 0 94752 112 94864 0 FreeSans 448 0 0 0 Tile_X0Y11_C_config_C_bit2
port 675 nsew signal output
flabel metal3 s 0 95648 112 95760 0 FreeSans 448 0 0 0 Tile_X0Y11_C_config_C_bit3
port 676 nsew signal output
flabel metal3 s 0 84000 112 84112 0 FreeSans 448 0 0 0 Tile_X0Y11_D_I_top
port 677 nsew signal output
flabel metal3 s 0 83104 112 83216 0 FreeSans 448 0 0 0 Tile_X0Y11_D_O_top
port 678 nsew signal input
flabel metal3 s 0 84896 112 85008 0 FreeSans 448 0 0 0 Tile_X0Y11_D_T_top
port 679 nsew signal output
flabel metal3 s 0 96544 112 96656 0 FreeSans 448 0 0 0 Tile_X0Y11_D_config_C_bit0
port 680 nsew signal output
flabel metal3 s 0 97440 112 97552 0 FreeSans 448 0 0 0 Tile_X0Y11_D_config_C_bit1
port 681 nsew signal output
flabel metal3 s 0 98336 112 98448 0 FreeSans 448 0 0 0 Tile_X0Y11_D_config_C_bit2
port 682 nsew signal output
flabel metal3 s 0 99232 112 99344 0 FreeSans 448 0 0 0 Tile_X0Y11_D_config_C_bit3
port 683 nsew signal output
flabel metal3 s 0 18480 112 18592 0 FreeSans 448 0 0 0 Tile_X0Y12_A_I_top
port 684 nsew signal output
flabel metal3 s 0 17584 112 17696 0 FreeSans 448 0 0 0 Tile_X0Y12_A_O_top
port 685 nsew signal input
flabel metal3 s 0 19376 112 19488 0 FreeSans 448 0 0 0 Tile_X0Y12_A_T_top
port 686 nsew signal output
flabel metal3 s 0 28336 112 28448 0 FreeSans 448 0 0 0 Tile_X0Y12_A_config_C_bit0
port 687 nsew signal output
flabel metal3 s 0 29232 112 29344 0 FreeSans 448 0 0 0 Tile_X0Y12_A_config_C_bit1
port 688 nsew signal output
flabel metal3 s 0 30128 112 30240 0 FreeSans 448 0 0 0 Tile_X0Y12_A_config_C_bit2
port 689 nsew signal output
flabel metal3 s 0 31024 112 31136 0 FreeSans 448 0 0 0 Tile_X0Y12_A_config_C_bit3
port 690 nsew signal output
flabel metal3 s 0 21168 112 21280 0 FreeSans 448 0 0 0 Tile_X0Y12_B_I_top
port 691 nsew signal output
flabel metal3 s 0 20272 112 20384 0 FreeSans 448 0 0 0 Tile_X0Y12_B_O_top
port 692 nsew signal input
flabel metal3 s 0 22064 112 22176 0 FreeSans 448 0 0 0 Tile_X0Y12_B_T_top
port 693 nsew signal output
flabel metal3 s 0 31920 112 32032 0 FreeSans 448 0 0 0 Tile_X0Y12_B_config_C_bit0
port 694 nsew signal output
flabel metal3 s 0 32816 112 32928 0 FreeSans 448 0 0 0 Tile_X0Y12_B_config_C_bit1
port 695 nsew signal output
flabel metal3 s 0 33712 112 33824 0 FreeSans 448 0 0 0 Tile_X0Y12_B_config_C_bit2
port 696 nsew signal output
flabel metal3 s 0 34608 112 34720 0 FreeSans 448 0 0 0 Tile_X0Y12_B_config_C_bit3
port 697 nsew signal output
flabel metal3 s 0 23856 112 23968 0 FreeSans 448 0 0 0 Tile_X0Y12_C_I_top
port 698 nsew signal output
flabel metal3 s 0 22960 112 23072 0 FreeSans 448 0 0 0 Tile_X0Y12_C_O_top
port 699 nsew signal input
flabel metal3 s 0 24752 112 24864 0 FreeSans 448 0 0 0 Tile_X0Y12_C_T_top
port 700 nsew signal output
flabel metal3 s 0 35504 112 35616 0 FreeSans 448 0 0 0 Tile_X0Y12_C_config_C_bit0
port 701 nsew signal output
flabel metal3 s 0 36400 112 36512 0 FreeSans 448 0 0 0 Tile_X0Y12_C_config_C_bit1
port 702 nsew signal output
flabel metal3 s 0 37296 112 37408 0 FreeSans 448 0 0 0 Tile_X0Y12_C_config_C_bit2
port 703 nsew signal output
flabel metal3 s 0 38192 112 38304 0 FreeSans 448 0 0 0 Tile_X0Y12_C_config_C_bit3
port 704 nsew signal output
flabel metal3 s 0 26544 112 26656 0 FreeSans 448 0 0 0 Tile_X0Y12_D_I_top
port 705 nsew signal output
flabel metal3 s 0 25648 112 25760 0 FreeSans 448 0 0 0 Tile_X0Y12_D_O_top
port 706 nsew signal input
flabel metal3 s 0 27440 112 27552 0 FreeSans 448 0 0 0 Tile_X0Y12_D_T_top
port 707 nsew signal output
flabel metal3 s 0 39088 112 39200 0 FreeSans 448 0 0 0 Tile_X0Y12_D_config_C_bit0
port 708 nsew signal output
flabel metal3 s 0 39984 112 40096 0 FreeSans 448 0 0 0 Tile_X0Y12_D_config_C_bit1
port 709 nsew signal output
flabel metal3 s 0 40880 112 40992 0 FreeSans 448 0 0 0 Tile_X0Y12_D_config_C_bit2
port 710 nsew signal output
flabel metal3 s 0 41776 112 41888 0 FreeSans 448 0 0 0 Tile_X0Y12_D_config_C_bit3
port 711 nsew signal output
flabel metal3 s 0 650496 112 650608 0 FreeSans 448 0 0 0 Tile_X0Y1_A_I_top
port 712 nsew signal output
flabel metal3 s 0 649600 112 649712 0 FreeSans 448 0 0 0 Tile_X0Y1_A_O_top
port 713 nsew signal input
flabel metal3 s 0 651392 112 651504 0 FreeSans 448 0 0 0 Tile_X0Y1_A_T_top
port 714 nsew signal output
flabel metal3 s 0 660352 112 660464 0 FreeSans 448 0 0 0 Tile_X0Y1_A_config_C_bit0
port 715 nsew signal output
flabel metal3 s 0 661248 112 661360 0 FreeSans 448 0 0 0 Tile_X0Y1_A_config_C_bit1
port 716 nsew signal output
flabel metal3 s 0 662144 112 662256 0 FreeSans 448 0 0 0 Tile_X0Y1_A_config_C_bit2
port 717 nsew signal output
flabel metal3 s 0 663040 112 663152 0 FreeSans 448 0 0 0 Tile_X0Y1_A_config_C_bit3
port 718 nsew signal output
flabel metal3 s 0 653184 112 653296 0 FreeSans 448 0 0 0 Tile_X0Y1_B_I_top
port 719 nsew signal output
flabel metal3 s 0 652288 112 652400 0 FreeSans 448 0 0 0 Tile_X0Y1_B_O_top
port 720 nsew signal input
flabel metal3 s 0 654080 112 654192 0 FreeSans 448 0 0 0 Tile_X0Y1_B_T_top
port 721 nsew signal output
flabel metal3 s 0 663936 112 664048 0 FreeSans 448 0 0 0 Tile_X0Y1_B_config_C_bit0
port 722 nsew signal output
flabel metal3 s 0 664832 112 664944 0 FreeSans 448 0 0 0 Tile_X0Y1_B_config_C_bit1
port 723 nsew signal output
flabel metal3 s 0 665728 112 665840 0 FreeSans 448 0 0 0 Tile_X0Y1_B_config_C_bit2
port 724 nsew signal output
flabel metal3 s 0 666624 112 666736 0 FreeSans 448 0 0 0 Tile_X0Y1_B_config_C_bit3
port 725 nsew signal output
flabel metal3 s 0 655872 112 655984 0 FreeSans 448 0 0 0 Tile_X0Y1_C_I_top
port 726 nsew signal output
flabel metal3 s 0 654976 112 655088 0 FreeSans 448 0 0 0 Tile_X0Y1_C_O_top
port 727 nsew signal input
flabel metal3 s 0 656768 112 656880 0 FreeSans 448 0 0 0 Tile_X0Y1_C_T_top
port 728 nsew signal output
flabel metal3 s 0 667520 112 667632 0 FreeSans 448 0 0 0 Tile_X0Y1_C_config_C_bit0
port 729 nsew signal output
flabel metal3 s 0 668416 112 668528 0 FreeSans 448 0 0 0 Tile_X0Y1_C_config_C_bit1
port 730 nsew signal output
flabel metal3 s 0 669312 112 669424 0 FreeSans 448 0 0 0 Tile_X0Y1_C_config_C_bit2
port 731 nsew signal output
flabel metal3 s 0 670208 112 670320 0 FreeSans 448 0 0 0 Tile_X0Y1_C_config_C_bit3
port 732 nsew signal output
flabel metal3 s 0 658560 112 658672 0 FreeSans 448 0 0 0 Tile_X0Y1_D_I_top
port 733 nsew signal output
flabel metal3 s 0 657664 112 657776 0 FreeSans 448 0 0 0 Tile_X0Y1_D_O_top
port 734 nsew signal input
flabel metal3 s 0 659456 112 659568 0 FreeSans 448 0 0 0 Tile_X0Y1_D_T_top
port 735 nsew signal output
flabel metal3 s 0 671104 112 671216 0 FreeSans 448 0 0 0 Tile_X0Y1_D_config_C_bit0
port 736 nsew signal output
flabel metal3 s 0 672000 112 672112 0 FreeSans 448 0 0 0 Tile_X0Y1_D_config_C_bit1
port 737 nsew signal output
flabel metal3 s 0 672896 112 673008 0 FreeSans 448 0 0 0 Tile_X0Y1_D_config_C_bit2
port 738 nsew signal output
flabel metal3 s 0 673792 112 673904 0 FreeSans 448 0 0 0 Tile_X0Y1_D_config_C_bit3
port 739 nsew signal output
flabel metal3 s 0 593040 112 593152 0 FreeSans 448 0 0 0 Tile_X0Y2_A_I_top
port 740 nsew signal output
flabel metal3 s 0 592144 112 592256 0 FreeSans 448 0 0 0 Tile_X0Y2_A_O_top
port 741 nsew signal input
flabel metal3 s 0 593936 112 594048 0 FreeSans 448 0 0 0 Tile_X0Y2_A_T_top
port 742 nsew signal output
flabel metal3 s 0 602896 112 603008 0 FreeSans 448 0 0 0 Tile_X0Y2_A_config_C_bit0
port 743 nsew signal output
flabel metal3 s 0 603792 112 603904 0 FreeSans 448 0 0 0 Tile_X0Y2_A_config_C_bit1
port 744 nsew signal output
flabel metal3 s 0 604688 112 604800 0 FreeSans 448 0 0 0 Tile_X0Y2_A_config_C_bit2
port 745 nsew signal output
flabel metal3 s 0 605584 112 605696 0 FreeSans 448 0 0 0 Tile_X0Y2_A_config_C_bit3
port 746 nsew signal output
flabel metal3 s 0 595728 112 595840 0 FreeSans 448 0 0 0 Tile_X0Y2_B_I_top
port 747 nsew signal output
flabel metal3 s 0 594832 112 594944 0 FreeSans 448 0 0 0 Tile_X0Y2_B_O_top
port 748 nsew signal input
flabel metal3 s 0 596624 112 596736 0 FreeSans 448 0 0 0 Tile_X0Y2_B_T_top
port 749 nsew signal output
flabel metal3 s 0 606480 112 606592 0 FreeSans 448 0 0 0 Tile_X0Y2_B_config_C_bit0
port 750 nsew signal output
flabel metal3 s 0 607376 112 607488 0 FreeSans 448 0 0 0 Tile_X0Y2_B_config_C_bit1
port 751 nsew signal output
flabel metal3 s 0 608272 112 608384 0 FreeSans 448 0 0 0 Tile_X0Y2_B_config_C_bit2
port 752 nsew signal output
flabel metal3 s 0 609168 112 609280 0 FreeSans 448 0 0 0 Tile_X0Y2_B_config_C_bit3
port 753 nsew signal output
flabel metal3 s 0 598416 112 598528 0 FreeSans 448 0 0 0 Tile_X0Y2_C_I_top
port 754 nsew signal output
flabel metal3 s 0 597520 112 597632 0 FreeSans 448 0 0 0 Tile_X0Y2_C_O_top
port 755 nsew signal input
flabel metal3 s 0 599312 112 599424 0 FreeSans 448 0 0 0 Tile_X0Y2_C_T_top
port 756 nsew signal output
flabel metal3 s 0 610064 112 610176 0 FreeSans 448 0 0 0 Tile_X0Y2_C_config_C_bit0
port 757 nsew signal output
flabel metal3 s 0 610960 112 611072 0 FreeSans 448 0 0 0 Tile_X0Y2_C_config_C_bit1
port 758 nsew signal output
flabel metal3 s 0 611856 112 611968 0 FreeSans 448 0 0 0 Tile_X0Y2_C_config_C_bit2
port 759 nsew signal output
flabel metal3 s 0 612752 112 612864 0 FreeSans 448 0 0 0 Tile_X0Y2_C_config_C_bit3
port 760 nsew signal output
flabel metal3 s 0 601104 112 601216 0 FreeSans 448 0 0 0 Tile_X0Y2_D_I_top
port 761 nsew signal output
flabel metal3 s 0 600208 112 600320 0 FreeSans 448 0 0 0 Tile_X0Y2_D_O_top
port 762 nsew signal input
flabel metal3 s 0 602000 112 602112 0 FreeSans 448 0 0 0 Tile_X0Y2_D_T_top
port 763 nsew signal output
flabel metal3 s 0 613648 112 613760 0 FreeSans 448 0 0 0 Tile_X0Y2_D_config_C_bit0
port 764 nsew signal output
flabel metal3 s 0 614544 112 614656 0 FreeSans 448 0 0 0 Tile_X0Y2_D_config_C_bit1
port 765 nsew signal output
flabel metal3 s 0 615440 112 615552 0 FreeSans 448 0 0 0 Tile_X0Y2_D_config_C_bit2
port 766 nsew signal output
flabel metal3 s 0 616336 112 616448 0 FreeSans 448 0 0 0 Tile_X0Y2_D_config_C_bit3
port 767 nsew signal output
flabel metal3 s 0 535584 112 535696 0 FreeSans 448 0 0 0 Tile_X0Y3_A_I_top
port 768 nsew signal output
flabel metal3 s 0 534688 112 534800 0 FreeSans 448 0 0 0 Tile_X0Y3_A_O_top
port 769 nsew signal input
flabel metal3 s 0 536480 112 536592 0 FreeSans 448 0 0 0 Tile_X0Y3_A_T_top
port 770 nsew signal output
flabel metal3 s 0 545440 112 545552 0 FreeSans 448 0 0 0 Tile_X0Y3_A_config_C_bit0
port 771 nsew signal output
flabel metal3 s 0 546336 112 546448 0 FreeSans 448 0 0 0 Tile_X0Y3_A_config_C_bit1
port 772 nsew signal output
flabel metal3 s 0 547232 112 547344 0 FreeSans 448 0 0 0 Tile_X0Y3_A_config_C_bit2
port 773 nsew signal output
flabel metal3 s 0 548128 112 548240 0 FreeSans 448 0 0 0 Tile_X0Y3_A_config_C_bit3
port 774 nsew signal output
flabel metal3 s 0 538272 112 538384 0 FreeSans 448 0 0 0 Tile_X0Y3_B_I_top
port 775 nsew signal output
flabel metal3 s 0 537376 112 537488 0 FreeSans 448 0 0 0 Tile_X0Y3_B_O_top
port 776 nsew signal input
flabel metal3 s 0 539168 112 539280 0 FreeSans 448 0 0 0 Tile_X0Y3_B_T_top
port 777 nsew signal output
flabel metal3 s 0 549024 112 549136 0 FreeSans 448 0 0 0 Tile_X0Y3_B_config_C_bit0
port 778 nsew signal output
flabel metal3 s 0 549920 112 550032 0 FreeSans 448 0 0 0 Tile_X0Y3_B_config_C_bit1
port 779 nsew signal output
flabel metal3 s 0 550816 112 550928 0 FreeSans 448 0 0 0 Tile_X0Y3_B_config_C_bit2
port 780 nsew signal output
flabel metal3 s 0 551712 112 551824 0 FreeSans 448 0 0 0 Tile_X0Y3_B_config_C_bit3
port 781 nsew signal output
flabel metal3 s 0 540960 112 541072 0 FreeSans 448 0 0 0 Tile_X0Y3_C_I_top
port 782 nsew signal output
flabel metal3 s 0 540064 112 540176 0 FreeSans 448 0 0 0 Tile_X0Y3_C_O_top
port 783 nsew signal input
flabel metal3 s 0 541856 112 541968 0 FreeSans 448 0 0 0 Tile_X0Y3_C_T_top
port 784 nsew signal output
flabel metal3 s 0 552608 112 552720 0 FreeSans 448 0 0 0 Tile_X0Y3_C_config_C_bit0
port 785 nsew signal output
flabel metal3 s 0 553504 112 553616 0 FreeSans 448 0 0 0 Tile_X0Y3_C_config_C_bit1
port 786 nsew signal output
flabel metal3 s 0 554400 112 554512 0 FreeSans 448 0 0 0 Tile_X0Y3_C_config_C_bit2
port 787 nsew signal output
flabel metal3 s 0 555296 112 555408 0 FreeSans 448 0 0 0 Tile_X0Y3_C_config_C_bit3
port 788 nsew signal output
flabel metal3 s 0 543648 112 543760 0 FreeSans 448 0 0 0 Tile_X0Y3_D_I_top
port 789 nsew signal output
flabel metal3 s 0 542752 112 542864 0 FreeSans 448 0 0 0 Tile_X0Y3_D_O_top
port 790 nsew signal input
flabel metal3 s 0 544544 112 544656 0 FreeSans 448 0 0 0 Tile_X0Y3_D_T_top
port 791 nsew signal output
flabel metal3 s 0 556192 112 556304 0 FreeSans 448 0 0 0 Tile_X0Y3_D_config_C_bit0
port 792 nsew signal output
flabel metal3 s 0 557088 112 557200 0 FreeSans 448 0 0 0 Tile_X0Y3_D_config_C_bit1
port 793 nsew signal output
flabel metal3 s 0 557984 112 558096 0 FreeSans 448 0 0 0 Tile_X0Y3_D_config_C_bit2
port 794 nsew signal output
flabel metal3 s 0 558880 112 558992 0 FreeSans 448 0 0 0 Tile_X0Y3_D_config_C_bit3
port 795 nsew signal output
flabel metal3 s 0 478128 112 478240 0 FreeSans 448 0 0 0 Tile_X0Y4_A_I_top
port 796 nsew signal output
flabel metal3 s 0 477232 112 477344 0 FreeSans 448 0 0 0 Tile_X0Y4_A_O_top
port 797 nsew signal input
flabel metal3 s 0 479024 112 479136 0 FreeSans 448 0 0 0 Tile_X0Y4_A_T_top
port 798 nsew signal output
flabel metal3 s 0 487984 112 488096 0 FreeSans 448 0 0 0 Tile_X0Y4_A_config_C_bit0
port 799 nsew signal output
flabel metal3 s 0 488880 112 488992 0 FreeSans 448 0 0 0 Tile_X0Y4_A_config_C_bit1
port 800 nsew signal output
flabel metal3 s 0 489776 112 489888 0 FreeSans 448 0 0 0 Tile_X0Y4_A_config_C_bit2
port 801 nsew signal output
flabel metal3 s 0 490672 112 490784 0 FreeSans 448 0 0 0 Tile_X0Y4_A_config_C_bit3
port 802 nsew signal output
flabel metal3 s 0 480816 112 480928 0 FreeSans 448 0 0 0 Tile_X0Y4_B_I_top
port 803 nsew signal output
flabel metal3 s 0 479920 112 480032 0 FreeSans 448 0 0 0 Tile_X0Y4_B_O_top
port 804 nsew signal input
flabel metal3 s 0 481712 112 481824 0 FreeSans 448 0 0 0 Tile_X0Y4_B_T_top
port 805 nsew signal output
flabel metal3 s 0 491568 112 491680 0 FreeSans 448 0 0 0 Tile_X0Y4_B_config_C_bit0
port 806 nsew signal output
flabel metal3 s 0 492464 112 492576 0 FreeSans 448 0 0 0 Tile_X0Y4_B_config_C_bit1
port 807 nsew signal output
flabel metal3 s 0 493360 112 493472 0 FreeSans 448 0 0 0 Tile_X0Y4_B_config_C_bit2
port 808 nsew signal output
flabel metal3 s 0 494256 112 494368 0 FreeSans 448 0 0 0 Tile_X0Y4_B_config_C_bit3
port 809 nsew signal output
flabel metal3 s 0 483504 112 483616 0 FreeSans 448 0 0 0 Tile_X0Y4_C_I_top
port 810 nsew signal output
flabel metal3 s 0 482608 112 482720 0 FreeSans 448 0 0 0 Tile_X0Y4_C_O_top
port 811 nsew signal input
flabel metal3 s 0 484400 112 484512 0 FreeSans 448 0 0 0 Tile_X0Y4_C_T_top
port 812 nsew signal output
flabel metal3 s 0 495152 112 495264 0 FreeSans 448 0 0 0 Tile_X0Y4_C_config_C_bit0
port 813 nsew signal output
flabel metal3 s 0 496048 112 496160 0 FreeSans 448 0 0 0 Tile_X0Y4_C_config_C_bit1
port 814 nsew signal output
flabel metal3 s 0 496944 112 497056 0 FreeSans 448 0 0 0 Tile_X0Y4_C_config_C_bit2
port 815 nsew signal output
flabel metal3 s 0 497840 112 497952 0 FreeSans 448 0 0 0 Tile_X0Y4_C_config_C_bit3
port 816 nsew signal output
flabel metal3 s 0 486192 112 486304 0 FreeSans 448 0 0 0 Tile_X0Y4_D_I_top
port 817 nsew signal output
flabel metal3 s 0 485296 112 485408 0 FreeSans 448 0 0 0 Tile_X0Y4_D_O_top
port 818 nsew signal input
flabel metal3 s 0 487088 112 487200 0 FreeSans 448 0 0 0 Tile_X0Y4_D_T_top
port 819 nsew signal output
flabel metal3 s 0 498736 112 498848 0 FreeSans 448 0 0 0 Tile_X0Y4_D_config_C_bit0
port 820 nsew signal output
flabel metal3 s 0 499632 112 499744 0 FreeSans 448 0 0 0 Tile_X0Y4_D_config_C_bit1
port 821 nsew signal output
flabel metal3 s 0 500528 112 500640 0 FreeSans 448 0 0 0 Tile_X0Y4_D_config_C_bit2
port 822 nsew signal output
flabel metal3 s 0 501424 112 501536 0 FreeSans 448 0 0 0 Tile_X0Y4_D_config_C_bit3
port 823 nsew signal output
flabel metal3 s 0 420672 112 420784 0 FreeSans 448 0 0 0 Tile_X0Y5_A_I_top
port 824 nsew signal output
flabel metal3 s 0 419776 112 419888 0 FreeSans 448 0 0 0 Tile_X0Y5_A_O_top
port 825 nsew signal input
flabel metal3 s 0 421568 112 421680 0 FreeSans 448 0 0 0 Tile_X0Y5_A_T_top
port 826 nsew signal output
flabel metal3 s 0 430528 112 430640 0 FreeSans 448 0 0 0 Tile_X0Y5_A_config_C_bit0
port 827 nsew signal output
flabel metal3 s 0 431424 112 431536 0 FreeSans 448 0 0 0 Tile_X0Y5_A_config_C_bit1
port 828 nsew signal output
flabel metal3 s 0 432320 112 432432 0 FreeSans 448 0 0 0 Tile_X0Y5_A_config_C_bit2
port 829 nsew signal output
flabel metal3 s 0 433216 112 433328 0 FreeSans 448 0 0 0 Tile_X0Y5_A_config_C_bit3
port 830 nsew signal output
flabel metal3 s 0 423360 112 423472 0 FreeSans 448 0 0 0 Tile_X0Y5_B_I_top
port 831 nsew signal output
flabel metal3 s 0 422464 112 422576 0 FreeSans 448 0 0 0 Tile_X0Y5_B_O_top
port 832 nsew signal input
flabel metal3 s 0 424256 112 424368 0 FreeSans 448 0 0 0 Tile_X0Y5_B_T_top
port 833 nsew signal output
flabel metal3 s 0 434112 112 434224 0 FreeSans 448 0 0 0 Tile_X0Y5_B_config_C_bit0
port 834 nsew signal output
flabel metal3 s 0 435008 112 435120 0 FreeSans 448 0 0 0 Tile_X0Y5_B_config_C_bit1
port 835 nsew signal output
flabel metal3 s 0 435904 112 436016 0 FreeSans 448 0 0 0 Tile_X0Y5_B_config_C_bit2
port 836 nsew signal output
flabel metal3 s 0 436800 112 436912 0 FreeSans 448 0 0 0 Tile_X0Y5_B_config_C_bit3
port 837 nsew signal output
flabel metal3 s 0 426048 112 426160 0 FreeSans 448 0 0 0 Tile_X0Y5_C_I_top
port 838 nsew signal output
flabel metal3 s 0 425152 112 425264 0 FreeSans 448 0 0 0 Tile_X0Y5_C_O_top
port 839 nsew signal input
flabel metal3 s 0 426944 112 427056 0 FreeSans 448 0 0 0 Tile_X0Y5_C_T_top
port 840 nsew signal output
flabel metal3 s 0 437696 112 437808 0 FreeSans 448 0 0 0 Tile_X0Y5_C_config_C_bit0
port 841 nsew signal output
flabel metal3 s 0 438592 112 438704 0 FreeSans 448 0 0 0 Tile_X0Y5_C_config_C_bit1
port 842 nsew signal output
flabel metal3 s 0 439488 112 439600 0 FreeSans 448 0 0 0 Tile_X0Y5_C_config_C_bit2
port 843 nsew signal output
flabel metal3 s 0 440384 112 440496 0 FreeSans 448 0 0 0 Tile_X0Y5_C_config_C_bit3
port 844 nsew signal output
flabel metal3 s 0 428736 112 428848 0 FreeSans 448 0 0 0 Tile_X0Y5_D_I_top
port 845 nsew signal output
flabel metal3 s 0 427840 112 427952 0 FreeSans 448 0 0 0 Tile_X0Y5_D_O_top
port 846 nsew signal input
flabel metal3 s 0 429632 112 429744 0 FreeSans 448 0 0 0 Tile_X0Y5_D_T_top
port 847 nsew signal output
flabel metal3 s 0 441280 112 441392 0 FreeSans 448 0 0 0 Tile_X0Y5_D_config_C_bit0
port 848 nsew signal output
flabel metal3 s 0 442176 112 442288 0 FreeSans 448 0 0 0 Tile_X0Y5_D_config_C_bit1
port 849 nsew signal output
flabel metal3 s 0 443072 112 443184 0 FreeSans 448 0 0 0 Tile_X0Y5_D_config_C_bit2
port 850 nsew signal output
flabel metal3 s 0 443968 112 444080 0 FreeSans 448 0 0 0 Tile_X0Y5_D_config_C_bit3
port 851 nsew signal output
flabel metal3 s 0 363216 112 363328 0 FreeSans 448 0 0 0 Tile_X0Y6_A_I_top
port 852 nsew signal output
flabel metal3 s 0 362320 112 362432 0 FreeSans 448 0 0 0 Tile_X0Y6_A_O_top
port 853 nsew signal input
flabel metal3 s 0 364112 112 364224 0 FreeSans 448 0 0 0 Tile_X0Y6_A_T_top
port 854 nsew signal output
flabel metal3 s 0 373072 112 373184 0 FreeSans 448 0 0 0 Tile_X0Y6_A_config_C_bit0
port 855 nsew signal output
flabel metal3 s 0 373968 112 374080 0 FreeSans 448 0 0 0 Tile_X0Y6_A_config_C_bit1
port 856 nsew signal output
flabel metal3 s 0 374864 112 374976 0 FreeSans 448 0 0 0 Tile_X0Y6_A_config_C_bit2
port 857 nsew signal output
flabel metal3 s 0 375760 112 375872 0 FreeSans 448 0 0 0 Tile_X0Y6_A_config_C_bit3
port 858 nsew signal output
flabel metal3 s 0 365904 112 366016 0 FreeSans 448 0 0 0 Tile_X0Y6_B_I_top
port 859 nsew signal output
flabel metal3 s 0 365008 112 365120 0 FreeSans 448 0 0 0 Tile_X0Y6_B_O_top
port 860 nsew signal input
flabel metal3 s 0 366800 112 366912 0 FreeSans 448 0 0 0 Tile_X0Y6_B_T_top
port 861 nsew signal output
flabel metal3 s 0 376656 112 376768 0 FreeSans 448 0 0 0 Tile_X0Y6_B_config_C_bit0
port 862 nsew signal output
flabel metal3 s 0 377552 112 377664 0 FreeSans 448 0 0 0 Tile_X0Y6_B_config_C_bit1
port 863 nsew signal output
flabel metal3 s 0 378448 112 378560 0 FreeSans 448 0 0 0 Tile_X0Y6_B_config_C_bit2
port 864 nsew signal output
flabel metal3 s 0 379344 112 379456 0 FreeSans 448 0 0 0 Tile_X0Y6_B_config_C_bit3
port 865 nsew signal output
flabel metal3 s 0 368592 112 368704 0 FreeSans 448 0 0 0 Tile_X0Y6_C_I_top
port 866 nsew signal output
flabel metal3 s 0 367696 112 367808 0 FreeSans 448 0 0 0 Tile_X0Y6_C_O_top
port 867 nsew signal input
flabel metal3 s 0 369488 112 369600 0 FreeSans 448 0 0 0 Tile_X0Y6_C_T_top
port 868 nsew signal output
flabel metal3 s 0 380240 112 380352 0 FreeSans 448 0 0 0 Tile_X0Y6_C_config_C_bit0
port 869 nsew signal output
flabel metal3 s 0 381136 112 381248 0 FreeSans 448 0 0 0 Tile_X0Y6_C_config_C_bit1
port 870 nsew signal output
flabel metal3 s 0 382032 112 382144 0 FreeSans 448 0 0 0 Tile_X0Y6_C_config_C_bit2
port 871 nsew signal output
flabel metal3 s 0 382928 112 383040 0 FreeSans 448 0 0 0 Tile_X0Y6_C_config_C_bit3
port 872 nsew signal output
flabel metal3 s 0 371280 112 371392 0 FreeSans 448 0 0 0 Tile_X0Y6_D_I_top
port 873 nsew signal output
flabel metal3 s 0 370384 112 370496 0 FreeSans 448 0 0 0 Tile_X0Y6_D_O_top
port 874 nsew signal input
flabel metal3 s 0 372176 112 372288 0 FreeSans 448 0 0 0 Tile_X0Y6_D_T_top
port 875 nsew signal output
flabel metal3 s 0 383824 112 383936 0 FreeSans 448 0 0 0 Tile_X0Y6_D_config_C_bit0
port 876 nsew signal output
flabel metal3 s 0 384720 112 384832 0 FreeSans 448 0 0 0 Tile_X0Y6_D_config_C_bit1
port 877 nsew signal output
flabel metal3 s 0 385616 112 385728 0 FreeSans 448 0 0 0 Tile_X0Y6_D_config_C_bit2
port 878 nsew signal output
flabel metal3 s 0 386512 112 386624 0 FreeSans 448 0 0 0 Tile_X0Y6_D_config_C_bit3
port 879 nsew signal output
flabel metal3 s 0 305760 112 305872 0 FreeSans 448 0 0 0 Tile_X0Y7_A_I_top
port 880 nsew signal output
flabel metal3 s 0 304864 112 304976 0 FreeSans 448 0 0 0 Tile_X0Y7_A_O_top
port 881 nsew signal input
flabel metal3 s 0 306656 112 306768 0 FreeSans 448 0 0 0 Tile_X0Y7_A_T_top
port 882 nsew signal output
flabel metal3 s 0 315616 112 315728 0 FreeSans 448 0 0 0 Tile_X0Y7_A_config_C_bit0
port 883 nsew signal output
flabel metal3 s 0 316512 112 316624 0 FreeSans 448 0 0 0 Tile_X0Y7_A_config_C_bit1
port 884 nsew signal output
flabel metal3 s 0 317408 112 317520 0 FreeSans 448 0 0 0 Tile_X0Y7_A_config_C_bit2
port 885 nsew signal output
flabel metal3 s 0 318304 112 318416 0 FreeSans 448 0 0 0 Tile_X0Y7_A_config_C_bit3
port 886 nsew signal output
flabel metal3 s 0 308448 112 308560 0 FreeSans 448 0 0 0 Tile_X0Y7_B_I_top
port 887 nsew signal output
flabel metal3 s 0 307552 112 307664 0 FreeSans 448 0 0 0 Tile_X0Y7_B_O_top
port 888 nsew signal input
flabel metal3 s 0 309344 112 309456 0 FreeSans 448 0 0 0 Tile_X0Y7_B_T_top
port 889 nsew signal output
flabel metal3 s 0 319200 112 319312 0 FreeSans 448 0 0 0 Tile_X0Y7_B_config_C_bit0
port 890 nsew signal output
flabel metal3 s 0 320096 112 320208 0 FreeSans 448 0 0 0 Tile_X0Y7_B_config_C_bit1
port 891 nsew signal output
flabel metal3 s 0 320992 112 321104 0 FreeSans 448 0 0 0 Tile_X0Y7_B_config_C_bit2
port 892 nsew signal output
flabel metal3 s 0 321888 112 322000 0 FreeSans 448 0 0 0 Tile_X0Y7_B_config_C_bit3
port 893 nsew signal output
flabel metal3 s 0 311136 112 311248 0 FreeSans 448 0 0 0 Tile_X0Y7_C_I_top
port 894 nsew signal output
flabel metal3 s 0 310240 112 310352 0 FreeSans 448 0 0 0 Tile_X0Y7_C_O_top
port 895 nsew signal input
flabel metal3 s 0 312032 112 312144 0 FreeSans 448 0 0 0 Tile_X0Y7_C_T_top
port 896 nsew signal output
flabel metal3 s 0 322784 112 322896 0 FreeSans 448 0 0 0 Tile_X0Y7_C_config_C_bit0
port 897 nsew signal output
flabel metal3 s 0 323680 112 323792 0 FreeSans 448 0 0 0 Tile_X0Y7_C_config_C_bit1
port 898 nsew signal output
flabel metal3 s 0 324576 112 324688 0 FreeSans 448 0 0 0 Tile_X0Y7_C_config_C_bit2
port 899 nsew signal output
flabel metal3 s 0 325472 112 325584 0 FreeSans 448 0 0 0 Tile_X0Y7_C_config_C_bit3
port 900 nsew signal output
flabel metal3 s 0 313824 112 313936 0 FreeSans 448 0 0 0 Tile_X0Y7_D_I_top
port 901 nsew signal output
flabel metal3 s 0 312928 112 313040 0 FreeSans 448 0 0 0 Tile_X0Y7_D_O_top
port 902 nsew signal input
flabel metal3 s 0 314720 112 314832 0 FreeSans 448 0 0 0 Tile_X0Y7_D_T_top
port 903 nsew signal output
flabel metal3 s 0 326368 112 326480 0 FreeSans 448 0 0 0 Tile_X0Y7_D_config_C_bit0
port 904 nsew signal output
flabel metal3 s 0 327264 112 327376 0 FreeSans 448 0 0 0 Tile_X0Y7_D_config_C_bit1
port 905 nsew signal output
flabel metal3 s 0 328160 112 328272 0 FreeSans 448 0 0 0 Tile_X0Y7_D_config_C_bit2
port 906 nsew signal output
flabel metal3 s 0 329056 112 329168 0 FreeSans 448 0 0 0 Tile_X0Y7_D_config_C_bit3
port 907 nsew signal output
flabel metal3 s 0 248304 112 248416 0 FreeSans 448 0 0 0 Tile_X0Y8_A_I_top
port 908 nsew signal output
flabel metal3 s 0 247408 112 247520 0 FreeSans 448 0 0 0 Tile_X0Y8_A_O_top
port 909 nsew signal input
flabel metal3 s 0 249200 112 249312 0 FreeSans 448 0 0 0 Tile_X0Y8_A_T_top
port 910 nsew signal output
flabel metal3 s 0 258160 112 258272 0 FreeSans 448 0 0 0 Tile_X0Y8_A_config_C_bit0
port 911 nsew signal output
flabel metal3 s 0 259056 112 259168 0 FreeSans 448 0 0 0 Tile_X0Y8_A_config_C_bit1
port 912 nsew signal output
flabel metal3 s 0 259952 112 260064 0 FreeSans 448 0 0 0 Tile_X0Y8_A_config_C_bit2
port 913 nsew signal output
flabel metal3 s 0 260848 112 260960 0 FreeSans 448 0 0 0 Tile_X0Y8_A_config_C_bit3
port 914 nsew signal output
flabel metal3 s 0 250992 112 251104 0 FreeSans 448 0 0 0 Tile_X0Y8_B_I_top
port 915 nsew signal output
flabel metal3 s 0 250096 112 250208 0 FreeSans 448 0 0 0 Tile_X0Y8_B_O_top
port 916 nsew signal input
flabel metal3 s 0 251888 112 252000 0 FreeSans 448 0 0 0 Tile_X0Y8_B_T_top
port 917 nsew signal output
flabel metal3 s 0 261744 112 261856 0 FreeSans 448 0 0 0 Tile_X0Y8_B_config_C_bit0
port 918 nsew signal output
flabel metal3 s 0 262640 112 262752 0 FreeSans 448 0 0 0 Tile_X0Y8_B_config_C_bit1
port 919 nsew signal output
flabel metal3 s 0 263536 112 263648 0 FreeSans 448 0 0 0 Tile_X0Y8_B_config_C_bit2
port 920 nsew signal output
flabel metal3 s 0 264432 112 264544 0 FreeSans 448 0 0 0 Tile_X0Y8_B_config_C_bit3
port 921 nsew signal output
flabel metal3 s 0 253680 112 253792 0 FreeSans 448 0 0 0 Tile_X0Y8_C_I_top
port 922 nsew signal output
flabel metal3 s 0 252784 112 252896 0 FreeSans 448 0 0 0 Tile_X0Y8_C_O_top
port 923 nsew signal input
flabel metal3 s 0 254576 112 254688 0 FreeSans 448 0 0 0 Tile_X0Y8_C_T_top
port 924 nsew signal output
flabel metal3 s 0 265328 112 265440 0 FreeSans 448 0 0 0 Tile_X0Y8_C_config_C_bit0
port 925 nsew signal output
flabel metal3 s 0 266224 112 266336 0 FreeSans 448 0 0 0 Tile_X0Y8_C_config_C_bit1
port 926 nsew signal output
flabel metal3 s 0 267120 112 267232 0 FreeSans 448 0 0 0 Tile_X0Y8_C_config_C_bit2
port 927 nsew signal output
flabel metal3 s 0 268016 112 268128 0 FreeSans 448 0 0 0 Tile_X0Y8_C_config_C_bit3
port 928 nsew signal output
flabel metal3 s 0 256368 112 256480 0 FreeSans 448 0 0 0 Tile_X0Y8_D_I_top
port 929 nsew signal output
flabel metal3 s 0 255472 112 255584 0 FreeSans 448 0 0 0 Tile_X0Y8_D_O_top
port 930 nsew signal input
flabel metal3 s 0 257264 112 257376 0 FreeSans 448 0 0 0 Tile_X0Y8_D_T_top
port 931 nsew signal output
flabel metal3 s 0 268912 112 269024 0 FreeSans 448 0 0 0 Tile_X0Y8_D_config_C_bit0
port 932 nsew signal output
flabel metal3 s 0 269808 112 269920 0 FreeSans 448 0 0 0 Tile_X0Y8_D_config_C_bit1
port 933 nsew signal output
flabel metal3 s 0 270704 112 270816 0 FreeSans 448 0 0 0 Tile_X0Y8_D_config_C_bit2
port 934 nsew signal output
flabel metal3 s 0 271600 112 271712 0 FreeSans 448 0 0 0 Tile_X0Y8_D_config_C_bit3
port 935 nsew signal output
flabel metal3 s 0 190848 112 190960 0 FreeSans 448 0 0 0 Tile_X0Y9_A_I_top
port 936 nsew signal output
flabel metal3 s 0 189952 112 190064 0 FreeSans 448 0 0 0 Tile_X0Y9_A_O_top
port 937 nsew signal input
flabel metal3 s 0 191744 112 191856 0 FreeSans 448 0 0 0 Tile_X0Y9_A_T_top
port 938 nsew signal output
flabel metal3 s 0 200704 112 200816 0 FreeSans 448 0 0 0 Tile_X0Y9_A_config_C_bit0
port 939 nsew signal output
flabel metal3 s 0 201600 112 201712 0 FreeSans 448 0 0 0 Tile_X0Y9_A_config_C_bit1
port 940 nsew signal output
flabel metal3 s 0 202496 112 202608 0 FreeSans 448 0 0 0 Tile_X0Y9_A_config_C_bit2
port 941 nsew signal output
flabel metal3 s 0 203392 112 203504 0 FreeSans 448 0 0 0 Tile_X0Y9_A_config_C_bit3
port 942 nsew signal output
flabel metal3 s 0 193536 112 193648 0 FreeSans 448 0 0 0 Tile_X0Y9_B_I_top
port 943 nsew signal output
flabel metal3 s 0 192640 112 192752 0 FreeSans 448 0 0 0 Tile_X0Y9_B_O_top
port 944 nsew signal input
flabel metal3 s 0 194432 112 194544 0 FreeSans 448 0 0 0 Tile_X0Y9_B_T_top
port 945 nsew signal output
flabel metal3 s 0 204288 112 204400 0 FreeSans 448 0 0 0 Tile_X0Y9_B_config_C_bit0
port 946 nsew signal output
flabel metal3 s 0 205184 112 205296 0 FreeSans 448 0 0 0 Tile_X0Y9_B_config_C_bit1
port 947 nsew signal output
flabel metal3 s 0 206080 112 206192 0 FreeSans 448 0 0 0 Tile_X0Y9_B_config_C_bit2
port 948 nsew signal output
flabel metal3 s 0 206976 112 207088 0 FreeSans 448 0 0 0 Tile_X0Y9_B_config_C_bit3
port 949 nsew signal output
flabel metal3 s 0 196224 112 196336 0 FreeSans 448 0 0 0 Tile_X0Y9_C_I_top
port 950 nsew signal output
flabel metal3 s 0 195328 112 195440 0 FreeSans 448 0 0 0 Tile_X0Y9_C_O_top
port 951 nsew signal input
flabel metal3 s 0 197120 112 197232 0 FreeSans 448 0 0 0 Tile_X0Y9_C_T_top
port 952 nsew signal output
flabel metal3 s 0 207872 112 207984 0 FreeSans 448 0 0 0 Tile_X0Y9_C_config_C_bit0
port 953 nsew signal output
flabel metal3 s 0 208768 112 208880 0 FreeSans 448 0 0 0 Tile_X0Y9_C_config_C_bit1
port 954 nsew signal output
flabel metal3 s 0 209664 112 209776 0 FreeSans 448 0 0 0 Tile_X0Y9_C_config_C_bit2
port 955 nsew signal output
flabel metal3 s 0 210560 112 210672 0 FreeSans 448 0 0 0 Tile_X0Y9_C_config_C_bit3
port 956 nsew signal output
flabel metal3 s 0 198912 112 199024 0 FreeSans 448 0 0 0 Tile_X0Y9_D_I_top
port 957 nsew signal output
flabel metal3 s 0 198016 112 198128 0 FreeSans 448 0 0 0 Tile_X0Y9_D_O_top
port 958 nsew signal input
flabel metal3 s 0 199808 112 199920 0 FreeSans 448 0 0 0 Tile_X0Y9_D_T_top
port 959 nsew signal output
flabel metal3 s 0 211456 112 211568 0 FreeSans 448 0 0 0 Tile_X0Y9_D_config_C_bit0
port 960 nsew signal output
flabel metal3 s 0 212352 112 212464 0 FreeSans 448 0 0 0 Tile_X0Y9_D_config_C_bit1
port 961 nsew signal output
flabel metal3 s 0 213248 112 213360 0 FreeSans 448 0 0 0 Tile_X0Y9_D_config_C_bit2
port 962 nsew signal output
flabel metal3 s 0 214144 112 214256 0 FreeSans 448 0 0 0 Tile_X0Y9_D_config_C_bit3
port 963 nsew signal output
flabel metal2 s 42112 0 42224 112 0 FreeSans 448 0 0 0 Tile_X1Y13_BOOT_top
port 964 nsew signal output
flabel metal2 s 32032 0 32144 112 0 FreeSans 448 0 0 0 Tile_X1Y13_CONFIGURED_top
port 965 nsew signal input
flabel metal2 s 30016 0 30128 112 0 FreeSans 448 0 0 0 Tile_X1Y13_RESET_top
port 966 nsew signal input
flabel metal2 s 34048 0 34160 112 0 FreeSans 448 0 0 0 Tile_X1Y13_SLOT_top0
port 967 nsew signal output
flabel metal2 s 36064 0 36176 112 0 FreeSans 448 0 0 0 Tile_X1Y13_SLOT_top1
port 968 nsew signal output
flabel metal2 s 38080 0 38192 112 0 FreeSans 448 0 0 0 Tile_X1Y13_SLOT_top2
port 969 nsew signal output
flabel metal2 s 40096 0 40208 112 0 FreeSans 448 0 0 0 Tile_X1Y13_SLOT_top3
port 970 nsew signal output
flabel metal3 s 464800 150192 464912 150304 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM0
port 971 nsew signal output
flabel metal3 s 464800 151088 464912 151200 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM1
port 972 nsew signal output
flabel metal3 s 464800 151984 464912 152096 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM2
port 973 nsew signal output
flabel metal3 s 464800 152880 464912 152992 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM3
port 974 nsew signal output
flabel metal3 s 464800 153776 464912 153888 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM4
port 975 nsew signal output
flabel metal3 s 464800 154672 464912 154784 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM5
port 976 nsew signal output
flabel metal3 s 464800 155568 464912 155680 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM6
port 977 nsew signal output
flabel metal3 s 464800 156464 464912 156576 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM7
port 978 nsew signal output
flabel metal3 s 464800 157360 464912 157472 0 FreeSans 448 0 0 0 Tile_X8Y10_A_SRAM8
port 979 nsew signal output
flabel metal3 s 464800 141232 464912 141344 0 FreeSans 448 0 0 0 Tile_X8Y10_CEN_SRAM
port 980 nsew signal output
flabel metal3 s 464800 165424 464912 165536 0 FreeSans 448 0 0 0 Tile_X8Y10_CLK_SRAM
port 981 nsew signal output
flabel metal3 s 464800 140336 464912 140448 0 FreeSans 448 0 0 0 Tile_X8Y10_CONFIGURED_top
port 982 nsew signal input
flabel metal3 s 464800 158256 464912 158368 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM0
port 983 nsew signal output
flabel metal3 s 464800 159152 464912 159264 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM1
port 984 nsew signal output
flabel metal3 s 464800 160048 464912 160160 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM2
port 985 nsew signal output
flabel metal3 s 464800 160944 464912 161056 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM3
port 986 nsew signal output
flabel metal3 s 464800 161840 464912 161952 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM4
port 987 nsew signal output
flabel metal3 s 464800 162736 464912 162848 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM5
port 988 nsew signal output
flabel metal3 s 464800 163632 464912 163744 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM6
port 989 nsew signal output
flabel metal3 s 464800 164528 464912 164640 0 FreeSans 448 0 0 0 Tile_X8Y10_D_SRAM7
port 990 nsew signal output
flabel metal3 s 464800 142128 464912 142240 0 FreeSans 448 0 0 0 Tile_X8Y10_GWEN_SRAM
port 991 nsew signal output
flabel metal3 s 464800 133168 464912 133280 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM0
port 992 nsew signal input
flabel metal3 s 464800 134064 464912 134176 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM1
port 993 nsew signal input
flabel metal3 s 464800 134960 464912 135072 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM2
port 994 nsew signal input
flabel metal3 s 464800 135856 464912 135968 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM3
port 995 nsew signal input
flabel metal3 s 464800 136752 464912 136864 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM4
port 996 nsew signal input
flabel metal3 s 464800 137648 464912 137760 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM5
port 997 nsew signal input
flabel metal3 s 464800 138544 464912 138656 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM6
port 998 nsew signal input
flabel metal3 s 464800 139440 464912 139552 0 FreeSans 448 0 0 0 Tile_X8Y10_Q_SRAM7
port 999 nsew signal input
flabel metal3 s 464800 143024 464912 143136 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM0
port 1000 nsew signal output
flabel metal3 s 464800 143920 464912 144032 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM1
port 1001 nsew signal output
flabel metal3 s 464800 144816 464912 144928 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM2
port 1002 nsew signal output
flabel metal3 s 464800 145712 464912 145824 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM3
port 1003 nsew signal output
flabel metal3 s 464800 146608 464912 146720 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM4
port 1004 nsew signal output
flabel metal3 s 464800 147504 464912 147616 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM5
port 1005 nsew signal output
flabel metal3 s 464800 148400 464912 148512 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM6
port 1006 nsew signal output
flabel metal3 s 464800 149296 464912 149408 0 FreeSans 448 0 0 0 Tile_X8Y10_WEN_SRAM7
port 1007 nsew signal output
flabel metal3 s 464800 35280 464912 35392 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM0
port 1008 nsew signal output
flabel metal3 s 464800 36176 464912 36288 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM1
port 1009 nsew signal output
flabel metal3 s 464800 37072 464912 37184 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM2
port 1010 nsew signal output
flabel metal3 s 464800 37968 464912 38080 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM3
port 1011 nsew signal output
flabel metal3 s 464800 38864 464912 38976 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM4
port 1012 nsew signal output
flabel metal3 s 464800 39760 464912 39872 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM5
port 1013 nsew signal output
flabel metal3 s 464800 40656 464912 40768 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM6
port 1014 nsew signal output
flabel metal3 s 464800 41552 464912 41664 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM7
port 1015 nsew signal output
flabel metal3 s 464800 42448 464912 42560 0 FreeSans 448 0 0 0 Tile_X8Y12_A_SRAM8
port 1016 nsew signal output
flabel metal3 s 464800 26320 464912 26432 0 FreeSans 448 0 0 0 Tile_X8Y12_CEN_SRAM
port 1017 nsew signal output
flabel metal3 s 464800 50512 464912 50624 0 FreeSans 448 0 0 0 Tile_X8Y12_CLK_SRAM
port 1018 nsew signal output
flabel metal3 s 464800 25424 464912 25536 0 FreeSans 448 0 0 0 Tile_X8Y12_CONFIGURED_top
port 1019 nsew signal input
flabel metal3 s 464800 43344 464912 43456 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM0
port 1020 nsew signal output
flabel metal3 s 464800 44240 464912 44352 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM1
port 1021 nsew signal output
flabel metal3 s 464800 45136 464912 45248 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM2
port 1022 nsew signal output
flabel metal3 s 464800 46032 464912 46144 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM3
port 1023 nsew signal output
flabel metal3 s 464800 46928 464912 47040 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM4
port 1024 nsew signal output
flabel metal3 s 464800 47824 464912 47936 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM5
port 1025 nsew signal output
flabel metal3 s 464800 48720 464912 48832 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM6
port 1026 nsew signal output
flabel metal3 s 464800 49616 464912 49728 0 FreeSans 448 0 0 0 Tile_X8Y12_D_SRAM7
port 1027 nsew signal output
flabel metal3 s 464800 27216 464912 27328 0 FreeSans 448 0 0 0 Tile_X8Y12_GWEN_SRAM
port 1028 nsew signal output
flabel metal3 s 464800 18256 464912 18368 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM0
port 1029 nsew signal input
flabel metal3 s 464800 19152 464912 19264 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM1
port 1030 nsew signal input
flabel metal3 s 464800 20048 464912 20160 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM2
port 1031 nsew signal input
flabel metal3 s 464800 20944 464912 21056 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM3
port 1032 nsew signal input
flabel metal3 s 464800 21840 464912 21952 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM4
port 1033 nsew signal input
flabel metal3 s 464800 22736 464912 22848 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM5
port 1034 nsew signal input
flabel metal3 s 464800 23632 464912 23744 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM6
port 1035 nsew signal input
flabel metal3 s 464800 24528 464912 24640 0 FreeSans 448 0 0 0 Tile_X8Y12_Q_SRAM7
port 1036 nsew signal input
flabel metal3 s 464800 28112 464912 28224 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM0
port 1037 nsew signal output
flabel metal3 s 464800 29008 464912 29120 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM1
port 1038 nsew signal output
flabel metal3 s 464800 29904 464912 30016 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM2
port 1039 nsew signal output
flabel metal3 s 464800 30800 464912 30912 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM3
port 1040 nsew signal output
flabel metal3 s 464800 31696 464912 31808 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM4
port 1041 nsew signal output
flabel metal3 s 464800 32592 464912 32704 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM5
port 1042 nsew signal output
flabel metal3 s 464800 33488 464912 33600 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM6
port 1043 nsew signal output
flabel metal3 s 464800 34384 464912 34496 0 FreeSans 448 0 0 0 Tile_X8Y12_WEN_SRAM7
port 1044 nsew signal output
flabel metal3 s 464800 609840 464912 609952 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM0
port 1045 nsew signal output
flabel metal3 s 464800 610736 464912 610848 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM1
port 1046 nsew signal output
flabel metal3 s 464800 611632 464912 611744 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM2
port 1047 nsew signal output
flabel metal3 s 464800 612528 464912 612640 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM3
port 1048 nsew signal output
flabel metal3 s 464800 613424 464912 613536 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM4
port 1049 nsew signal output
flabel metal3 s 464800 614320 464912 614432 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM5
port 1050 nsew signal output
flabel metal3 s 464800 615216 464912 615328 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM6
port 1051 nsew signal output
flabel metal3 s 464800 616112 464912 616224 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM7
port 1052 nsew signal output
flabel metal3 s 464800 617008 464912 617120 0 FreeSans 448 0 0 0 Tile_X8Y2_A_SRAM8
port 1053 nsew signal output
flabel metal3 s 464800 600880 464912 600992 0 FreeSans 448 0 0 0 Tile_X8Y2_CEN_SRAM
port 1054 nsew signal output
flabel metal3 s 464800 625072 464912 625184 0 FreeSans 448 0 0 0 Tile_X8Y2_CLK_SRAM
port 1055 nsew signal output
flabel metal3 s 464800 599984 464912 600096 0 FreeSans 448 0 0 0 Tile_X8Y2_CONFIGURED_top
port 1056 nsew signal input
flabel metal3 s 464800 617904 464912 618016 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM0
port 1057 nsew signal output
flabel metal3 s 464800 618800 464912 618912 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM1
port 1058 nsew signal output
flabel metal3 s 464800 619696 464912 619808 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM2
port 1059 nsew signal output
flabel metal3 s 464800 620592 464912 620704 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM3
port 1060 nsew signal output
flabel metal3 s 464800 621488 464912 621600 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM4
port 1061 nsew signal output
flabel metal3 s 464800 622384 464912 622496 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM5
port 1062 nsew signal output
flabel metal3 s 464800 623280 464912 623392 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM6
port 1063 nsew signal output
flabel metal3 s 464800 624176 464912 624288 0 FreeSans 448 0 0 0 Tile_X8Y2_D_SRAM7
port 1064 nsew signal output
flabel metal3 s 464800 601776 464912 601888 0 FreeSans 448 0 0 0 Tile_X8Y2_GWEN_SRAM
port 1065 nsew signal output
flabel metal3 s 464800 592816 464912 592928 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM0
port 1066 nsew signal input
flabel metal3 s 464800 593712 464912 593824 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM1
port 1067 nsew signal input
flabel metal3 s 464800 594608 464912 594720 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM2
port 1068 nsew signal input
flabel metal3 s 464800 595504 464912 595616 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM3
port 1069 nsew signal input
flabel metal3 s 464800 596400 464912 596512 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM4
port 1070 nsew signal input
flabel metal3 s 464800 597296 464912 597408 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM5
port 1071 nsew signal input
flabel metal3 s 464800 598192 464912 598304 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM6
port 1072 nsew signal input
flabel metal3 s 464800 599088 464912 599200 0 FreeSans 448 0 0 0 Tile_X8Y2_Q_SRAM7
port 1073 nsew signal input
flabel metal3 s 464800 602672 464912 602784 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM0
port 1074 nsew signal output
flabel metal3 s 464800 603568 464912 603680 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM1
port 1075 nsew signal output
flabel metal3 s 464800 604464 464912 604576 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM2
port 1076 nsew signal output
flabel metal3 s 464800 605360 464912 605472 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM3
port 1077 nsew signal output
flabel metal3 s 464800 606256 464912 606368 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM4
port 1078 nsew signal output
flabel metal3 s 464800 607152 464912 607264 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM5
port 1079 nsew signal output
flabel metal3 s 464800 608048 464912 608160 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM6
port 1080 nsew signal output
flabel metal3 s 464800 608944 464912 609056 0 FreeSans 448 0 0 0 Tile_X8Y2_WEN_SRAM7
port 1081 nsew signal output
flabel metal3 s 464800 494928 464912 495040 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM0
port 1082 nsew signal output
flabel metal3 s 464800 495824 464912 495936 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM1
port 1083 nsew signal output
flabel metal3 s 464800 496720 464912 496832 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM2
port 1084 nsew signal output
flabel metal3 s 464800 497616 464912 497728 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM3
port 1085 nsew signal output
flabel metal3 s 464800 498512 464912 498624 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM4
port 1086 nsew signal output
flabel metal3 s 464800 499408 464912 499520 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM5
port 1087 nsew signal output
flabel metal3 s 464800 500304 464912 500416 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM6
port 1088 nsew signal output
flabel metal3 s 464800 501200 464912 501312 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM7
port 1089 nsew signal output
flabel metal3 s 464800 502096 464912 502208 0 FreeSans 448 0 0 0 Tile_X8Y4_A_SRAM8
port 1090 nsew signal output
flabel metal3 s 464800 485968 464912 486080 0 FreeSans 448 0 0 0 Tile_X8Y4_CEN_SRAM
port 1091 nsew signal output
flabel metal3 s 464800 510160 464912 510272 0 FreeSans 448 0 0 0 Tile_X8Y4_CLK_SRAM
port 1092 nsew signal output
flabel metal3 s 464800 485072 464912 485184 0 FreeSans 448 0 0 0 Tile_X8Y4_CONFIGURED_top
port 1093 nsew signal input
flabel metal3 s 464800 502992 464912 503104 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM0
port 1094 nsew signal output
flabel metal3 s 464800 503888 464912 504000 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM1
port 1095 nsew signal output
flabel metal3 s 464800 504784 464912 504896 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM2
port 1096 nsew signal output
flabel metal3 s 464800 505680 464912 505792 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM3
port 1097 nsew signal output
flabel metal3 s 464800 506576 464912 506688 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM4
port 1098 nsew signal output
flabel metal3 s 464800 507472 464912 507584 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM5
port 1099 nsew signal output
flabel metal3 s 464800 508368 464912 508480 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM6
port 1100 nsew signal output
flabel metal3 s 464800 509264 464912 509376 0 FreeSans 448 0 0 0 Tile_X8Y4_D_SRAM7
port 1101 nsew signal output
flabel metal3 s 464800 486864 464912 486976 0 FreeSans 448 0 0 0 Tile_X8Y4_GWEN_SRAM
port 1102 nsew signal output
flabel metal3 s 464800 477904 464912 478016 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM0
port 1103 nsew signal input
flabel metal3 s 464800 478800 464912 478912 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM1
port 1104 nsew signal input
flabel metal3 s 464800 479696 464912 479808 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM2
port 1105 nsew signal input
flabel metal3 s 464800 480592 464912 480704 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM3
port 1106 nsew signal input
flabel metal3 s 464800 481488 464912 481600 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM4
port 1107 nsew signal input
flabel metal3 s 464800 482384 464912 482496 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM5
port 1108 nsew signal input
flabel metal3 s 464800 483280 464912 483392 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM6
port 1109 nsew signal input
flabel metal3 s 464800 484176 464912 484288 0 FreeSans 448 0 0 0 Tile_X8Y4_Q_SRAM7
port 1110 nsew signal input
flabel metal3 s 464800 487760 464912 487872 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM0
port 1111 nsew signal output
flabel metal3 s 464800 488656 464912 488768 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM1
port 1112 nsew signal output
flabel metal3 s 464800 489552 464912 489664 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM2
port 1113 nsew signal output
flabel metal3 s 464800 490448 464912 490560 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM3
port 1114 nsew signal output
flabel metal3 s 464800 491344 464912 491456 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM4
port 1115 nsew signal output
flabel metal3 s 464800 492240 464912 492352 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM5
port 1116 nsew signal output
flabel metal3 s 464800 493136 464912 493248 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM6
port 1117 nsew signal output
flabel metal3 s 464800 494032 464912 494144 0 FreeSans 448 0 0 0 Tile_X8Y4_WEN_SRAM7
port 1118 nsew signal output
flabel metal3 s 464800 380016 464912 380128 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM0
port 1119 nsew signal output
flabel metal3 s 464800 380912 464912 381024 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM1
port 1120 nsew signal output
flabel metal3 s 464800 381808 464912 381920 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM2
port 1121 nsew signal output
flabel metal3 s 464800 382704 464912 382816 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM3
port 1122 nsew signal output
flabel metal3 s 464800 383600 464912 383712 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM4
port 1123 nsew signal output
flabel metal3 s 464800 384496 464912 384608 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM5
port 1124 nsew signal output
flabel metal3 s 464800 385392 464912 385504 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM6
port 1125 nsew signal output
flabel metal3 s 464800 386288 464912 386400 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM7
port 1126 nsew signal output
flabel metal3 s 464800 387184 464912 387296 0 FreeSans 448 0 0 0 Tile_X8Y6_A_SRAM8
port 1127 nsew signal output
flabel metal3 s 464800 371056 464912 371168 0 FreeSans 448 0 0 0 Tile_X8Y6_CEN_SRAM
port 1128 nsew signal output
flabel metal3 s 464800 395248 464912 395360 0 FreeSans 448 0 0 0 Tile_X8Y6_CLK_SRAM
port 1129 nsew signal output
flabel metal3 s 464800 370160 464912 370272 0 FreeSans 448 0 0 0 Tile_X8Y6_CONFIGURED_top
port 1130 nsew signal input
flabel metal3 s 464800 388080 464912 388192 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM0
port 1131 nsew signal output
flabel metal3 s 464800 388976 464912 389088 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM1
port 1132 nsew signal output
flabel metal3 s 464800 389872 464912 389984 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM2
port 1133 nsew signal output
flabel metal3 s 464800 390768 464912 390880 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM3
port 1134 nsew signal output
flabel metal3 s 464800 391664 464912 391776 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM4
port 1135 nsew signal output
flabel metal3 s 464800 392560 464912 392672 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM5
port 1136 nsew signal output
flabel metal3 s 464800 393456 464912 393568 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM6
port 1137 nsew signal output
flabel metal3 s 464800 394352 464912 394464 0 FreeSans 448 0 0 0 Tile_X8Y6_D_SRAM7
port 1138 nsew signal output
flabel metal3 s 464800 371952 464912 372064 0 FreeSans 448 0 0 0 Tile_X8Y6_GWEN_SRAM
port 1139 nsew signal output
flabel metal3 s 464800 362992 464912 363104 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM0
port 1140 nsew signal input
flabel metal3 s 464800 363888 464912 364000 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM1
port 1141 nsew signal input
flabel metal3 s 464800 364784 464912 364896 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM2
port 1142 nsew signal input
flabel metal3 s 464800 365680 464912 365792 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM3
port 1143 nsew signal input
flabel metal3 s 464800 366576 464912 366688 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM4
port 1144 nsew signal input
flabel metal3 s 464800 367472 464912 367584 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM5
port 1145 nsew signal input
flabel metal3 s 464800 368368 464912 368480 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM6
port 1146 nsew signal input
flabel metal3 s 464800 369264 464912 369376 0 FreeSans 448 0 0 0 Tile_X8Y6_Q_SRAM7
port 1147 nsew signal input
flabel metal3 s 464800 372848 464912 372960 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM0
port 1148 nsew signal output
flabel metal3 s 464800 373744 464912 373856 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM1
port 1149 nsew signal output
flabel metal3 s 464800 374640 464912 374752 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM2
port 1150 nsew signal output
flabel metal3 s 464800 375536 464912 375648 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM3
port 1151 nsew signal output
flabel metal3 s 464800 376432 464912 376544 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM4
port 1152 nsew signal output
flabel metal3 s 464800 377328 464912 377440 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM5
port 1153 nsew signal output
flabel metal3 s 464800 378224 464912 378336 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM6
port 1154 nsew signal output
flabel metal3 s 464800 379120 464912 379232 0 FreeSans 448 0 0 0 Tile_X8Y6_WEN_SRAM7
port 1155 nsew signal output
flabel metal3 s 464800 265104 464912 265216 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM0
port 1156 nsew signal output
flabel metal3 s 464800 266000 464912 266112 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM1
port 1157 nsew signal output
flabel metal3 s 464800 266896 464912 267008 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM2
port 1158 nsew signal output
flabel metal3 s 464800 267792 464912 267904 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM3
port 1159 nsew signal output
flabel metal3 s 464800 268688 464912 268800 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM4
port 1160 nsew signal output
flabel metal3 s 464800 269584 464912 269696 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM5
port 1161 nsew signal output
flabel metal3 s 464800 270480 464912 270592 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM6
port 1162 nsew signal output
flabel metal3 s 464800 271376 464912 271488 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM7
port 1163 nsew signal output
flabel metal3 s 464800 272272 464912 272384 0 FreeSans 448 0 0 0 Tile_X8Y8_A_SRAM8
port 1164 nsew signal output
flabel metal3 s 464800 256144 464912 256256 0 FreeSans 448 0 0 0 Tile_X8Y8_CEN_SRAM
port 1165 nsew signal output
flabel metal3 s 464800 280336 464912 280448 0 FreeSans 448 0 0 0 Tile_X8Y8_CLK_SRAM
port 1166 nsew signal output
flabel metal3 s 464800 255248 464912 255360 0 FreeSans 448 0 0 0 Tile_X8Y8_CONFIGURED_top
port 1167 nsew signal input
flabel metal3 s 464800 273168 464912 273280 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM0
port 1168 nsew signal output
flabel metal3 s 464800 274064 464912 274176 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM1
port 1169 nsew signal output
flabel metal3 s 464800 274960 464912 275072 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM2
port 1170 nsew signal output
flabel metal3 s 464800 275856 464912 275968 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM3
port 1171 nsew signal output
flabel metal3 s 464800 276752 464912 276864 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM4
port 1172 nsew signal output
flabel metal3 s 464800 277648 464912 277760 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM5
port 1173 nsew signal output
flabel metal3 s 464800 278544 464912 278656 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM6
port 1174 nsew signal output
flabel metal3 s 464800 279440 464912 279552 0 FreeSans 448 0 0 0 Tile_X8Y8_D_SRAM7
port 1175 nsew signal output
flabel metal3 s 464800 257040 464912 257152 0 FreeSans 448 0 0 0 Tile_X8Y8_GWEN_SRAM
port 1176 nsew signal output
flabel metal3 s 464800 248080 464912 248192 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM0
port 1177 nsew signal input
flabel metal3 s 464800 248976 464912 249088 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM1
port 1178 nsew signal input
flabel metal3 s 464800 249872 464912 249984 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM2
port 1179 nsew signal input
flabel metal3 s 464800 250768 464912 250880 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM3
port 1180 nsew signal input
flabel metal3 s 464800 251664 464912 251776 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM4
port 1181 nsew signal input
flabel metal3 s 464800 252560 464912 252672 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM5
port 1182 nsew signal input
flabel metal3 s 464800 253456 464912 253568 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM6
port 1183 nsew signal input
flabel metal3 s 464800 254352 464912 254464 0 FreeSans 448 0 0 0 Tile_X8Y8_Q_SRAM7
port 1184 nsew signal input
flabel metal3 s 464800 257936 464912 258048 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM0
port 1185 nsew signal output
flabel metal3 s 464800 258832 464912 258944 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM1
port 1186 nsew signal output
flabel metal3 s 464800 259728 464912 259840 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM2
port 1187 nsew signal output
flabel metal3 s 464800 260624 464912 260736 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM3
port 1188 nsew signal output
flabel metal3 s 464800 261520 464912 261632 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM4
port 1189 nsew signal output
flabel metal3 s 464800 262416 464912 262528 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM5
port 1190 nsew signal output
flabel metal3 s 464800 263312 464912 263424 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM6
port 1191 nsew signal output
flabel metal3 s 464800 264208 464912 264320 0 FreeSans 448 0 0 0 Tile_X8Y8_WEN_SRAM7
port 1192 nsew signal output
flabel metal2 s 784 0 896 112 0 FreeSans 448 0 0 0 UserCLK
port 1193 nsew signal input
flabel metal4 s 3888 130256 4208 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 130256 24208 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 72800 4208 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 72800 24208 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 15344 4208 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 15344 24208 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 647360 4208 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 647360 24208 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 589904 4208 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 589904 24208 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 532448 4208 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 532448 24208 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 474992 4208 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 474992 24208 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 417536 4208 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 417536 24208 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 360080 4208 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 360080 24208 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 302624 4208 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 302624 24208 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 245168 4208 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 245168 24208 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 3888 187712 4208 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 23888 187712 24208 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 704816 32768 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 704816 52768 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 704816 72768 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 130256 32768 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 130256 52768 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 130256 72768 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 72800 32768 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 72800 52768 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 72800 72768 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 15344 32768 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 15344 52768 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 15344 72768 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 1120 32768 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 1120 52768 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 1120 72768 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 647360 32768 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 647360 52768 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 647360 72768 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 589904 32768 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 589904 52768 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 589904 72768 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 532448 32768 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 532448 52768 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 532448 72768 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 474992 32768 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 474992 52768 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 474992 72768 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 417536 32768 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 417536 52768 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 417536 72768 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 360080 32768 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 360080 52768 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 360080 72768 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 302624 32768 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 302624 52768 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 302624 72768 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 245168 32768 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 245168 52768 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 245168 72768 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 32448 187712 32768 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 52448 187712 52768 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 72448 187712 72768 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 704816 90224 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 704816 110224 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 704816 130224 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 130256 90224 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 130256 110224 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 130256 130224 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 72800 90224 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 72800 110224 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 72800 130224 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 15344 90224 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 15344 110224 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 15344 130224 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 1120 90224 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 1120 110224 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 1120 130224 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 647360 90224 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 647360 110224 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 647360 130224 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 589904 90224 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 589904 110224 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 589904 130224 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 532448 90224 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 532448 110224 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 532448 130224 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 474992 90224 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 474992 110224 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 474992 130224 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 417536 90224 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 417536 110224 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 417536 130224 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 360080 90224 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 360080 110224 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 360080 130224 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 302624 90224 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 302624 110224 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 302624 130224 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 245168 90224 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 245168 110224 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 245168 130224 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 89904 187712 90224 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 109904 187712 110224 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 129904 187712 130224 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 704816 147680 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 704816 167680 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 704816 187680 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 130256 147680 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 130256 167680 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 130256 187680 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 72800 147680 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 72800 167680 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 72800 187680 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 15344 147680 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 15344 167680 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 15344 187680 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 1120 147680 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 1120 167680 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 1120 187680 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 647360 147680 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 647360 167680 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 647360 187680 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 589904 147680 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 589904 167680 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 589904 187680 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 532448 147680 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 532448 167680 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 532448 187680 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 474992 147680 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 474992 167680 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 474992 187680 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 417536 147680 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 417536 167680 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 417536 187680 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 360080 147680 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 360080 167680 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 360080 187680 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 302624 147680 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 302624 167680 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 302624 187680 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 245168 147680 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 245168 167680 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 245168 187680 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 147360 187712 147680 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 167360 187712 167680 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 187360 187712 187680 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 704816 205136 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 704816 225136 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 704816 245136 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 130256 205136 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 130256 225136 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 130256 245136 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 72800 205136 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 72800 225136 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 72800 245136 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 15344 205136 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 15344 225136 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 15344 245136 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 1120 205136 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 1120 225136 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 1120 245136 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 647360 205136 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 647360 225136 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 647360 245136 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 589904 205136 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 589904 225136 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 589904 245136 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 532448 205136 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 532448 225136 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 532448 245136 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 474992 205136 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 474992 225136 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 474992 245136 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 417536 205136 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 417536 225136 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 417536 245136 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 360080 205136 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 360080 225136 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 360080 245136 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 302624 205136 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 302624 225136 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 302624 245136 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 245168 205136 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 245168 225136 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 245168 245136 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 204816 187712 205136 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 224816 187712 225136 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 244816 187712 245136 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 704816 269536 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 704816 289536 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 704816 309536 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 130256 269536 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 130256 289536 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 130256 309536 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 72800 269536 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 72800 289536 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 72800 309536 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 15344 269536 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 15344 289536 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 15344 309536 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 1120 269536 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 1120 289536 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 1120 309536 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 647360 269536 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 647360 289536 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 647360 309536 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 589904 269536 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 589904 289536 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 589904 309536 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 532448 269536 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 532448 289536 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 532448 309536 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 474992 269536 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 474992 289536 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 474992 309536 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 417536 269536 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 417536 289536 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 417536 309536 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 360080 269536 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 360080 289536 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 360080 309536 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 302624 269536 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 302624 289536 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 302624 309536 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 245168 269536 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 245168 289536 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 245168 309536 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 269216 187712 269536 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 289216 187712 289536 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 309216 187712 309536 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 704816 326992 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 704816 346992 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 704816 366992 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 15344 326992 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 15344 346992 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 15344 366992 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 1120 326992 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 1120 346992 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 1120 366992 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 589904 326992 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 589904 346992 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 589904 366992 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 474992 326992 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 474992 346992 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 474992 366992 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 360080 326992 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 360080 346992 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 360080 366992 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 245168 326992 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 245168 346992 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 245168 366992 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 326672 130256 326992 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 346672 130256 346992 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 366672 130256 366992 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 704816 379744 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 704816 399744 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 704816 419744 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 130256 379744 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 130256 399744 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 130256 419744 187712 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 72800 379744 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 72800 399744 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 72800 419744 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 15344 379744 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 15344 399744 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 15344 419744 72800 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 1120 379744 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 1120 399744 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 1120 419744 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 647360 379744 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 647360 399744 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 647360 419744 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 589904 379744 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 589904 399744 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 589904 419744 647360 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 532448 379744 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 532448 399744 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 532448 419744 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 474992 379744 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 474992 399744 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 474992 419744 532448 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 417536 379744 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 417536 399744 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 417536 419744 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 360080 379744 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 360080 399744 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 360080 419744 417536 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 302624 379744 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 302624 399744 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 302624 419744 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 245168 379744 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 245168 399744 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 245168 419744 302624 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 379424 187712 379744 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 399424 187712 399744 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 419424 187712 419744 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 704816 437200 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 704816 457200 719040 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 15344 437200 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 15344 457200 130256 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 1120 437200 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 1120 457200 15344 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 589904 437200 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 589904 457200 704816 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 474992 437200 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 474992 457200 589904 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 360080 437200 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 360080 457200 474992 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 245168 437200 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 245168 457200 360080 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 436880 130256 437200 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 456880 130256 457200 245168 0 FreeSans 1472 90 0 0 VDD
port 1194 nsew power bidirectional
flabel metal4 s 4548 130256 4868 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 130256 24868 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 72800 4868 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 72800 24868 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 15344 4868 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 15344 24868 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 647360 4868 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 647360 24868 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 589904 4868 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 589904 24868 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 532448 4868 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 532448 24868 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 474992 4868 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 474992 24868 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 417536 4868 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 417536 24868 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 360080 4868 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 360080 24868 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 302624 4868 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 302624 24868 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 245168 4868 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 245168 24868 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 4548 187712 4868 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 24548 187712 24868 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 704816 33428 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 704816 53428 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 704816 73428 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 130256 33428 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 130256 53428 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 130256 73428 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 72800 33428 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 72800 53428 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 72800 73428 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 15344 33428 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 15344 53428 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 15344 73428 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 1120 33428 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 1120 53428 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 1120 73428 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 647360 33428 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 647360 53428 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 647360 73428 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 589904 33428 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 589904 53428 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 589904 73428 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 532448 33428 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 532448 53428 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 532448 73428 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 474992 33428 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 474992 53428 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 474992 73428 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 417536 33428 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 417536 53428 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 417536 73428 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 360080 33428 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 360080 53428 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 360080 73428 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 302624 33428 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 302624 53428 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 302624 73428 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 245168 33428 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 245168 53428 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 245168 73428 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 33108 187712 33428 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 53108 187712 53428 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 73108 187712 73428 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 704816 90884 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 704816 110884 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 704816 130884 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 130256 90884 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 130256 110884 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 130256 130884 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 72800 90884 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 72800 110884 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 72800 130884 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 15344 90884 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 15344 110884 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 15344 130884 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 1120 90884 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 1120 110884 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 1120 130884 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 647360 90884 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 647360 110884 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 647360 130884 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 589904 90884 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 589904 110884 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 589904 130884 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 532448 90884 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 532448 110884 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 532448 130884 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 474992 90884 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 474992 110884 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 474992 130884 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 417536 90884 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 417536 110884 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 417536 130884 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 360080 90884 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 360080 110884 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 360080 130884 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 302624 90884 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 302624 110884 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 302624 130884 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 245168 90884 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 245168 110884 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 245168 130884 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 90564 187712 90884 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 110564 187712 110884 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 130564 187712 130884 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 704816 148340 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 704816 168340 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 704816 188340 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 130256 148340 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 130256 168340 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 130256 188340 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 72800 148340 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 72800 168340 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 72800 188340 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 15344 148340 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 15344 168340 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 15344 188340 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 1120 148340 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 1120 168340 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 1120 188340 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 647360 148340 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 647360 168340 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 647360 188340 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 589904 148340 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 589904 168340 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 589904 188340 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 532448 148340 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 532448 168340 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 532448 188340 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 474992 148340 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 474992 168340 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 474992 188340 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 417536 148340 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 417536 168340 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 417536 188340 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 360080 148340 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 360080 168340 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 360080 188340 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 302624 148340 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 302624 168340 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 302624 188340 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 245168 148340 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 245168 168340 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 245168 188340 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 148020 187712 148340 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 168020 187712 168340 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 188020 187712 188340 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 704816 205796 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 704816 225796 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 704816 245796 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 130256 205796 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 130256 225796 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 130256 245796 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 72800 205796 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 72800 225796 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 72800 245796 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 15344 205796 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 15344 225796 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 15344 245796 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 1120 205796 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 1120 225796 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 1120 245796 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 647360 205796 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 647360 225796 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 647360 245796 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 589904 205796 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 589904 225796 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 589904 245796 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 532448 205796 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 532448 225796 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 532448 245796 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 474992 205796 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 474992 225796 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 474992 245796 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 417536 205796 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 417536 225796 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 417536 245796 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 360080 205796 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 360080 225796 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 360080 245796 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 302624 205796 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 302624 225796 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 302624 245796 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 245168 205796 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 245168 225796 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 245168 245796 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 205476 187712 205796 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 225476 187712 225796 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 245476 187712 245796 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 704816 270196 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 704816 290196 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 704816 310196 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 130256 270196 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 130256 290196 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 130256 310196 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 72800 270196 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 72800 290196 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 72800 310196 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 15344 270196 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 15344 290196 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 15344 310196 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 1120 270196 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 1120 290196 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 1120 310196 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 647360 270196 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 647360 290196 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 647360 310196 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 589904 270196 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 589904 290196 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 589904 310196 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 532448 270196 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 532448 290196 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 532448 310196 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 474992 270196 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 474992 290196 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 474992 310196 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 417536 270196 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 417536 290196 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 417536 310196 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 360080 270196 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 360080 290196 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 360080 310196 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 302624 270196 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 302624 290196 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 302624 310196 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 245168 270196 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 245168 290196 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 245168 310196 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 269876 187712 270196 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 289876 187712 290196 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 309876 187712 310196 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 704816 327652 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 704816 347652 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 704816 367652 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 15344 327652 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 15344 347652 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 15344 367652 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 1120 327652 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 1120 347652 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 1120 367652 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 589904 327652 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 589904 347652 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 589904 367652 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 474992 327652 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 474992 347652 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 474992 367652 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 360080 327652 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 360080 347652 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 360080 367652 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 245168 327652 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 245168 347652 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 245168 367652 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 327332 130256 327652 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 347332 130256 347652 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 367332 130256 367652 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 704816 380404 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 704816 400404 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 704816 420404 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 130256 380404 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 130256 400404 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 130256 420404 187712 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 72800 380404 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 72800 400404 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 72800 420404 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 15344 380404 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 15344 400404 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 15344 420404 72800 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 1120 380404 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 1120 400404 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 1120 420404 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 647360 380404 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 647360 400404 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 647360 420404 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 589904 380404 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 589904 400404 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 589904 420404 647360 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 532448 380404 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 532448 400404 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 532448 420404 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 474992 380404 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 474992 400404 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 474992 420404 532448 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 417536 380404 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 417536 400404 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 417536 420404 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 360080 380404 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 360080 400404 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 360080 420404 417536 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 302624 380404 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 302624 400404 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 302624 420404 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 245168 380404 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 245168 400404 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 245168 420404 302624 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 380084 187712 380404 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 400084 187712 400404 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 420084 187712 420404 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 704816 437860 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 704816 457860 719040 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 15344 437860 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 15344 457860 130256 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 1120 437860 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 1120 457860 15344 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 589904 437860 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 589904 457860 704816 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 474992 437860 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 474992 457860 589904 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 360080 437860 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 360080 457860 474992 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 245168 437860 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 245168 457860 360080 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 437540 130256 437860 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
flabel metal4 s 457540 130256 457860 245168 0 FreeSans 1472 90 0 0 VSS
port 1195 nsew ground bidirectional
rlabel metal4 457040 187712 457040 187712 0 VDD
rlabel metal4 457700 187712 457700 187712 0 VSS
rlabel metal3 28056 704788 28056 704788 0 FrameData[0]
rlabel metal3 112 563416 112 563416 0 FrameData[100]
rlabel metal3 112 564312 112 564312 0 FrameData[101]
rlabel metal3 112 565208 112 565208 0 FrameData[102]
rlabel metal3 112 566104 112 566104 0 FrameData[103]
rlabel metal3 112 567000 112 567000 0 FrameData[104]
rlabel metal3 112 567896 112 567896 0 FrameData[105]
rlabel metal3 112 568792 112 568792 0 FrameData[106]
rlabel metal3 112 569688 112 569688 0 FrameData[107]
rlabel metal3 112 570584 112 570584 0 FrameData[108]
rlabel metal3 112 571480 112 571480 0 FrameData[109]
rlabel metal3 14392 709352 14392 709352 0 FrameData[10]
rlabel metal3 112 572376 112 572376 0 FrameData[110]
rlabel metal3 112 573272 112 573272 0 FrameData[111]
rlabel metal3 112 574168 112 574168 0 FrameData[112]
rlabel metal3 112 575064 112 575064 0 FrameData[113]
rlabel metal3 112 575960 112 575960 0 FrameData[114]
rlabel metal3 112 576856 112 576856 0 FrameData[115]
rlabel metal3 112 577752 112 577752 0 FrameData[116]
rlabel metal3 112 578648 112 578648 0 FrameData[117]
rlabel metal3 112 579544 112 579544 0 FrameData[118]
rlabel metal3 112 580440 112 580440 0 FrameData[119]
rlabel metal3 14392 709800 14392 709800 0 FrameData[11]
rlabel metal3 112 581336 112 581336 0 FrameData[120]
rlabel metal3 112 582232 112 582232 0 FrameData[121]
rlabel metal3 112 583128 112 583128 0 FrameData[122]
rlabel metal3 112 584024 112 584024 0 FrameData[123]
rlabel metal3 112 584920 112 584920 0 FrameData[124]
rlabel metal3 112 585816 112 585816 0 FrameData[125]
rlabel metal3 112 586712 112 586712 0 FrameData[126]
rlabel metal3 112 587608 112 587608 0 FrameData[127]
rlabel metal3 112 502376 112 502376 0 FrameData[128]
rlabel metal3 112 503272 112 503272 0 FrameData[129]
rlabel metal3 14392 710248 14392 710248 0 FrameData[12]
rlabel metal3 112 504168 112 504168 0 FrameData[130]
rlabel metal3 112 505064 112 505064 0 FrameData[131]
rlabel metal3 112 505960 112 505960 0 FrameData[132]
rlabel metal3 112 506856 112 506856 0 FrameData[133]
rlabel metal3 112 507752 112 507752 0 FrameData[134]
rlabel metal3 112 508648 112 508648 0 FrameData[135]
rlabel metal3 112 509544 112 509544 0 FrameData[136]
rlabel metal3 112 510440 112 510440 0 FrameData[137]
rlabel metal3 112 511336 112 511336 0 FrameData[138]
rlabel metal3 112 512232 112 512232 0 FrameData[139]
rlabel metal3 14392 710696 14392 710696 0 FrameData[13]
rlabel metal3 112 513128 112 513128 0 FrameData[140]
rlabel metal3 112 514024 112 514024 0 FrameData[141]
rlabel metal3 112 514920 112 514920 0 FrameData[142]
rlabel metal3 112 515816 112 515816 0 FrameData[143]
rlabel metal3 112 516712 112 516712 0 FrameData[144]
rlabel metal3 112 517608 112 517608 0 FrameData[145]
rlabel metal3 112 518504 112 518504 0 FrameData[146]
rlabel metal3 112 519400 112 519400 0 FrameData[147]
rlabel metal3 112 520296 112 520296 0 FrameData[148]
rlabel metal3 112 521192 112 521192 0 FrameData[149]
rlabel metal3 14392 711144 14392 711144 0 FrameData[14]
rlabel metal3 112 522088 112 522088 0 FrameData[150]
rlabel metal3 112 522984 112 522984 0 FrameData[151]
rlabel metal3 112 523880 112 523880 0 FrameData[152]
rlabel metal3 112 524776 112 524776 0 FrameData[153]
rlabel metal3 112 525672 112 525672 0 FrameData[154]
rlabel metal3 112 526568 112 526568 0 FrameData[155]
rlabel metal3 112 527464 112 527464 0 FrameData[156]
rlabel metal3 112 528360 112 528360 0 FrameData[157]
rlabel metal3 112 529256 112 529256 0 FrameData[158]
rlabel metal3 112 530152 112 530152 0 FrameData[159]
rlabel metal3 14392 711592 14392 711592 0 FrameData[15]
rlabel metal3 112 444920 112 444920 0 FrameData[160]
rlabel metal3 112 445816 112 445816 0 FrameData[161]
rlabel metal3 112 446712 112 446712 0 FrameData[162]
rlabel metal3 112 447608 112 447608 0 FrameData[163]
rlabel metal3 112 448504 112 448504 0 FrameData[164]
rlabel metal3 112 449400 112 449400 0 FrameData[165]
rlabel metal3 112 450296 112 450296 0 FrameData[166]
rlabel metal3 112 451192 112 451192 0 FrameData[167]
rlabel metal3 112 452088 112 452088 0 FrameData[168]
rlabel metal3 112 452984 112 452984 0 FrameData[169]
rlabel metal3 14392 712040 14392 712040 0 FrameData[16]
rlabel metal3 112 453880 112 453880 0 FrameData[170]
rlabel metal3 112 454776 112 454776 0 FrameData[171]
rlabel metal3 112 455672 112 455672 0 FrameData[172]
rlabel metal3 112 456568 112 456568 0 FrameData[173]
rlabel metal3 112 457464 112 457464 0 FrameData[174]
rlabel metal3 112 458360 112 458360 0 FrameData[175]
rlabel metal3 112 459256 112 459256 0 FrameData[176]
rlabel metal3 112 460152 112 460152 0 FrameData[177]
rlabel metal3 112 461048 112 461048 0 FrameData[178]
rlabel metal3 112 461944 112 461944 0 FrameData[179]
rlabel metal3 14392 712488 14392 712488 0 FrameData[17]
rlabel metal3 112 462840 112 462840 0 FrameData[180]
rlabel metal3 112 463736 112 463736 0 FrameData[181]
rlabel metal3 112 464632 112 464632 0 FrameData[182]
rlabel metal3 112 465528 112 465528 0 FrameData[183]
rlabel metal3 112 466424 112 466424 0 FrameData[184]
rlabel metal3 112 467320 112 467320 0 FrameData[185]
rlabel metal3 112 468216 112 468216 0 FrameData[186]
rlabel metal3 112 469112 112 469112 0 FrameData[187]
rlabel metal3 112 470008 112 470008 0 FrameData[188]
rlabel metal3 112 470904 112 470904 0 FrameData[189]
rlabel metal3 14392 712936 14392 712936 0 FrameData[18]
rlabel metal3 112 471800 112 471800 0 FrameData[190]
rlabel metal3 112 472696 112 472696 0 FrameData[191]
rlabel metal3 112 387464 112 387464 0 FrameData[192]
rlabel metal3 112 388360 112 388360 0 FrameData[193]
rlabel metal3 112 389256 112 389256 0 FrameData[194]
rlabel metal3 112 390152 112 390152 0 FrameData[195]
rlabel metal3 112 391048 112 391048 0 FrameData[196]
rlabel metal3 112 391944 112 391944 0 FrameData[197]
rlabel metal3 112 392840 112 392840 0 FrameData[198]
rlabel metal3 112 393736 112 393736 0 FrameData[199]
rlabel metal3 14392 713384 14392 713384 0 FrameData[19]
rlabel metal3 14392 705320 14392 705320 0 FrameData[1]
rlabel metal3 112 394632 112 394632 0 FrameData[200]
rlabel metal3 112 395528 112 395528 0 FrameData[201]
rlabel metal3 112 396424 112 396424 0 FrameData[202]
rlabel metal3 112 397320 112 397320 0 FrameData[203]
rlabel metal3 112 398216 112 398216 0 FrameData[204]
rlabel metal3 112 399112 112 399112 0 FrameData[205]
rlabel metal3 112 400008 112 400008 0 FrameData[206]
rlabel metal3 112 400904 112 400904 0 FrameData[207]
rlabel metal3 112 401800 112 401800 0 FrameData[208]
rlabel metal3 112 402696 112 402696 0 FrameData[209]
rlabel metal3 14392 713832 14392 713832 0 FrameData[20]
rlabel metal3 112 403592 112 403592 0 FrameData[210]
rlabel metal3 112 404488 112 404488 0 FrameData[211]
rlabel metal3 112 405384 112 405384 0 FrameData[212]
rlabel metal3 112 406280 112 406280 0 FrameData[213]
rlabel metal3 112 407176 112 407176 0 FrameData[214]
rlabel metal3 112 408072 112 408072 0 FrameData[215]
rlabel metal3 112 408968 112 408968 0 FrameData[216]
rlabel metal3 112 409864 112 409864 0 FrameData[217]
rlabel metal3 112 410760 112 410760 0 FrameData[218]
rlabel metal3 112 411656 112 411656 0 FrameData[219]
rlabel metal3 14392 714280 14392 714280 0 FrameData[21]
rlabel metal3 112 412552 112 412552 0 FrameData[220]
rlabel metal3 112 413448 112 413448 0 FrameData[221]
rlabel metal3 112 414344 112 414344 0 FrameData[222]
rlabel metal3 112 415240 112 415240 0 FrameData[223]
rlabel metal3 112 330008 112 330008 0 FrameData[224]
rlabel metal3 112 330904 112 330904 0 FrameData[225]
rlabel metal3 112 331800 112 331800 0 FrameData[226]
rlabel metal3 112 332696 112 332696 0 FrameData[227]
rlabel metal3 112 333592 112 333592 0 FrameData[228]
rlabel metal3 112 334488 112 334488 0 FrameData[229]
rlabel metal3 14392 714728 14392 714728 0 FrameData[22]
rlabel metal3 112 335384 112 335384 0 FrameData[230]
rlabel metal3 112 336280 112 336280 0 FrameData[231]
rlabel metal3 112 337176 112 337176 0 FrameData[232]
rlabel metal3 112 338072 112 338072 0 FrameData[233]
rlabel metal3 112 338968 112 338968 0 FrameData[234]
rlabel metal3 112 339864 112 339864 0 FrameData[235]
rlabel metal3 112 340760 112 340760 0 FrameData[236]
rlabel metal3 112 341656 112 341656 0 FrameData[237]
rlabel metal3 112 342552 112 342552 0 FrameData[238]
rlabel metal3 112 343448 112 343448 0 FrameData[239]
rlabel metal3 14392 715176 14392 715176 0 FrameData[23]
rlabel metal3 112 344344 112 344344 0 FrameData[240]
rlabel metal3 112 345240 112 345240 0 FrameData[241]
rlabel metal3 112 346136 112 346136 0 FrameData[242]
rlabel metal3 112 347032 112 347032 0 FrameData[243]
rlabel metal3 112 347928 112 347928 0 FrameData[244]
rlabel metal3 112 348824 112 348824 0 FrameData[245]
rlabel metal3 112 349720 112 349720 0 FrameData[246]
rlabel metal3 112 350616 112 350616 0 FrameData[247]
rlabel metal3 112 351512 112 351512 0 FrameData[248]
rlabel metal3 112 352408 112 352408 0 FrameData[249]
rlabel metal3 14392 715624 14392 715624 0 FrameData[24]
rlabel metal3 112 353304 112 353304 0 FrameData[250]
rlabel metal3 112 354200 112 354200 0 FrameData[251]
rlabel metal3 112 355096 112 355096 0 FrameData[252]
rlabel metal3 112 355992 112 355992 0 FrameData[253]
rlabel metal3 112 356888 112 356888 0 FrameData[254]
rlabel metal3 112 357784 112 357784 0 FrameData[255]
rlabel metal3 112 272552 112 272552 0 FrameData[256]
rlabel metal3 112 273448 112 273448 0 FrameData[257]
rlabel metal3 112 274344 112 274344 0 FrameData[258]
rlabel metal3 112 275240 112 275240 0 FrameData[259]
rlabel metal3 14392 716072 14392 716072 0 FrameData[25]
rlabel metal3 112 276136 112 276136 0 FrameData[260]
rlabel metal3 112 277032 112 277032 0 FrameData[261]
rlabel metal3 112 277928 112 277928 0 FrameData[262]
rlabel metal3 112 278824 112 278824 0 FrameData[263]
rlabel metal3 112 279720 112 279720 0 FrameData[264]
rlabel metal3 112 280616 112 280616 0 FrameData[265]
rlabel metal3 112 281512 112 281512 0 FrameData[266]
rlabel metal3 112 282408 112 282408 0 FrameData[267]
rlabel metal3 112 283304 112 283304 0 FrameData[268]
rlabel metal3 112 284200 112 284200 0 FrameData[269]
rlabel metal3 14392 716520 14392 716520 0 FrameData[26]
rlabel metal3 112 285096 112 285096 0 FrameData[270]
rlabel metal3 112 285992 112 285992 0 FrameData[271]
rlabel metal3 112 286888 112 286888 0 FrameData[272]
rlabel metal3 112 287784 112 287784 0 FrameData[273]
rlabel metal3 112 288680 112 288680 0 FrameData[274]
rlabel metal3 112 289576 112 289576 0 FrameData[275]
rlabel metal3 112 290472 112 290472 0 FrameData[276]
rlabel metal3 112 291368 112 291368 0 FrameData[277]
rlabel metal3 112 292264 112 292264 0 FrameData[278]
rlabel metal3 112 293160 112 293160 0 FrameData[279]
rlabel metal3 14392 716968 14392 716968 0 FrameData[27]
rlabel metal3 112 294056 112 294056 0 FrameData[280]
rlabel metal3 112 294952 112 294952 0 FrameData[281]
rlabel metal3 112 295848 112 295848 0 FrameData[282]
rlabel metal3 112 296744 112 296744 0 FrameData[283]
rlabel metal3 112 297640 112 297640 0 FrameData[284]
rlabel metal3 112 298536 112 298536 0 FrameData[285]
rlabel metal3 112 299432 112 299432 0 FrameData[286]
rlabel metal3 112 300328 112 300328 0 FrameData[287]
rlabel metal3 112 215096 112 215096 0 FrameData[288]
rlabel metal3 112 215992 112 215992 0 FrameData[289]
rlabel metal3 966 717416 966 717416 0 FrameData[28]
rlabel metal3 112 216888 112 216888 0 FrameData[290]
rlabel metal3 112 217784 112 217784 0 FrameData[291]
rlabel metal3 112 218680 112 218680 0 FrameData[292]
rlabel metal3 112 219576 112 219576 0 FrameData[293]
rlabel metal3 112 220472 112 220472 0 FrameData[294]
rlabel metal3 112 221368 112 221368 0 FrameData[295]
rlabel metal3 112 222264 112 222264 0 FrameData[296]
rlabel metal3 112 223160 112 223160 0 FrameData[297]
rlabel metal3 112 224056 112 224056 0 FrameData[298]
rlabel metal3 112 224952 112 224952 0 FrameData[299]
rlabel metal3 14392 717864 14392 717864 0 FrameData[29]
rlabel metal3 14392 705768 14392 705768 0 FrameData[2]
rlabel metal3 112 225848 112 225848 0 FrameData[300]
rlabel metal3 112 226744 112 226744 0 FrameData[301]
rlabel metal3 112 227640 112 227640 0 FrameData[302]
rlabel metal3 112 228536 112 228536 0 FrameData[303]
rlabel metal3 112 229432 112 229432 0 FrameData[304]
rlabel metal3 112 230328 112 230328 0 FrameData[305]
rlabel metal3 112 231224 112 231224 0 FrameData[306]
rlabel metal3 112 232120 112 232120 0 FrameData[307]
rlabel metal3 112 233016 112 233016 0 FrameData[308]
rlabel metal3 112 233912 112 233912 0 FrameData[309]
rlabel metal3 14392 718312 14392 718312 0 FrameData[30]
rlabel metal3 112 234808 112 234808 0 FrameData[310]
rlabel metal3 112 235704 112 235704 0 FrameData[311]
rlabel metal3 112 236600 112 236600 0 FrameData[312]
rlabel metal3 112 237496 112 237496 0 FrameData[313]
rlabel metal3 112 238392 112 238392 0 FrameData[314]
rlabel metal3 112 239288 112 239288 0 FrameData[315]
rlabel metal3 112 240184 112 240184 0 FrameData[316]
rlabel metal3 112 241080 112 241080 0 FrameData[317]
rlabel metal3 112 241976 112 241976 0 FrameData[318]
rlabel metal3 112 242872 112 242872 0 FrameData[319]
rlabel metal3 14392 718760 14392 718760 0 FrameData[31]
rlabel metal3 112 157640 112 157640 0 FrameData[320]
rlabel metal3 112 158536 112 158536 0 FrameData[321]
rlabel metal3 112 159432 112 159432 0 FrameData[322]
rlabel metal3 112 160328 112 160328 0 FrameData[323]
rlabel metal3 112 161224 112 161224 0 FrameData[324]
rlabel metal3 112 162120 112 162120 0 FrameData[325]
rlabel metal3 112 163016 112 163016 0 FrameData[326]
rlabel metal3 112 163912 112 163912 0 FrameData[327]
rlabel metal3 112 164808 112 164808 0 FrameData[328]
rlabel metal3 112 165704 112 165704 0 FrameData[329]
rlabel metal3 112 674744 112 674744 0 FrameData[32]
rlabel metal3 112 166600 112 166600 0 FrameData[330]
rlabel metal3 112 167496 112 167496 0 FrameData[331]
rlabel metal3 112 168392 112 168392 0 FrameData[332]
rlabel metal3 112 169288 112 169288 0 FrameData[333]
rlabel metal3 112 170184 112 170184 0 FrameData[334]
rlabel metal3 112 171080 112 171080 0 FrameData[335]
rlabel metal3 112 171976 112 171976 0 FrameData[336]
rlabel metal3 112 172872 112 172872 0 FrameData[337]
rlabel metal3 112 173768 112 173768 0 FrameData[338]
rlabel metal3 112 174664 112 174664 0 FrameData[339]
rlabel metal3 112 675640 112 675640 0 FrameData[33]
rlabel metal3 112 175560 112 175560 0 FrameData[340]
rlabel metal3 112 176456 112 176456 0 FrameData[341]
rlabel metal3 112 177352 112 177352 0 FrameData[342]
rlabel metal3 112 178248 112 178248 0 FrameData[343]
rlabel metal3 112 179144 112 179144 0 FrameData[344]
rlabel metal3 112 180040 112 180040 0 FrameData[345]
rlabel metal3 112 180936 112 180936 0 FrameData[346]
rlabel metal3 112 181832 112 181832 0 FrameData[347]
rlabel metal3 112 182728 112 182728 0 FrameData[348]
rlabel metal3 112 183624 112 183624 0 FrameData[349]
rlabel metal3 112 676536 112 676536 0 FrameData[34]
rlabel metal3 112 184520 112 184520 0 FrameData[350]
rlabel metal3 112 185416 112 185416 0 FrameData[351]
rlabel metal3 112 100184 112 100184 0 FrameData[352]
rlabel metal3 112 101080 112 101080 0 FrameData[353]
rlabel metal3 112 101976 112 101976 0 FrameData[354]
rlabel metal3 112 102872 112 102872 0 FrameData[355]
rlabel metal3 112 103768 112 103768 0 FrameData[356]
rlabel metal3 112 104664 112 104664 0 FrameData[357]
rlabel metal3 112 105560 112 105560 0 FrameData[358]
rlabel metal3 112 106456 112 106456 0 FrameData[359]
rlabel metal3 112 677432 112 677432 0 FrameData[35]
rlabel metal3 112 107352 112 107352 0 FrameData[360]
rlabel metal3 112 108248 112 108248 0 FrameData[361]
rlabel metal3 112 109144 112 109144 0 FrameData[362]
rlabel metal3 112 110040 112 110040 0 FrameData[363]
rlabel metal3 112 110936 112 110936 0 FrameData[364]
rlabel metal3 112 111832 112 111832 0 FrameData[365]
rlabel metal3 112 112728 112 112728 0 FrameData[366]
rlabel metal3 112 113624 112 113624 0 FrameData[367]
rlabel metal3 112 114520 112 114520 0 FrameData[368]
rlabel metal3 112 115416 112 115416 0 FrameData[369]
rlabel metal3 112 678328 112 678328 0 FrameData[36]
rlabel metal3 112 116312 112 116312 0 FrameData[370]
rlabel metal3 112 117208 112 117208 0 FrameData[371]
rlabel metal3 112 118104 112 118104 0 FrameData[372]
rlabel metal3 112 119000 112 119000 0 FrameData[373]
rlabel metal3 112 119896 112 119896 0 FrameData[374]
rlabel metal3 112 120792 112 120792 0 FrameData[375]
rlabel metal3 112 121688 112 121688 0 FrameData[376]
rlabel metal3 112 122584 112 122584 0 FrameData[377]
rlabel metal3 112 123480 112 123480 0 FrameData[378]
rlabel metal3 112 124376 112 124376 0 FrameData[379]
rlabel metal3 112 679224 112 679224 0 FrameData[37]
rlabel metal3 112 125272 112 125272 0 FrameData[380]
rlabel metal3 112 126168 112 126168 0 FrameData[381]
rlabel metal3 112 127064 112 127064 0 FrameData[382]
rlabel metal3 112 127960 112 127960 0 FrameData[383]
rlabel metal3 112 42728 112 42728 0 FrameData[384]
rlabel metal3 112 43624 112 43624 0 FrameData[385]
rlabel metal3 112 44520 112 44520 0 FrameData[386]
rlabel metal3 112 45416 112 45416 0 FrameData[387]
rlabel metal3 112 46312 112 46312 0 FrameData[388]
rlabel metal3 112 47208 112 47208 0 FrameData[389]
rlabel metal3 112 680120 112 680120 0 FrameData[38]
rlabel metal3 112 48104 112 48104 0 FrameData[390]
rlabel metal3 112 49000 112 49000 0 FrameData[391]
rlabel metal3 112 49896 112 49896 0 FrameData[392]
rlabel metal3 112 50792 112 50792 0 FrameData[393]
rlabel metal3 112 51688 112 51688 0 FrameData[394]
rlabel metal3 112 52584 112 52584 0 FrameData[395]
rlabel metal3 112 53480 112 53480 0 FrameData[396]
rlabel metal3 112 54376 112 54376 0 FrameData[397]
rlabel metal3 112 55272 112 55272 0 FrameData[398]
rlabel metal3 112 56168 112 56168 0 FrameData[399]
rlabel metal3 112 681016 112 681016 0 FrameData[39]
rlabel metal3 14392 706216 14392 706216 0 FrameData[3]
rlabel metal3 112 57064 112 57064 0 FrameData[400]
rlabel metal3 112 57960 112 57960 0 FrameData[401]
rlabel metal3 112 58856 112 58856 0 FrameData[402]
rlabel metal3 112 59752 112 59752 0 FrameData[403]
rlabel metal3 112 60648 112 60648 0 FrameData[404]
rlabel metal3 112 61544 112 61544 0 FrameData[405]
rlabel metal3 112 62440 112 62440 0 FrameData[406]
rlabel metal3 112 63336 112 63336 0 FrameData[407]
rlabel metal3 112 64232 112 64232 0 FrameData[408]
rlabel metal3 112 65128 112 65128 0 FrameData[409]
rlabel metal3 112 681912 112 681912 0 FrameData[40]
rlabel metal3 112 66024 112 66024 0 FrameData[410]
rlabel metal3 112 66920 112 66920 0 FrameData[411]
rlabel metal3 112 67816 112 67816 0 FrameData[412]
rlabel metal3 112 68712 112 68712 0 FrameData[413]
rlabel metal3 112 69608 112 69608 0 FrameData[414]
rlabel metal3 112 70504 112 70504 0 FrameData[415]
rlabel metal3 28728 966 28728 966 0 FrameData[416]
rlabel metal3 28056 1260 28056 1260 0 FrameData[417]
rlabel metal3 14392 2072 14392 2072 0 FrameData[418]
rlabel metal3 14392 2520 14392 2520 0 FrameData[419]
rlabel metal3 112 682808 112 682808 0 FrameData[41]
rlabel metal3 14392 2968 14392 2968 0 FrameData[420]
rlabel metal3 14392 3416 14392 3416 0 FrameData[421]
rlabel metal3 14392 3864 14392 3864 0 FrameData[422]
rlabel metal3 14392 4312 14392 4312 0 FrameData[423]
rlabel metal3 14392 4760 14392 4760 0 FrameData[424]
rlabel metal3 14392 5208 14392 5208 0 FrameData[425]
rlabel metal3 14392 5656 14392 5656 0 FrameData[426]
rlabel metal3 14392 6104 14392 6104 0 FrameData[427]
rlabel metal3 14392 6552 14392 6552 0 FrameData[428]
rlabel metal3 14392 7000 14392 7000 0 FrameData[429]
rlabel metal3 112 683704 112 683704 0 FrameData[42]
rlabel metal3 14392 7448 14392 7448 0 FrameData[430]
rlabel metal3 14392 7896 14392 7896 0 FrameData[431]
rlabel metal3 14392 8344 14392 8344 0 FrameData[432]
rlabel metal3 14392 8792 14392 8792 0 FrameData[433]
rlabel metal3 14392 9240 14392 9240 0 FrameData[434]
rlabel metal3 14392 9688 14392 9688 0 FrameData[435]
rlabel metal3 14392 10136 14392 10136 0 FrameData[436]
rlabel metal3 14392 10584 14392 10584 0 FrameData[437]
rlabel metal3 14392 11032 14392 11032 0 FrameData[438]
rlabel metal3 14392 11480 14392 11480 0 FrameData[439]
rlabel metal3 112 684600 112 684600 0 FrameData[43]
rlabel metal3 14392 11928 14392 11928 0 FrameData[440]
rlabel metal3 14392 12376 14392 12376 0 FrameData[441]
rlabel metal3 14392 12824 14392 12824 0 FrameData[442]
rlabel metal3 14392 13272 14392 13272 0 FrameData[443]
rlabel metal3 14392 13720 14392 13720 0 FrameData[444]
rlabel metal3 14392 14168 14392 14168 0 FrameData[445]
rlabel metal3 14392 14616 14392 14616 0 FrameData[446]
rlabel metal3 14392 15064 14392 15064 0 FrameData[447]
rlabel metal3 112 685496 112 685496 0 FrameData[44]
rlabel metal3 112 686392 112 686392 0 FrameData[45]
rlabel metal3 112 687288 112 687288 0 FrameData[46]
rlabel metal3 112 688184 112 688184 0 FrameData[47]
rlabel metal3 112 689080 112 689080 0 FrameData[48]
rlabel metal3 112 689976 112 689976 0 FrameData[49]
rlabel metal3 14392 706664 14392 706664 0 FrameData[4]
rlabel metal3 112 690872 112 690872 0 FrameData[50]
rlabel metal3 112 691768 112 691768 0 FrameData[51]
rlabel metal3 112 692664 112 692664 0 FrameData[52]
rlabel metal3 112 693560 112 693560 0 FrameData[53]
rlabel metal3 112 694456 112 694456 0 FrameData[54]
rlabel metal3 112 695352 112 695352 0 FrameData[55]
rlabel metal3 112 696248 112 696248 0 FrameData[56]
rlabel metal3 112 697144 112 697144 0 FrameData[57]
rlabel metal3 112 698040 112 698040 0 FrameData[58]
rlabel metal3 112 698936 112 698936 0 FrameData[59]
rlabel metal3 14392 707112 14392 707112 0 FrameData[5]
rlabel metal3 112 699832 112 699832 0 FrameData[60]
rlabel metal3 112 700728 112 700728 0 FrameData[61]
rlabel metal3 112 701624 112 701624 0 FrameData[62]
rlabel metal3 112 702520 112 702520 0 FrameData[63]
rlabel metal3 112 617288 112 617288 0 FrameData[64]
rlabel metal3 112 618184 112 618184 0 FrameData[65]
rlabel metal3 112 619080 112 619080 0 FrameData[66]
rlabel metal3 112 619976 112 619976 0 FrameData[67]
rlabel metal3 112 620872 112 620872 0 FrameData[68]
rlabel metal3 112 621768 112 621768 0 FrameData[69]
rlabel metal3 14392 707560 14392 707560 0 FrameData[6]
rlabel metal3 112 622664 112 622664 0 FrameData[70]
rlabel metal3 112 623560 112 623560 0 FrameData[71]
rlabel metal3 112 624456 112 624456 0 FrameData[72]
rlabel metal3 112 625352 112 625352 0 FrameData[73]
rlabel metal3 112 626248 112 626248 0 FrameData[74]
rlabel metal3 112 627144 112 627144 0 FrameData[75]
rlabel metal3 112 628040 112 628040 0 FrameData[76]
rlabel metal3 112 628936 112 628936 0 FrameData[77]
rlabel metal3 112 629832 112 629832 0 FrameData[78]
rlabel metal3 112 630728 112 630728 0 FrameData[79]
rlabel metal3 14392 708008 14392 708008 0 FrameData[7]
rlabel metal3 112 631624 112 631624 0 FrameData[80]
rlabel metal3 112 632520 112 632520 0 FrameData[81]
rlabel metal3 112 633416 112 633416 0 FrameData[82]
rlabel metal3 112 634312 112 634312 0 FrameData[83]
rlabel metal3 112 635208 112 635208 0 FrameData[84]
rlabel metal3 112 636104 112 636104 0 FrameData[85]
rlabel metal3 112 637000 112 637000 0 FrameData[86]
rlabel metal3 112 637896 112 637896 0 FrameData[87]
rlabel metal3 112 638792 112 638792 0 FrameData[88]
rlabel metal3 112 639688 112 639688 0 FrameData[89]
rlabel metal3 14392 708456 14392 708456 0 FrameData[8]
rlabel metal3 112 640584 112 640584 0 FrameData[90]
rlabel metal3 112 641480 112 641480 0 FrameData[91]
rlabel metal3 112 642376 112 642376 0 FrameData[92]
rlabel metal3 112 643272 112 643272 0 FrameData[93]
rlabel metal3 112 644168 112 644168 0 FrameData[94]
rlabel metal3 112 645064 112 645064 0 FrameData[95]
rlabel metal3 112 559832 112 559832 0 FrameData[96]
rlabel metal3 112 560728 112 560728 0 FrameData[97]
rlabel metal3 112 561624 112 561624 0 FrameData[98]
rlabel metal3 112 562520 112 562520 0 FrameData[99]
rlabel metal3 14392 708904 14392 708904 0 FrameData[9]
rlabel metal2 2184 7714 2184 7714 0 FrameStrobe[0]
rlabel metal2 269976 602 269976 602 0 FrameStrobe[100]
rlabel metal2 272664 602 272664 602 0 FrameStrobe[101]
rlabel metal2 275352 602 275352 602 0 FrameStrobe[102]
rlabel metal2 278040 602 278040 602 0 FrameStrobe[103]
rlabel metal2 280728 602 280728 602 0 FrameStrobe[104]
rlabel metal2 283416 602 283416 602 0 FrameStrobe[105]
rlabel metal2 286104 602 286104 602 0 FrameStrobe[106]
rlabel metal2 288792 602 288792 602 0 FrameStrobe[107]
rlabel metal2 291480 602 291480 602 0 FrameStrobe[108]
rlabel metal2 294168 602 294168 602 0 FrameStrobe[109]
rlabel metal2 15624 7714 15624 7714 0 FrameStrobe[10]
rlabel metal2 296856 602 296856 602 0 FrameStrobe[110]
rlabel metal2 299544 602 299544 602 0 FrameStrobe[111]
rlabel metal2 302232 602 302232 602 0 FrameStrobe[112]
rlabel metal2 304920 602 304920 602 0 FrameStrobe[113]
rlabel metal2 307608 602 307608 602 0 FrameStrobe[114]
rlabel metal2 310296 602 310296 602 0 FrameStrobe[115]
rlabel metal2 312984 602 312984 602 0 FrameStrobe[116]
rlabel metal2 315672 602 315672 602 0 FrameStrobe[117]
rlabel metal2 318360 602 318360 602 0 FrameStrobe[118]
rlabel metal2 321048 602 321048 602 0 FrameStrobe[119]
rlabel metal2 16968 7714 16968 7714 0 FrameStrobe[11]
rlabel metal2 326984 602 326984 602 0 FrameStrobe[120]
rlabel metal2 329448 602 329448 602 0 FrameStrobe[121]
rlabel metal2 331912 602 331912 602 0 FrameStrobe[122]
rlabel metal2 334376 602 334376 602 0 FrameStrobe[123]
rlabel metal2 336840 602 336840 602 0 FrameStrobe[124]
rlabel metal2 339304 602 339304 602 0 FrameStrobe[125]
rlabel metal2 341768 602 341768 602 0 FrameStrobe[126]
rlabel metal2 344232 602 344232 602 0 FrameStrobe[127]
rlabel metal2 346696 602 346696 602 0 FrameStrobe[128]
rlabel metal2 349160 602 349160 602 0 FrameStrobe[129]
rlabel metal2 18312 7714 18312 7714 0 FrameStrobe[12]
rlabel metal2 351624 602 351624 602 0 FrameStrobe[130]
rlabel metal2 354088 602 354088 602 0 FrameStrobe[131]
rlabel metal2 356552 602 356552 602 0 FrameStrobe[132]
rlabel metal2 359016 602 359016 602 0 FrameStrobe[133]
rlabel metal2 361480 602 361480 602 0 FrameStrobe[134]
rlabel metal2 363944 602 363944 602 0 FrameStrobe[135]
rlabel metal2 366408 602 366408 602 0 FrameStrobe[136]
rlabel metal2 368872 602 368872 602 0 FrameStrobe[137]
rlabel metal2 371336 602 371336 602 0 FrameStrobe[138]
rlabel metal2 373800 602 373800 602 0 FrameStrobe[139]
rlabel metal2 19656 7714 19656 7714 0 FrameStrobe[13]
rlabel metal2 380184 602 380184 602 0 FrameStrobe[140]
rlabel metal2 382872 602 382872 602 0 FrameStrobe[141]
rlabel metal2 385560 602 385560 602 0 FrameStrobe[142]
rlabel metal2 388248 602 388248 602 0 FrameStrobe[143]
rlabel metal2 390936 602 390936 602 0 FrameStrobe[144]
rlabel metal2 393624 602 393624 602 0 FrameStrobe[145]
rlabel metal2 396312 602 396312 602 0 FrameStrobe[146]
rlabel metal2 399000 602 399000 602 0 FrameStrobe[147]
rlabel metal2 401688 602 401688 602 0 FrameStrobe[148]
rlabel metal2 404376 602 404376 602 0 FrameStrobe[149]
rlabel metal2 21000 7714 21000 7714 0 FrameStrobe[14]
rlabel metal2 407064 602 407064 602 0 FrameStrobe[150]
rlabel metal2 409752 602 409752 602 0 FrameStrobe[151]
rlabel metal2 412440 602 412440 602 0 FrameStrobe[152]
rlabel metal2 415128 602 415128 602 0 FrameStrobe[153]
rlabel metal2 417816 602 417816 602 0 FrameStrobe[154]
rlabel metal2 420504 602 420504 602 0 FrameStrobe[155]
rlabel metal2 423192 602 423192 602 0 FrameStrobe[156]
rlabel metal2 425880 602 425880 602 0 FrameStrobe[157]
rlabel metal2 428568 602 428568 602 0 FrameStrobe[158]
rlabel metal2 431256 602 431256 602 0 FrameStrobe[159]
rlabel metal2 22344 7714 22344 7714 0 FrameStrobe[15]
rlabel metal2 436744 602 436744 602 0 FrameStrobe[160]
rlabel metal2 438088 602 438088 602 0 FrameStrobe[161]
rlabel metal2 439432 602 439432 602 0 FrameStrobe[162]
rlabel metal2 440776 602 440776 602 0 FrameStrobe[163]
rlabel metal2 442120 602 442120 602 0 FrameStrobe[164]
rlabel metal2 443464 602 443464 602 0 FrameStrobe[165]
rlabel metal2 444808 602 444808 602 0 FrameStrobe[166]
rlabel metal2 446152 602 446152 602 0 FrameStrobe[167]
rlabel metal2 448280 126 448280 126 0 FrameStrobe[168]
rlabel metal2 448840 602 448840 602 0 FrameStrobe[169]
rlabel metal2 23688 7714 23688 7714 0 FrameStrobe[16]
rlabel metal2 450184 602 450184 602 0 FrameStrobe[170]
rlabel metal2 451528 602 451528 602 0 FrameStrobe[171]
rlabel metal2 452872 602 452872 602 0 FrameStrobe[172]
rlabel metal2 454216 602 454216 602 0 FrameStrobe[173]
rlabel metal2 455560 602 455560 602 0 FrameStrobe[174]
rlabel metal2 456904 602 456904 602 0 FrameStrobe[175]
rlabel metal2 458248 602 458248 602 0 FrameStrobe[176]
rlabel metal2 459592 602 459592 602 0 FrameStrobe[177]
rlabel metal2 460936 602 460936 602 0 FrameStrobe[178]
rlabel metal2 462280 602 462280 602 0 FrameStrobe[179]
rlabel metal2 25032 7714 25032 7714 0 FrameStrobe[17]
rlabel metal2 26376 7714 26376 7714 0 FrameStrobe[18]
rlabel metal2 27720 7714 27720 7714 0 FrameStrobe[19]
rlabel metal2 3528 7714 3528 7714 0 FrameStrobe[1]
rlabel metal2 46200 602 46200 602 0 FrameStrobe[20]
rlabel metal2 48216 602 48216 602 0 FrameStrobe[21]
rlabel metal2 50232 602 50232 602 0 FrameStrobe[22]
rlabel metal2 52248 602 52248 602 0 FrameStrobe[23]
rlabel metal2 54264 602 54264 602 0 FrameStrobe[24]
rlabel metal2 56280 602 56280 602 0 FrameStrobe[25]
rlabel metal2 58296 602 58296 602 0 FrameStrobe[26]
rlabel metal2 60312 602 60312 602 0 FrameStrobe[27]
rlabel metal2 62328 602 62328 602 0 FrameStrobe[28]
rlabel metal2 64344 602 64344 602 0 FrameStrobe[29]
rlabel metal2 4872 7714 4872 7714 0 FrameStrobe[2]
rlabel metal2 66360 602 66360 602 0 FrameStrobe[30]
rlabel metal2 68376 602 68376 602 0 FrameStrobe[31]
rlabel metal2 70392 602 70392 602 0 FrameStrobe[32]
rlabel metal2 72408 602 72408 602 0 FrameStrobe[33]
rlabel metal2 74424 602 74424 602 0 FrameStrobe[34]
rlabel metal2 76440 602 76440 602 0 FrameStrobe[35]
rlabel metal2 78456 602 78456 602 0 FrameStrobe[36]
rlabel metal2 80472 602 80472 602 0 FrameStrobe[37]
rlabel metal2 82488 602 82488 602 0 FrameStrobe[38]
rlabel metal2 84504 602 84504 602 0 FrameStrobe[39]
rlabel metal2 6216 7714 6216 7714 0 FrameStrobe[3]
rlabel metal2 90664 602 90664 602 0 FrameStrobe[40]
rlabel metal2 93352 602 93352 602 0 FrameStrobe[41]
rlabel metal2 96040 602 96040 602 0 FrameStrobe[42]
rlabel metal2 98728 602 98728 602 0 FrameStrobe[43]
rlabel metal2 101416 602 101416 602 0 FrameStrobe[44]
rlabel metal2 104104 602 104104 602 0 FrameStrobe[45]
rlabel metal2 106792 602 106792 602 0 FrameStrobe[46]
rlabel metal2 109480 602 109480 602 0 FrameStrobe[47]
rlabel metal2 112168 602 112168 602 0 FrameStrobe[48]
rlabel metal2 114856 602 114856 602 0 FrameStrobe[49]
rlabel metal2 7560 7714 7560 7714 0 FrameStrobe[4]
rlabel metal2 117544 602 117544 602 0 FrameStrobe[50]
rlabel metal2 120232 602 120232 602 0 FrameStrobe[51]
rlabel metal2 122920 602 122920 602 0 FrameStrobe[52]
rlabel metal2 125608 602 125608 602 0 FrameStrobe[53]
rlabel metal2 128296 602 128296 602 0 FrameStrobe[54]
rlabel metal2 130984 602 130984 602 0 FrameStrobe[55]
rlabel metal2 133672 602 133672 602 0 FrameStrobe[56]
rlabel metal2 136360 602 136360 602 0 FrameStrobe[57]
rlabel metal2 139048 602 139048 602 0 FrameStrobe[58]
rlabel metal2 141736 602 141736 602 0 FrameStrobe[59]
rlabel metal2 8904 7714 8904 7714 0 FrameStrobe[5]
rlabel metal2 148120 602 148120 602 0 FrameStrobe[60]
rlabel metal2 150808 602 150808 602 0 FrameStrobe[61]
rlabel metal2 153496 602 153496 602 0 FrameStrobe[62]
rlabel metal2 156184 602 156184 602 0 FrameStrobe[63]
rlabel metal2 158872 602 158872 602 0 FrameStrobe[64]
rlabel metal2 161560 602 161560 602 0 FrameStrobe[65]
rlabel metal2 164248 602 164248 602 0 FrameStrobe[66]
rlabel metal2 166936 602 166936 602 0 FrameStrobe[67]
rlabel metal2 169624 602 169624 602 0 FrameStrobe[68]
rlabel metal2 172312 602 172312 602 0 FrameStrobe[69]
rlabel metal2 10248 7714 10248 7714 0 FrameStrobe[6]
rlabel metal2 175000 602 175000 602 0 FrameStrobe[70]
rlabel metal2 177688 602 177688 602 0 FrameStrobe[71]
rlabel metal2 180376 602 180376 602 0 FrameStrobe[72]
rlabel metal2 183064 602 183064 602 0 FrameStrobe[73]
rlabel metal2 185752 602 185752 602 0 FrameStrobe[74]
rlabel metal2 188440 602 188440 602 0 FrameStrobe[75]
rlabel metal2 191128 602 191128 602 0 FrameStrobe[76]
rlabel metal2 193816 602 193816 602 0 FrameStrobe[77]
rlabel metal2 196504 602 196504 602 0 FrameStrobe[78]
rlabel metal2 199192 602 199192 602 0 FrameStrobe[79]
rlabel metal2 11592 7714 11592 7714 0 FrameStrobe[7]
rlabel metal2 206920 602 206920 602 0 FrameStrobe[80]
rlabel metal2 209832 602 209832 602 0 FrameStrobe[81]
rlabel metal2 212744 602 212744 602 0 FrameStrobe[82]
rlabel metal2 215656 602 215656 602 0 FrameStrobe[83]
rlabel metal2 218568 602 218568 602 0 FrameStrobe[84]
rlabel metal2 221480 602 221480 602 0 FrameStrobe[85]
rlabel metal2 224392 602 224392 602 0 FrameStrobe[86]
rlabel metal2 227304 602 227304 602 0 FrameStrobe[87]
rlabel metal2 230216 602 230216 602 0 FrameStrobe[88]
rlabel metal2 233128 602 233128 602 0 FrameStrobe[89]
rlabel metal2 12936 7714 12936 7714 0 FrameStrobe[8]
rlabel metal2 236040 602 236040 602 0 FrameStrobe[90]
rlabel metal2 238952 602 238952 602 0 FrameStrobe[91]
rlabel metal2 241864 602 241864 602 0 FrameStrobe[92]
rlabel metal2 244776 602 244776 602 0 FrameStrobe[93]
rlabel metal2 247688 602 247688 602 0 FrameStrobe[94]
rlabel metal2 250600 602 250600 602 0 FrameStrobe[95]
rlabel metal2 253512 602 253512 602 0 FrameStrobe[96]
rlabel metal2 256424 602 256424 602 0 FrameStrobe[97]
rlabel metal2 259336 602 259336 602 0 FrameStrobe[98]
rlabel metal2 262248 602 262248 602 0 FrameStrobe[99]
rlabel metal2 14280 7714 14280 7714 0 FrameStrobe[9]
rlabel metal3 112 133448 112 133448 0 Tile_X0Y10_A_I_top
rlabel metal3 112 132552 112 132552 0 Tile_X0Y10_A_O_top
rlabel metal3 112 134344 112 134344 0 Tile_X0Y10_A_T_top
rlabel metal3 112 143304 112 143304 0 Tile_X0Y10_A_config_C_bit0
rlabel metal3 112 144200 112 144200 0 Tile_X0Y10_A_config_C_bit1
rlabel metal3 112 145096 112 145096 0 Tile_X0Y10_A_config_C_bit2
rlabel metal3 112 145992 112 145992 0 Tile_X0Y10_A_config_C_bit3
rlabel metal3 112 136136 112 136136 0 Tile_X0Y10_B_I_top
rlabel metal3 112 135240 112 135240 0 Tile_X0Y10_B_O_top
rlabel metal3 112 137032 112 137032 0 Tile_X0Y10_B_T_top
rlabel metal3 112 146888 112 146888 0 Tile_X0Y10_B_config_C_bit0
rlabel metal3 112 147784 112 147784 0 Tile_X0Y10_B_config_C_bit1
rlabel metal3 112 148680 112 148680 0 Tile_X0Y10_B_config_C_bit2
rlabel metal3 112 149576 112 149576 0 Tile_X0Y10_B_config_C_bit3
rlabel metal3 112 138824 112 138824 0 Tile_X0Y10_C_I_top
rlabel metal3 112 137928 112 137928 0 Tile_X0Y10_C_O_top
rlabel metal3 112 139720 112 139720 0 Tile_X0Y10_C_T_top
rlabel metal3 112 150472 112 150472 0 Tile_X0Y10_C_config_C_bit0
rlabel metal3 112 151368 112 151368 0 Tile_X0Y10_C_config_C_bit1
rlabel metal3 112 152264 112 152264 0 Tile_X0Y10_C_config_C_bit2
rlabel metal3 112 153160 112 153160 0 Tile_X0Y10_C_config_C_bit3
rlabel metal3 112 141512 112 141512 0 Tile_X0Y10_D_I_top
rlabel metal3 112 140616 112 140616 0 Tile_X0Y10_D_O_top
rlabel metal3 112 142408 112 142408 0 Tile_X0Y10_D_T_top
rlabel metal3 112 154056 112 154056 0 Tile_X0Y10_D_config_C_bit0
rlabel metal3 112 154952 112 154952 0 Tile_X0Y10_D_config_C_bit1
rlabel metal3 112 155848 112 155848 0 Tile_X0Y10_D_config_C_bit2
rlabel metal3 112 156744 112 156744 0 Tile_X0Y10_D_config_C_bit3
rlabel metal3 112 75992 112 75992 0 Tile_X0Y11_A_I_top
rlabel metal3 112 75096 112 75096 0 Tile_X0Y11_A_O_top
rlabel metal3 112 76888 112 76888 0 Tile_X0Y11_A_T_top
rlabel metal3 112 85848 112 85848 0 Tile_X0Y11_A_config_C_bit0
rlabel metal3 112 86744 112 86744 0 Tile_X0Y11_A_config_C_bit1
rlabel metal3 112 87640 112 87640 0 Tile_X0Y11_A_config_C_bit2
rlabel metal3 112 88536 112 88536 0 Tile_X0Y11_A_config_C_bit3
rlabel metal3 112 78680 112 78680 0 Tile_X0Y11_B_I_top
rlabel metal3 112 77784 112 77784 0 Tile_X0Y11_B_O_top
rlabel metal3 112 79576 112 79576 0 Tile_X0Y11_B_T_top
rlabel metal3 112 89432 112 89432 0 Tile_X0Y11_B_config_C_bit0
rlabel metal3 112 90328 112 90328 0 Tile_X0Y11_B_config_C_bit1
rlabel metal3 112 91224 112 91224 0 Tile_X0Y11_B_config_C_bit2
rlabel metal3 112 92120 112 92120 0 Tile_X0Y11_B_config_C_bit3
rlabel metal3 112 81368 112 81368 0 Tile_X0Y11_C_I_top
rlabel metal3 112 80472 112 80472 0 Tile_X0Y11_C_O_top
rlabel metal3 112 82264 112 82264 0 Tile_X0Y11_C_T_top
rlabel metal3 112 93016 112 93016 0 Tile_X0Y11_C_config_C_bit0
rlabel metal3 112 93912 112 93912 0 Tile_X0Y11_C_config_C_bit1
rlabel metal3 112 94808 112 94808 0 Tile_X0Y11_C_config_C_bit2
rlabel metal3 112 95704 112 95704 0 Tile_X0Y11_C_config_C_bit3
rlabel metal3 112 84056 112 84056 0 Tile_X0Y11_D_I_top
rlabel metal3 112 83160 112 83160 0 Tile_X0Y11_D_O_top
rlabel metal3 112 84952 112 84952 0 Tile_X0Y11_D_T_top
rlabel metal3 112 96600 112 96600 0 Tile_X0Y11_D_config_C_bit0
rlabel metal3 112 97496 112 97496 0 Tile_X0Y11_D_config_C_bit1
rlabel metal3 112 98392 112 98392 0 Tile_X0Y11_D_config_C_bit2
rlabel metal3 112 99288 112 99288 0 Tile_X0Y11_D_config_C_bit3
rlabel metal3 112 18536 112 18536 0 Tile_X0Y12_A_I_top
rlabel metal3 112 17640 112 17640 0 Tile_X0Y12_A_O_top
rlabel metal3 112 19432 112 19432 0 Tile_X0Y12_A_T_top
rlabel metal3 112 28392 112 28392 0 Tile_X0Y12_A_config_C_bit0
rlabel metal3 112 29288 112 29288 0 Tile_X0Y12_A_config_C_bit1
rlabel metal3 112 30184 112 30184 0 Tile_X0Y12_A_config_C_bit2
rlabel metal3 112 31080 112 31080 0 Tile_X0Y12_A_config_C_bit3
rlabel metal3 112 21224 112 21224 0 Tile_X0Y12_B_I_top
rlabel metal3 112 20328 112 20328 0 Tile_X0Y12_B_O_top
rlabel metal3 112 22120 112 22120 0 Tile_X0Y12_B_T_top
rlabel metal3 112 31976 112 31976 0 Tile_X0Y12_B_config_C_bit0
rlabel metal3 112 32872 112 32872 0 Tile_X0Y12_B_config_C_bit1
rlabel metal3 112 33768 112 33768 0 Tile_X0Y12_B_config_C_bit2
rlabel metal3 112 34664 112 34664 0 Tile_X0Y12_B_config_C_bit3
rlabel metal3 112 23912 112 23912 0 Tile_X0Y12_C_I_top
rlabel metal3 112 23016 112 23016 0 Tile_X0Y12_C_O_top
rlabel metal3 112 24808 112 24808 0 Tile_X0Y12_C_T_top
rlabel metal3 112 35560 112 35560 0 Tile_X0Y12_C_config_C_bit0
rlabel metal3 112 36456 112 36456 0 Tile_X0Y12_C_config_C_bit1
rlabel metal3 112 37352 112 37352 0 Tile_X0Y12_C_config_C_bit2
rlabel metal3 112 38248 112 38248 0 Tile_X0Y12_C_config_C_bit3
rlabel metal3 112 26600 112 26600 0 Tile_X0Y12_D_I_top
rlabel metal3 112 25704 112 25704 0 Tile_X0Y12_D_O_top
rlabel metal3 112 27496 112 27496 0 Tile_X0Y12_D_T_top
rlabel metal3 112 39144 112 39144 0 Tile_X0Y12_D_config_C_bit0
rlabel metal3 112 40040 112 40040 0 Tile_X0Y12_D_config_C_bit1
rlabel metal3 112 40936 112 40936 0 Tile_X0Y12_D_config_C_bit2
rlabel metal3 112 41832 112 41832 0 Tile_X0Y12_D_config_C_bit3
rlabel metal3 112 650552 112 650552 0 Tile_X0Y1_A_I_top
rlabel metal3 112 649656 112 649656 0 Tile_X0Y1_A_O_top
rlabel metal3 112 651448 112 651448 0 Tile_X0Y1_A_T_top
rlabel metal3 112 660408 112 660408 0 Tile_X0Y1_A_config_C_bit0
rlabel metal3 112 661304 112 661304 0 Tile_X0Y1_A_config_C_bit1
rlabel metal3 112 662200 112 662200 0 Tile_X0Y1_A_config_C_bit2
rlabel metal3 112 663096 112 663096 0 Tile_X0Y1_A_config_C_bit3
rlabel metal3 112 653240 112 653240 0 Tile_X0Y1_B_I_top
rlabel metal3 112 652344 112 652344 0 Tile_X0Y1_B_O_top
rlabel metal3 112 654136 112 654136 0 Tile_X0Y1_B_T_top
rlabel metal3 112 663992 112 663992 0 Tile_X0Y1_B_config_C_bit0
rlabel metal3 112 664888 112 664888 0 Tile_X0Y1_B_config_C_bit1
rlabel metal3 112 665784 112 665784 0 Tile_X0Y1_B_config_C_bit2
rlabel metal3 112 666680 112 666680 0 Tile_X0Y1_B_config_C_bit3
rlabel metal3 112 655928 112 655928 0 Tile_X0Y1_C_I_top
rlabel metal3 112 655032 112 655032 0 Tile_X0Y1_C_O_top
rlabel metal3 112 656824 112 656824 0 Tile_X0Y1_C_T_top
rlabel metal3 112 667576 112 667576 0 Tile_X0Y1_C_config_C_bit0
rlabel metal3 112 668472 112 668472 0 Tile_X0Y1_C_config_C_bit1
rlabel metal3 112 669368 112 669368 0 Tile_X0Y1_C_config_C_bit2
rlabel metal3 112 670264 112 670264 0 Tile_X0Y1_C_config_C_bit3
rlabel metal3 112 658616 112 658616 0 Tile_X0Y1_D_I_top
rlabel metal3 112 657720 112 657720 0 Tile_X0Y1_D_O_top
rlabel metal3 112 659512 112 659512 0 Tile_X0Y1_D_T_top
rlabel metal3 112 671160 112 671160 0 Tile_X0Y1_D_config_C_bit0
rlabel metal3 112 672056 112 672056 0 Tile_X0Y1_D_config_C_bit1
rlabel metal3 112 672952 112 672952 0 Tile_X0Y1_D_config_C_bit2
rlabel metal3 112 673848 112 673848 0 Tile_X0Y1_D_config_C_bit3
rlabel metal3 112 593096 112 593096 0 Tile_X0Y2_A_I_top
rlabel metal3 112 592200 112 592200 0 Tile_X0Y2_A_O_top
rlabel metal3 112 593992 112 593992 0 Tile_X0Y2_A_T_top
rlabel metal3 112 602952 112 602952 0 Tile_X0Y2_A_config_C_bit0
rlabel metal3 112 603848 112 603848 0 Tile_X0Y2_A_config_C_bit1
rlabel metal3 112 604744 112 604744 0 Tile_X0Y2_A_config_C_bit2
rlabel metal3 112 605640 112 605640 0 Tile_X0Y2_A_config_C_bit3
rlabel metal3 112 595784 112 595784 0 Tile_X0Y2_B_I_top
rlabel metal3 112 594888 112 594888 0 Tile_X0Y2_B_O_top
rlabel metal3 112 596680 112 596680 0 Tile_X0Y2_B_T_top
rlabel metal3 112 606536 112 606536 0 Tile_X0Y2_B_config_C_bit0
rlabel metal3 112 607432 112 607432 0 Tile_X0Y2_B_config_C_bit1
rlabel metal3 112 608328 112 608328 0 Tile_X0Y2_B_config_C_bit2
rlabel metal3 112 609224 112 609224 0 Tile_X0Y2_B_config_C_bit3
rlabel metal3 112 598472 112 598472 0 Tile_X0Y2_C_I_top
rlabel metal3 112 597576 112 597576 0 Tile_X0Y2_C_O_top
rlabel metal3 112 599368 112 599368 0 Tile_X0Y2_C_T_top
rlabel metal3 112 610120 112 610120 0 Tile_X0Y2_C_config_C_bit0
rlabel metal3 112 611016 112 611016 0 Tile_X0Y2_C_config_C_bit1
rlabel metal3 112 611912 112 611912 0 Tile_X0Y2_C_config_C_bit2
rlabel metal3 112 612808 112 612808 0 Tile_X0Y2_C_config_C_bit3
rlabel metal3 112 601160 112 601160 0 Tile_X0Y2_D_I_top
rlabel metal3 112 600264 112 600264 0 Tile_X0Y2_D_O_top
rlabel metal3 112 602056 112 602056 0 Tile_X0Y2_D_T_top
rlabel metal3 112 613704 112 613704 0 Tile_X0Y2_D_config_C_bit0
rlabel metal3 112 614600 112 614600 0 Tile_X0Y2_D_config_C_bit1
rlabel metal3 112 615496 112 615496 0 Tile_X0Y2_D_config_C_bit2
rlabel metal3 112 616392 112 616392 0 Tile_X0Y2_D_config_C_bit3
rlabel metal3 112 535640 112 535640 0 Tile_X0Y3_A_I_top
rlabel metal3 112 534744 112 534744 0 Tile_X0Y3_A_O_top
rlabel metal3 112 536536 112 536536 0 Tile_X0Y3_A_T_top
rlabel metal3 112 545496 112 545496 0 Tile_X0Y3_A_config_C_bit0
rlabel metal3 112 546392 112 546392 0 Tile_X0Y3_A_config_C_bit1
rlabel metal3 112 547288 112 547288 0 Tile_X0Y3_A_config_C_bit2
rlabel metal3 112 548184 112 548184 0 Tile_X0Y3_A_config_C_bit3
rlabel metal3 112 538328 112 538328 0 Tile_X0Y3_B_I_top
rlabel metal3 112 537432 112 537432 0 Tile_X0Y3_B_O_top
rlabel metal3 112 539224 112 539224 0 Tile_X0Y3_B_T_top
rlabel metal3 112 549080 112 549080 0 Tile_X0Y3_B_config_C_bit0
rlabel metal3 112 549976 112 549976 0 Tile_X0Y3_B_config_C_bit1
rlabel metal3 112 550872 112 550872 0 Tile_X0Y3_B_config_C_bit2
rlabel metal3 112 551768 112 551768 0 Tile_X0Y3_B_config_C_bit3
rlabel metal3 112 541016 112 541016 0 Tile_X0Y3_C_I_top
rlabel metal3 112 540120 112 540120 0 Tile_X0Y3_C_O_top
rlabel metal3 112 541912 112 541912 0 Tile_X0Y3_C_T_top
rlabel metal3 112 552664 112 552664 0 Tile_X0Y3_C_config_C_bit0
rlabel metal3 112 553560 112 553560 0 Tile_X0Y3_C_config_C_bit1
rlabel metal3 112 554456 112 554456 0 Tile_X0Y3_C_config_C_bit2
rlabel metal3 112 555352 112 555352 0 Tile_X0Y3_C_config_C_bit3
rlabel metal3 112 543704 112 543704 0 Tile_X0Y3_D_I_top
rlabel metal3 112 542808 112 542808 0 Tile_X0Y3_D_O_top
rlabel metal3 112 544600 112 544600 0 Tile_X0Y3_D_T_top
rlabel metal3 112 556248 112 556248 0 Tile_X0Y3_D_config_C_bit0
rlabel metal3 112 557144 112 557144 0 Tile_X0Y3_D_config_C_bit1
rlabel metal3 112 558040 112 558040 0 Tile_X0Y3_D_config_C_bit2
rlabel metal3 112 558936 112 558936 0 Tile_X0Y3_D_config_C_bit3
rlabel metal3 112 478184 112 478184 0 Tile_X0Y4_A_I_top
rlabel metal3 112 477288 112 477288 0 Tile_X0Y4_A_O_top
rlabel metal3 112 479080 112 479080 0 Tile_X0Y4_A_T_top
rlabel metal3 112 488040 112 488040 0 Tile_X0Y4_A_config_C_bit0
rlabel metal3 112 488936 112 488936 0 Tile_X0Y4_A_config_C_bit1
rlabel metal3 112 489832 112 489832 0 Tile_X0Y4_A_config_C_bit2
rlabel metal3 112 490728 112 490728 0 Tile_X0Y4_A_config_C_bit3
rlabel metal3 112 480872 112 480872 0 Tile_X0Y4_B_I_top
rlabel metal3 112 479976 112 479976 0 Tile_X0Y4_B_O_top
rlabel metal3 112 481768 112 481768 0 Tile_X0Y4_B_T_top
rlabel metal3 112 491624 112 491624 0 Tile_X0Y4_B_config_C_bit0
rlabel metal3 112 492520 112 492520 0 Tile_X0Y4_B_config_C_bit1
rlabel metal3 112 493416 112 493416 0 Tile_X0Y4_B_config_C_bit2
rlabel metal3 112 494312 112 494312 0 Tile_X0Y4_B_config_C_bit3
rlabel metal3 112 483560 112 483560 0 Tile_X0Y4_C_I_top
rlabel metal3 112 482664 112 482664 0 Tile_X0Y4_C_O_top
rlabel metal3 112 484456 112 484456 0 Tile_X0Y4_C_T_top
rlabel metal3 112 495208 112 495208 0 Tile_X0Y4_C_config_C_bit0
rlabel metal3 112 496104 112 496104 0 Tile_X0Y4_C_config_C_bit1
rlabel metal3 112 497000 112 497000 0 Tile_X0Y4_C_config_C_bit2
rlabel metal3 112 497896 112 497896 0 Tile_X0Y4_C_config_C_bit3
rlabel metal3 112 486248 112 486248 0 Tile_X0Y4_D_I_top
rlabel metal3 112 485352 112 485352 0 Tile_X0Y4_D_O_top
rlabel metal3 112 487144 112 487144 0 Tile_X0Y4_D_T_top
rlabel metal3 112 498792 112 498792 0 Tile_X0Y4_D_config_C_bit0
rlabel metal3 112 499688 112 499688 0 Tile_X0Y4_D_config_C_bit1
rlabel metal3 112 500584 112 500584 0 Tile_X0Y4_D_config_C_bit2
rlabel metal3 112 501480 112 501480 0 Tile_X0Y4_D_config_C_bit3
rlabel metal3 112 420728 112 420728 0 Tile_X0Y5_A_I_top
rlabel metal3 112 419832 112 419832 0 Tile_X0Y5_A_O_top
rlabel metal3 112 421624 112 421624 0 Tile_X0Y5_A_T_top
rlabel metal3 112 430584 112 430584 0 Tile_X0Y5_A_config_C_bit0
rlabel metal3 112 431480 112 431480 0 Tile_X0Y5_A_config_C_bit1
rlabel metal3 112 432376 112 432376 0 Tile_X0Y5_A_config_C_bit2
rlabel metal3 112 433272 112 433272 0 Tile_X0Y5_A_config_C_bit3
rlabel metal3 112 423416 112 423416 0 Tile_X0Y5_B_I_top
rlabel metal3 112 422520 112 422520 0 Tile_X0Y5_B_O_top
rlabel metal3 112 424312 112 424312 0 Tile_X0Y5_B_T_top
rlabel metal3 112 434168 112 434168 0 Tile_X0Y5_B_config_C_bit0
rlabel metal3 112 435064 112 435064 0 Tile_X0Y5_B_config_C_bit1
rlabel metal3 112 435960 112 435960 0 Tile_X0Y5_B_config_C_bit2
rlabel metal3 112 436856 112 436856 0 Tile_X0Y5_B_config_C_bit3
rlabel metal3 112 426104 112 426104 0 Tile_X0Y5_C_I_top
rlabel metal3 112 425208 112 425208 0 Tile_X0Y5_C_O_top
rlabel metal3 112 427000 112 427000 0 Tile_X0Y5_C_T_top
rlabel metal3 112 437752 112 437752 0 Tile_X0Y5_C_config_C_bit0
rlabel metal3 112 438648 112 438648 0 Tile_X0Y5_C_config_C_bit1
rlabel metal3 112 439544 112 439544 0 Tile_X0Y5_C_config_C_bit2
rlabel metal3 112 440440 112 440440 0 Tile_X0Y5_C_config_C_bit3
rlabel metal3 112 428792 112 428792 0 Tile_X0Y5_D_I_top
rlabel metal3 112 427896 112 427896 0 Tile_X0Y5_D_O_top
rlabel metal3 112 429688 112 429688 0 Tile_X0Y5_D_T_top
rlabel metal3 112 441336 112 441336 0 Tile_X0Y5_D_config_C_bit0
rlabel metal3 112 442232 112 442232 0 Tile_X0Y5_D_config_C_bit1
rlabel metal3 112 443128 112 443128 0 Tile_X0Y5_D_config_C_bit2
rlabel metal3 112 444024 112 444024 0 Tile_X0Y5_D_config_C_bit3
rlabel metal3 112 363272 112 363272 0 Tile_X0Y6_A_I_top
rlabel metal3 112 362376 112 362376 0 Tile_X0Y6_A_O_top
rlabel metal3 112 364168 112 364168 0 Tile_X0Y6_A_T_top
rlabel metal3 112 373128 112 373128 0 Tile_X0Y6_A_config_C_bit0
rlabel metal3 112 374024 112 374024 0 Tile_X0Y6_A_config_C_bit1
rlabel metal3 112 374920 112 374920 0 Tile_X0Y6_A_config_C_bit2
rlabel metal3 112 375816 112 375816 0 Tile_X0Y6_A_config_C_bit3
rlabel metal3 112 365960 112 365960 0 Tile_X0Y6_B_I_top
rlabel metal3 112 365064 112 365064 0 Tile_X0Y6_B_O_top
rlabel metal3 112 366856 112 366856 0 Tile_X0Y6_B_T_top
rlabel metal3 112 376712 112 376712 0 Tile_X0Y6_B_config_C_bit0
rlabel metal3 112 377608 112 377608 0 Tile_X0Y6_B_config_C_bit1
rlabel metal3 112 378504 112 378504 0 Tile_X0Y6_B_config_C_bit2
rlabel metal3 112 379400 112 379400 0 Tile_X0Y6_B_config_C_bit3
rlabel metal3 112 368648 112 368648 0 Tile_X0Y6_C_I_top
rlabel metal3 112 367752 112 367752 0 Tile_X0Y6_C_O_top
rlabel metal3 112 369544 112 369544 0 Tile_X0Y6_C_T_top
rlabel metal3 112 380296 112 380296 0 Tile_X0Y6_C_config_C_bit0
rlabel metal3 112 381192 112 381192 0 Tile_X0Y6_C_config_C_bit1
rlabel metal3 112 382088 112 382088 0 Tile_X0Y6_C_config_C_bit2
rlabel metal3 112 382984 112 382984 0 Tile_X0Y6_C_config_C_bit3
rlabel metal3 112 371336 112 371336 0 Tile_X0Y6_D_I_top
rlabel metal3 112 370440 112 370440 0 Tile_X0Y6_D_O_top
rlabel metal3 112 372232 112 372232 0 Tile_X0Y6_D_T_top
rlabel metal3 112 383880 112 383880 0 Tile_X0Y6_D_config_C_bit0
rlabel metal3 112 384776 112 384776 0 Tile_X0Y6_D_config_C_bit1
rlabel metal3 112 385672 112 385672 0 Tile_X0Y6_D_config_C_bit2
rlabel metal3 112 386568 112 386568 0 Tile_X0Y6_D_config_C_bit3
rlabel metal3 112 305816 112 305816 0 Tile_X0Y7_A_I_top
rlabel metal3 112 304920 112 304920 0 Tile_X0Y7_A_O_top
rlabel metal3 112 306712 112 306712 0 Tile_X0Y7_A_T_top
rlabel metal3 112 315672 112 315672 0 Tile_X0Y7_A_config_C_bit0
rlabel metal3 112 316568 112 316568 0 Tile_X0Y7_A_config_C_bit1
rlabel metal3 112 317464 112 317464 0 Tile_X0Y7_A_config_C_bit2
rlabel metal3 112 318360 112 318360 0 Tile_X0Y7_A_config_C_bit3
rlabel metal3 112 308504 112 308504 0 Tile_X0Y7_B_I_top
rlabel metal3 112 307608 112 307608 0 Tile_X0Y7_B_O_top
rlabel metal3 112 309400 112 309400 0 Tile_X0Y7_B_T_top
rlabel metal3 112 319256 112 319256 0 Tile_X0Y7_B_config_C_bit0
rlabel metal3 112 320152 112 320152 0 Tile_X0Y7_B_config_C_bit1
rlabel metal3 112 321048 112 321048 0 Tile_X0Y7_B_config_C_bit2
rlabel metal3 112 321944 112 321944 0 Tile_X0Y7_B_config_C_bit3
rlabel metal3 112 311192 112 311192 0 Tile_X0Y7_C_I_top
rlabel metal3 112 310296 112 310296 0 Tile_X0Y7_C_O_top
rlabel metal3 112 312088 112 312088 0 Tile_X0Y7_C_T_top
rlabel metal3 112 322840 112 322840 0 Tile_X0Y7_C_config_C_bit0
rlabel metal3 112 323736 112 323736 0 Tile_X0Y7_C_config_C_bit1
rlabel metal3 112 324632 112 324632 0 Tile_X0Y7_C_config_C_bit2
rlabel metal3 112 325528 112 325528 0 Tile_X0Y7_C_config_C_bit3
rlabel metal3 112 313880 112 313880 0 Tile_X0Y7_D_I_top
rlabel metal3 112 312984 112 312984 0 Tile_X0Y7_D_O_top
rlabel metal3 112 314776 112 314776 0 Tile_X0Y7_D_T_top
rlabel metal3 112 326424 112 326424 0 Tile_X0Y7_D_config_C_bit0
rlabel metal3 112 327320 112 327320 0 Tile_X0Y7_D_config_C_bit1
rlabel metal3 112 328216 112 328216 0 Tile_X0Y7_D_config_C_bit2
rlabel metal3 112 329112 112 329112 0 Tile_X0Y7_D_config_C_bit3
rlabel metal3 112 248360 112 248360 0 Tile_X0Y8_A_I_top
rlabel metal3 112 247464 112 247464 0 Tile_X0Y8_A_O_top
rlabel metal3 112 249256 112 249256 0 Tile_X0Y8_A_T_top
rlabel metal3 112 258216 112 258216 0 Tile_X0Y8_A_config_C_bit0
rlabel metal3 112 259112 112 259112 0 Tile_X0Y8_A_config_C_bit1
rlabel metal3 112 260008 112 260008 0 Tile_X0Y8_A_config_C_bit2
rlabel metal3 112 260904 112 260904 0 Tile_X0Y8_A_config_C_bit3
rlabel metal3 112 251048 112 251048 0 Tile_X0Y8_B_I_top
rlabel metal3 112 250152 112 250152 0 Tile_X0Y8_B_O_top
rlabel metal3 112 251944 112 251944 0 Tile_X0Y8_B_T_top
rlabel metal3 112 261800 112 261800 0 Tile_X0Y8_B_config_C_bit0
rlabel metal3 112 262696 112 262696 0 Tile_X0Y8_B_config_C_bit1
rlabel metal3 112 263592 112 263592 0 Tile_X0Y8_B_config_C_bit2
rlabel metal3 112 264488 112 264488 0 Tile_X0Y8_B_config_C_bit3
rlabel metal3 112 253736 112 253736 0 Tile_X0Y8_C_I_top
rlabel metal3 112 252840 112 252840 0 Tile_X0Y8_C_O_top
rlabel metal3 112 254632 112 254632 0 Tile_X0Y8_C_T_top
rlabel metal3 112 265384 112 265384 0 Tile_X0Y8_C_config_C_bit0
rlabel metal3 112 266280 112 266280 0 Tile_X0Y8_C_config_C_bit1
rlabel metal3 112 267176 112 267176 0 Tile_X0Y8_C_config_C_bit2
rlabel metal3 112 268072 112 268072 0 Tile_X0Y8_C_config_C_bit3
rlabel metal3 112 256424 112 256424 0 Tile_X0Y8_D_I_top
rlabel metal3 112 255528 112 255528 0 Tile_X0Y8_D_O_top
rlabel metal3 112 257320 112 257320 0 Tile_X0Y8_D_T_top
rlabel metal3 112 268968 112 268968 0 Tile_X0Y8_D_config_C_bit0
rlabel metal3 112 269864 112 269864 0 Tile_X0Y8_D_config_C_bit1
rlabel metal3 112 270760 112 270760 0 Tile_X0Y8_D_config_C_bit2
rlabel metal3 112 271656 112 271656 0 Tile_X0Y8_D_config_C_bit3
rlabel metal3 112 190904 112 190904 0 Tile_X0Y9_A_I_top
rlabel metal3 112 190008 112 190008 0 Tile_X0Y9_A_O_top
rlabel metal3 112 191800 112 191800 0 Tile_X0Y9_A_T_top
rlabel metal3 112 200760 112 200760 0 Tile_X0Y9_A_config_C_bit0
rlabel metal3 112 201656 112 201656 0 Tile_X0Y9_A_config_C_bit1
rlabel metal3 112 202552 112 202552 0 Tile_X0Y9_A_config_C_bit2
rlabel metal3 112 203448 112 203448 0 Tile_X0Y9_A_config_C_bit3
rlabel metal3 112 193592 112 193592 0 Tile_X0Y9_B_I_top
rlabel metal3 112 192696 112 192696 0 Tile_X0Y9_B_O_top
rlabel metal3 112 194488 112 194488 0 Tile_X0Y9_B_T_top
rlabel metal3 112 204344 112 204344 0 Tile_X0Y9_B_config_C_bit0
rlabel metal3 112 205240 112 205240 0 Tile_X0Y9_B_config_C_bit1
rlabel metal3 112 206136 112 206136 0 Tile_X0Y9_B_config_C_bit2
rlabel metal3 112 207032 112 207032 0 Tile_X0Y9_B_config_C_bit3
rlabel metal3 112 196280 112 196280 0 Tile_X0Y9_C_I_top
rlabel metal3 112 195384 112 195384 0 Tile_X0Y9_C_O_top
rlabel metal3 112 197176 112 197176 0 Tile_X0Y9_C_T_top
rlabel metal3 112 207928 112 207928 0 Tile_X0Y9_C_config_C_bit0
rlabel metal3 112 208824 112 208824 0 Tile_X0Y9_C_config_C_bit1
rlabel metal3 112 209720 112 209720 0 Tile_X0Y9_C_config_C_bit2
rlabel metal3 112 210616 112 210616 0 Tile_X0Y9_C_config_C_bit3
rlabel metal3 112 198968 112 198968 0 Tile_X0Y9_D_I_top
rlabel metal3 112 198072 112 198072 0 Tile_X0Y9_D_O_top
rlabel metal3 112 199864 112 199864 0 Tile_X0Y9_D_T_top
rlabel metal3 112 211512 112 211512 0 Tile_X0Y9_D_config_C_bit0
rlabel metal3 112 212408 112 212408 0 Tile_X0Y9_D_config_C_bit1
rlabel metal3 112 213304 112 213304 0 Tile_X0Y9_D_config_C_bit2
rlabel metal3 112 214200 112 214200 0 Tile_X0Y9_D_config_C_bit3
rlabel metal2 42168 602 42168 602 0 Tile_X1Y13_BOOT_top
rlabel metal2 32088 602 32088 602 0 Tile_X1Y13_CONFIGURED_top
rlabel metal2 30072 602 30072 602 0 Tile_X1Y13_RESET_top
rlabel metal2 34104 602 34104 602 0 Tile_X1Y13_SLOT_top0
rlabel metal2 36120 602 36120 602 0 Tile_X1Y13_SLOT_top1
rlabel metal2 38136 602 38136 602 0 Tile_X1Y13_SLOT_top2
rlabel metal2 40152 602 40152 602 0 Tile_X1Y13_SLOT_top3
rlabel metal3 464814 150248 464814 150248 0 Tile_X8Y10_A_SRAM0
rlabel metal3 464814 151144 464814 151144 0 Tile_X8Y10_A_SRAM1
rlabel metal3 464814 152040 464814 152040 0 Tile_X8Y10_A_SRAM2
rlabel metal3 464814 152936 464814 152936 0 Tile_X8Y10_A_SRAM3
rlabel metal3 464814 153832 464814 153832 0 Tile_X8Y10_A_SRAM4
rlabel metal3 464814 154728 464814 154728 0 Tile_X8Y10_A_SRAM5
rlabel metal3 464814 155624 464814 155624 0 Tile_X8Y10_A_SRAM6
rlabel metal3 464814 156520 464814 156520 0 Tile_X8Y10_A_SRAM7
rlabel metal3 464814 157416 464814 157416 0 Tile_X8Y10_A_SRAM8
rlabel metal3 464814 141288 464814 141288 0 Tile_X8Y10_CEN_SRAM
rlabel metal3 464814 165480 464814 165480 0 Tile_X8Y10_CLK_SRAM
rlabel metal3 464814 140392 464814 140392 0 Tile_X8Y10_CONFIGURED_top
rlabel metal3 464814 158312 464814 158312 0 Tile_X8Y10_D_SRAM0
rlabel metal3 464814 159208 464814 159208 0 Tile_X8Y10_D_SRAM1
rlabel metal3 464814 160104 464814 160104 0 Tile_X8Y10_D_SRAM2
rlabel metal3 464814 161000 464814 161000 0 Tile_X8Y10_D_SRAM3
rlabel metal3 464814 161896 464814 161896 0 Tile_X8Y10_D_SRAM4
rlabel metal3 464814 162792 464814 162792 0 Tile_X8Y10_D_SRAM5
rlabel metal3 464814 163688 464814 163688 0 Tile_X8Y10_D_SRAM6
rlabel metal3 464814 164584 464814 164584 0 Tile_X8Y10_D_SRAM7
rlabel metal3 464814 142184 464814 142184 0 Tile_X8Y10_GWEN_SRAM
rlabel metal3 464814 133224 464814 133224 0 Tile_X8Y10_Q_SRAM0
rlabel metal3 464814 134120 464814 134120 0 Tile_X8Y10_Q_SRAM1
rlabel metal3 464814 135016 464814 135016 0 Tile_X8Y10_Q_SRAM2
rlabel metal3 464814 135912 464814 135912 0 Tile_X8Y10_Q_SRAM3
rlabel metal3 464814 136808 464814 136808 0 Tile_X8Y10_Q_SRAM4
rlabel metal3 464814 137704 464814 137704 0 Tile_X8Y10_Q_SRAM5
rlabel metal3 464814 138600 464814 138600 0 Tile_X8Y10_Q_SRAM6
rlabel metal3 464814 139496 464814 139496 0 Tile_X8Y10_Q_SRAM7
rlabel metal3 464814 143080 464814 143080 0 Tile_X8Y10_WEN_SRAM0
rlabel metal3 464814 143976 464814 143976 0 Tile_X8Y10_WEN_SRAM1
rlabel metal3 464814 144872 464814 144872 0 Tile_X8Y10_WEN_SRAM2
rlabel metal3 464814 145768 464814 145768 0 Tile_X8Y10_WEN_SRAM3
rlabel metal3 464814 146664 464814 146664 0 Tile_X8Y10_WEN_SRAM4
rlabel metal3 464814 147560 464814 147560 0 Tile_X8Y10_WEN_SRAM5
rlabel metal3 464814 148456 464814 148456 0 Tile_X8Y10_WEN_SRAM6
rlabel metal3 464814 149352 464814 149352 0 Tile_X8Y10_WEN_SRAM7
rlabel metal3 464814 35336 464814 35336 0 Tile_X8Y12_A_SRAM0
rlabel metal3 464814 36232 464814 36232 0 Tile_X8Y12_A_SRAM1
rlabel metal3 464814 37128 464814 37128 0 Tile_X8Y12_A_SRAM2
rlabel metal3 464814 38024 464814 38024 0 Tile_X8Y12_A_SRAM3
rlabel metal3 464814 38920 464814 38920 0 Tile_X8Y12_A_SRAM4
rlabel metal3 464814 39816 464814 39816 0 Tile_X8Y12_A_SRAM5
rlabel metal3 464814 40712 464814 40712 0 Tile_X8Y12_A_SRAM6
rlabel metal3 464814 41608 464814 41608 0 Tile_X8Y12_A_SRAM7
rlabel metal3 464814 42504 464814 42504 0 Tile_X8Y12_A_SRAM8
rlabel metal3 464814 26376 464814 26376 0 Tile_X8Y12_CEN_SRAM
rlabel metal3 464814 50568 464814 50568 0 Tile_X8Y12_CLK_SRAM
rlabel metal3 464814 25480 464814 25480 0 Tile_X8Y12_CONFIGURED_top
rlabel metal3 464814 43400 464814 43400 0 Tile_X8Y12_D_SRAM0
rlabel metal3 464814 44296 464814 44296 0 Tile_X8Y12_D_SRAM1
rlabel metal3 464814 45192 464814 45192 0 Tile_X8Y12_D_SRAM2
rlabel metal3 464814 46088 464814 46088 0 Tile_X8Y12_D_SRAM3
rlabel metal3 464814 46984 464814 46984 0 Tile_X8Y12_D_SRAM4
rlabel metal3 464814 47880 464814 47880 0 Tile_X8Y12_D_SRAM5
rlabel metal3 464814 48776 464814 48776 0 Tile_X8Y12_D_SRAM6
rlabel metal3 464814 49672 464814 49672 0 Tile_X8Y12_D_SRAM7
rlabel metal3 464814 27272 464814 27272 0 Tile_X8Y12_GWEN_SRAM
rlabel metal3 464814 18312 464814 18312 0 Tile_X8Y12_Q_SRAM0
rlabel metal3 464814 19208 464814 19208 0 Tile_X8Y12_Q_SRAM1
rlabel metal3 464814 20104 464814 20104 0 Tile_X8Y12_Q_SRAM2
rlabel metal3 464814 21000 464814 21000 0 Tile_X8Y12_Q_SRAM3
rlabel metal3 464814 21896 464814 21896 0 Tile_X8Y12_Q_SRAM4
rlabel metal3 464814 22792 464814 22792 0 Tile_X8Y12_Q_SRAM5
rlabel metal3 464814 23688 464814 23688 0 Tile_X8Y12_Q_SRAM6
rlabel metal3 464814 24584 464814 24584 0 Tile_X8Y12_Q_SRAM7
rlabel metal3 464814 28168 464814 28168 0 Tile_X8Y12_WEN_SRAM0
rlabel metal3 464814 29064 464814 29064 0 Tile_X8Y12_WEN_SRAM1
rlabel metal3 464814 29960 464814 29960 0 Tile_X8Y12_WEN_SRAM2
rlabel metal3 464814 30856 464814 30856 0 Tile_X8Y12_WEN_SRAM3
rlabel metal3 464814 31752 464814 31752 0 Tile_X8Y12_WEN_SRAM4
rlabel metal3 464814 32648 464814 32648 0 Tile_X8Y12_WEN_SRAM5
rlabel metal3 464814 33544 464814 33544 0 Tile_X8Y12_WEN_SRAM6
rlabel metal3 464814 34440 464814 34440 0 Tile_X8Y12_WEN_SRAM7
rlabel metal3 464814 609896 464814 609896 0 Tile_X8Y2_A_SRAM0
rlabel metal3 464814 610792 464814 610792 0 Tile_X8Y2_A_SRAM1
rlabel metal3 464814 611688 464814 611688 0 Tile_X8Y2_A_SRAM2
rlabel metal3 464814 612584 464814 612584 0 Tile_X8Y2_A_SRAM3
rlabel metal3 464814 613480 464814 613480 0 Tile_X8Y2_A_SRAM4
rlabel metal3 464814 614376 464814 614376 0 Tile_X8Y2_A_SRAM5
rlabel metal3 464814 615272 464814 615272 0 Tile_X8Y2_A_SRAM6
rlabel metal3 464814 616168 464814 616168 0 Tile_X8Y2_A_SRAM7
rlabel metal3 464814 617064 464814 617064 0 Tile_X8Y2_A_SRAM8
rlabel metal3 464814 600936 464814 600936 0 Tile_X8Y2_CEN_SRAM
rlabel metal3 464814 625128 464814 625128 0 Tile_X8Y2_CLK_SRAM
rlabel metal3 464814 600040 464814 600040 0 Tile_X8Y2_CONFIGURED_top
rlabel metal3 464814 617960 464814 617960 0 Tile_X8Y2_D_SRAM0
rlabel metal3 464814 618856 464814 618856 0 Tile_X8Y2_D_SRAM1
rlabel metal3 464814 619752 464814 619752 0 Tile_X8Y2_D_SRAM2
rlabel metal3 464814 620648 464814 620648 0 Tile_X8Y2_D_SRAM3
rlabel metal3 464814 621544 464814 621544 0 Tile_X8Y2_D_SRAM4
rlabel metal3 464814 622440 464814 622440 0 Tile_X8Y2_D_SRAM5
rlabel metal3 464814 623336 464814 623336 0 Tile_X8Y2_D_SRAM6
rlabel metal3 464814 624232 464814 624232 0 Tile_X8Y2_D_SRAM7
rlabel metal3 464814 601832 464814 601832 0 Tile_X8Y2_GWEN_SRAM
rlabel metal3 464814 592872 464814 592872 0 Tile_X8Y2_Q_SRAM0
rlabel metal3 464814 593768 464814 593768 0 Tile_X8Y2_Q_SRAM1
rlabel metal3 464814 594664 464814 594664 0 Tile_X8Y2_Q_SRAM2
rlabel metal3 464814 595560 464814 595560 0 Tile_X8Y2_Q_SRAM3
rlabel metal3 464814 596456 464814 596456 0 Tile_X8Y2_Q_SRAM4
rlabel metal3 464814 597352 464814 597352 0 Tile_X8Y2_Q_SRAM5
rlabel metal3 464814 598248 464814 598248 0 Tile_X8Y2_Q_SRAM6
rlabel metal3 464814 599144 464814 599144 0 Tile_X8Y2_Q_SRAM7
rlabel metal3 464814 602728 464814 602728 0 Tile_X8Y2_WEN_SRAM0
rlabel metal3 464814 603624 464814 603624 0 Tile_X8Y2_WEN_SRAM1
rlabel metal3 464814 604520 464814 604520 0 Tile_X8Y2_WEN_SRAM2
rlabel metal3 464814 605416 464814 605416 0 Tile_X8Y2_WEN_SRAM3
rlabel metal3 464814 606312 464814 606312 0 Tile_X8Y2_WEN_SRAM4
rlabel metal3 464814 607208 464814 607208 0 Tile_X8Y2_WEN_SRAM5
rlabel metal3 464814 608104 464814 608104 0 Tile_X8Y2_WEN_SRAM6
rlabel metal3 464814 609000 464814 609000 0 Tile_X8Y2_WEN_SRAM7
rlabel metal3 464814 494984 464814 494984 0 Tile_X8Y4_A_SRAM0
rlabel metal3 464814 495880 464814 495880 0 Tile_X8Y4_A_SRAM1
rlabel metal3 464814 496776 464814 496776 0 Tile_X8Y4_A_SRAM2
rlabel metal3 464814 497672 464814 497672 0 Tile_X8Y4_A_SRAM3
rlabel metal3 464814 498568 464814 498568 0 Tile_X8Y4_A_SRAM4
rlabel metal3 464814 499464 464814 499464 0 Tile_X8Y4_A_SRAM5
rlabel metal3 464814 500360 464814 500360 0 Tile_X8Y4_A_SRAM6
rlabel metal3 464814 501256 464814 501256 0 Tile_X8Y4_A_SRAM7
rlabel metal3 464814 502152 464814 502152 0 Tile_X8Y4_A_SRAM8
rlabel metal3 464814 486024 464814 486024 0 Tile_X8Y4_CEN_SRAM
rlabel metal3 464814 510216 464814 510216 0 Tile_X8Y4_CLK_SRAM
rlabel metal3 464814 485128 464814 485128 0 Tile_X8Y4_CONFIGURED_top
rlabel metal3 464814 503048 464814 503048 0 Tile_X8Y4_D_SRAM0
rlabel metal3 464814 503944 464814 503944 0 Tile_X8Y4_D_SRAM1
rlabel metal3 464814 504840 464814 504840 0 Tile_X8Y4_D_SRAM2
rlabel metal3 464814 505736 464814 505736 0 Tile_X8Y4_D_SRAM3
rlabel metal3 464814 506632 464814 506632 0 Tile_X8Y4_D_SRAM4
rlabel metal3 464814 507528 464814 507528 0 Tile_X8Y4_D_SRAM5
rlabel metal3 464814 508424 464814 508424 0 Tile_X8Y4_D_SRAM6
rlabel metal3 464814 509320 464814 509320 0 Tile_X8Y4_D_SRAM7
rlabel metal3 464814 486920 464814 486920 0 Tile_X8Y4_GWEN_SRAM
rlabel metal3 464814 477960 464814 477960 0 Tile_X8Y4_Q_SRAM0
rlabel metal3 464814 478856 464814 478856 0 Tile_X8Y4_Q_SRAM1
rlabel metal3 464814 479752 464814 479752 0 Tile_X8Y4_Q_SRAM2
rlabel metal3 464814 480648 464814 480648 0 Tile_X8Y4_Q_SRAM3
rlabel metal3 464814 481544 464814 481544 0 Tile_X8Y4_Q_SRAM4
rlabel metal3 464814 482440 464814 482440 0 Tile_X8Y4_Q_SRAM5
rlabel metal3 464814 483336 464814 483336 0 Tile_X8Y4_Q_SRAM6
rlabel metal3 464814 484232 464814 484232 0 Tile_X8Y4_Q_SRAM7
rlabel metal3 464814 487816 464814 487816 0 Tile_X8Y4_WEN_SRAM0
rlabel metal3 464814 488712 464814 488712 0 Tile_X8Y4_WEN_SRAM1
rlabel metal3 464814 489608 464814 489608 0 Tile_X8Y4_WEN_SRAM2
rlabel metal3 464814 490504 464814 490504 0 Tile_X8Y4_WEN_SRAM3
rlabel metal3 464814 491400 464814 491400 0 Tile_X8Y4_WEN_SRAM4
rlabel metal3 464814 492296 464814 492296 0 Tile_X8Y4_WEN_SRAM5
rlabel metal3 464814 493192 464814 493192 0 Tile_X8Y4_WEN_SRAM6
rlabel metal3 464814 494088 464814 494088 0 Tile_X8Y4_WEN_SRAM7
rlabel metal3 464814 380072 464814 380072 0 Tile_X8Y6_A_SRAM0
rlabel metal3 464814 380968 464814 380968 0 Tile_X8Y6_A_SRAM1
rlabel metal3 464814 381864 464814 381864 0 Tile_X8Y6_A_SRAM2
rlabel metal3 464814 382760 464814 382760 0 Tile_X8Y6_A_SRAM3
rlabel metal3 464814 383656 464814 383656 0 Tile_X8Y6_A_SRAM4
rlabel metal3 464814 384552 464814 384552 0 Tile_X8Y6_A_SRAM5
rlabel metal3 464814 385448 464814 385448 0 Tile_X8Y6_A_SRAM6
rlabel metal3 464814 386344 464814 386344 0 Tile_X8Y6_A_SRAM7
rlabel metal3 464814 387240 464814 387240 0 Tile_X8Y6_A_SRAM8
rlabel metal3 464814 371112 464814 371112 0 Tile_X8Y6_CEN_SRAM
rlabel metal3 464814 395304 464814 395304 0 Tile_X8Y6_CLK_SRAM
rlabel metal3 464814 370216 464814 370216 0 Tile_X8Y6_CONFIGURED_top
rlabel metal3 464814 388136 464814 388136 0 Tile_X8Y6_D_SRAM0
rlabel metal3 464814 389032 464814 389032 0 Tile_X8Y6_D_SRAM1
rlabel metal3 464814 389928 464814 389928 0 Tile_X8Y6_D_SRAM2
rlabel metal3 464814 390824 464814 390824 0 Tile_X8Y6_D_SRAM3
rlabel metal3 464814 391720 464814 391720 0 Tile_X8Y6_D_SRAM4
rlabel metal3 464814 392616 464814 392616 0 Tile_X8Y6_D_SRAM5
rlabel metal3 464814 393512 464814 393512 0 Tile_X8Y6_D_SRAM6
rlabel metal3 464814 394408 464814 394408 0 Tile_X8Y6_D_SRAM7
rlabel metal3 464814 372008 464814 372008 0 Tile_X8Y6_GWEN_SRAM
rlabel metal3 464814 363048 464814 363048 0 Tile_X8Y6_Q_SRAM0
rlabel metal3 464814 363944 464814 363944 0 Tile_X8Y6_Q_SRAM1
rlabel metal3 464814 364840 464814 364840 0 Tile_X8Y6_Q_SRAM2
rlabel metal3 464814 365736 464814 365736 0 Tile_X8Y6_Q_SRAM3
rlabel metal3 464814 366632 464814 366632 0 Tile_X8Y6_Q_SRAM4
rlabel metal3 464814 367528 464814 367528 0 Tile_X8Y6_Q_SRAM5
rlabel metal3 464814 368424 464814 368424 0 Tile_X8Y6_Q_SRAM6
rlabel metal3 464814 369320 464814 369320 0 Tile_X8Y6_Q_SRAM7
rlabel metal3 464814 372904 464814 372904 0 Tile_X8Y6_WEN_SRAM0
rlabel metal3 464814 373800 464814 373800 0 Tile_X8Y6_WEN_SRAM1
rlabel metal3 464814 374696 464814 374696 0 Tile_X8Y6_WEN_SRAM2
rlabel metal3 464814 375592 464814 375592 0 Tile_X8Y6_WEN_SRAM3
rlabel metal3 464814 376488 464814 376488 0 Tile_X8Y6_WEN_SRAM4
rlabel metal3 464814 377384 464814 377384 0 Tile_X8Y6_WEN_SRAM5
rlabel metal3 464814 378280 464814 378280 0 Tile_X8Y6_WEN_SRAM6
rlabel metal3 464814 379176 464814 379176 0 Tile_X8Y6_WEN_SRAM7
rlabel metal3 464814 265160 464814 265160 0 Tile_X8Y8_A_SRAM0
rlabel metal3 464814 266056 464814 266056 0 Tile_X8Y8_A_SRAM1
rlabel metal3 464814 266952 464814 266952 0 Tile_X8Y8_A_SRAM2
rlabel metal3 464814 267848 464814 267848 0 Tile_X8Y8_A_SRAM3
rlabel metal3 464814 268744 464814 268744 0 Tile_X8Y8_A_SRAM4
rlabel metal3 464814 269640 464814 269640 0 Tile_X8Y8_A_SRAM5
rlabel metal3 464814 270536 464814 270536 0 Tile_X8Y8_A_SRAM6
rlabel metal3 464814 271432 464814 271432 0 Tile_X8Y8_A_SRAM7
rlabel metal3 464814 272328 464814 272328 0 Tile_X8Y8_A_SRAM8
rlabel metal3 464814 256200 464814 256200 0 Tile_X8Y8_CEN_SRAM
rlabel metal3 464814 280392 464814 280392 0 Tile_X8Y8_CLK_SRAM
rlabel metal3 464814 255304 464814 255304 0 Tile_X8Y8_CONFIGURED_top
rlabel metal3 464814 273224 464814 273224 0 Tile_X8Y8_D_SRAM0
rlabel metal3 464814 274120 464814 274120 0 Tile_X8Y8_D_SRAM1
rlabel metal3 464814 275016 464814 275016 0 Tile_X8Y8_D_SRAM2
rlabel metal3 464814 275912 464814 275912 0 Tile_X8Y8_D_SRAM3
rlabel metal3 464814 276808 464814 276808 0 Tile_X8Y8_D_SRAM4
rlabel metal3 464814 277704 464814 277704 0 Tile_X8Y8_D_SRAM5
rlabel metal3 464814 278600 464814 278600 0 Tile_X8Y8_D_SRAM6
rlabel metal3 464814 279496 464814 279496 0 Tile_X8Y8_D_SRAM7
rlabel metal3 464814 257096 464814 257096 0 Tile_X8Y8_GWEN_SRAM
rlabel metal3 464814 248136 464814 248136 0 Tile_X8Y8_Q_SRAM0
rlabel metal3 464814 249032 464814 249032 0 Tile_X8Y8_Q_SRAM1
rlabel metal3 464814 249928 464814 249928 0 Tile_X8Y8_Q_SRAM2
rlabel metal3 464814 250824 464814 250824 0 Tile_X8Y8_Q_SRAM3
rlabel metal3 464814 251720 464814 251720 0 Tile_X8Y8_Q_SRAM4
rlabel metal3 464814 252616 464814 252616 0 Tile_X8Y8_Q_SRAM5
rlabel metal3 464814 253512 464814 253512 0 Tile_X8Y8_Q_SRAM6
rlabel metal3 464814 254408 464814 254408 0 Tile_X8Y8_Q_SRAM7
rlabel metal3 464814 257992 464814 257992 0 Tile_X8Y8_WEN_SRAM0
rlabel metal3 464814 258888 464814 258888 0 Tile_X8Y8_WEN_SRAM1
rlabel metal3 464814 259784 464814 259784 0 Tile_X8Y8_WEN_SRAM2
rlabel metal3 464814 260680 464814 260680 0 Tile_X8Y8_WEN_SRAM3
rlabel metal3 464814 261576 464814 261576 0 Tile_X8Y8_WEN_SRAM4
rlabel metal3 464814 262472 464814 262472 0 Tile_X8Y8_WEN_SRAM5
rlabel metal3 464814 263368 464814 263368 0 Tile_X8Y8_WEN_SRAM6
rlabel metal3 464814 264264 464814 264264 0 Tile_X8Y8_WEN_SRAM7
rlabel metal2 44212 1036 44212 1036 0 UserCLK
<< properties >>
string FIXED_BBOX 0 0 464912 719152
<< end >>
