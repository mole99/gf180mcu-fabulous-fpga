// Copyright 2025 Leo Moser
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

(* blackbox, keep *)
module OBI_PERIPHERAL (
    output REQ,
    output WE,
    
    output BE0,
    output BE1,
    output BE2,
    output BE3,
    
    output ADDR0,
    output ADDR1,
    output ADDR2,
    output ADDR3,
    output ADDR4,
    output ADDR5,
    output ADDR6,
    output ADDR7,
    output ADDR8,
    output ADDR9,
    output ADDR10,
    output ADDR11,
    output ADDR12,
    output ADDR13,
    output ADDR14,
    output ADDR15,
    output ADDR16,
    output ADDR17,
    output ADDR18,
    output ADDR19,
    output ADDR20,
    output ADDR21,
    output ADDR22,
    output ADDR23,

    output WDATA0,
    output WDATA1,
    output WDATA2,
    output WDATA3,
    output WDATA4,
    output WDATA5,
    output WDATA6,
    output WDATA7,
    output WDATA8,
    output WDATA9,
    output WDATA10,
    output WDATA11,
    output WDATA12,
    output WDATA13,
    output WDATA14,
    output WDATA15,
    output WDATA16,
    output WDATA17,
    output WDATA18,
    output WDATA19,
    output WDATA20,
    output WDATA21,
    output WDATA22,
    output WDATA23,
    output WDATA24,
    output WDATA25,
    output WDATA26,
    output WDATA27,
    output WDATA28,
    output WDATA29,
    output WDATA30,
    output WDATA31,
    
    input  GNT,
    input  RVALID,
    
    input  RDATA0,
    input  RDATA1,
    input  RDATA2,
    input  RDATA3,
    input  RDATA4,
    input  RDATA5,
    input  RDATA6,
    input  RDATA7,
    input  RDATA8,
    input  RDATA9,
    input  RDATA10,
    input  RDATA11,
    input  RDATA12,
    input  RDATA13,
    input  RDATA14,
    input  RDATA15,
    input  RDATA16,
    input  RDATA17,
    input  RDATA18,
    input  RDATA19,
    input  RDATA20,
    input  RDATA21,
    input  RDATA22,
    input  RDATA23,
    input  RDATA24,
    input  RDATA25,
    input  RDATA26,
    input  RDATA27,
    input  RDATA28,
    input  RDATA29,
    input  RDATA30,
    input  RDATA31
);

endmodule

(* blackbox, keep *)
module CUSTOM_INSTRUCTION (
    input  ISSUE_READY,
    input  ISSUE_ACCEPT,
    output ISSUE_VALID,
    
    output ISSUE_INSTR0,
    output ISSUE_INSTR1,
    output ISSUE_INSTR2,
    output ISSUE_INSTR3,
    output ISSUE_INSTR4,
    output ISSUE_INSTR5,
    output ISSUE_INSTR6,
    output ISSUE_INSTR7,
    output ISSUE_INSTR8,
    output ISSUE_INSTR9,
    output ISSUE_INSTR10,
    output ISSUE_INSTR11,
    output ISSUE_INSTR12,
    output ISSUE_INSTR13,
    output ISSUE_INSTR14,
    output ISSUE_INSTR15,
    output ISSUE_INSTR16,
    output ISSUE_INSTR17,
    output ISSUE_INSTR18,
    output ISSUE_INSTR19,
    output ISSUE_INSTR20,
    output ISSUE_INSTR21,
    output ISSUE_INSTR22,
    output ISSUE_INSTR23,
    output ISSUE_INSTR24,
    output ISSUE_INSTR25,
    output ISSUE_INSTR26,
    output ISSUE_INSTR27,
    output ISSUE_INSTR28,
    output ISSUE_INSTR29,
    output ISSUE_INSTR30,
    output ISSUE_INSTR31,

    output ISSUE_OPA0,
    output ISSUE_OPA1,
    output ISSUE_OPA2,
    output ISSUE_OPA3,
    output ISSUE_OPA4,
    output ISSUE_OPA5,
    output ISSUE_OPA6,
    output ISSUE_OPA7,
    output ISSUE_OPA8,
    output ISSUE_OPA9,
    output ISSUE_OPA10,
    output ISSUE_OPA11,
    output ISSUE_OPA12,
    output ISSUE_OPA13,
    output ISSUE_OPA14,
    output ISSUE_OPA15,
    output ISSUE_OPA16,
    output ISSUE_OPA17,
    output ISSUE_OPA18,
    output ISSUE_OPA19,
    output ISSUE_OPA20,
    output ISSUE_OPA21,
    output ISSUE_OPA22,
    output ISSUE_OPA23,
    output ISSUE_OPA24,
    output ISSUE_OPA25,
    output ISSUE_OPA26,
    output ISSUE_OPA27,
    output ISSUE_OPA28,
    output ISSUE_OPA29,
    output ISSUE_OPA30,
    output ISSUE_OPA31,
    
    output ISSUE_OPB0,
    output ISSUE_OPB1,
    output ISSUE_OPB2,
    output ISSUE_OPB3,
    output ISSUE_OPB4,
    output ISSUE_OPB5,
    output ISSUE_OPB6,
    output ISSUE_OPB7,
    output ISSUE_OPB8,
    output ISSUE_OPB9,
    output ISSUE_OPB10,
    output ISSUE_OPB11,
    output ISSUE_OPB12,
    output ISSUE_OPB13,
    output ISSUE_OPB14,
    output ISSUE_OPB15,
    output ISSUE_OPB16,
    output ISSUE_OPB17,
    output ISSUE_OPB18,
    output ISSUE_OPB19,
    output ISSUE_OPB20,
    output ISSUE_OPB21,
    output ISSUE_OPB22,
    output ISSUE_OPB23,
    output ISSUE_OPB24,
    output ISSUE_OPB25,
    output ISSUE_OPB26,
    output ISSUE_OPB27,
    output ISSUE_OPB28,
    output ISSUE_OPB29,
    output ISSUE_OPB30,
    output ISSUE_OPB31,
    
    output ISSUE_ID0,
    output ISSUE_ID1,
    output ISSUE_ID2,
    output ISSUE_ID3,
    
    input  RESULT_VALID,

    input RESULT_ID0,
    input RESULT_ID1,
    input RESULT_ID2,
    input RESULT_ID3,

    input RESULT_RD0,
    input RESULT_RD1,
    input RESULT_RD2,
    input RESULT_RD3,
    input RESULT_RD4,

    input RESULT0,
    input RESULT1,
    input RESULT2,
    input RESULT3,
    input RESULT4,
    input RESULT5,
    input RESULT6,
    input RESULT7,
    input RESULT8,
    input RESULT9,
    input RESULT10,
    input RESULT11,
    input RESULT12,
    input RESULT13,
    input RESULT14,
    input RESULT15,
    input RESULT16,
    input RESULT17,
    input RESULT18,
    input RESULT19,
    input RESULT20,
    input RESULT21,
    input RESULT22,
    input RESULT23,
    input RESULT24,
    input RESULT25,
    input RESULT26,
    input RESULT27,
    input RESULT28,
    input RESULT29,
    input RESULT30,
    input RESULT31
);

endmodule

(* blackbox *)
module IHP_BRAM_1024x16 (
    input  A_ADDR0,
    input  A_ADDR1,
    input  A_ADDR2,
    input  A_ADDR3,
    input  A_ADDR4,
    input  A_ADDR5,
    input  A_ADDR6,
    input  A_ADDR7,
    input  A_ADDR8,
    input  A_ADDR9,

    input  A_BM0,
    input  A_BM1,
    input  A_BM2,
    input  A_BM3,
    input  A_BM4,
    input  A_BM5,
    input  A_BM6,
    input  A_BM7,
    input  A_BM8,
    input  A_BM9,
    input  A_BM10,
    input  A_BM11,
    input  A_BM12,
    input  A_BM13,
    input  A_BM14,
    input  A_BM15,

    input  A_DIN0,
    input  A_DIN1,
    input  A_DIN2,
    input  A_DIN3,
    input  A_DIN4,
    input  A_DIN5,
    input  A_DIN6,
    input  A_DIN7,
    input  A_DIN8,
    input  A_DIN9,
    input  A_DIN10,
    input  A_DIN11,
    input  A_DIN12,
    input  A_DIN13,
    input  A_DIN14,
    input  A_DIN15,

    input  A_WEN,
    input  A_MEN,
    input  A_REN,

    output A_DOUT0,
    output A_DOUT1,
    output A_DOUT2,
    output A_DOUT3,
    output A_DOUT4,
    output A_DOUT5,
    output A_DOUT6,
    output A_DOUT7,
    output A_DOUT8,
    output A_DOUT9,
    output A_DOUT10,
    output A_DOUT11,
    output A_DOUT12,
    output A_DOUT13,
    output A_DOUT14,
    output A_DOUT15,

    input  B_ADDR0,
    input  B_ADDR1,
    input  B_ADDR2,
    input  B_ADDR3,
    input  B_ADDR4,
    input  B_ADDR5,
    input  B_ADDR6,
    input  B_ADDR7,
    input  B_ADDR8,
    input  B_ADDR9,

    input  B_BM0,
    input  B_BM1,
    input  B_BM2,
    input  B_BM3,
    input  B_BM4,
    input  B_BM5,
    input  B_BM6,
    input  B_BM7,
    input  B_BM8,
    input  B_BM9,
    input  B_BM10,
    input  B_BM11,
    input  B_BM12,
    input  B_BM13,
    input  B_BM14,
    input  B_BM15,

    input  B_DIN0,
    input  B_DIN1,
    input  B_DIN2,
    input  B_DIN3,
    input  B_DIN4,
    input  B_DIN5,
    input  B_DIN6,
    input  B_DIN7,
    input  B_DIN8,
    input  B_DIN9,
    input  B_DIN10,
    input  B_DIN11,
    input  B_DIN12,
    input  B_DIN13,
    input  B_DIN14,
    input  B_DIN15,

    input  B_WEN,
    input  B_MEN,
    input  B_REN,

    output B_DOUT0,
    output B_DOUT1,
    output B_DOUT2,
    output B_DOUT3,
    output B_DOUT4,
    output B_DOUT5,
    output B_DOUT6,
    output B_DOUT7,
    output B_DOUT8,
    output B_DOUT9,
    output B_DOUT10,
    output B_DOUT11,
    output B_DOUT12,
    output B_DOUT13,
    output B_DOUT14,
    output B_DOUT15
);

endmodule

(* blackbox *)
module IHP_SRAM_1024x32 (
    input  A_ADDR0,
    input  A_ADDR1,
    input  A_ADDR2,
    input  A_ADDR3,
    input  A_ADDR4,
    input  A_ADDR5,
    input  A_ADDR6,
    input  A_ADDR7,
    input  A_ADDR8,
    input  A_ADDR9,

    input  A_BM0,
    input  A_BM1,
    input  A_BM2,
    input  A_BM3,
    input  A_BM4,
    input  A_BM5,
    input  A_BM6,
    input  A_BM7,
    input  A_BM8,
    input  A_BM9,
    input  A_BM10,
    input  A_BM11,
    input  A_BM12,
    input  A_BM13,
    input  A_BM14,
    input  A_BM15,
    input  A_BM16,
    input  A_BM17,
    input  A_BM18,
    input  A_BM19,
    input  A_BM20,
    input  A_BM21,
    input  A_BM22,
    input  A_BM23,
    input  A_BM24,
    input  A_BM25,
    input  A_BM26,
    input  A_BM27,
    input  A_BM28,
    input  A_BM29,
    input  A_BM30,
    input  A_BM31,

    input  A_DIN0,
    input  A_DIN1,
    input  A_DIN2,
    input  A_DIN3,
    input  A_DIN4,
    input  A_DIN5,
    input  A_DIN6,
    input  A_DIN7,
    input  A_DIN8,
    input  A_DIN9,
    input  A_DIN10,
    input  A_DIN11,
    input  A_DIN12,
    input  A_DIN13,
    input  A_DIN14,
    input  A_DIN15,
    input  A_DIN16,
    input  A_DIN17,
    input  A_DIN18,
    input  A_DIN19,
    input  A_DIN20,
    input  A_DIN21,
    input  A_DIN22,
    input  A_DIN23,
    input  A_DIN24,
    input  A_DIN25,
    input  A_DIN26,
    input  A_DIN27,
    input  A_DIN28,
    input  A_DIN29,
    input  A_DIN30,
    input  A_DIN31,

    input  A_WEN,
    input  A_MEN,
    input  A_REN,

    output A_DOUT0,
    output A_DOUT1,
    output A_DOUT2,
    output A_DOUT3,
    output A_DOUT4,
    output A_DOUT5,
    output A_DOUT6,
    output A_DOUT7,
    output A_DOUT8,
    output A_DOUT9,
    output A_DOUT10,
    output A_DOUT11,
    output A_DOUT12,
    output A_DOUT13,
    output A_DOUT14,
    output A_DOUT15,
    output A_DOUT16,
    output A_DOUT17,
    output A_DOUT18,
    output A_DOUT19,
    output A_DOUT20,
    output A_DOUT21,
    output A_DOUT22,
    output A_DOUT23,
    output A_DOUT24,
    output A_DOUT25,
    output A_DOUT26,
    output A_DOUT27,
    output A_DOUT28,
    output A_DOUT29,
    output A_DOUT30,
    output A_DOUT31
);

endmodule

(* blackbox, keep *)
module WARMBOOT (
    input  SLOT0,
    input  SLOT1,
    input  SLOT2,
    input  SLOT3,
    input  BOOT,
    output RESET
);

endmodule

(* blackbox, keep *)
module CPU_IRQ (
    input  IRQ0,
    input  IRQ1,
    input  IRQ2,
    input  IRQ3
);

endmodule

(* blackbox *)
module MULADD #(
    parameter A_reg=0,
    parameter B_reg=0,
    parameter C_reg=0,
    parameter signExtension=0,
    parameter ACC=0,
    parameter ACCout=0
)(
    input A0,
    input A1,
    input A2,
    input A3,
    input A4,
    input A5,
    input A6,
    input A7,
    
    input B0,
    input B1,
    input B2,
    input B3,
    input B4,
    input B5,
    input B6,
    input B7,
    
    input C0,
    input C1,
    input C2,
    input C3,
    input C4,
    input C5,
    input C6,
    input C7,
    input C8,
    input C9,
    input C10,
    input C11,
    input C12,
    input C13,
    input C14,
    input C15,
    input C16,
    input C17,
    input C18,
    input C19,
    
    input clr,
    
    output Q0,
    output Q1,
    output Q2,
    output Q3,
    output Q4,
    output Q5,
    output Q6,
    output Q7,
    output Q8,
    output Q9,
    output Q10,
    output Q11,
    output Q12,
    output Q13,
    output Q14,
    output Q15,
    output Q16,
    output Q17,
    output Q18,
    output Q19
);

endmodule
