// Copyright 2025 Leo Moser
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module OBI_PERIPHERAL_wrapper (
    output        REQ,
    output        WE,
    output [3: 0] BE,
    output [23:0] ADDR,
    output [31:0] WDATA,
    
    input         GNT,
    input         RVALID,
    input  [31:0] RDATA,
);

    OBI_PERIPHERAL i_OBI_PERIPHERAL (
        .REQ    (REQ),
        .WE     (WE),

        .BE0    (BE[0]),
        .BE1    (BE[1]),
        .BE2    (BE[2]),
        .BE3    (BE[3]),

        .ADDR0    (ADDR[0]),
        .ADDR1    (ADDR[1]),
        .ADDR2    (ADDR[2]),
        .ADDR3    (ADDR[3]),
        .ADDR4    (ADDR[4]),
        .ADDR5    (ADDR[5]),
        .ADDR6    (ADDR[6]),
        .ADDR7    (ADDR[7]),
        .ADDR8    (ADDR[8]),
        .ADDR9    (ADDR[9]),
        .ADDR10    (ADDR[10]),
        .ADDR11    (ADDR[11]),
        .ADDR12    (ADDR[12]),
        .ADDR13    (ADDR[13]),
        .ADDR14    (ADDR[14]),
        .ADDR15    (ADDR[15]),
        .ADDR16    (ADDR[16]),
        .ADDR17    (ADDR[17]),
        .ADDR18    (ADDR[18]),
        .ADDR19    (ADDR[19]),
        .ADDR20    (ADDR[20]),
        .ADDR21    (ADDR[21]),
        .ADDR22    (ADDR[22]),
        .ADDR23    (ADDR[23]),
        
        .WDATA0    (WDATA[0]),
        .WDATA1    (WDATA[1]),
        .WDATA2    (WDATA[2]),
        .WDATA3    (WDATA[3]),
        .WDATA4    (WDATA[4]),
        .WDATA5    (WDATA[5]),
        .WDATA6    (WDATA[6]),
        .WDATA7    (WDATA[7]),
        .WDATA8    (WDATA[8]),
        .WDATA9    (WDATA[9]),
        .WDATA10    (WDATA[10]),
        .WDATA11    (WDATA[11]),
        .WDATA12    (WDATA[12]),
        .WDATA13    (WDATA[13]),
        .WDATA14    (WDATA[14]),
        .WDATA15    (WDATA[15]),
        .WDATA16    (WDATA[16]),
        .WDATA17    (WDATA[17]),
        .WDATA18    (WDATA[18]),
        .WDATA19    (WDATA[19]),
        .WDATA20    (WDATA[20]),
        .WDATA21    (WDATA[21]),
        .WDATA22    (WDATA[22]),
        .WDATA23    (WDATA[23]),
        .WDATA24    (WDATA[24]),
        .WDATA25    (WDATA[25]),
        .WDATA26    (WDATA[26]),
        .WDATA27    (WDATA[27]),
        .WDATA28    (WDATA[28]),
        .WDATA29    (WDATA[29]),
        .WDATA30    (WDATA[30]),
        .WDATA31    (WDATA[31]),

        .GNT        (GNT),
        .RVALID     (RVALID),

        .RDATA0    (RDATA[0]),
        .RDATA1    (RDATA[1]),
        .RDATA2    (RDATA[2]),
        .RDATA3    (RDATA[3]),
        .RDATA4    (RDATA[4]),
        .RDATA5    (RDATA[5]),
        .RDATA6    (RDATA[6]),
        .RDATA7    (RDATA[7]),
        .RDATA8    (RDATA[8]),
        .RDATA9    (RDATA[9]),
        .RDATA10    (RDATA[10]),
        .RDATA11    (RDATA[11]),
        .RDATA12    (RDATA[12]),
        .RDATA13    (RDATA[13]),
        .RDATA14    (RDATA[14]),
        .RDATA15    (RDATA[15]),
        .RDATA16    (RDATA[16]),
        .RDATA17    (RDATA[17]),
        .RDATA18    (RDATA[18]),
        .RDATA19    (RDATA[19]),
        .RDATA20    (RDATA[20]),
        .RDATA21    (RDATA[21]),
        .RDATA22    (RDATA[22]),
        .RDATA23    (RDATA[23]),
        .RDATA24    (RDATA[24]),
        .RDATA25    (RDATA[25]),
        .RDATA26    (RDATA[26]),
        .RDATA27    (RDATA[27]),
        .RDATA28    (RDATA[28]),
        .RDATA29    (RDATA[29]),
        .RDATA30    (RDATA[30]),
        .RDATA31    (RDATA[31])
    );

endmodule

module CUSTOM_INSTRUCTION_wrapper (
    input         ISSUE_READY,
    input         ISSUE_ACCEPT,
    output        ISSUE_VALID,
    output [31:0] ISSUE_INSTR,
    output [31:0] ISSUE_OPA,
    output [31:0] ISSUE_OPB,
    output [ 3:0] ISSUE_ID,
    
    input         RESULT_VALID,
    input  [ 3:0] RESULT_ID,
    input  [ 4:0] RESULT_RD,
    input  [31:0] RESULT
);

    CUSTOM_INSTRUCTION i_CUSTOM_INSTRUCTION (
        .ISSUE_READY    (ISSUE_READY),
        .ISSUE_ACCEPT   (ISSUE_ACCEPT),
        .ISSUE_VALID    (ISSUE_VALID),

        .ISSUE_INSTR0    (ISSUE_INSTR[0]),
        .ISSUE_INSTR1    (ISSUE_INSTR[1]),
        .ISSUE_INSTR2    (ISSUE_INSTR[2]),
        .ISSUE_INSTR3    (ISSUE_INSTR[3]),
        .ISSUE_INSTR4    (ISSUE_INSTR[4]),
        .ISSUE_INSTR5    (ISSUE_INSTR[5]),
        .ISSUE_INSTR6    (ISSUE_INSTR[6]),
        .ISSUE_INSTR7    (ISSUE_INSTR[7]),
        .ISSUE_INSTR8    (ISSUE_INSTR[8]),
        .ISSUE_INSTR9    (ISSUE_INSTR[9]),
        .ISSUE_INSTR10    (ISSUE_INSTR[10]),
        .ISSUE_INSTR11    (ISSUE_INSTR[11]),
        .ISSUE_INSTR12    (ISSUE_INSTR[12]),
        .ISSUE_INSTR13    (ISSUE_INSTR[13]),
        .ISSUE_INSTR14    (ISSUE_INSTR[14]),
        .ISSUE_INSTR15    (ISSUE_INSTR[15]),
        .ISSUE_INSTR16    (ISSUE_INSTR[16]),
        .ISSUE_INSTR17    (ISSUE_INSTR[17]),
        .ISSUE_INSTR18    (ISSUE_INSTR[18]),
        .ISSUE_INSTR19    (ISSUE_INSTR[19]),
        .ISSUE_INSTR20    (ISSUE_INSTR[20]),
        .ISSUE_INSTR21    (ISSUE_INSTR[21]),
        .ISSUE_INSTR22    (ISSUE_INSTR[22]),
        .ISSUE_INSTR23    (ISSUE_INSTR[23]),
        .ISSUE_INSTR24    (ISSUE_INSTR[24]),
        .ISSUE_INSTR25    (ISSUE_INSTR[25]),
        .ISSUE_INSTR26    (ISSUE_INSTR[26]),
        .ISSUE_INSTR27    (ISSUE_INSTR[27]),
        .ISSUE_INSTR28    (ISSUE_INSTR[28]),
        .ISSUE_INSTR29    (ISSUE_INSTR[29]),
        .ISSUE_INSTR30    (ISSUE_INSTR[30]),
        .ISSUE_INSTR31    (ISSUE_INSTR[31]),

        .ISSUE_OPA0    (ISSUE_OPA[0]),
        .ISSUE_OPA1    (ISSUE_OPA[1]),
        .ISSUE_OPA2    (ISSUE_OPA[2]),
        .ISSUE_OPA3    (ISSUE_OPA[3]),
        .ISSUE_OPA4    (ISSUE_OPA[4]),
        .ISSUE_OPA5    (ISSUE_OPA[5]),
        .ISSUE_OPA6    (ISSUE_OPA[6]),
        .ISSUE_OPA7    (ISSUE_OPA[7]),
        .ISSUE_OPA8    (ISSUE_OPA[8]),
        .ISSUE_OPA9    (ISSUE_OPA[9]),
        .ISSUE_OPA10    (ISSUE_OPA[10]),
        .ISSUE_OPA11    (ISSUE_OPA[11]),
        .ISSUE_OPA12    (ISSUE_OPA[12]),
        .ISSUE_OPA13    (ISSUE_OPA[13]),
        .ISSUE_OPA14    (ISSUE_OPA[14]),
        .ISSUE_OPA15    (ISSUE_OPA[15]),
        .ISSUE_OPA16    (ISSUE_OPA[16]),
        .ISSUE_OPA17    (ISSUE_OPA[17]),
        .ISSUE_OPA18    (ISSUE_OPA[18]),
        .ISSUE_OPA19    (ISSUE_OPA[19]),
        .ISSUE_OPA20    (ISSUE_OPA[20]),
        .ISSUE_OPA21    (ISSUE_OPA[21]),
        .ISSUE_OPA22    (ISSUE_OPA[22]),
        .ISSUE_OPA23    (ISSUE_OPA[23]),
        .ISSUE_OPA24    (ISSUE_OPA[24]),
        .ISSUE_OPA25    (ISSUE_OPA[25]),
        .ISSUE_OPA26    (ISSUE_OPA[26]),
        .ISSUE_OPA27    (ISSUE_OPA[27]),
        .ISSUE_OPA28    (ISSUE_OPA[28]),
        .ISSUE_OPA29    (ISSUE_OPA[29]),
        .ISSUE_OPA30    (ISSUE_OPA[30]),
        .ISSUE_OPA31    (ISSUE_OPA[31]),

        .ISSUE_OPB0    (ISSUE_OPB[0]),
        .ISSUE_OPB1    (ISSUE_OPB[1]),
        .ISSUE_OPB2    (ISSUE_OPB[2]),
        .ISSUE_OPB3    (ISSUE_OPB[3]),
        .ISSUE_OPB4    (ISSUE_OPB[4]),
        .ISSUE_OPB5    (ISSUE_OPB[5]),
        .ISSUE_OPB6    (ISSUE_OPB[6]),
        .ISSUE_OPB7    (ISSUE_OPB[7]),
        .ISSUE_OPB8    (ISSUE_OPB[8]),
        .ISSUE_OPB9    (ISSUE_OPB[9]),
        .ISSUE_OPB10    (ISSUE_OPB[10]),
        .ISSUE_OPB11    (ISSUE_OPB[11]),
        .ISSUE_OPB12    (ISSUE_OPB[12]),
        .ISSUE_OPB13    (ISSUE_OPB[13]),
        .ISSUE_OPB14    (ISSUE_OPB[14]),
        .ISSUE_OPB15    (ISSUE_OPB[15]),
        .ISSUE_OPB16    (ISSUE_OPB[16]),
        .ISSUE_OPB17    (ISSUE_OPB[17]),
        .ISSUE_OPB18    (ISSUE_OPB[18]),
        .ISSUE_OPB19    (ISSUE_OPB[19]),
        .ISSUE_OPB20    (ISSUE_OPB[20]),
        .ISSUE_OPB21    (ISSUE_OPB[21]),
        .ISSUE_OPB22    (ISSUE_OPB[22]),
        .ISSUE_OPB23    (ISSUE_OPB[23]),
        .ISSUE_OPB24    (ISSUE_OPB[24]),
        .ISSUE_OPB25    (ISSUE_OPB[25]),
        .ISSUE_OPB26    (ISSUE_OPB[26]),
        .ISSUE_OPB27    (ISSUE_OPB[27]),
        .ISSUE_OPB28    (ISSUE_OPB[28]),
        .ISSUE_OPB29    (ISSUE_OPB[29]),
        .ISSUE_OPB30    (ISSUE_OPB[30]),
        .ISSUE_OPB31    (ISSUE_OPB[31]),

        .ISSUE_ID0    (ISSUE_ID[0]),
        .ISSUE_ID1    (ISSUE_ID[1]),
        .ISSUE_ID2    (ISSUE_ID[2]),
        .ISSUE_ID3    (ISSUE_ID[3]),
        
        .RESULT_VALID   (RESULT_VALID),
        
        .RESULT_ID0    (RESULT_ID[0]),
        .RESULT_ID1    (RESULT_ID[1]),
        .RESULT_ID2    (RESULT_ID[2]),
        .RESULT_ID3    (RESULT_ID[3]),

        .RESULT_RD0    (RESULT_RD[0]),
        .RESULT_RD1    (RESULT_RD[1]),
        .RESULT_RD2    (RESULT_RD[2]),
        .RESULT_RD3    (RESULT_RD[3]),
        .RESULT_RD4    (RESULT_RD[4]),

        .RESULT0    (RESULT[0]),
        .RESULT1    (RESULT[1]),
        .RESULT2    (RESULT[2]),
        .RESULT3    (RESULT[3]),
        .RESULT4    (RESULT[4]),
        .RESULT5    (RESULT[5]),
        .RESULT6    (RESULT[6]),
        .RESULT7    (RESULT[7]),
        .RESULT8    (RESULT[8]),
        .RESULT9    (RESULT[9]),
        .RESULT10    (RESULT[10]),
        .RESULT11    (RESULT[11]),
        .RESULT12    (RESULT[12]),
        .RESULT13    (RESULT[13]),
        .RESULT14    (RESULT[14]),
        .RESULT15    (RESULT[15]),
        .RESULT16    (RESULT[16]),
        .RESULT17    (RESULT[17]),
        .RESULT18    (RESULT[18]),
        .RESULT19    (RESULT[19]),
        .RESULT20    (RESULT[20]),
        .RESULT21    (RESULT[21]),
        .RESULT22    (RESULT[22]),
        .RESULT23    (RESULT[23]),
        .RESULT24    (RESULT[24]),
        .RESULT25    (RESULT[25]),
        .RESULT26    (RESULT[26]),
        .RESULT27    (RESULT[27]),
        .RESULT28    (RESULT[28]),
        .RESULT29    (RESULT[29]),
        .RESULT30    (RESULT[30]),
        .RESULT31    (RESULT[31])
    );

endmodule

module IHP_BRAM_1024x16_wrapper (
    input  [ 9:0] A_ADDR,
    input  [16:0] A_BM,
    input  [16:0] A_DIN,
    input         A_WEN,
    input         A_MEN,
    input         A_REN,
    output [16:0] A_DOUT,

    input  [ 9:0] B_ADDR,
    input  [16:0] B_BM,
    input  [16:0] B_DIN,
    input         B_WEN,
    input         B_MEN,
    input         B_REN,
    output [16:0] B_DOUT
);
    IHP_BRAM_1024x16 i_IHP_BRAM_1024x16 (
        .A_ADDR0 (A_ADDR[0]),
        .A_ADDR1 (A_ADDR[1]),
        .A_ADDR2 (A_ADDR[2]),
        .A_ADDR3 (A_ADDR[3]),
        .A_ADDR4 (A_ADDR[4]),
        .A_ADDR5 (A_ADDR[5]),
        .A_ADDR6 (A_ADDR[6]),
        .A_ADDR7 (A_ADDR[7]),
        .A_ADDR8 (A_ADDR[8]),
        .A_ADDR9 (A_ADDR[9]),

        .A_BM0 (A_BM[0]),
        .A_BM1 (A_BM[1]),
        .A_BM2 (A_BM[2]),
        .A_BM3 (A_BM[3]),
        .A_BM4 (A_BM[4]),
        .A_BM5 (A_BM[5]),
        .A_BM6 (A_BM[6]),
        .A_BM7 (A_BM[7]),
        .A_BM8 (A_BM[8]),
        .A_BM9 (A_BM[9]),
        .A_BM10 (A_BM[10]),
        .A_BM11 (A_BM[11]),
        .A_BM12 (A_BM[12]),
        .A_BM13 (A_BM[13]),
        .A_BM14 (A_BM[14]),
        .A_BM15 (A_BM[15]),

        .A_DIN0 (A_DIN[0]),
        .A_DIN1 (A_DIN[1]),
        .A_DIN2 (A_DIN[2]),
        .A_DIN3 (A_DIN[3]),
        .A_DIN4 (A_DIN[4]),
        .A_DIN5 (A_DIN[5]),
        .A_DIN6 (A_DIN[6]),
        .A_DIN7 (A_DIN[7]),
        .A_DIN8 (A_DIN[8]),
        .A_DIN9 (A_DIN[9]),
        .A_DIN10 (A_DIN[10]),
        .A_DIN11 (A_DIN[11]),
        .A_DIN12 (A_DIN[12]),
        .A_DIN13 (A_DIN[13]),
        .A_DIN14 (A_DIN[14]),
        .A_DIN15 (A_DIN[15]),

        .A_WEN (A_WEN),
        .A_MEN (A_MEN),
        .A_REN (A_REN),

        .A_DOUT0 (A_DOUT[0]),
        .A_DOUT1 (A_DOUT[1]),
        .A_DOUT2 (A_DOUT[2]),
        .A_DOUT3 (A_DOUT[3]),
        .A_DOUT4 (A_DOUT[4]),
        .A_DOUT5 (A_DOUT[5]),
        .A_DOUT6 (A_DOUT[6]),
        .A_DOUT7 (A_DOUT[7]),
        .A_DOUT8 (A_DOUT[8]),
        .A_DOUT9 (A_DOUT[9]),
        .A_DOUT10 (A_DOUT[10]),
        .A_DOUT11 (A_DOUT[11]),
        .A_DOUT12 (A_DOUT[12]),
        .A_DOUT13 (A_DOUT[13]),
        .A_DOUT14 (A_DOUT[14]),
        .A_DOUT15 (A_DOUT[15]),

        .B_ADDR0 (B_ADDR[0]),
        .B_ADDR1 (B_ADDR[1]),
        .B_ADDR2 (B_ADDR[2]),
        .B_ADDR3 (B_ADDR[3]),
        .B_ADDR4 (B_ADDR[4]),
        .B_ADDR5 (B_ADDR[5]),
        .B_ADDR6 (B_ADDR[6]),
        .B_ADDR7 (B_ADDR[7]),
        .B_ADDR8 (B_ADDR[8]),
        .B_ADDR9 (B_ADDR[9]),

        .B_BM0 (B_BM[0]),
        .B_BM1 (B_BM[1]),
        .B_BM2 (B_BM[2]),
        .B_BM3 (B_BM[3]),
        .B_BM4 (B_BM[4]),
        .B_BM5 (B_BM[5]),
        .B_BM6 (B_BM[6]),
        .B_BM7 (B_BM[7]),
        .B_BM8 (B_BM[8]),
        .B_BM9 (B_BM[9]),
        .B_BM10 (B_BM[10]),
        .B_BM11 (B_BM[11]),
        .B_BM12 (B_BM[12]),
        .B_BM13 (B_BM[13]),
        .B_BM14 (B_BM[14]),
        .B_BM15 (B_BM[15]),

        .B_DIN0 (B_DIN[0]),
        .B_DIN1 (B_DIN[1]),
        .B_DIN2 (B_DIN[2]),
        .B_DIN3 (B_DIN[3]),
        .B_DIN4 (B_DIN[4]),
        .B_DIN5 (B_DIN[5]),
        .B_DIN6 (B_DIN[6]),
        .B_DIN7 (B_DIN[7]),
        .B_DIN8 (B_DIN[8]),
        .B_DIN9 (B_DIN[9]),
        .B_DIN10 (B_DIN[10]),
        .B_DIN11 (B_DIN[11]),
        .B_DIN12 (B_DIN[12]),
        .B_DIN13 (B_DIN[13]),
        .B_DIN14 (B_DIN[14]),
        .B_DIN15 (B_DIN[15]),

        .B_WEN (B_WEN),
        .B_MEN (B_MEN),
        .B_REN (B_REN),

        .B_DOUT0 (B_DOUT[0]),
        .B_DOUT1 (B_DOUT[1]),
        .B_DOUT2 (B_DOUT[2]),
        .B_DOUT3 (B_DOUT[3]),
        .B_DOUT4 (B_DOUT[4]),
        .B_DOUT5 (B_DOUT[5]),
        .B_DOUT6 (B_DOUT[6]),
        .B_DOUT7 (B_DOUT[7]),
        .B_DOUT8 (B_DOUT[8]),
        .B_DOUT9 (B_DOUT[9]),
        .B_DOUT10 (B_DOUT[10]),
        .B_DOUT11 (B_DOUT[11]),
        .B_DOUT12 (B_DOUT[12]),
        .B_DOUT13 (B_DOUT[13]),
        .B_DOUT14 (B_DOUT[14]),
        .B_DOUT15 (B_DOUT[15])
    );

endmodule

module IHP_SRAM_1024x32_wrapper (
    input  [ 9:0] A_ADDR,
    input  [31:0] A_BM,
    input  [31:0] A_DIN,
    input         A_WEN,
    input         A_MEN,
    input         A_REN,
    output [31:0] A_DOUT
);
    IHP_SRAM_1024x32 i_IHP_SRAM_1024x32 (
        .A_ADDR0 (A_ADDR[0]),
        .A_ADDR1 (A_ADDR[1]),
        .A_ADDR2 (A_ADDR[2]),
        .A_ADDR3 (A_ADDR[3]),
        .A_ADDR4 (A_ADDR[4]),
        .A_ADDR5 (A_ADDR[5]),
        .A_ADDR6 (A_ADDR[6]),
        .A_ADDR7 (A_ADDR[7]),
        .A_ADDR8 (A_ADDR[8]),
        .A_ADDR9 (A_ADDR[9]),

        .A_BM0 (A_BM[0]),
        .A_BM1 (A_BM[1]),
        .A_BM2 (A_BM[2]),
        .A_BM3 (A_BM[3]),
        .A_BM4 (A_BM[4]),
        .A_BM5 (A_BM[5]),
        .A_BM6 (A_BM[6]),
        .A_BM7 (A_BM[7]),
        .A_BM8 (A_BM[8]),
        .A_BM9 (A_BM[9]),
        .A_BM10 (A_BM[10]),
        .A_BM11 (A_BM[11]),
        .A_BM12 (A_BM[12]),
        .A_BM13 (A_BM[13]),
        .A_BM14 (A_BM[14]),
        .A_BM15 (A_BM[15]),
        .A_BM16 (A_BM[16]),
        .A_BM17 (A_BM[17]),
        .A_BM18 (A_BM[18]),
        .A_BM19 (A_BM[19]),
        .A_BM20 (A_BM[20]),
        .A_BM21 (A_BM[21]),
        .A_BM22 (A_BM[22]),
        .A_BM23 (A_BM[23]),
        .A_BM24 (A_BM[24]),
        .A_BM25 (A_BM[25]),
        .A_BM26 (A_BM[26]),
        .A_BM27 (A_BM[27]),
        .A_BM28 (A_BM[28]),
        .A_BM29 (A_BM[29]),
        .A_BM30 (A_BM[30]),
        .A_BM31 (A_BM[31]),

        .A_DIN0 (A_DIN[0]),
        .A_DIN1 (A_DIN[1]),
        .A_DIN2 (A_DIN[2]),
        .A_DIN3 (A_DIN[3]),
        .A_DIN4 (A_DIN[4]),
        .A_DIN5 (A_DIN[5]),
        .A_DIN6 (A_DIN[6]),
        .A_DIN7 (A_DIN[7]),
        .A_DIN8 (A_DIN[8]),
        .A_DIN9 (A_DIN[9]),
        .A_DIN10 (A_DIN[10]),
        .A_DIN11 (A_DIN[11]),
        .A_DIN12 (A_DIN[12]),
        .A_DIN13 (A_DIN[13]),
        .A_DIN14 (A_DIN[14]),
        .A_DIN15 (A_DIN[15]),
        .A_DIN16 (A_DIN[16]),
        .A_DIN17 (A_DIN[17]),
        .A_DIN18 (A_DIN[18]),
        .A_DIN19 (A_DIN[19]),
        .A_DIN20 (A_DIN[20]),
        .A_DIN21 (A_DIN[21]),
        .A_DIN22 (A_DIN[22]),
        .A_DIN23 (A_DIN[23]),
        .A_DIN24 (A_DIN[24]),
        .A_DIN25 (A_DIN[25]),
        .A_DIN26 (A_DIN[26]),
        .A_DIN27 (A_DIN[27]),
        .A_DIN28 (A_DIN[28]),
        .A_DIN29 (A_DIN[29]),
        .A_DIN30 (A_DIN[30]),
        .A_DIN31 (A_DIN[31]),

        .A_WEN (A_WEN),
        .A_MEN (A_MEN),
        .A_REN (A_REN),

        .A_DOUT0 (A_DOUT[0]),
        .A_DOUT1 (A_DOUT[1]),
        .A_DOUT2 (A_DOUT[2]),
        .A_DOUT3 (A_DOUT[3]),
        .A_DOUT4 (A_DOUT[4]),
        .A_DOUT5 (A_DOUT[5]),
        .A_DOUT6 (A_DOUT[6]),
        .A_DOUT7 (A_DOUT[7]),
        .A_DOUT8 (A_DOUT[8]),
        .A_DOUT9 (A_DOUT[9]),
        .A_DOUT10 (A_DOUT[10]),
        .A_DOUT11 (A_DOUT[11]),
        .A_DOUT12 (A_DOUT[12]),
        .A_DOUT13 (A_DOUT[13]),
        .A_DOUT14 (A_DOUT[14]),
        .A_DOUT15 (A_DOUT[15]),
        .A_DOUT16 (A_DOUT[16]),
        .A_DOUT17 (A_DOUT[17]),
        .A_DOUT18 (A_DOUT[18]),
        .A_DOUT19 (A_DOUT[19]),
        .A_DOUT20 (A_DOUT[20]),
        .A_DOUT21 (A_DOUT[21]),
        .A_DOUT22 (A_DOUT[22]),
        .A_DOUT23 (A_DOUT[23]),
        .A_DOUT24 (A_DOUT[24]),
        .A_DOUT25 (A_DOUT[25]),
        .A_DOUT26 (A_DOUT[26]),
        .A_DOUT27 (A_DOUT[27]),
        .A_DOUT28 (A_DOUT[28]),
        .A_DOUT29 (A_DOUT[29]),
        .A_DOUT30 (A_DOUT[30]),
        .A_DOUT31 (A_DOUT[31])
    );

endmodule

module WARMBOOT_wrapper (
    input  [3:0] SLOT,
    input        BOOT,
    output       RESET
);

    WARMBOOT i_WARMBOOT (
        .SLOT0  (SLOT[0]),
        .SLOT1  (SLOT[1]),
        .SLOT2  (SLOT[2]),
        .SLOT3  (SLOT[3]),
        .BOOT   (BOOT),
        .RESET  (RESET)
    );

endmodule

module CPU_IRQ_wrapper (
    input  [3:0] IRQ,
);

    CPU_IRQ i_CPU_IRQ (
        .IRQ0   (IRQ[0]),
        .IRQ1   (IRQ[1]),
        .IRQ2   (IRQ[2]),
        .IRQ3   (IRQ[3])
    );

endmodule

module MULADD_wrapper #(
    parameter A_reg=0,
    parameter B_reg=0,
    parameter C_reg=0,
    parameter signExtension=0,
    parameter ACC=0,
    parameter ACCout=0
) (
    input [7:0] A,
    input [7:0] B,
    input [19:0] C,
    input clr,
    
    output [19:0] Q
);

    MULADD #(
        .A_reg  (A_reg),
        .B_reg  (B_reg),
        .C_reg  (C_reg),
        
        .signExtension  (signExtension),
        .ACC            (ACC),
        .ACCout         (ACCout),
    ) muladd (
        .A0 (A[0]),
        .A1 (A[1]),
        .A2 (A[2]),
        .A3 (A[3]),
        .A4 (A[4]),
        .A5 (A[5]),
        .A6 (A[6]),
        .A7 (A[7]),

        .B0 (B[0]),
        .B1 (B[1]),
        .B2 (B[2]),
        .B3 (B[3]),
        .B4 (B[4]),
        .B5 (B[5]),
        .B6 (B[6]),
        .B7 (B[7]),
        
        .C0 (C[0]),
        .C1 (C[1]),
        .C2 (C[2]),
        .C3 (C[3]),
        .C4 (C[4]),
        .C5 (C[5]),
        .C6 (C[6]),
        .C7 (C[7]),
        .C8 (C[8]),
        .C9 (C[9]),
        .C10 (C[10]),
        .C11 (C[11]),
        .C12 (C[12]),
        .C13 (C[13]),
        .C14 (C[14]),
        .C15 (C[15]),
        .C16 (C[16]),
        .C17 (C[17]),
        .C18 (C[18]),
        .C19 (C[19]),
        
        .clr (clr),
        
        .Q0 (Q[0]),
        .Q1 (Q[1]),
        .Q2 (Q[2]),
        .Q3 (Q[3]),
        .Q4 (Q[4]),
        .Q5 (Q[5]),
        .Q6 (Q[6]),
        .Q7 (Q[7]),
        .Q8 (Q[8]),
        .Q9 (Q[9]),
        .Q10 (Q[10]),
        .Q11 (Q[11]),
        .Q12 (Q[12]),
        .Q13 (Q[13]),
        .Q14 (Q[14]),
        .Q15 (Q[15]),
        .Q16 (Q[16]),
        .Q17 (Q[17]),
        .Q18 (Q[18]),
        .Q19 (Q[19])
    );

endmodule
